magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 558 203
rect 31 -17 65 21
<< locali >>
rect 390 401 446 471
rect 342 367 446 401
rect 18 195 84 265
rect 120 199 205 265
rect 239 199 291 265
rect 342 199 387 367
rect 482 333 530 467
rect 421 299 530 333
rect 120 53 159 199
rect 239 132 273 199
rect 421 165 455 299
rect 489 199 537 265
rect 193 53 273 132
rect 307 131 530 165
rect 307 51 341 131
rect 481 59 530 131
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 19 299 85 527
rect 120 349 154 461
rect 188 383 240 527
rect 274 435 340 469
rect 274 349 308 435
rect 120 315 308 349
rect 19 17 85 161
rect 381 17 447 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 193 53 273 132 6 A1
port 1 nsew signal input
rlabel locali s 239 132 273 199 6 A1
port 1 nsew signal input
rlabel locali s 239 199 291 265 6 A1
port 1 nsew signal input
rlabel locali s 120 53 159 199 6 A2
port 2 nsew signal input
rlabel locali s 120 199 205 265 6 A2
port 2 nsew signal input
rlabel locali s 18 195 84 265 6 A3
port 3 nsew signal input
rlabel locali s 342 199 387 367 6 B1
port 4 nsew signal input
rlabel locali s 342 367 446 401 6 B1
port 4 nsew signal input
rlabel locali s 390 401 446 471 6 B1
port 4 nsew signal input
rlabel locali s 489 199 537 265 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 31 -17 65 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 558 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 481 59 530 131 6 Y
port 10 nsew signal output
rlabel locali s 307 51 341 131 6 Y
port 10 nsew signal output
rlabel locali s 307 131 530 165 6 Y
port 10 nsew signal output
rlabel locali s 421 165 455 299 6 Y
port 10 nsew signal output
rlabel locali s 421 299 530 333 6 Y
port 10 nsew signal output
rlabel locali s 482 333 530 467 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3719530
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3713376
<< end >>
