/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/cap_vpp_04p4x04p6_m1m2_noshield/sky130_fd_pr__cap_vpp_04p4x04p6_m1m2_noshield_o2.spice