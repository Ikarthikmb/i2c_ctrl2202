magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect 4335 3660 4829 3776
rect 3699 3502 4829 3660
rect 3699 3336 4943 3502
<< pwell >>
rect 577 923 991 1175
rect 293 97 1611 749
rect 299 70 1611 97
rect 299 -16 1646 70
<< mvnmos >>
rect 656 949 756 1149
rect 812 949 912 1149
rect 372 123 472 723
rect 528 123 628 723
rect 684 123 784 723
rect 840 123 940 723
rect 996 123 1096 723
rect 1152 123 1252 723
rect 1432 123 1532 723
<< mvpmos >>
rect 3818 3510 4018 3594
rect 4074 3510 4274 3594
rect 4454 3510 4554 3710
rect 4610 3510 4710 3710
<< mvndiff >>
rect 603 1131 656 1149
rect 603 1097 611 1131
rect 645 1097 656 1131
rect 603 1063 656 1097
rect 603 1029 611 1063
rect 645 1029 656 1063
rect 603 995 656 1029
rect 603 961 611 995
rect 645 961 656 995
rect 603 949 656 961
rect 756 1131 812 1149
rect 756 1097 767 1131
rect 801 1097 812 1131
rect 756 1063 812 1097
rect 756 1029 767 1063
rect 801 1029 812 1063
rect 756 995 812 1029
rect 756 961 767 995
rect 801 961 812 995
rect 756 949 812 961
rect 912 1131 965 1149
rect 912 1097 923 1131
rect 957 1097 965 1131
rect 912 1063 965 1097
rect 912 1029 923 1063
rect 957 1029 965 1063
rect 912 995 965 1029
rect 912 961 923 995
rect 957 961 965 995
rect 912 949 965 961
rect 319 645 372 723
rect 319 611 327 645
rect 361 611 372 645
rect 319 577 372 611
rect 319 543 327 577
rect 361 543 372 577
rect 319 509 372 543
rect 319 475 327 509
rect 361 475 372 509
rect 319 441 372 475
rect 319 407 327 441
rect 361 407 372 441
rect 319 373 372 407
rect 319 339 327 373
rect 361 339 372 373
rect 319 305 372 339
rect 319 271 327 305
rect 361 271 372 305
rect 319 237 372 271
rect 319 203 327 237
rect 361 203 372 237
rect 319 169 372 203
rect 319 135 327 169
rect 361 135 372 169
rect 319 123 372 135
rect 472 645 528 723
rect 472 611 483 645
rect 517 611 528 645
rect 472 577 528 611
rect 472 543 483 577
rect 517 543 528 577
rect 472 509 528 543
rect 472 475 483 509
rect 517 475 528 509
rect 472 441 528 475
rect 472 407 483 441
rect 517 407 528 441
rect 472 373 528 407
rect 472 339 483 373
rect 517 339 528 373
rect 472 305 528 339
rect 472 271 483 305
rect 517 271 528 305
rect 472 237 528 271
rect 472 203 483 237
rect 517 203 528 237
rect 472 169 528 203
rect 472 135 483 169
rect 517 135 528 169
rect 472 123 528 135
rect 628 645 684 723
rect 628 611 639 645
rect 673 611 684 645
rect 628 577 684 611
rect 628 543 639 577
rect 673 543 684 577
rect 628 509 684 543
rect 628 475 639 509
rect 673 475 684 509
rect 628 441 684 475
rect 628 407 639 441
rect 673 407 684 441
rect 628 373 684 407
rect 628 339 639 373
rect 673 339 684 373
rect 628 305 684 339
rect 628 271 639 305
rect 673 271 684 305
rect 628 237 684 271
rect 628 203 639 237
rect 673 203 684 237
rect 628 169 684 203
rect 628 135 639 169
rect 673 135 684 169
rect 628 123 684 135
rect 784 645 840 723
rect 784 611 795 645
rect 829 611 840 645
rect 784 577 840 611
rect 784 543 795 577
rect 829 543 840 577
rect 784 509 840 543
rect 784 475 795 509
rect 829 475 840 509
rect 784 441 840 475
rect 784 407 795 441
rect 829 407 840 441
rect 784 373 840 407
rect 784 339 795 373
rect 829 339 840 373
rect 784 305 840 339
rect 784 271 795 305
rect 829 271 840 305
rect 784 237 840 271
rect 784 203 795 237
rect 829 203 840 237
rect 784 169 840 203
rect 784 135 795 169
rect 829 135 840 169
rect 784 123 840 135
rect 940 645 996 723
rect 940 611 951 645
rect 985 611 996 645
rect 940 577 996 611
rect 940 543 951 577
rect 985 543 996 577
rect 940 509 996 543
rect 940 475 951 509
rect 985 475 996 509
rect 940 441 996 475
rect 940 407 951 441
rect 985 407 996 441
rect 940 373 996 407
rect 940 339 951 373
rect 985 339 996 373
rect 940 305 996 339
rect 940 271 951 305
rect 985 271 996 305
rect 940 237 996 271
rect 940 203 951 237
rect 985 203 996 237
rect 940 169 996 203
rect 940 135 951 169
rect 985 135 996 169
rect 940 123 996 135
rect 1096 645 1152 723
rect 1096 611 1107 645
rect 1141 611 1152 645
rect 1096 577 1152 611
rect 1096 543 1107 577
rect 1141 543 1152 577
rect 1096 509 1152 543
rect 1096 475 1107 509
rect 1141 475 1152 509
rect 1096 441 1152 475
rect 1096 407 1107 441
rect 1141 407 1152 441
rect 1096 373 1152 407
rect 1096 339 1107 373
rect 1141 339 1152 373
rect 1096 305 1152 339
rect 1096 271 1107 305
rect 1141 271 1152 305
rect 1096 237 1152 271
rect 1096 203 1107 237
rect 1141 203 1152 237
rect 1096 169 1152 203
rect 1096 135 1107 169
rect 1141 135 1152 169
rect 1096 123 1152 135
rect 1252 645 1305 723
rect 1252 611 1263 645
rect 1297 611 1305 645
rect 1252 577 1305 611
rect 1252 543 1263 577
rect 1297 543 1305 577
rect 1252 509 1305 543
rect 1252 475 1263 509
rect 1297 475 1305 509
rect 1252 441 1305 475
rect 1252 407 1263 441
rect 1297 407 1305 441
rect 1252 373 1305 407
rect 1252 339 1263 373
rect 1297 339 1305 373
rect 1252 305 1305 339
rect 1252 271 1263 305
rect 1297 271 1305 305
rect 1252 237 1305 271
rect 1252 203 1263 237
rect 1297 203 1305 237
rect 1252 169 1305 203
rect 1252 135 1263 169
rect 1297 135 1305 169
rect 1252 123 1305 135
rect 1379 645 1432 723
rect 1379 611 1387 645
rect 1421 611 1432 645
rect 1379 577 1432 611
rect 1379 543 1387 577
rect 1421 543 1432 577
rect 1379 509 1432 543
rect 1379 475 1387 509
rect 1421 475 1432 509
rect 1379 441 1432 475
rect 1379 407 1387 441
rect 1421 407 1432 441
rect 1379 373 1432 407
rect 1379 339 1387 373
rect 1421 339 1432 373
rect 1379 305 1432 339
rect 1379 271 1387 305
rect 1421 271 1432 305
rect 1379 237 1432 271
rect 1379 203 1387 237
rect 1421 203 1432 237
rect 1379 169 1432 203
rect 1379 135 1387 169
rect 1421 135 1432 169
rect 1379 123 1432 135
rect 1532 645 1585 723
rect 1532 611 1543 645
rect 1577 611 1585 645
rect 1532 577 1585 611
rect 1532 543 1543 577
rect 1577 543 1585 577
rect 1532 509 1585 543
rect 1532 475 1543 509
rect 1577 475 1585 509
rect 1532 441 1585 475
rect 1532 407 1543 441
rect 1577 407 1585 441
rect 1532 373 1585 407
rect 1532 339 1543 373
rect 1577 339 1585 373
rect 1532 305 1585 339
rect 1532 271 1543 305
rect 1577 271 1585 305
rect 1532 237 1585 271
rect 1532 203 1543 237
rect 1577 203 1585 237
rect 1532 169 1585 203
rect 1532 135 1543 169
rect 1577 135 1585 169
rect 1532 123 1585 135
<< mvpdiff >>
rect 4401 3698 4454 3710
rect 4401 3664 4409 3698
rect 4443 3664 4454 3698
rect 4401 3630 4454 3664
rect 4401 3596 4409 3630
rect 4443 3596 4454 3630
rect 3765 3556 3818 3594
rect 3765 3522 3773 3556
rect 3807 3522 3818 3556
rect 3765 3510 3818 3522
rect 4018 3556 4074 3594
rect 4018 3522 4029 3556
rect 4063 3522 4074 3556
rect 4018 3510 4074 3522
rect 4274 3556 4327 3594
rect 4274 3522 4285 3556
rect 4319 3522 4327 3556
rect 4274 3510 4327 3522
rect 4401 3562 4454 3596
rect 4401 3528 4409 3562
rect 4443 3528 4454 3562
rect 4401 3510 4454 3528
rect 4554 3698 4610 3710
rect 4554 3664 4565 3698
rect 4599 3664 4610 3698
rect 4554 3630 4610 3664
rect 4554 3596 4565 3630
rect 4599 3596 4610 3630
rect 4554 3562 4610 3596
rect 4554 3528 4565 3562
rect 4599 3528 4610 3562
rect 4554 3510 4610 3528
rect 4710 3698 4763 3710
rect 4710 3664 4721 3698
rect 4755 3664 4763 3698
rect 4710 3630 4763 3664
rect 4710 3596 4721 3630
rect 4755 3596 4763 3630
rect 4710 3562 4763 3596
rect 4710 3528 4721 3562
rect 4755 3528 4763 3562
rect 4710 3510 4763 3528
<< mvndiffc >>
rect 611 1097 645 1131
rect 611 1029 645 1063
rect 611 961 645 995
rect 767 1097 801 1131
rect 767 1029 801 1063
rect 767 961 801 995
rect 923 1097 957 1131
rect 923 1029 957 1063
rect 923 961 957 995
rect 327 611 361 645
rect 327 543 361 577
rect 327 475 361 509
rect 327 407 361 441
rect 327 339 361 373
rect 327 271 361 305
rect 327 203 361 237
rect 327 135 361 169
rect 483 611 517 645
rect 483 543 517 577
rect 483 475 517 509
rect 483 407 517 441
rect 483 339 517 373
rect 483 271 517 305
rect 483 203 517 237
rect 483 135 517 169
rect 639 611 673 645
rect 639 543 673 577
rect 639 475 673 509
rect 639 407 673 441
rect 639 339 673 373
rect 639 271 673 305
rect 639 203 673 237
rect 639 135 673 169
rect 795 611 829 645
rect 795 543 829 577
rect 795 475 829 509
rect 795 407 829 441
rect 795 339 829 373
rect 795 271 829 305
rect 795 203 829 237
rect 795 135 829 169
rect 951 611 985 645
rect 951 543 985 577
rect 951 475 985 509
rect 951 407 985 441
rect 951 339 985 373
rect 951 271 985 305
rect 951 203 985 237
rect 951 135 985 169
rect 1107 611 1141 645
rect 1107 543 1141 577
rect 1107 475 1141 509
rect 1107 407 1141 441
rect 1107 339 1141 373
rect 1107 271 1141 305
rect 1107 203 1141 237
rect 1107 135 1141 169
rect 1263 611 1297 645
rect 1263 543 1297 577
rect 1263 475 1297 509
rect 1263 407 1297 441
rect 1263 339 1297 373
rect 1263 271 1297 305
rect 1263 203 1297 237
rect 1263 135 1297 169
rect 1387 611 1421 645
rect 1387 543 1421 577
rect 1387 475 1421 509
rect 1387 407 1421 441
rect 1387 339 1421 373
rect 1387 271 1421 305
rect 1387 203 1421 237
rect 1387 135 1421 169
rect 1543 611 1577 645
rect 1543 543 1577 577
rect 1543 475 1577 509
rect 1543 407 1577 441
rect 1543 339 1577 373
rect 1543 271 1577 305
rect 1543 203 1577 237
rect 1543 135 1577 169
<< mvpdiffc >>
rect 4409 3664 4443 3698
rect 4409 3596 4443 3630
rect 3773 3522 3807 3556
rect 4029 3522 4063 3556
rect 4285 3522 4319 3556
rect 4409 3528 4443 3562
rect 4565 3664 4599 3698
rect 4565 3596 4599 3630
rect 4565 3528 4599 3562
rect 4721 3664 4755 3698
rect 4721 3596 4755 3630
rect 4721 3528 4755 3562
<< psubdiff >>
rect 325 10 349 44
rect 383 10 421 44
rect 455 10 493 44
rect 527 10 565 44
rect 599 10 637 44
rect 671 10 709 44
rect 743 10 781 44
rect 815 10 852 44
rect 886 10 923 44
rect 957 10 994 44
rect 1028 10 1065 44
rect 1099 10 1136 44
rect 1170 10 1207 44
rect 1241 10 1278 44
rect 1312 10 1349 44
rect 1383 10 1420 44
rect 1454 10 1491 44
rect 1525 10 1562 44
rect 1596 10 1620 44
<< mvnsubdiff >>
rect 3765 3402 3799 3436
rect 3833 3402 3871 3436
rect 3905 3402 3943 3436
rect 3977 3402 4015 3436
rect 4049 3402 4087 3436
rect 4121 3402 4159 3436
rect 4193 3402 4231 3436
rect 4265 3402 4303 3436
rect 4337 3402 4375 3436
rect 4409 3402 4447 3436
rect 4481 3402 4519 3436
rect 4553 3402 4591 3436
rect 4625 3402 4663 3436
rect 4697 3402 4736 3436
rect 4770 3402 4809 3436
rect 4843 3402 4877 3436
<< psubdiffcont >>
rect 349 10 383 44
rect 421 10 455 44
rect 493 10 527 44
rect 565 10 599 44
rect 637 10 671 44
rect 709 10 743 44
rect 781 10 815 44
rect 852 10 886 44
rect 923 10 957 44
rect 994 10 1028 44
rect 1065 10 1099 44
rect 1136 10 1170 44
rect 1207 10 1241 44
rect 1278 10 1312 44
rect 1349 10 1383 44
rect 1420 10 1454 44
rect 1491 10 1525 44
rect 1562 10 1596 44
<< mvnsubdiffcont >>
rect 3799 3402 3833 3436
rect 3871 3402 3905 3436
rect 3943 3402 3977 3436
rect 4015 3402 4049 3436
rect 4087 3402 4121 3436
rect 4159 3402 4193 3436
rect 4231 3402 4265 3436
rect 4303 3402 4337 3436
rect 4375 3402 4409 3436
rect 4447 3402 4481 3436
rect 4519 3402 4553 3436
rect 4591 3402 4625 3436
rect 4663 3402 4697 3436
rect 4736 3402 4770 3436
rect 4809 3402 4843 3436
<< poly >>
rect 4454 3792 4710 3808
rect 4454 3758 4470 3792
rect 4504 3758 4565 3792
rect 4599 3758 4660 3792
rect 4694 3758 4710 3792
rect 4454 3742 4710 3758
rect 4454 3710 4554 3742
rect 4610 3710 4710 3742
rect 3818 3676 4018 3692
rect 3818 3642 3834 3676
rect 3868 3642 3968 3676
rect 4002 3642 4018 3676
rect 3818 3594 4018 3642
rect 4074 3676 4274 3692
rect 4074 3642 4090 3676
rect 4124 3642 4224 3676
rect 4258 3642 4274 3676
rect 4074 3594 4274 3642
rect 3818 3478 4018 3510
rect 4074 3478 4274 3510
rect 4454 3478 4554 3510
rect 4610 3478 4710 3510
rect 656 1149 756 1175
rect 812 1149 912 1175
rect 656 923 756 949
rect 622 907 756 923
rect 622 873 638 907
rect 672 873 706 907
rect 740 873 756 907
rect 622 857 756 873
rect 812 923 912 949
rect 812 907 946 923
rect 812 873 828 907
rect 862 873 896 907
rect 930 873 946 907
rect 812 857 946 873
rect 372 799 784 815
rect 372 765 388 799
rect 422 765 458 799
rect 492 765 527 799
rect 561 765 596 799
rect 630 765 665 799
rect 699 765 734 799
rect 768 765 784 799
rect 372 749 784 765
rect 372 723 472 749
rect 528 723 628 749
rect 684 723 784 749
rect 840 799 1252 815
rect 840 765 856 799
rect 890 765 925 799
rect 959 765 994 799
rect 1028 765 1063 799
rect 1097 765 1132 799
rect 1166 765 1202 799
rect 1236 765 1252 799
rect 840 749 1252 765
rect 840 723 940 749
rect 996 723 1096 749
rect 1152 723 1252 749
rect 1432 799 1566 815
rect 1432 765 1448 799
rect 1482 765 1516 799
rect 1550 765 1566 799
rect 1432 749 1566 765
rect 1432 723 1532 749
rect 372 97 472 123
rect 528 97 628 123
rect 684 97 784 123
rect 840 97 940 123
rect 996 97 1096 123
rect 1152 97 1252 123
rect 1432 97 1532 123
<< polycont >>
rect 4470 3758 4504 3792
rect 4565 3758 4599 3792
rect 4660 3758 4694 3792
rect 3834 3642 3868 3676
rect 3968 3642 4002 3676
rect 4090 3642 4124 3676
rect 4224 3642 4258 3676
rect 638 873 672 907
rect 706 873 740 907
rect 828 873 862 907
rect 896 873 930 907
rect 388 765 422 799
rect 458 765 492 799
rect 527 765 561 799
rect 596 765 630 799
rect 665 765 699 799
rect 734 765 768 799
rect 856 765 890 799
rect 925 765 959 799
rect 994 765 1028 799
rect 1063 765 1097 799
rect 1132 765 1166 799
rect 1202 765 1236 799
rect 1448 765 1482 799
rect 1516 765 1550 799
<< locali >>
rect 3818 3792 4710 3838
rect 3818 3758 4470 3792
rect 4504 3758 4565 3792
rect 4599 3758 4660 3792
rect 4694 3758 4710 3792
rect 3818 3750 4375 3758
rect 3818 3716 3833 3750
rect 3867 3716 3905 3750
rect 3939 3723 4375 3750
rect 3939 3716 4018 3723
rect 3818 3676 4018 3716
rect 3708 3642 3746 3676
rect 3818 3642 3834 3676
rect 3868 3642 3968 3676
rect 4002 3642 4018 3676
rect 4074 3642 4090 3676
rect 4137 3642 4175 3676
rect 4209 3642 4224 3676
rect 4258 3642 4274 3676
rect 3674 3572 3784 3642
rect 3674 3556 3807 3572
rect 3674 3522 3773 3556
rect 3674 3506 3807 3522
rect 4308 3572 4375 3723
rect 4029 3508 4063 3522
rect 4285 3556 4375 3572
rect 4319 3522 4375 3556
rect 4285 3506 4375 3522
rect 4409 3698 4443 3714
rect 4565 3712 4599 3714
rect 4562 3698 4600 3712
rect 4562 3678 4565 3698
rect 4409 3630 4443 3664
rect 4409 3580 4443 3596
rect 4409 3508 4443 3528
rect 4599 3678 4600 3698
rect 4721 3698 4755 3714
rect 4565 3630 4599 3664
rect 4565 3562 4599 3596
rect 4565 3512 4599 3528
rect 4721 3630 4755 3664
rect 4721 3580 4755 3596
rect 4721 3508 4755 3528
rect 3765 3402 3766 3436
rect 3833 3402 3838 3436
rect 3905 3402 3910 3436
rect 3977 3402 3982 3436
rect 4049 3402 4054 3436
rect 4121 3402 4126 3436
rect 4193 3402 4198 3436
rect 4265 3402 4271 3436
rect 4337 3402 4344 3436
rect 4409 3402 4417 3436
rect 4481 3402 4490 3436
rect 4553 3402 4563 3436
rect 4625 3402 4636 3436
rect 4697 3402 4709 3436
rect 4770 3402 4782 3436
rect 4843 3402 4877 3436
rect 611 1131 645 1147
rect 611 1087 645 1097
rect 611 1015 645 1029
rect 611 945 645 961
rect 767 1145 801 1147
rect 767 1131 771 1145
rect 801 1097 805 1111
rect 767 1073 805 1097
rect 767 1063 771 1073
rect 923 1131 957 1147
rect 923 1078 957 1097
rect 923 1063 924 1078
rect 767 995 801 1029
rect 767 945 801 961
rect 957 1029 958 1044
rect 923 1006 958 1029
rect 923 995 924 1006
rect 923 945 957 961
rect 622 901 638 907
rect 672 901 706 907
rect 622 873 633 901
rect 672 873 705 901
rect 740 873 756 907
rect 812 901 828 907
rect 812 873 826 901
rect 862 873 896 907
rect 930 901 946 907
rect 932 873 946 901
rect 667 867 705 873
rect 860 867 898 873
rect 372 765 388 799
rect 422 765 458 799
rect 492 765 510 799
rect 561 765 582 799
rect 630 765 665 799
rect 699 765 734 799
rect 768 765 784 799
rect 840 765 856 799
rect 897 765 925 799
rect 969 765 994 799
rect 1028 765 1063 799
rect 1097 765 1132 799
rect 1166 765 1202 799
rect 1236 765 1252 799
rect 1432 765 1448 799
rect 1482 765 1516 799
rect 1577 765 1615 799
rect 327 645 361 661
rect 327 577 361 611
rect 325 543 327 570
rect 483 645 517 661
rect 483 577 517 611
rect 361 543 363 570
rect 325 536 363 543
rect 639 645 673 661
rect 639 577 673 611
rect 327 509 361 536
rect 483 509 517 543
rect 635 543 639 570
rect 795 645 829 661
rect 795 577 829 611
rect 635 536 673 543
rect 951 645 985 661
rect 951 577 985 611
rect 639 509 673 536
rect 327 441 361 475
rect 517 475 522 496
rect 484 462 522 475
rect 795 509 829 543
rect 949 543 951 570
rect 1107 645 1141 661
rect 1107 577 1141 611
rect 985 543 987 570
rect 949 536 987 543
rect 1263 645 1297 661
rect 1263 577 1297 611
rect 327 373 361 407
rect 327 305 361 339
rect 327 237 361 271
rect 327 169 361 203
rect 327 119 361 135
rect 483 441 517 462
rect 483 373 517 407
rect 483 305 517 339
rect 483 237 517 271
rect 483 169 517 203
rect 483 119 517 135
rect 639 441 673 475
rect 794 475 795 496
rect 951 509 985 536
rect 829 475 832 496
rect 794 462 832 475
rect 1107 509 1141 543
rect 1260 543 1263 570
rect 1387 645 1421 661
rect 1387 577 1421 611
rect 1297 543 1298 570
rect 1260 536 1298 543
rect 1263 509 1297 536
rect 639 373 673 407
rect 639 305 673 339
rect 639 237 673 271
rect 639 169 673 203
rect 639 119 673 135
rect 795 441 829 462
rect 795 373 829 407
rect 795 305 829 339
rect 795 237 829 271
rect 795 169 829 203
rect 795 119 829 135
rect 951 441 985 475
rect 1075 475 1107 496
rect 1075 462 1113 475
rect 1387 509 1421 543
rect 951 373 985 407
rect 951 305 985 339
rect 951 237 985 271
rect 951 169 985 203
rect 951 119 985 135
rect 1107 441 1141 462
rect 1107 373 1141 407
rect 1107 305 1141 339
rect 1107 237 1141 271
rect 1107 169 1141 203
rect 1107 119 1141 135
rect 1263 441 1297 475
rect 1385 475 1387 496
rect 1543 645 1577 661
rect 1543 577 1577 611
rect 1543 509 1577 543
rect 1421 475 1423 496
rect 1385 462 1423 475
rect 1263 373 1297 407
rect 1263 305 1297 339
rect 1263 237 1297 271
rect 1263 169 1297 203
rect 1263 119 1297 135
rect 1387 441 1421 462
rect 1387 373 1421 407
rect 1387 305 1421 339
rect 1387 237 1421 271
rect 1387 169 1421 203
rect 1387 119 1421 135
rect 1543 441 1577 475
rect 1543 373 1577 407
rect 1543 305 1577 339
rect 1543 237 1577 271
rect 1543 189 1577 203
rect 1543 117 1577 135
rect 325 10 346 44
rect 383 10 419 44
rect 455 10 492 44
rect 527 10 565 44
rect 599 10 637 44
rect 672 10 709 44
rect 744 10 781 44
rect 816 10 852 44
rect 888 10 923 44
rect 960 10 994 44
rect 1032 10 1065 44
rect 1104 10 1136 44
rect 1176 10 1207 44
rect 1248 10 1278 44
rect 1320 10 1349 44
rect 1392 10 1420 44
rect 1464 10 1491 44
rect 1536 10 1562 44
rect 1596 10 1620 44
<< viali >>
rect 3833 3716 3867 3750
rect 3905 3716 3939 3750
rect 3674 3642 3708 3676
rect 3746 3642 3780 3676
rect 4103 3642 4124 3676
rect 4124 3642 4137 3676
rect 4175 3642 4209 3676
rect 4029 3556 4063 3580
rect 4029 3546 4063 3556
rect 4029 3474 4063 3508
rect 4528 3678 4562 3712
rect 4409 3562 4443 3580
rect 4409 3546 4443 3562
rect 4600 3678 4634 3712
rect 4721 3562 4755 3580
rect 4721 3546 4755 3562
rect 4409 3474 4443 3508
rect 4721 3474 4755 3508
rect 3766 3402 3799 3436
rect 3799 3402 3800 3436
rect 3838 3402 3871 3436
rect 3871 3402 3872 3436
rect 3910 3402 3943 3436
rect 3943 3402 3944 3436
rect 3982 3402 4015 3436
rect 4015 3402 4016 3436
rect 4054 3402 4087 3436
rect 4087 3402 4088 3436
rect 4126 3402 4159 3436
rect 4159 3402 4160 3436
rect 4198 3402 4231 3436
rect 4231 3402 4232 3436
rect 4271 3402 4303 3436
rect 4303 3402 4305 3436
rect 4344 3402 4375 3436
rect 4375 3402 4378 3436
rect 4417 3402 4447 3436
rect 4447 3402 4451 3436
rect 4490 3402 4519 3436
rect 4519 3402 4524 3436
rect 4563 3402 4591 3436
rect 4591 3402 4597 3436
rect 4636 3402 4663 3436
rect 4663 3402 4670 3436
rect 4709 3402 4736 3436
rect 4736 3402 4743 3436
rect 4782 3402 4809 3436
rect 4809 3402 4816 3436
rect 611 1063 645 1087
rect 611 1053 645 1063
rect 611 995 645 1015
rect 611 981 645 995
rect 771 1131 805 1145
rect 771 1111 801 1131
rect 801 1111 805 1131
rect 771 1063 805 1073
rect 771 1039 801 1063
rect 801 1039 805 1063
rect 924 1063 958 1078
rect 924 1044 957 1063
rect 957 1044 958 1063
rect 924 995 958 1006
rect 924 972 957 995
rect 957 972 958 995
rect 633 873 638 901
rect 638 873 667 901
rect 705 873 706 901
rect 706 873 739 901
rect 826 873 828 901
rect 828 873 860 901
rect 898 873 930 901
rect 930 873 932 901
rect 633 867 667 873
rect 705 867 739 873
rect 826 867 860 873
rect 898 867 932 873
rect 510 765 527 799
rect 527 765 544 799
rect 582 765 596 799
rect 596 765 616 799
rect 863 765 890 799
rect 890 765 897 799
rect 935 765 959 799
rect 959 765 969 799
rect 1543 765 1550 799
rect 1550 765 1577 799
rect 1615 765 1649 799
rect 291 536 325 570
rect 363 536 397 570
rect 601 536 635 570
rect 673 536 707 570
rect 450 475 483 496
rect 483 475 484 496
rect 450 462 484 475
rect 522 462 556 496
rect 915 536 949 570
rect 987 536 1021 570
rect 760 462 794 496
rect 832 462 866 496
rect 1226 536 1260 570
rect 1298 536 1332 570
rect 1041 462 1075 496
rect 1113 475 1141 496
rect 1141 475 1147 496
rect 1113 462 1147 475
rect 1351 462 1385 496
rect 1423 462 1457 496
rect 1543 169 1577 189
rect 1543 155 1577 169
rect 1543 83 1577 117
rect 346 10 349 44
rect 349 10 380 44
rect 419 10 421 44
rect 421 10 453 44
rect 492 10 493 44
rect 493 10 526 44
rect 565 10 599 44
rect 638 10 671 44
rect 671 10 672 44
rect 710 10 743 44
rect 743 10 744 44
rect 782 10 815 44
rect 815 10 816 44
rect 854 10 886 44
rect 886 10 888 44
rect 926 10 957 44
rect 957 10 960 44
rect 998 10 1028 44
rect 1028 10 1032 44
rect 1070 10 1099 44
rect 1099 10 1104 44
rect 1142 10 1170 44
rect 1170 10 1176 44
rect 1214 10 1241 44
rect 1241 10 1248 44
rect 1286 10 1312 44
rect 1312 10 1320 44
rect 1358 10 1383 44
rect 1383 10 1392 44
rect 1430 10 1454 44
rect 1454 10 1464 44
rect 1502 10 1525 44
rect 1525 10 1536 44
<< metal1 >>
rect 3224 3816 4646 3822
rect 3276 3788 4646 3816
rect 3224 3752 3276 3764
tri 4469 3756 4501 3788 ne
rect 4501 3756 4646 3788
tri 3815 3750 3821 3756 se
rect 3821 3750 3951 3756
tri 3809 3744 3815 3750 se
rect 3815 3744 3833 3750
rect 3224 3694 3276 3700
rect 3320 3738 3833 3744
rect 3372 3716 3833 3738
rect 3867 3716 3905 3750
rect 3939 3716 3951 3750
tri 4501 3741 4516 3756 ne
rect 3372 3710 3951 3716
rect 4516 3712 4646 3756
rect 3320 3674 3372 3686
rect 3320 3616 3372 3622
rect 3409 3676 4221 3682
rect 3461 3642 3674 3676
rect 3708 3642 3746 3676
rect 3780 3642 4103 3676
rect 4137 3642 4175 3676
rect 4209 3642 4221 3676
rect 4516 3678 4528 3712
rect 4562 3678 4600 3712
rect 4634 3678 4646 3712
rect 4516 3672 4646 3678
rect 3461 3636 4221 3642
rect 3409 3612 3461 3624
rect 3409 3554 3461 3560
rect 4023 3580 4761 3592
rect 4023 3546 4029 3580
rect 4063 3546 4409 3580
rect 4443 3546 4721 3580
rect 4755 3546 4761 3580
rect 4023 3508 4761 3546
rect 4023 3474 4029 3508
rect 4063 3474 4409 3508
rect 4443 3474 4721 3508
rect 4755 3474 4761 3508
rect 4023 3442 4761 3474
rect 3754 3436 4828 3442
rect 3754 3402 3766 3436
rect 3800 3402 3838 3436
rect 3872 3402 3910 3436
rect 3944 3402 3982 3436
rect 4016 3402 4054 3436
rect 4088 3402 4126 3436
rect 4160 3402 4198 3436
rect 4232 3402 4271 3436
rect 4305 3402 4344 3436
rect 4378 3402 4417 3436
rect 4451 3402 4490 3436
rect 4524 3402 4563 3436
rect 4597 3402 4636 3436
rect 4670 3402 4709 3436
rect 4743 3402 4782 3436
rect 4816 3402 4828 3436
rect 3754 3396 4828 3402
rect 3224 1760 3276 1766
tri 3190 1666 3224 1700 se
rect 3224 1696 3276 1708
rect 605 1644 3224 1666
rect 605 1638 3276 1644
rect 3320 1700 3372 1706
tri 3318 1638 3320 1640 se
rect 3320 1638 3372 1648
rect 605 1087 651 1638
tri 651 1605 684 1638 nw
tri 3286 1606 3318 1638 se
rect 3318 1636 3372 1638
rect 3318 1606 3320 1636
rect 923 1584 3320 1606
rect 923 1578 3372 1584
rect 605 1053 611 1087
rect 645 1053 651 1087
rect 605 1015 651 1053
rect 765 1145 811 1157
rect 765 1111 771 1145
rect 805 1111 811 1145
rect 765 1073 811 1111
rect 923 1090 957 1578
tri 957 1544 991 1578 nw
tri 3309 1374 3333 1398 se
rect 3333 1374 3339 1398
rect 1191 1346 3339 1374
rect 3391 1346 3403 1398
rect 3455 1346 3461 1398
rect 765 1039 771 1073
rect 805 1039 811 1073
rect 765 1027 811 1039
rect 918 1078 964 1090
rect 918 1044 924 1078
rect 958 1044 964 1078
rect 605 981 611 1015
rect 645 981 651 1015
rect 918 1006 964 1044
rect 918 994 924 1006
rect 605 969 651 981
rect 697 972 924 994
rect 958 972 964 1006
rect 697 960 964 972
rect 697 907 751 960
tri 751 922 789 960 nw
rect 621 901 751 907
rect 621 867 633 901
rect 667 867 705 901
rect 739 867 751 901
rect 621 861 751 867
rect 814 901 944 907
rect 814 867 826 901
rect 860 867 898 901
rect 932 867 944 901
rect 814 861 944 867
rect 498 799 628 805
rect 498 765 510 799
rect 544 765 582 799
rect 616 765 628 799
rect 498 759 628 765
rect 705 576 751 861
rect 851 799 981 805
rect 851 765 863 799
rect 897 765 935 799
rect 969 765 981 799
rect 851 759 981 765
rect 1191 576 1237 1346
tri 1237 1312 1271 1346 nw
rect 1531 799 1661 805
rect 1531 765 1543 799
rect 1577 765 1615 799
rect 1649 765 1661 799
rect 1531 759 1661 765
rect 279 570 751 576
rect 279 536 291 570
rect 325 536 363 570
rect 397 536 601 570
rect 635 536 673 570
rect 707 536 751 570
rect 279 530 751 536
rect 903 570 1344 576
rect 903 536 915 570
rect 949 536 987 570
rect 1021 536 1226 570
rect 1260 536 1298 570
rect 1332 536 1344 570
rect 903 530 1344 536
rect 438 496 1469 502
rect 438 462 450 496
rect 484 462 522 496
rect 556 462 760 496
rect 794 462 832 496
rect 866 462 1041 496
rect 1075 462 1113 496
rect 1147 462 1351 496
rect 1385 462 1423 496
rect 1457 462 1469 496
rect 438 456 1469 462
rect 334 189 1583 201
rect 334 155 1543 189
rect 1577 155 1583 189
rect 334 117 1583 155
rect 334 83 1543 117
rect 1577 83 1583 117
rect 334 44 1583 83
rect 334 10 346 44
rect 380 10 419 44
rect 453 10 492 44
rect 526 10 565 44
rect 599 10 638 44
rect 672 10 710 44
rect 744 10 782 44
rect 816 10 854 44
rect 888 10 926 44
rect 960 10 998 44
rect 1032 10 1070 44
rect 1104 10 1142 44
rect 1176 10 1214 44
rect 1248 10 1286 44
rect 1320 10 1358 44
rect 1392 10 1430 44
rect 1464 10 1502 44
rect 1536 10 1583 44
rect 334 4 1583 10
<< via1 >>
rect 3224 3764 3276 3816
rect 3224 3700 3276 3752
rect 3320 3686 3372 3738
rect 3320 3622 3372 3674
rect 3409 3624 3461 3676
rect 3409 3560 3461 3612
rect 3224 1708 3276 1760
rect 3224 1644 3276 1696
rect 3320 1648 3372 1700
rect 3320 1584 3372 1636
rect 3339 1346 3391 1398
rect 3403 1346 3455 1398
<< metal2 >>
rect 3224 3816 3276 3822
rect 3224 3752 3276 3764
rect 3224 1760 3276 3700
rect 3224 1696 3276 1708
rect 3224 1638 3276 1644
rect 3320 3738 3372 3744
rect 3320 3674 3372 3686
rect 3320 1700 3372 3622
rect 3320 1636 3372 1648
rect 3320 1578 3372 1584
rect 3409 3676 3461 3682
rect 3409 3612 3461 3624
tri 3375 1398 3409 1432 se
rect 3409 1398 3461 3560
rect 3333 1346 3339 1398
rect 3391 1346 3403 1398
rect 3455 1346 3461 1398
use sky130_fd_pr__nfet_01v8__example_55959141808568  sky130_fd_pr__nfet_01v8__example_55959141808568_0
timestamp 1644511149
transform -1 0 1532 0 1 123
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_0
timestamp 1644511149
transform -1 0 784 0 1 123
box -28 0 440 267
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_1
timestamp 1644511149
transform 1 0 840 0 1 123
box -28 0 440 267
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_0
timestamp 1644511149
transform 1 0 812 0 1 949
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_1
timestamp 1644511149
transform -1 0 756 0 1 949
box -28 0 128 97
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_0
timestamp 1644511149
transform -1 0 4018 0 1 3510
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_1
timestamp 1644511149
transform 1 0 4074 0 1 3510
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808567  sky130_fd_pr__pfet_01v8__example_55959141808567_0
timestamp 1644511149
transform -1 0 4710 0 -1 3710
box -28 0 284 97
<< labels >>
flabel metal1 s 4568 3462 4596 3490 3 FreeSans 520 180 0 0 VPWR_HV
port 1 nsew
flabel metal1 s 894 771 922 799 3 FreeSans 520 0 0 0 IN
port 2 nsew
flabel metal1 s 1452 126 1480 154 3 FreeSans 520 0 0 0 VGND
port 3 nsew
flabel metal1 s 848 866 876 894 3 FreeSans 520 0 0 0 RST_H
port 4 nsew
flabel metal1 s 1583 768 1611 796 3 FreeSans 520 0 0 0 HLD_H_N
port 5 nsew
flabel metal1 s 552 770 580 798 3 FreeSans 520 0 0 0 IN_B
port 6 nsew
flabel metal1 s 614 1026 642 1054 3 FreeSans 520 0 0 0 OUT_H_N
port 7 nsew
flabel metal1 s 776 1123 804 1151 3 FreeSans 520 0 0 0 VGND
port 3 nsew
<< properties >>
string GDS_END 8176984
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8157906
<< end >>
