magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -66 377 162 897
<< pwell >>
rect -26 -43 122 43
<< obsli1 >>
rect 0 797 31 831
rect 65 797 96 831
rect 0 -17 31 17
rect 65 -17 96 17
<< obsli1c >>
rect 31 797 65 831
rect 31 -17 65 17
<< metal1 >>
rect 0 831 96 837
rect 0 797 31 831
rect 65 797 96 831
rect 0 791 96 797
rect 0 689 96 763
rect 0 51 96 125
rect 0 17 96 23
rect 0 -17 31 17
rect 65 -17 96 17
rect 0 -23 96 -17
<< labels >>
rlabel metal1 s 0 51 96 125 6 VGND
port 1 nsew ground bidirectional
rlabel metal1 s 0 -23 96 23 8 VNB
port 2 nsew ground bidirectional
rlabel pwell s -26 -43 122 43 8 VNB
port 2 nsew ground bidirectional
rlabel metal1 s 0 791 96 837 6 VPB
port 3 nsew power bidirectional
rlabel nwell s -66 377 162 897 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 689 96 763 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 96 814
string LEFclass CORE SPACER
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 1242032
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 1239652
<< end >>
