magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 1 21 551 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 155 47 185 177
rect 351 47 381 177
rect 423 47 453 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 351 297 381 497
rect 435 297 465 497
<< ndiff >>
rect 27 119 79 177
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 47 155 177
rect 185 101 237 177
rect 185 67 195 101
rect 229 67 237 101
rect 185 47 237 67
rect 299 101 351 177
rect 299 67 307 101
rect 341 67 351 101
rect 299 47 351 67
rect 381 47 423 177
rect 453 97 525 177
rect 453 63 477 97
rect 511 63 525 97
rect 453 47 525 63
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 409 163 497
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 485 245 497
rect 193 451 203 485
rect 237 451 245 485
rect 193 297 245 451
rect 299 485 351 497
rect 299 451 307 485
rect 341 451 351 485
rect 299 297 351 451
rect 381 417 435 497
rect 381 383 391 417
rect 425 383 435 417
rect 381 297 435 383
rect 465 489 525 497
rect 465 455 475 489
rect 509 455 525 489
rect 465 421 525 455
rect 465 387 475 421
rect 509 387 525 421
rect 465 297 525 387
<< ndiffc >>
rect 35 85 69 119
rect 195 67 229 101
rect 307 67 341 101
rect 477 63 511 97
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 375 153 409
rect 203 451 237 485
rect 307 451 341 485
rect 391 383 425 417
rect 475 455 509 489
rect 475 387 509 421
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 351 497 381 523
rect 435 497 465 523
rect 79 265 109 297
rect 163 265 193 297
rect 351 265 381 297
rect 435 265 465 297
rect 55 249 109 265
rect 55 215 65 249
rect 99 215 109 249
rect 55 199 109 215
rect 79 177 109 199
rect 155 249 213 265
rect 155 215 169 249
rect 203 215 213 249
rect 155 199 213 215
rect 304 249 381 265
rect 304 215 318 249
rect 352 215 381 249
rect 304 199 381 215
rect 155 177 185 199
rect 351 177 381 199
rect 423 249 477 265
rect 423 215 433 249
rect 467 215 477 249
rect 423 199 477 215
rect 423 177 453 199
rect 79 21 109 47
rect 155 21 185 47
rect 351 21 381 47
rect 423 21 453 47
<< polycont >>
rect 65 215 99 249
rect 169 215 203 249
rect 318 215 352 249
rect 433 215 467 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 19 485 253 493
rect 19 451 35 485
rect 69 459 203 485
rect 69 451 85 459
rect 187 451 203 459
rect 237 451 253 485
rect 287 485 362 527
rect 287 451 307 485
rect 341 451 362 485
rect 472 489 525 527
rect 472 455 475 489
rect 509 455 525 489
rect 19 417 85 451
rect 19 383 35 417
rect 69 383 85 417
rect 19 349 85 383
rect 119 417 165 425
rect 391 417 425 433
rect 119 409 242 417
rect 153 407 242 409
rect 153 383 391 407
rect 153 375 425 383
rect 119 367 425 375
rect 472 421 525 455
rect 472 387 475 421
rect 509 387 525 421
rect 472 371 525 387
rect 119 359 295 367
rect 19 315 35 349
rect 69 325 85 349
rect 323 325 535 333
rect 69 315 535 325
rect 19 299 535 315
rect 19 289 368 299
rect 25 249 115 255
rect 25 215 65 249
rect 99 215 115 249
rect 153 249 248 255
rect 153 215 169 249
rect 203 215 248 249
rect 25 153 115 215
rect 198 135 248 215
rect 298 249 368 255
rect 298 215 318 249
rect 352 215 368 249
rect 402 249 467 265
rect 402 215 433 249
rect 298 135 340 215
rect 402 199 467 215
rect 501 165 535 299
rect 389 131 535 165
rect 19 85 35 119
rect 69 85 109 119
rect 389 101 425 131
rect 19 17 109 85
rect 164 67 195 101
rect 229 67 307 101
rect 341 67 425 101
rect 164 51 425 67
rect 461 63 477 97
rect 511 63 527 97
rect 461 17 527 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 214 153 248 187 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 306 153 340 187 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 402 221 436 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 306 221 340 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 306 289 340 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a22oi_1
rlabel metal1 s 0 -48 552 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 4085032
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4079418
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 13.800 0.000 
<< end >>
