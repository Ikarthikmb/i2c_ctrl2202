magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< obsli1 >>
rect 0 4544 4498 4610
rect 0 66 28 4516
rect 56 94 84 4544
rect 112 66 140 4516
rect 168 94 196 4544
rect 224 66 252 4516
rect 280 94 308 4544
rect 336 66 364 4516
rect 392 94 420 4544
rect 448 66 476 4516
rect 504 94 532 4544
rect 560 66 588 4516
rect 616 94 644 4544
rect 672 66 700 4516
rect 728 94 756 4544
rect 784 66 812 4516
rect 840 94 868 4544
rect 896 66 924 4516
rect 952 94 980 4544
rect 1008 66 1036 4516
rect 1064 94 1092 4544
rect 1120 66 1148 4516
rect 1176 94 1204 4544
rect 1232 66 1260 4516
rect 1288 94 1316 4544
rect 1344 66 1372 4516
rect 1400 94 1428 4544
rect 1456 66 1484 4516
rect 1512 94 1540 4544
rect 1568 66 1596 4516
rect 1624 94 1652 4544
rect 1680 66 1708 4516
rect 1736 94 1764 4544
rect 1792 66 1820 4516
rect 1848 94 1876 4544
rect 1904 66 1932 4516
rect 1960 94 1988 4544
rect 2016 66 2044 4516
rect 2072 94 2100 4544
rect 2128 66 2156 4516
rect 2184 94 2212 4544
rect 2240 66 2268 4516
rect 2296 94 2324 4544
rect 2352 66 2380 4516
rect 2408 94 2436 4544
rect 2464 66 2492 4516
rect 2520 94 2548 4544
rect 2576 66 2604 4516
rect 2632 94 2660 4544
rect 2688 66 2716 4516
rect 2744 94 2772 4544
rect 2800 66 2828 4516
rect 2856 94 2884 4544
rect 2912 66 2940 4516
rect 2968 94 2996 4544
rect 3024 66 3052 4516
rect 3080 94 3108 4544
rect 3136 66 3164 4516
rect 3192 94 3220 4544
rect 3248 66 3276 4516
rect 3304 94 3332 4544
rect 3360 66 3388 4516
rect 3416 94 3444 4544
rect 3472 66 3500 4516
rect 3528 94 3556 4544
rect 3584 66 3612 4516
rect 3640 94 3668 4544
rect 3696 66 3724 4516
rect 3752 94 3780 4544
rect 3808 66 3836 4516
rect 3864 94 3892 4544
rect 3920 66 3948 4516
rect 3976 94 4004 4544
rect 4032 66 4060 4516
rect 4088 94 4116 4544
rect 4144 66 4172 4516
rect 4200 94 4228 4544
rect 4256 66 4284 4516
rect 4312 94 4340 4544
rect 4368 66 4396 4516
rect 4424 94 4498 4544
rect 0 0 4498 66
<< obsm1 >>
rect 0 4544 4498 4610
rect 0 94 28 4544
rect 56 66 84 4516
rect 112 94 140 4544
rect 168 66 196 4516
rect 224 94 252 4544
rect 280 66 308 4516
rect 336 94 364 4544
rect 392 66 420 4516
rect 448 94 476 4544
rect 504 66 532 4516
rect 560 94 588 4544
rect 616 66 644 4516
rect 672 94 700 4544
rect 728 66 756 4516
rect 784 94 812 4544
rect 840 66 868 4516
rect 896 94 924 4544
rect 952 66 980 4516
rect 1008 94 1036 4544
rect 1064 66 1092 4516
rect 1120 94 1148 4544
rect 1176 66 1204 4516
rect 1232 94 1260 4544
rect 1288 66 1316 4516
rect 1344 94 1372 4544
rect 1400 66 1428 4516
rect 1456 94 1484 4544
rect 1512 66 1540 4516
rect 1568 94 1596 4544
rect 1624 66 1652 4516
rect 1680 94 1708 4544
rect 1736 66 1764 4516
rect 1792 94 1820 4544
rect 1848 66 1876 4516
rect 1904 94 1932 4544
rect 1960 66 1988 4516
rect 2016 94 2044 4544
rect 2072 66 2100 4516
rect 2128 94 2156 4544
rect 2184 66 2212 4516
rect 2240 94 2268 4544
rect 2296 66 2324 4516
rect 2352 94 2380 4544
rect 2408 66 2436 4516
rect 2464 94 2492 4544
rect 2520 66 2548 4516
rect 2576 94 2604 4544
rect 2632 66 2660 4516
rect 2688 94 2716 4544
rect 2744 66 2772 4516
rect 2800 94 2828 4544
rect 2856 66 2884 4516
rect 2912 94 2940 4544
rect 2968 66 2996 4516
rect 3024 94 3052 4544
rect 3080 66 3108 4516
rect 3136 94 3164 4544
rect 3192 66 3220 4516
rect 3248 94 3276 4544
rect 3304 66 3332 4516
rect 3360 94 3388 4544
rect 3416 66 3444 4516
rect 3472 94 3500 4544
rect 3528 66 3556 4516
rect 3584 94 3612 4544
rect 3640 66 3668 4516
rect 3696 94 3724 4544
rect 3752 66 3780 4516
rect 3808 94 3836 4544
rect 3864 66 3892 4516
rect 3920 94 3948 4544
rect 3976 66 4004 4516
rect 4032 94 4060 4544
rect 4088 66 4116 4516
rect 4144 94 4172 4544
rect 4200 66 4228 4516
rect 4256 94 4284 4544
rect 4312 66 4340 4516
rect 4368 94 4396 4544
rect 4424 66 4498 4516
rect 0 0 4498 66
<< obsm2 >>
rect 0 66 28 4610
rect 56 4544 196 4610
rect 56 94 84 4544
rect 112 66 140 4516
rect 0 0 140 66
rect 168 0 196 4544
rect 224 66 252 4610
rect 280 4544 420 4610
rect 280 94 308 4544
rect 336 66 364 4516
rect 224 0 364 66
rect 392 0 420 4544
rect 448 66 476 4610
rect 504 4544 644 4610
rect 504 94 532 4544
rect 560 66 588 4516
rect 448 0 588 66
rect 616 0 644 4544
rect 672 66 700 4610
rect 728 4544 868 4610
rect 728 94 756 4544
rect 784 66 812 4516
rect 672 0 812 66
rect 840 0 868 4544
rect 896 66 924 4610
rect 952 4544 1092 4610
rect 952 94 980 4544
rect 1008 66 1036 4516
rect 896 0 1036 66
rect 1064 0 1092 4544
rect 1120 66 1148 4610
rect 1176 4544 1316 4610
rect 1176 94 1204 4544
rect 1232 66 1260 4516
rect 1120 0 1260 66
rect 1288 0 1316 4544
rect 1344 66 1372 4610
rect 1400 4544 1540 4610
rect 1400 94 1428 4544
rect 1456 66 1484 4516
rect 1344 0 1484 66
rect 1512 0 1540 4544
rect 1568 66 1596 4610
rect 1624 4544 1764 4610
rect 1624 94 1652 4544
rect 1680 66 1708 4516
rect 1568 0 1708 66
rect 1736 0 1764 4544
rect 1792 66 1820 4610
rect 1848 4544 1988 4610
rect 1848 94 1876 4544
rect 1904 66 1932 4516
rect 1792 0 1932 66
rect 1960 0 1988 4544
rect 2016 66 2044 4610
rect 2072 4544 2212 4610
rect 2072 94 2100 4544
rect 2128 66 2156 4516
rect 2016 0 2156 66
rect 2184 0 2212 4544
rect 2240 66 2268 4610
rect 2296 4544 2436 4610
rect 2296 94 2324 4544
rect 2352 66 2380 4516
rect 2240 0 2380 66
rect 2408 0 2436 4544
rect 2464 66 2492 4610
rect 2520 4544 2660 4610
rect 2520 94 2548 4544
rect 2576 66 2604 4516
rect 2464 0 2604 66
rect 2632 0 2660 4544
rect 2688 66 2716 4610
rect 2744 4544 2884 4610
rect 2744 94 2772 4544
rect 2800 66 2828 4516
rect 2688 0 2828 66
rect 2856 0 2884 4544
rect 2912 66 2940 4610
rect 2968 4544 3108 4610
rect 2968 94 2996 4544
rect 3024 66 3052 4516
rect 2912 0 3052 66
rect 3080 0 3108 4544
rect 3136 66 3164 4610
rect 3192 4544 3332 4610
rect 3192 94 3220 4544
rect 3248 66 3276 4516
rect 3136 0 3276 66
rect 3304 0 3332 4544
rect 3360 66 3388 4610
rect 3416 4544 3556 4610
rect 3416 94 3444 4544
rect 3472 66 3500 4516
rect 3360 0 3500 66
rect 3528 0 3556 4544
rect 3584 66 3612 4610
rect 3640 4544 3780 4610
rect 3640 94 3668 4544
rect 3696 66 3724 4516
rect 3584 0 3724 66
rect 3752 0 3780 4544
rect 3808 66 3836 4610
rect 3864 4544 4004 4610
rect 3864 94 3892 4544
rect 3920 66 3948 4516
rect 3808 0 3948 66
rect 3976 0 4004 4544
rect 4032 66 4060 4610
rect 4088 4544 4498 4610
rect 4088 94 4116 4544
rect 4144 66 4172 4516
rect 4032 0 4172 66
rect 4200 0 4228 4544
rect 4256 66 4284 4516
rect 4312 94 4340 4544
rect 4368 66 4396 4516
rect 4424 94 4498 4544
rect 4256 0 4498 66
<< obsm3 >>
rect 0 4544 4498 4610
rect 0 126 60 4544
rect 120 66 180 4484
rect 240 126 300 4544
rect 360 66 420 4484
rect 480 126 540 4544
rect 600 66 660 4484
rect 720 126 780 4544
rect 840 66 900 4484
rect 960 126 1020 4544
rect 1080 66 1140 4484
rect 1200 126 1260 4544
rect 1320 66 1380 4484
rect 1440 126 1500 4544
rect 1560 66 1620 4484
rect 1680 126 1740 4544
rect 1800 66 1860 4484
rect 1920 126 1980 4544
rect 2040 66 2100 4484
rect 2160 126 2220 4544
rect 2280 66 2340 4484
rect 2400 126 2460 4544
rect 2520 66 2580 4484
rect 2640 126 2700 4544
rect 2760 66 2820 4484
rect 2880 126 2940 4544
rect 3000 66 3060 4484
rect 3120 126 3180 4544
rect 3240 66 3300 4484
rect 3360 126 3420 4544
rect 3480 66 3540 4484
rect 3600 126 3660 4544
rect 3720 66 3780 4484
rect 3840 126 3900 4544
rect 3960 66 4020 4484
rect 4080 126 4140 4544
rect 4200 66 4260 4484
rect 4320 126 4498 4544
rect 0 0 4498 66
<< obsm4 >>
rect 0 4544 4498 4610
rect 0 66 60 4484
rect 120 4299 420 4544
rect 120 126 180 4299
rect 240 311 300 4239
rect 360 371 420 4299
rect 480 311 540 4484
rect 240 66 540 311
rect 600 126 660 4544
rect 720 66 780 4484
rect 840 126 900 4544
rect 960 66 1020 4484
rect 1080 126 1140 4544
rect 1200 66 1260 4484
rect 1320 126 1380 4544
rect 1440 66 1500 4484
rect 1560 4299 1860 4544
rect 1560 126 1620 4299
rect 1680 311 1740 4239
rect 1800 371 1860 4299
rect 1920 311 1980 4484
rect 1680 66 1980 311
rect 2040 126 2100 4544
rect 2160 66 2220 4484
rect 2280 126 2340 4544
rect 2400 66 2460 4484
rect 2520 126 2580 4544
rect 2640 66 2700 4484
rect 2760 126 2820 4544
rect 2880 66 2940 4484
rect 3000 4299 3300 4544
rect 3000 126 3060 4299
rect 3120 311 3180 4239
rect 3240 371 3300 4299
rect 3360 311 3420 4484
rect 3120 66 3420 311
rect 3480 126 3540 4544
rect 3600 66 3660 4484
rect 3720 126 3780 4544
rect 3840 66 3900 4484
rect 3960 126 4020 4544
rect 4080 66 4140 4484
rect 4200 126 4260 4544
rect 4320 66 4498 4484
rect 0 0 4498 66
<< obsm5 >>
rect 0 4275 4498 4610
rect 0 655 320 4275
rect 640 335 960 3955
rect 1280 655 1600 4275
rect 1920 335 2240 3955
rect 2560 655 2880 4275
rect 3200 335 3520 3955
rect 3840 655 4498 4275
rect 0 0 4498 335
<< properties >>
string FIXED_BBOX 0 0 4498 4610
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1231494
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 1168706
<< end >>
