magic
tech sky130B
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_0
timestamp 1644511149
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_1
timestamp 1644511149
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_2
timestamp 1644511149
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_3
timestamp 1644511149
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_4
timestamp 1644511149
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_5
timestamp 1644511149
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808202  sky130_fd_pr__hvdfl1sd2__example_55959141808202_6
timestamp 1644511149
transform 1 0 1036 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808194  sky130_fd_pr__hvdfl1sd__example_55959141808194_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808194  sky130_fd_pr__hvdfl1sd__example_55959141808194_1
timestamp 1644511149
transform 1 0 1192 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 1220 471 1220 471 0 FreeSans 300 0 0 0 S
flabel comment s 1064 471 1064 471 0 FreeSans 300 0 0 0 D
flabel comment s 908 471 908 471 0 FreeSans 300 0 0 0 S
flabel comment s 752 471 752 471 0 FreeSans 300 0 0 0 D
flabel comment s 596 471 596 471 0 FreeSans 300 0 0 0 S
flabel comment s 440 471 440 471 0 FreeSans 300 0 0 0 D
flabel comment s 284 471 284 471 0 FreeSans 300 0 0 0 S
flabel comment s 128 471 128 471 0 FreeSans 300 0 0 0 D
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7340162
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7335482
<< end >>
