magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 31 21 762 203
rect 31 17 63 21
rect 29 -17 63 17
<< locali >>
rect 17 199 83 257
rect 299 265 363 341
rect 185 215 251 257
rect 287 215 363 265
rect 401 257 476 341
rect 678 375 811 493
rect 401 215 498 257
rect 536 215 626 257
rect 761 181 811 375
rect 674 53 811 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 48 325 108 493
rect 147 359 197 527
rect 315 409 476 493
rect 231 375 544 409
rect 231 325 265 375
rect 48 291 265 325
rect 117 165 151 291
rect 510 325 544 375
rect 578 359 644 527
rect 510 291 694 325
rect 660 257 694 291
rect 660 215 727 257
rect 49 129 151 165
rect 232 147 572 181
rect 232 129 309 147
rect 49 51 115 129
rect 149 61 386 95
rect 438 17 472 111
rect 506 54 572 147
rect 606 17 640 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 536 215 626 257 6 A1
port 1 nsew signal input
rlabel locali s 401 215 498 257 6 A2
port 2 nsew signal input
rlabel locali s 401 257 476 341 6 A2
port 2 nsew signal input
rlabel locali s 185 215 251 257 6 B1
port 3 nsew signal input
rlabel locali s 287 215 363 265 6 B2
port 4 nsew signal input
rlabel locali s 299 265 363 341 6 B2
port 4 nsew signal input
rlabel locali s 17 199 83 257 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 7 nsew ground bidirectional
rlabel pwell s 31 17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 31 21 762 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 674 53 811 181 6 X
port 10 nsew signal output
rlabel locali s 761 181 811 375 6 X
port 10 nsew signal output
rlabel locali s 678 375 811 493 6 X
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 810304
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 803074
<< end >>
