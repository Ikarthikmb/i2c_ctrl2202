magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< pwell >>
rect -13 -26 73 8246
rect 258 570 279 619
rect 467 -26 553 8246
<< locali >>
rect 13 0 47 8220
rect 493 0 527 8220
<< metal1 >>
rect 14 8213 526 8220
rect 14 8161 44 8213
rect 96 8161 284 8213
rect 336 8161 364 8213
rect 416 8161 444 8213
rect 496 8161 526 8213
rect 14 8154 526 8161
rect 14 126 46 8154
rect 74 66 106 8094
rect 134 126 166 8154
rect 194 66 226 8094
rect 254 126 286 8154
rect 314 66 346 8094
rect 374 126 406 8154
rect 434 66 466 8094
rect 494 126 526 8154
rect 60 59 480 66
rect 60 7 84 59
rect 136 7 164 59
rect 216 7 244 59
rect 296 7 324 59
rect 376 7 404 59
rect 456 7 480 59
rect 60 0 480 7
<< via1 >>
rect 44 8161 96 8213
rect 284 8161 336 8213
rect 364 8161 416 8213
rect 444 8161 496 8213
rect 84 7 136 59
rect 164 7 216 59
rect 244 7 296 59
rect 324 7 376 59
rect 404 7 456 59
<< metal2 >>
rect 14 8215 166 8220
rect 14 8159 42 8215
rect 98 8159 166 8215
rect 14 8154 166 8159
rect 14 126 46 8154
rect 74 66 106 8094
rect 134 126 166 8154
rect 194 66 226 8220
rect 254 8215 526 8220
rect 254 8159 282 8215
rect 338 8159 362 8215
rect 418 8159 442 8215
rect 498 8159 526 8215
rect 254 8154 526 8159
rect 254 126 286 8154
rect 314 66 346 8094
rect 374 126 406 8154
rect 434 66 466 8094
rect 494 126 526 8154
rect 60 61 480 66
rect 60 5 82 61
rect 138 5 162 61
rect 218 5 242 61
rect 298 5 322 61
rect 378 5 402 61
rect 458 5 480 61
rect 60 0 480 5
<< via2 >>
rect 42 8213 98 8215
rect 42 8161 44 8213
rect 44 8161 96 8213
rect 96 8161 98 8213
rect 42 8159 98 8161
rect 282 8213 338 8215
rect 282 8161 284 8213
rect 284 8161 336 8213
rect 336 8161 338 8213
rect 282 8159 338 8161
rect 362 8213 418 8215
rect 362 8161 364 8213
rect 364 8161 416 8213
rect 416 8161 418 8213
rect 362 8159 418 8161
rect 442 8213 498 8215
rect 442 8161 444 8213
rect 444 8161 496 8213
rect 496 8161 498 8213
rect 442 8159 498 8161
rect 82 59 138 61
rect 82 7 84 59
rect 84 7 136 59
rect 136 7 138 59
rect 82 5 138 7
rect 162 59 218 61
rect 162 7 164 59
rect 164 7 216 59
rect 216 7 218 59
rect 162 5 218 7
rect 242 59 298 61
rect 242 7 244 59
rect 244 7 296 59
rect 296 7 298 59
rect 242 5 298 7
rect 322 59 378 61
rect 322 7 324 59
rect 324 7 376 59
rect 376 7 378 59
rect 322 5 378 7
rect 402 59 458 61
rect 402 7 404 59
rect 404 7 456 59
rect 456 7 458 59
rect 402 5 458 7
<< metal3 >>
rect 0 8219 540 8220
rect 0 8155 38 8219
rect 102 8155 118 8219
rect 182 8155 198 8219
rect 262 8155 278 8219
rect 342 8155 358 8219
rect 422 8155 438 8219
rect 502 8155 540 8219
rect 0 8154 540 8155
rect 0 126 60 8154
rect 120 66 180 8094
rect 240 126 300 8154
rect 360 66 420 8094
rect 480 126 540 8154
rect 60 65 480 66
rect 60 1 78 65
rect 142 1 158 65
rect 222 1 238 65
rect 302 1 318 65
rect 382 1 398 65
rect 462 1 480 65
rect 60 0 480 1
<< via3 >>
rect 38 8215 102 8219
rect 38 8159 42 8215
rect 42 8159 98 8215
rect 98 8159 102 8215
rect 38 8155 102 8159
rect 118 8155 182 8219
rect 198 8155 262 8219
rect 278 8215 342 8219
rect 278 8159 282 8215
rect 282 8159 338 8215
rect 338 8159 342 8215
rect 278 8155 342 8159
rect 358 8215 422 8219
rect 358 8159 362 8215
rect 362 8159 418 8215
rect 418 8159 422 8215
rect 358 8155 422 8159
rect 438 8215 502 8219
rect 438 8159 442 8215
rect 442 8159 498 8215
rect 498 8159 502 8215
rect 438 8155 502 8159
rect 78 61 142 65
rect 78 5 82 61
rect 82 5 138 61
rect 138 5 142 61
rect 78 1 142 5
rect 158 61 222 65
rect 158 5 162 61
rect 162 5 218 61
rect 218 5 222 61
rect 158 1 222 5
rect 238 61 302 65
rect 238 5 242 61
rect 242 5 298 61
rect 298 5 302 61
rect 238 1 302 5
rect 318 61 382 65
rect 318 5 322 61
rect 322 5 378 61
rect 378 5 382 61
rect 318 1 382 5
rect 398 61 462 65
rect 398 5 402 61
rect 402 5 458 61
rect 458 5 462 61
rect 398 1 462 5
<< metal4 >>
rect 0 8219 540 8220
rect 0 8155 38 8219
rect 102 8155 118 8219
rect 182 8155 198 8219
rect 262 8155 278 8219
rect 342 8155 358 8219
rect 422 8155 438 8219
rect 502 8155 540 8219
rect 0 8154 540 8155
rect 0 126 60 8154
rect 120 66 180 8094
rect 240 126 300 8154
rect 360 66 420 8094
rect 480 126 540 8154
rect 60 65 480 66
rect 60 1 78 65
rect 142 1 158 65
rect 222 1 238 65
rect 302 1 318 65
rect 382 1 398 65
rect 462 1 480 65
rect 60 0 480 1
<< labels >>
flabel metal2 s 141 268 160 288 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 288 19 324 55 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 258 570 279 619 0 FreeSans 400 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 30676
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 13348
string path 0.750 40.470 0.750 0.330 
<< end >>
