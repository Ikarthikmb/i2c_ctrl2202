magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -36 679 1916 1471
<< pwell >>
rect 1744 25 1846 159
<< psubdiff >>
rect 1770 109 1820 133
rect 1770 75 1778 109
rect 1812 75 1820 109
rect 1770 51 1820 75
<< nsubdiff >>
rect 1770 1339 1820 1363
rect 1770 1305 1778 1339
rect 1812 1305 1820 1339
rect 1770 1281 1820 1305
<< psubdiffcont >>
rect 1778 75 1812 109
<< nsubdiffcont >>
rect 1778 1305 1812 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 1880 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 490 1130 524 1397
rect 706 1130 740 1397
rect 922 1130 956 1397
rect 1138 1130 1172 1397
rect 1354 1130 1388 1397
rect 1570 1130 1604 1397
rect 1778 1339 1812 1397
rect 1778 1289 1812 1305
rect 64 724 98 740
rect 64 674 98 690
rect 920 724 954 1096
rect 920 690 971 724
rect 920 318 954 690
rect 62 17 96 218
rect 274 17 308 218
rect 490 17 524 218
rect 706 17 740 218
rect 922 17 956 218
rect 1138 17 1172 218
rect 1354 17 1388 218
rect 1570 17 1604 218
rect 1778 109 1812 125
rect 1778 17 1812 75
rect 0 -17 1880 17
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1644511149
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1644511149
transform 1 0 1770 0 1 1281
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1644511149
transform 1 0 1770 0 1 51
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m15_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m15_w2_000_sli_dli_da_p_0
timestamp 1644511149
transform 1 0 54 0 1 51
box -26 -26 1688 456
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m15_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m15_w2_000_sli_dli_da_p_0
timestamp 1644511149
transform 1 0 54 0 1 963
box -59 -56 1721 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 954 707 954 707 4 Z
port 2 nsew
rlabel locali s 940 0 940 0 4 gnd
port 3 nsew
rlabel locali s 940 1414 940 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 1880 1414
string GDS_END 388138
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 385372
<< end >>
