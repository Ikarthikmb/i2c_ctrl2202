/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/esd_rf_diode_pd2nw_11v0/sky130_fd_pr__esd_rf_diode_pd2nw_11v0_300.model.spice