magic
tech sky130B
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdfm1sd2__example_5595914180827  sky130_fd_pr__hvdfm1sd2__example_5595914180827_0
timestamp 1644511149
transform 1 0 160 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808233  sky130_fd_pr__hvdfm1sd__example_55959141808233_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_55959141808233  sky130_fd_pr__hvdfm1sd__example_55959141808233_1
timestamp 1644511149
transform 1 0 376 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 404 481 404 481 0 FreeSans 300 0 0 0 D
flabel comment s 188 481 188 481 0 FreeSans 300 0 0 0 S
flabel comment s -28 481 -28 481 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 27762128
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27760686
<< end >>
