/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/res_xhigh_po/sky130_fd_pr__res_xhigh_po_5p73.model.spice