/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/sky130A/libs.tech/ngspice/sky130_fd_pr__model__r+c.model.spice