magic
tech sky130B
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__dfl1sd__example_55959141808190  sky130_fd_pr__dfl1sd__example_55959141808190_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_55959141808190  sky130_fd_pr__dfl1sd__example_55959141808190_1
timestamp 1644511149
transform 1 0 160 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 188 471 188 471 0 FreeSans 300 0 0 0 D
flabel comment s -28 471 -28 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 3258494
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3257444
<< end >>
