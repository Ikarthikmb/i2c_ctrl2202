magic
tech sky130A
timestamp 1644511149
<< properties >>
string GDS_END 35982246
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35980194
<< end >>
