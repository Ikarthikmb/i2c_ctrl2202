magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 68 21 822 203
rect 29 -17 63 17
<< scnmos >>
rect 155 47 185 177
rect 264 47 294 177
rect 336 47 366 177
rect 451 47 481 177
rect 537 47 567 177
rect 623 47 653 177
rect 709 47 739 177
<< scpmoshvt >>
rect 155 297 185 497
rect 264 297 294 497
rect 350 297 380 497
rect 451 297 481 497
rect 537 297 567 497
rect 623 297 653 497
rect 709 297 739 497
<< ndiff >>
rect 94 161 155 177
rect 94 127 110 161
rect 144 127 155 161
rect 94 93 155 127
rect 94 59 110 93
rect 144 59 155 93
rect 94 47 155 59
rect 185 47 264 177
rect 294 47 336 177
rect 366 89 451 177
rect 366 55 397 89
rect 431 55 451 89
rect 366 47 451 55
rect 481 153 537 177
rect 481 119 492 153
rect 526 119 537 153
rect 481 47 537 119
rect 567 89 623 177
rect 567 55 578 89
rect 612 55 623 89
rect 567 47 623 55
rect 653 169 709 177
rect 653 135 664 169
rect 698 135 709 169
rect 653 101 709 135
rect 653 67 664 101
rect 698 67 709 101
rect 653 47 709 67
rect 739 89 796 177
rect 739 55 750 89
rect 784 55 796 89
rect 739 47 796 55
<< pdiff >>
rect 94 477 155 497
rect 94 443 110 477
rect 144 443 155 477
rect 94 409 155 443
rect 94 375 110 409
rect 144 375 155 409
rect 94 297 155 375
rect 185 489 264 497
rect 185 455 209 489
rect 243 455 264 489
rect 185 421 264 455
rect 185 387 209 421
rect 243 387 264 421
rect 185 297 264 387
rect 294 477 350 497
rect 294 443 305 477
rect 339 443 350 477
rect 294 409 350 443
rect 294 375 305 409
rect 339 375 350 409
rect 294 297 350 375
rect 380 489 451 497
rect 380 455 398 489
rect 432 455 451 489
rect 380 421 451 455
rect 380 387 398 421
rect 432 387 451 421
rect 380 297 451 387
rect 481 477 537 497
rect 481 443 492 477
rect 526 443 537 477
rect 481 409 537 443
rect 481 375 492 409
rect 526 375 537 409
rect 481 297 537 375
rect 567 489 623 497
rect 567 455 578 489
rect 612 455 623 489
rect 567 421 623 455
rect 567 387 578 421
rect 612 387 623 421
rect 567 297 623 387
rect 653 477 709 497
rect 653 443 664 477
rect 698 443 709 477
rect 653 409 709 443
rect 653 375 664 409
rect 698 375 709 409
rect 653 341 709 375
rect 653 307 664 341
rect 698 307 709 341
rect 653 297 709 307
rect 739 489 796 497
rect 739 455 750 489
rect 784 455 796 489
rect 739 421 796 455
rect 739 387 750 421
rect 784 387 796 421
rect 739 297 796 387
<< ndiffc >>
rect 110 127 144 161
rect 110 59 144 93
rect 397 55 431 89
rect 492 119 526 153
rect 578 55 612 89
rect 664 135 698 169
rect 664 67 698 101
rect 750 55 784 89
<< pdiffc >>
rect 110 443 144 477
rect 110 375 144 409
rect 209 455 243 489
rect 209 387 243 421
rect 305 443 339 477
rect 305 375 339 409
rect 398 455 432 489
rect 398 387 432 421
rect 492 443 526 477
rect 492 375 526 409
rect 578 455 612 489
rect 578 387 612 421
rect 664 443 698 477
rect 664 375 698 409
rect 664 307 698 341
rect 750 455 784 489
rect 750 387 784 421
<< poly >>
rect 155 497 185 523
rect 264 497 294 523
rect 350 497 380 523
rect 451 497 481 523
rect 537 497 567 523
rect 623 497 653 523
rect 709 497 739 523
rect 155 265 185 297
rect 264 265 294 297
rect 350 265 380 297
rect 451 265 481 297
rect 537 265 567 297
rect 623 265 653 297
rect 709 265 739 297
rect 131 249 185 265
rect 131 215 141 249
rect 175 215 185 249
rect 131 199 185 215
rect 227 249 294 265
rect 227 215 237 249
rect 271 215 294 249
rect 227 199 294 215
rect 155 177 185 199
rect 264 177 294 199
rect 336 249 390 265
rect 336 215 346 249
rect 380 215 390 249
rect 336 199 390 215
rect 451 249 739 265
rect 451 215 467 249
rect 501 215 535 249
rect 569 215 603 249
rect 637 215 671 249
rect 705 215 739 249
rect 451 199 739 215
rect 336 177 366 199
rect 451 177 481 199
rect 537 177 567 199
rect 623 177 653 199
rect 709 177 739 199
rect 155 21 185 47
rect 264 21 294 47
rect 336 21 366 47
rect 451 21 481 47
rect 537 21 567 47
rect 623 21 653 47
rect 709 21 739 47
<< polycont >>
rect 141 215 175 249
rect 237 215 271 249
rect 346 215 380 249
rect 467 215 501 249
rect 535 215 569 249
rect 603 215 637 249
rect 671 215 705 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 109 477 145 493
rect 23 268 73 467
rect 109 443 110 477
rect 144 443 145 477
rect 109 409 145 443
rect 109 375 110 409
rect 144 375 145 409
rect 179 489 269 527
rect 179 455 209 489
rect 243 455 269 489
rect 179 421 269 455
rect 179 387 209 421
rect 243 387 269 421
rect 304 477 340 493
rect 304 443 305 477
rect 339 443 340 477
rect 304 409 340 443
rect 109 350 145 375
rect 304 375 305 409
rect 339 375 340 409
rect 382 489 448 527
rect 382 455 398 489
rect 432 455 448 489
rect 382 421 448 455
rect 382 387 398 421
rect 432 387 448 421
rect 490 477 528 493
rect 490 443 492 477
rect 526 443 528 477
rect 490 409 528 443
rect 304 350 340 375
rect 490 375 492 409
rect 526 375 528 409
rect 562 489 628 527
rect 562 455 578 489
rect 612 455 628 489
rect 562 421 628 455
rect 562 387 578 421
rect 612 387 628 421
rect 662 477 700 493
rect 662 443 664 477
rect 698 443 700 477
rect 662 409 700 443
rect 490 352 528 375
rect 662 375 664 409
rect 698 375 700 409
rect 734 489 800 527
rect 734 455 750 489
rect 784 455 800 489
rect 734 421 800 455
rect 734 387 750 421
rect 784 387 800 421
rect 662 353 700 375
rect 662 352 811 353
rect 109 316 456 350
rect 414 271 456 316
rect 490 341 811 352
rect 490 307 664 341
rect 698 307 811 341
rect 23 249 175 268
rect 23 215 141 249
rect 23 199 175 215
rect 213 249 271 268
rect 213 215 237 249
rect 93 127 110 161
rect 144 127 160 161
rect 213 149 271 215
rect 305 249 380 265
rect 305 215 346 249
rect 305 199 380 215
rect 414 249 721 271
rect 414 215 467 249
rect 501 215 535 249
rect 569 215 603 249
rect 637 215 671 249
rect 705 215 721 249
rect 414 204 721 215
rect 414 161 456 204
rect 755 169 811 307
rect 93 113 160 127
rect 307 123 456 161
rect 490 153 664 169
rect 307 113 345 123
rect 93 93 345 113
rect 490 119 492 153
rect 526 135 664 153
rect 698 135 811 169
rect 526 123 811 135
rect 526 119 528 123
rect 490 103 528 119
rect 93 59 110 93
rect 144 75 345 93
rect 662 101 700 123
rect 144 59 160 75
rect 93 51 160 59
rect 381 55 397 89
rect 431 55 447 89
rect 381 17 447 55
rect 562 55 578 89
rect 612 55 628 89
rect 562 17 628 55
rect 662 67 664 101
rect 698 67 700 101
rect 662 51 700 67
rect 734 55 750 89
rect 784 55 800 89
rect 734 17 800 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 121 221 155 255 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 340 0 0 0 C
port 3 nsew signal input
flabel locali s 765 153 799 187 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 and3_4
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 3877458
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3870622
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
