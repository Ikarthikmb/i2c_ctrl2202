magic
tech sky130A
timestamp 1644511149
<< properties >>
string GDS_END 6765066
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6764678
<< end >>
