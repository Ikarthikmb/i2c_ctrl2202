magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< locali >>
rect 167 480 179 514
rect 213 480 251 514
rect 285 480 323 514
rect 357 480 369 514
rect 167 20 179 54
rect 213 20 251 54
rect 285 20 323 54
rect 357 20 369 54
<< viali >>
rect 179 480 213 514
rect 251 480 285 514
rect 323 480 357 514
rect 179 20 213 54
rect 251 20 285 54
rect 323 20 357 54
<< obsli1 >>
rect 48 392 82 402
rect 48 320 82 358
rect 48 248 82 286
rect 48 176 82 214
rect 48 132 82 142
rect 159 98 193 436
rect 251 98 285 436
rect 343 98 377 436
rect 454 392 488 402
rect 454 320 488 358
rect 454 248 488 286
rect 454 176 488 214
rect 454 132 488 142
<< obsli1c >>
rect 48 358 82 392
rect 48 286 82 320
rect 48 214 82 248
rect 48 142 82 176
rect 454 358 488 392
rect 454 286 488 320
rect 454 214 488 248
rect 454 142 488 176
<< metal1 >>
rect 167 514 369 534
rect 167 480 179 514
rect 213 480 251 514
rect 285 480 323 514
rect 357 480 369 514
rect 167 468 369 480
rect 36 392 94 420
rect 36 358 48 392
rect 82 358 94 392
rect 36 320 94 358
rect 36 286 48 320
rect 82 286 94 320
rect 36 248 94 286
rect 36 214 48 248
rect 82 214 94 248
rect 36 176 94 214
rect 36 142 48 176
rect 82 142 94 176
rect 36 114 94 142
rect 442 392 500 420
rect 442 358 454 392
rect 488 358 500 392
rect 442 320 500 358
rect 442 286 454 320
rect 488 286 500 320
rect 442 248 500 286
rect 442 214 454 248
rect 488 214 500 248
rect 442 176 500 214
rect 442 142 454 176
rect 488 142 500 176
rect 442 114 500 142
rect 167 54 369 66
rect 167 20 179 54
rect 213 20 251 54
rect 285 20 323 54
rect 357 20 369 54
rect 167 0 369 20
<< obsm1 >>
rect 150 114 202 420
rect 242 114 294 420
rect 334 114 386 420
<< metal2 >>
rect 10 292 526 420
rect 10 114 526 242
<< labels >>
rlabel metal1 s 442 114 500 420 6 BULK
port 1 nsew
rlabel metal1 s 36 114 94 420 6 BULK
port 1 nsew
rlabel metal2 s 10 292 526 420 6 DRAIN
port 2 nsew
rlabel viali s 323 480 357 514 6 GATE
port 3 nsew
rlabel viali s 323 20 357 54 6 GATE
port 3 nsew
rlabel viali s 251 480 285 514 6 GATE
port 3 nsew
rlabel viali s 251 20 285 54 6 GATE
port 3 nsew
rlabel viali s 179 480 213 514 6 GATE
port 3 nsew
rlabel viali s 179 20 213 54 6 GATE
port 3 nsew
rlabel locali s 167 480 369 514 6 GATE
port 3 nsew
rlabel locali s 167 20 369 54 6 GATE
port 3 nsew
rlabel metal1 s 167 468 369 534 6 GATE
port 3 nsew
rlabel metal1 s 167 0 369 66 6 GATE
port 3 nsew
rlabel metal2 s 10 114 526 242 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 536 534
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9346270
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9338618
<< end >>
