magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1970 582
<< pwell >>
rect 13 21 1919 203
rect 25 -17 59 21
<< locali >>
rect 811 345 861 423
rect 995 345 1029 423
rect 1163 345 1201 493
rect 1335 345 1369 493
rect 1503 345 1537 493
rect 1671 345 1705 493
rect 1839 345 1915 493
rect 811 297 1915 345
rect 17 211 355 263
rect 389 211 723 263
rect 761 211 1177 263
rect 1211 211 1539 263
rect 1573 211 1818 263
rect 1852 177 1915 297
rect 1579 131 1915 177
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 17 345 81 493
rect 119 379 185 527
rect 219 345 253 493
rect 287 379 353 527
rect 387 345 421 493
rect 455 459 1129 493
rect 455 379 521 459
rect 555 345 589 423
rect 623 379 689 459
rect 723 345 773 423
rect 17 297 773 345
rect 895 379 961 459
rect 1063 379 1129 459
rect 1235 379 1301 527
rect 1403 379 1469 527
rect 1571 379 1637 527
rect 1739 379 1805 527
rect 17 17 101 177
rect 135 131 1477 177
rect 135 51 169 131
rect 203 17 269 97
rect 303 51 337 131
rect 371 17 437 97
rect 471 51 505 131
rect 539 17 605 97
rect 639 51 673 131
rect 707 17 777 97
rect 811 51 845 131
rect 879 17 945 97
rect 979 51 1013 131
rect 1511 97 1545 177
rect 1047 17 1117 97
rect 1151 51 1915 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
<< metal1 >>
rect 0 561 1932 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1932 561
rect 0 496 1932 527
rect 0 17 1932 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1932 17
rect 0 -48 1932 -17
<< labels >>
rlabel locali s 17 211 355 263 6 A1
port 1 nsew signal input
rlabel locali s 389 211 723 263 6 A2
port 2 nsew signal input
rlabel locali s 761 211 1177 263 6 A3
port 3 nsew signal input
rlabel locali s 1211 211 1539 263 6 B1
port 4 nsew signal input
rlabel locali s 1573 211 1818 263 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 1932 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 25 -17 59 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 13 21 1919 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1970 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1932 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1579 131 1915 177 6 Y
port 10 nsew signal output
rlabel locali s 1852 177 1915 297 6 Y
port 10 nsew signal output
rlabel locali s 811 297 1915 345 6 Y
port 10 nsew signal output
rlabel locali s 1839 345 1915 493 6 Y
port 10 nsew signal output
rlabel locali s 1671 345 1705 493 6 Y
port 10 nsew signal output
rlabel locali s 1503 345 1537 493 6 Y
port 10 nsew signal output
rlabel locali s 1335 345 1369 493 6 Y
port 10 nsew signal output
rlabel locali s 1163 345 1201 493 6 Y
port 10 nsew signal output
rlabel locali s 995 345 1029 423 6 Y
port 10 nsew signal output
rlabel locali s 811 345 861 423 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1932 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 926530
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 910678
<< end >>
