magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1099 203
rect 30 -17 64 21
<< locali >>
rect 183 340 221 493
rect 355 340 391 493
rect 18 306 391 340
rect 18 161 64 306
rect 497 215 631 323
rect 696 299 1080 341
rect 696 198 757 299
rect 828 199 938 265
rect 1006 199 1080 299
rect 18 127 343 161
rect 119 123 343 127
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 83 374 149 527
rect 255 374 321 527
rect 427 451 497 527
rect 531 421 569 493
rect 603 455 737 527
rect 843 421 909 489
rect 531 417 909 421
rect 425 375 909 417
rect 1015 387 1087 527
rect 425 366 569 375
rect 425 267 463 366
rect 98 199 463 267
rect 423 174 463 199
rect 423 131 619 174
rect 655 123 1081 157
rect 655 97 721 123
rect 19 17 85 93
rect 191 17 257 89
rect 363 17 429 93
rect 467 51 721 97
rect 755 17 823 89
rect 929 17 995 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 1006 199 1080 299 6 A1
port 1 nsew signal input
rlabel locali s 696 198 757 299 6 A1
port 1 nsew signal input
rlabel locali s 696 299 1080 341 6 A1
port 1 nsew signal input
rlabel locali s 828 199 938 265 6 A2
port 2 nsew signal input
rlabel locali s 497 215 631 323 6 B1
port 3 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1099 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 119 123 343 127 6 X
port 8 nsew signal output
rlabel locali s 18 127 343 161 6 X
port 8 nsew signal output
rlabel locali s 18 161 64 306 6 X
port 8 nsew signal output
rlabel locali s 18 306 391 340 6 X
port 8 nsew signal output
rlabel locali s 355 340 391 493 6 X
port 8 nsew signal output
rlabel locali s 183 340 221 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1285428
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1277504
<< end >>
