magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1551 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 855 47 885 177
rect 939 47 969 177
rect 1023 47 1053 177
rect 1107 47 1137 177
rect 1191 47 1221 177
rect 1275 47 1305 177
rect 1359 47 1389 177
rect 1443 47 1473 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 855 297 885 497
rect 939 297 969 497
rect 1023 297 1053 497
rect 1107 297 1137 497
rect 1191 297 1221 497
rect 1275 297 1305 497
rect 1359 297 1389 497
rect 1443 297 1473 497
<< ndiff >>
rect 27 163 79 177
rect 27 129 35 163
rect 69 129 79 163
rect 27 95 79 129
rect 27 61 35 95
rect 69 61 79 95
rect 27 47 79 61
rect 109 95 163 177
rect 109 61 119 95
rect 153 61 163 95
rect 109 47 163 61
rect 193 163 247 177
rect 193 129 203 163
rect 237 129 247 163
rect 193 95 247 129
rect 193 61 203 95
rect 237 61 247 95
rect 193 47 247 61
rect 277 95 331 177
rect 277 61 287 95
rect 321 61 331 95
rect 277 47 331 61
rect 361 163 415 177
rect 361 129 371 163
rect 405 129 415 163
rect 361 95 415 129
rect 361 61 371 95
rect 405 61 415 95
rect 361 47 415 61
rect 445 163 499 177
rect 445 129 455 163
rect 489 129 499 163
rect 445 47 499 129
rect 529 95 583 177
rect 529 61 539 95
rect 573 61 583 95
rect 529 47 583 61
rect 613 163 667 177
rect 613 129 623 163
rect 657 129 667 163
rect 613 47 667 129
rect 697 95 749 177
rect 697 61 707 95
rect 741 61 749 95
rect 697 47 749 61
rect 803 95 855 177
rect 803 61 811 95
rect 845 61 855 95
rect 803 47 855 61
rect 885 163 939 177
rect 885 129 895 163
rect 929 129 939 163
rect 885 47 939 129
rect 969 95 1023 177
rect 969 61 979 95
rect 1013 61 1023 95
rect 969 47 1023 61
rect 1053 163 1107 177
rect 1053 129 1063 163
rect 1097 129 1107 163
rect 1053 47 1107 129
rect 1137 163 1191 177
rect 1137 129 1147 163
rect 1181 129 1191 163
rect 1137 95 1191 129
rect 1137 61 1147 95
rect 1181 61 1191 95
rect 1137 47 1191 61
rect 1221 95 1275 177
rect 1221 61 1231 95
rect 1265 61 1275 95
rect 1221 47 1275 61
rect 1305 163 1359 177
rect 1305 129 1315 163
rect 1349 129 1359 163
rect 1305 95 1359 129
rect 1305 61 1315 95
rect 1349 61 1359 95
rect 1305 47 1359 61
rect 1389 95 1443 177
rect 1389 61 1399 95
rect 1433 61 1443 95
rect 1389 47 1443 61
rect 1473 163 1525 177
rect 1473 129 1483 163
rect 1517 129 1525 163
rect 1473 95 1525 129
rect 1473 61 1483 95
rect 1517 61 1525 95
rect 1473 47 1525 61
<< pdiff >>
rect 27 481 79 497
rect 27 447 35 481
rect 69 447 79 481
rect 27 413 79 447
rect 27 379 35 413
rect 69 379 79 413
rect 27 345 79 379
rect 27 311 35 345
rect 69 311 79 345
rect 27 297 79 311
rect 109 409 163 497
rect 109 375 119 409
rect 153 375 163 409
rect 109 341 163 375
rect 109 307 119 341
rect 153 307 163 341
rect 109 297 163 307
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 409 331 497
rect 277 375 287 409
rect 321 375 331 409
rect 277 341 331 375
rect 277 307 287 341
rect 321 307 331 341
rect 277 297 331 307
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 409 415 443
rect 361 375 371 409
rect 405 375 415 409
rect 361 297 415 375
rect 445 409 499 497
rect 445 375 455 409
rect 489 375 499 409
rect 445 341 499 375
rect 445 307 455 341
rect 489 307 499 341
rect 445 297 499 307
rect 529 477 583 497
rect 529 443 539 477
rect 573 443 583 477
rect 529 409 583 443
rect 529 375 539 409
rect 573 375 583 409
rect 529 297 583 375
rect 613 409 667 497
rect 613 375 623 409
rect 657 375 667 409
rect 613 341 667 375
rect 613 307 623 341
rect 657 307 667 341
rect 613 297 667 307
rect 697 477 855 497
rect 697 443 707 477
rect 741 443 811 477
rect 845 443 855 477
rect 697 409 855 443
rect 697 375 707 409
rect 741 375 811 409
rect 845 375 855 409
rect 697 341 855 375
rect 697 307 707 341
rect 741 307 811 341
rect 845 307 855 341
rect 697 297 855 307
rect 885 477 939 497
rect 885 443 895 477
rect 929 443 939 477
rect 885 409 939 443
rect 885 375 895 409
rect 929 375 939 409
rect 885 297 939 375
rect 969 477 1023 497
rect 969 443 979 477
rect 1013 443 1023 477
rect 969 409 1023 443
rect 969 375 979 409
rect 1013 375 1023 409
rect 969 341 1023 375
rect 969 307 979 341
rect 1013 307 1023 341
rect 969 297 1023 307
rect 1053 477 1107 497
rect 1053 443 1063 477
rect 1097 443 1107 477
rect 1053 409 1107 443
rect 1053 375 1063 409
rect 1097 375 1107 409
rect 1053 297 1107 375
rect 1137 477 1191 497
rect 1137 443 1147 477
rect 1181 443 1191 477
rect 1137 409 1191 443
rect 1137 375 1147 409
rect 1181 375 1191 409
rect 1137 341 1191 375
rect 1137 307 1147 341
rect 1181 307 1191 341
rect 1137 297 1191 307
rect 1221 477 1275 497
rect 1221 443 1231 477
rect 1265 443 1275 477
rect 1221 409 1275 443
rect 1221 375 1231 409
rect 1265 375 1275 409
rect 1221 297 1275 375
rect 1305 477 1359 497
rect 1305 443 1315 477
rect 1349 443 1359 477
rect 1305 409 1359 443
rect 1305 375 1315 409
rect 1349 375 1359 409
rect 1305 341 1359 375
rect 1305 307 1315 341
rect 1349 307 1359 341
rect 1305 297 1359 307
rect 1389 477 1443 497
rect 1389 443 1399 477
rect 1433 443 1443 477
rect 1389 409 1443 443
rect 1389 375 1399 409
rect 1433 375 1443 409
rect 1389 297 1443 375
rect 1473 477 1533 497
rect 1473 443 1483 477
rect 1517 443 1533 477
rect 1473 409 1533 443
rect 1473 375 1483 409
rect 1517 375 1533 409
rect 1473 341 1533 375
rect 1473 307 1483 341
rect 1517 307 1533 341
rect 1473 297 1533 307
<< ndiffc >>
rect 35 129 69 163
rect 35 61 69 95
rect 119 61 153 95
rect 203 129 237 163
rect 203 61 237 95
rect 287 61 321 95
rect 371 129 405 163
rect 371 61 405 95
rect 455 129 489 163
rect 539 61 573 95
rect 623 129 657 163
rect 707 61 741 95
rect 811 61 845 95
rect 895 129 929 163
rect 979 61 1013 95
rect 1063 129 1097 163
rect 1147 129 1181 163
rect 1147 61 1181 95
rect 1231 61 1265 95
rect 1315 129 1349 163
rect 1315 61 1349 95
rect 1399 61 1433 95
rect 1483 129 1517 163
rect 1483 61 1517 95
<< pdiffc >>
rect 35 447 69 481
rect 35 379 69 413
rect 35 311 69 345
rect 119 375 153 409
rect 119 307 153 341
rect 203 443 237 477
rect 203 375 237 409
rect 287 375 321 409
rect 287 307 321 341
rect 371 443 405 477
rect 371 375 405 409
rect 455 375 489 409
rect 455 307 489 341
rect 539 443 573 477
rect 539 375 573 409
rect 623 375 657 409
rect 623 307 657 341
rect 707 443 741 477
rect 811 443 845 477
rect 707 375 741 409
rect 811 375 845 409
rect 707 307 741 341
rect 811 307 845 341
rect 895 443 929 477
rect 895 375 929 409
rect 979 443 1013 477
rect 979 375 1013 409
rect 979 307 1013 341
rect 1063 443 1097 477
rect 1063 375 1097 409
rect 1147 443 1181 477
rect 1147 375 1181 409
rect 1147 307 1181 341
rect 1231 443 1265 477
rect 1231 375 1265 409
rect 1315 443 1349 477
rect 1315 375 1349 409
rect 1315 307 1349 341
rect 1399 443 1433 477
rect 1399 375 1433 409
rect 1483 443 1517 477
rect 1483 375 1517 409
rect 1483 307 1517 341
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 855 497 885 523
rect 939 497 969 523
rect 1023 497 1053 523
rect 1107 497 1137 523
rect 1191 497 1221 523
rect 1275 497 1305 523
rect 1359 497 1389 523
rect 1443 497 1473 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 331 265 361 297
rect 79 249 361 265
rect 79 215 107 249
rect 141 215 175 249
rect 209 215 243 249
rect 277 215 311 249
rect 345 215 361 249
rect 79 199 361 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 331 177 361 199
rect 415 265 445 297
rect 499 265 529 297
rect 583 265 613 297
rect 667 265 697 297
rect 855 265 885 297
rect 939 265 969 297
rect 1023 265 1053 297
rect 1107 265 1137 297
rect 415 249 732 265
rect 415 215 546 249
rect 580 215 614 249
rect 648 215 682 249
rect 716 215 732 249
rect 415 199 732 215
rect 855 249 1137 265
rect 855 215 871 249
rect 905 215 939 249
rect 973 215 1007 249
rect 1041 215 1075 249
rect 1109 215 1137 249
rect 855 199 1137 215
rect 415 177 445 199
rect 499 177 529 199
rect 583 177 613 199
rect 667 177 697 199
rect 855 177 885 199
rect 939 177 969 199
rect 1023 177 1053 199
rect 1107 177 1137 199
rect 1191 265 1221 297
rect 1275 265 1305 297
rect 1359 265 1389 297
rect 1443 265 1473 297
rect 1191 249 1473 265
rect 1191 215 1207 249
rect 1241 215 1275 249
rect 1309 215 1343 249
rect 1377 215 1411 249
rect 1445 215 1473 249
rect 1191 199 1473 215
rect 1191 177 1221 199
rect 1275 177 1305 199
rect 1359 177 1389 199
rect 1443 177 1473 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 855 21 885 47
rect 939 21 969 47
rect 1023 21 1053 47
rect 1107 21 1137 47
rect 1191 21 1221 47
rect 1275 21 1305 47
rect 1359 21 1389 47
rect 1443 21 1473 47
<< polycont >>
rect 107 215 141 249
rect 175 215 209 249
rect 243 215 277 249
rect 311 215 345 249
rect 546 215 580 249
rect 614 215 648 249
rect 682 215 716 249
rect 871 215 905 249
rect 939 215 973 249
rect 1007 215 1041 249
rect 1075 215 1109 249
rect 1207 215 1241 249
rect 1275 215 1309 249
rect 1343 215 1377 249
rect 1411 215 1445 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 18 481 853 493
rect 18 447 35 481
rect 69 477 853 481
rect 69 459 203 477
rect 69 447 85 459
rect 18 413 85 447
rect 195 443 203 459
rect 237 459 371 477
rect 237 443 245 459
rect 18 379 35 413
rect 69 379 85 413
rect 18 345 85 379
rect 18 311 35 345
rect 69 311 85 345
rect 18 291 85 311
rect 119 409 161 425
rect 153 375 161 409
rect 119 341 161 375
rect 195 409 245 443
rect 363 443 371 459
rect 405 459 539 477
rect 405 443 413 459
rect 195 375 203 409
rect 237 375 245 409
rect 195 359 245 375
rect 279 409 329 425
rect 279 375 287 409
rect 321 375 329 409
rect 153 325 161 341
rect 279 341 329 375
rect 363 409 413 443
rect 531 443 539 459
rect 573 459 707 477
rect 573 443 581 459
rect 363 375 371 409
rect 405 375 413 409
rect 363 359 413 375
rect 447 409 497 425
rect 447 375 455 409
rect 489 375 497 409
rect 279 325 287 341
rect 153 307 287 325
rect 321 325 329 341
rect 447 341 497 375
rect 531 409 581 443
rect 699 443 707 459
rect 741 443 811 477
rect 845 443 853 477
rect 531 375 539 409
rect 573 375 581 409
rect 531 359 581 375
rect 615 409 665 425
rect 615 375 623 409
rect 657 375 665 409
rect 447 325 455 341
rect 321 307 455 325
rect 489 325 497 341
rect 615 341 665 375
rect 615 325 623 341
rect 489 307 623 325
rect 657 307 665 341
rect 119 289 665 307
rect 699 409 853 443
rect 699 375 707 409
rect 741 375 811 409
rect 845 375 853 409
rect 699 341 853 375
rect 887 477 937 527
rect 887 443 895 477
rect 929 443 937 477
rect 887 409 937 443
rect 887 375 895 409
rect 929 375 937 409
rect 887 359 937 375
rect 971 477 1021 493
rect 971 443 979 477
rect 1013 443 1021 477
rect 971 409 1021 443
rect 971 375 979 409
rect 1013 375 1021 409
rect 699 307 707 341
rect 741 307 811 341
rect 845 325 853 341
rect 971 341 1021 375
rect 1055 477 1105 527
rect 1055 443 1063 477
rect 1097 443 1105 477
rect 1055 409 1105 443
rect 1055 375 1063 409
rect 1097 375 1105 409
rect 1055 359 1105 375
rect 1139 477 1189 493
rect 1139 443 1147 477
rect 1181 443 1189 477
rect 1139 409 1189 443
rect 1139 375 1147 409
rect 1181 375 1189 409
rect 971 325 979 341
rect 845 307 979 325
rect 1013 325 1021 341
rect 1139 341 1189 375
rect 1223 477 1273 527
rect 1223 443 1231 477
rect 1265 443 1273 477
rect 1223 409 1273 443
rect 1223 375 1231 409
rect 1265 375 1273 409
rect 1223 359 1273 375
rect 1307 477 1357 493
rect 1307 443 1315 477
rect 1349 443 1357 477
rect 1307 409 1357 443
rect 1307 375 1315 409
rect 1349 375 1357 409
rect 1139 325 1147 341
rect 1013 307 1147 325
rect 1181 325 1189 341
rect 1307 341 1357 375
rect 1391 477 1441 527
rect 1391 443 1399 477
rect 1433 443 1441 477
rect 1391 409 1441 443
rect 1391 375 1399 409
rect 1433 375 1441 409
rect 1391 359 1441 375
rect 1475 477 1525 493
rect 1475 443 1483 477
rect 1517 443 1525 477
rect 1475 409 1525 443
rect 1475 375 1483 409
rect 1517 375 1525 409
rect 1307 325 1315 341
rect 1181 307 1315 325
rect 1349 325 1357 341
rect 1475 341 1525 375
rect 1475 325 1483 341
rect 1349 307 1483 325
rect 1517 307 1525 341
rect 699 291 1525 307
rect 18 249 379 255
rect 18 215 107 249
rect 141 215 175 249
rect 209 215 243 249
rect 277 215 311 249
rect 345 215 379 249
rect 19 163 405 181
rect 19 129 35 163
rect 69 145 203 163
rect 69 129 85 145
rect 19 95 85 129
rect 187 129 203 145
rect 237 145 371 163
rect 237 129 253 145
rect 19 61 35 95
rect 69 61 85 95
rect 19 51 85 61
rect 119 95 153 111
rect 119 17 153 61
rect 187 95 253 129
rect 355 129 371 145
rect 439 177 489 289
rect 523 249 808 255
rect 523 215 546 249
rect 580 215 614 249
rect 648 215 682 249
rect 716 215 808 249
rect 855 249 1137 257
rect 855 215 871 249
rect 905 215 939 249
rect 973 215 1007 249
rect 1041 215 1075 249
rect 1109 215 1137 249
rect 1182 249 1547 257
rect 1182 215 1207 249
rect 1241 215 1275 249
rect 1309 215 1343 249
rect 1377 215 1411 249
rect 1445 215 1547 249
rect 439 163 1113 177
rect 439 129 455 163
rect 489 129 623 163
rect 657 129 895 163
rect 929 129 1063 163
rect 1097 129 1113 163
rect 1147 163 1533 181
rect 1181 145 1315 163
rect 1181 129 1197 145
rect 187 61 203 95
rect 237 61 253 95
rect 187 51 253 61
rect 287 95 321 111
rect 287 17 321 61
rect 355 95 405 129
rect 1147 95 1197 129
rect 1299 129 1315 145
rect 1349 145 1483 163
rect 1349 129 1365 145
rect 355 61 371 95
rect 405 61 539 95
rect 573 61 707 95
rect 741 61 757 95
rect 355 51 757 61
rect 795 61 811 95
rect 845 61 979 95
rect 1013 61 1147 95
rect 1181 61 1197 95
rect 795 51 1197 61
rect 1231 95 1265 111
rect 1231 17 1265 61
rect 1299 95 1365 129
rect 1467 129 1483 145
rect 1517 129 1533 163
rect 1299 61 1315 95
rect 1349 61 1365 95
rect 1299 51 1365 61
rect 1399 95 1433 111
rect 1399 17 1433 61
rect 1467 95 1533 129
rect 1467 61 1483 95
rect 1517 61 1533 95
rect 1467 51 1533 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 1322 221 1356 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 400 180 0 0 B2
port 4 nsew signal input
flabel locali s 954 221 988 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 400 180 0 0 B1
port 3 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 400 180 0 0 Y
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a22oi_4
rlabel metal1 s 0 -48 1564 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 4110910
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4098918
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 39.100 0.000 
<< end >>
