magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< locali >>
rect 4094 50423 4122 50457
rect 86 50386 120 50402
rect 86 50336 120 50352
rect 70 50244 136 50278
rect 70 50052 136 50086
rect 86 49978 120 49994
rect 86 49928 120 49944
rect 4094 49873 4122 49907
rect 4094 49633 4122 49667
rect 86 49596 120 49612
rect 86 49546 120 49562
rect 70 49454 136 49488
rect 70 49262 136 49296
rect 86 49188 120 49204
rect 86 49138 120 49154
rect 4094 49083 4122 49117
rect 4094 48843 4122 48877
rect 86 48806 120 48822
rect 86 48756 120 48772
rect 70 48664 136 48698
rect 70 48472 136 48506
rect 86 48398 120 48414
rect 86 48348 120 48364
rect 4094 48293 4122 48327
rect 4094 48053 4122 48087
rect 86 48016 120 48032
rect 86 47966 120 47982
rect 70 47874 136 47908
rect 70 47682 136 47716
rect 86 47608 120 47624
rect 86 47558 120 47574
rect 4094 47503 4122 47537
rect 4094 47263 4122 47297
rect 86 47226 120 47242
rect 86 47176 120 47192
rect 70 47084 136 47118
rect 70 46892 136 46926
rect 86 46818 120 46834
rect 86 46768 120 46784
rect 4094 46713 4122 46747
rect 4094 46473 4122 46507
rect 86 46436 120 46452
rect 86 46386 120 46402
rect 70 46294 136 46328
rect 70 46102 136 46136
rect 86 46028 120 46044
rect 86 45978 120 45994
rect 4094 45923 4122 45957
rect 4094 45683 4122 45717
rect 86 45646 120 45662
rect 86 45596 120 45612
rect 70 45504 136 45538
rect 70 45312 136 45346
rect 86 45238 120 45254
rect 86 45188 120 45204
rect 4094 45133 4122 45167
rect 4094 44893 4122 44927
rect 86 44856 120 44872
rect 86 44806 120 44822
rect 70 44714 136 44748
rect 70 44522 136 44556
rect 86 44448 120 44464
rect 86 44398 120 44414
rect 4094 44343 4122 44377
rect 4094 44103 4122 44137
rect 86 44066 120 44082
rect 86 44016 120 44032
rect 70 43924 136 43958
rect 70 43732 136 43766
rect 86 43658 120 43674
rect 86 43608 120 43624
rect 4094 43553 4122 43587
rect 4094 43313 4122 43347
rect 86 43276 120 43292
rect 86 43226 120 43242
rect 70 43134 136 43168
rect 70 42942 136 42976
rect 86 42868 120 42884
rect 86 42818 120 42834
rect 4094 42763 4122 42797
rect 4094 42523 4122 42557
rect 86 42486 120 42502
rect 86 42436 120 42452
rect 70 42344 136 42378
rect 70 42152 136 42186
rect 86 42078 120 42094
rect 86 42028 120 42044
rect 4094 41973 4122 42007
rect 4094 41733 4122 41767
rect 86 41696 120 41712
rect 86 41646 120 41662
rect 70 41554 136 41588
rect 70 41362 136 41396
rect 86 41288 120 41304
rect 86 41238 120 41254
rect 4094 41183 4122 41217
rect 4094 40943 4122 40977
rect 86 40906 120 40922
rect 86 40856 120 40872
rect 70 40764 136 40798
rect 70 40572 136 40606
rect 86 40498 120 40514
rect 86 40448 120 40464
rect 4094 40393 4122 40427
rect 4094 40153 4122 40187
rect 86 40116 120 40132
rect 86 40066 120 40082
rect 70 39974 136 40008
rect 70 39782 136 39816
rect 86 39708 120 39724
rect 86 39658 120 39674
rect 4094 39603 4122 39637
rect 4094 39363 4122 39397
rect 86 39326 120 39342
rect 86 39276 120 39292
rect 70 39184 136 39218
rect 70 38992 136 39026
rect 86 38918 120 38934
rect 86 38868 120 38884
rect 4094 38813 4122 38847
rect 4094 38573 4122 38607
rect 86 38536 120 38552
rect 86 38486 120 38502
rect 70 38394 136 38428
rect 70 38202 136 38236
rect 86 38128 120 38144
rect 86 38078 120 38094
rect 4094 38023 4122 38057
rect 4094 37783 4122 37817
rect 86 37746 120 37762
rect 86 37696 120 37712
rect 70 37604 136 37638
rect 70 37412 136 37446
rect 86 37338 120 37354
rect 86 37288 120 37304
rect 4094 37233 4122 37267
rect 4094 36993 4122 37027
rect 86 36956 120 36972
rect 86 36906 120 36922
rect 70 36814 136 36848
rect 70 36622 136 36656
rect 86 36548 120 36564
rect 86 36498 120 36514
rect 4094 36443 4122 36477
rect 4094 36203 4122 36237
rect 86 36166 120 36182
rect 86 36116 120 36132
rect 70 36024 136 36058
rect 70 35832 136 35866
rect 86 35758 120 35774
rect 86 35708 120 35724
rect 4094 35653 4122 35687
rect 4094 35413 4122 35447
rect 86 35376 120 35392
rect 86 35326 120 35342
rect 70 35234 136 35268
rect 70 35042 136 35076
rect 86 34968 120 34984
rect 86 34918 120 34934
rect 4094 34863 4122 34897
rect 4094 34623 4122 34657
rect 86 34586 120 34602
rect 86 34536 120 34552
rect 70 34444 136 34478
rect 70 34252 136 34286
rect 86 34178 120 34194
rect 86 34128 120 34144
rect 4094 34073 4122 34107
rect 4094 33833 4122 33867
rect 86 33796 120 33812
rect 86 33746 120 33762
rect 70 33654 136 33688
rect 70 33462 136 33496
rect 86 33388 120 33404
rect 86 33338 120 33354
rect 4094 33283 4122 33317
rect 4094 33043 4122 33077
rect 86 33006 120 33022
rect 86 32956 120 32972
rect 70 32864 136 32898
rect 70 32672 136 32706
rect 86 32598 120 32614
rect 86 32548 120 32564
rect 4094 32493 4122 32527
rect 4094 32253 4122 32287
rect 86 32216 120 32232
rect 86 32166 120 32182
rect 70 32074 136 32108
rect 70 31882 136 31916
rect 86 31808 120 31824
rect 86 31758 120 31774
rect 4094 31703 4122 31737
rect 4094 31463 4122 31497
rect 86 31426 120 31442
rect 86 31376 120 31392
rect 70 31284 136 31318
rect 70 31092 136 31126
rect 86 31018 120 31034
rect 86 30968 120 30984
rect 4094 30913 4122 30947
rect 4094 30673 4122 30707
rect 86 30636 120 30652
rect 86 30586 120 30602
rect 70 30494 136 30528
rect 70 30302 136 30336
rect 86 30228 120 30244
rect 86 30178 120 30194
rect 4094 30123 4122 30157
rect 4094 29883 4122 29917
rect 86 29846 120 29862
rect 86 29796 120 29812
rect 70 29704 136 29738
rect 70 29512 136 29546
rect 86 29438 120 29454
rect 86 29388 120 29404
rect 4094 29333 4122 29367
rect 4094 29093 4122 29127
rect 86 29056 120 29072
rect 86 29006 120 29022
rect 70 28914 136 28948
rect 70 28722 136 28756
rect 86 28648 120 28664
rect 86 28598 120 28614
rect 4094 28543 4122 28577
rect 4094 28303 4122 28337
rect 86 28266 120 28282
rect 86 28216 120 28232
rect 70 28124 136 28158
rect 70 27932 136 27966
rect 86 27858 120 27874
rect 86 27808 120 27824
rect 4094 27753 4122 27787
rect 4094 27513 4122 27547
rect 86 27476 120 27492
rect 86 27426 120 27442
rect 70 27334 136 27368
rect 70 27142 136 27176
rect 86 27068 120 27084
rect 86 27018 120 27034
rect 4094 26963 4122 26997
rect 4094 26723 4122 26757
rect 86 26686 120 26702
rect 86 26636 120 26652
rect 70 26544 136 26578
rect 70 26352 136 26386
rect 86 26278 120 26294
rect 86 26228 120 26244
rect 4094 26173 4122 26207
rect 4094 25933 4122 25967
rect 86 25896 120 25912
rect 86 25846 120 25862
rect 70 25754 136 25788
rect 70 25562 136 25596
rect 86 25488 120 25504
rect 86 25438 120 25454
rect 4094 25383 4122 25417
rect 4094 25143 4122 25177
rect 86 25106 120 25122
rect 86 25056 120 25072
rect 70 24964 136 24998
rect 70 24772 136 24806
rect 86 24698 120 24714
rect 86 24648 120 24664
rect 4094 24593 4122 24627
rect 4094 24353 4122 24387
rect 86 24316 120 24332
rect 86 24266 120 24282
rect 70 24174 136 24208
rect 70 23982 136 24016
rect 86 23908 120 23924
rect 86 23858 120 23874
rect 4094 23803 4122 23837
rect 4094 23563 4122 23597
rect 86 23526 120 23542
rect 86 23476 120 23492
rect 70 23384 136 23418
rect 70 23192 136 23226
rect 86 23118 120 23134
rect 86 23068 120 23084
rect 4094 23013 4122 23047
rect 4094 22773 4122 22807
rect 86 22736 120 22752
rect 86 22686 120 22702
rect 70 22594 136 22628
rect 70 22402 136 22436
rect 86 22328 120 22344
rect 86 22278 120 22294
rect 4094 22223 4122 22257
rect 4094 21983 4122 22017
rect 86 21946 120 21962
rect 86 21896 120 21912
rect 70 21804 136 21838
rect 70 21612 136 21646
rect 86 21538 120 21554
rect 86 21488 120 21504
rect 4094 21433 4122 21467
rect 4094 21193 4122 21227
rect 86 21156 120 21172
rect 86 21106 120 21122
rect 70 21014 136 21048
rect 70 20822 136 20856
rect 86 20748 120 20764
rect 86 20698 120 20714
rect 4094 20643 4122 20677
rect 4094 20403 4122 20437
rect 86 20366 120 20382
rect 86 20316 120 20332
rect 70 20224 136 20258
rect 70 20032 136 20066
rect 86 19958 120 19974
rect 86 19908 120 19924
rect 4094 19853 4122 19887
rect 4094 19613 4122 19647
rect 86 19576 120 19592
rect 86 19526 120 19542
rect 70 19434 136 19468
rect 70 19242 136 19276
rect 86 19168 120 19184
rect 86 19118 120 19134
rect 4094 19063 4122 19097
rect 4094 18823 4122 18857
rect 86 18786 120 18802
rect 86 18736 120 18752
rect 70 18644 136 18678
rect 70 18452 136 18486
rect 86 18378 120 18394
rect 86 18328 120 18344
rect 4094 18273 4122 18307
rect 4094 18033 4122 18067
rect 86 17996 120 18012
rect 86 17946 120 17962
rect 70 17854 136 17888
rect 70 17662 136 17696
rect 86 17588 120 17604
rect 86 17538 120 17554
rect 4094 17483 4122 17517
rect 4094 17243 4122 17277
rect 86 17206 120 17222
rect 86 17156 120 17172
rect 70 17064 136 17098
rect 70 16872 136 16906
rect 86 16798 120 16814
rect 86 16748 120 16764
rect 4094 16693 4122 16727
rect 4094 16453 4122 16487
rect 86 16416 120 16432
rect 86 16366 120 16382
rect 70 16274 136 16308
rect 70 16082 136 16116
rect 86 16008 120 16024
rect 86 15958 120 15974
rect 4094 15903 4122 15937
rect 4094 15663 4122 15697
rect 86 15626 120 15642
rect 86 15576 120 15592
rect 70 15484 136 15518
rect 70 15292 136 15326
rect 86 15218 120 15234
rect 86 15168 120 15184
rect 4094 15113 4122 15147
rect 4094 14873 4122 14907
rect 86 14836 120 14852
rect 86 14786 120 14802
rect 70 14694 136 14728
rect 70 14502 136 14536
rect 86 14428 120 14444
rect 86 14378 120 14394
rect 4094 14323 4122 14357
rect 4094 14083 4122 14117
rect 86 14046 120 14062
rect 86 13996 120 14012
rect 70 13904 136 13938
rect 70 13712 136 13746
rect 86 13638 120 13654
rect 86 13588 120 13604
rect 4094 13533 4122 13567
rect 4094 13293 4122 13327
rect 86 13256 120 13272
rect 86 13206 120 13222
rect 70 13114 136 13148
rect 70 12922 136 12956
rect 86 12848 120 12864
rect 86 12798 120 12814
rect 4094 12743 4122 12777
rect 4094 12503 4122 12537
rect 86 12466 120 12482
rect 86 12416 120 12432
rect 70 12324 136 12358
rect 70 12132 136 12166
rect 86 12058 120 12074
rect 86 12008 120 12024
rect 4094 11953 4122 11987
rect 4094 11713 4122 11747
rect 86 11676 120 11692
rect 86 11626 120 11642
rect 70 11534 136 11568
rect 70 11342 136 11376
rect 86 11268 120 11284
rect 86 11218 120 11234
rect 4094 11163 4122 11197
rect 4094 10923 4122 10957
rect 86 10886 120 10902
rect 86 10836 120 10852
rect 70 10744 136 10778
rect 70 10552 136 10586
rect 86 10478 120 10494
rect 86 10428 120 10444
rect 4094 10373 4122 10407
rect 4094 10133 4122 10167
rect 86 10096 120 10112
rect 86 10046 120 10062
rect 70 9954 136 9988
rect 70 9762 136 9796
rect 86 9688 120 9704
rect 86 9638 120 9654
rect 4094 9583 4122 9617
rect 4094 9343 4122 9377
rect 86 9306 120 9322
rect 86 9256 120 9272
rect 70 9164 136 9198
rect 70 8972 136 9006
rect 86 8898 120 8914
rect 86 8848 120 8864
rect 4094 8793 4122 8827
rect 4094 8553 4122 8587
rect 86 8516 120 8532
rect 86 8466 120 8482
rect 70 8374 136 8408
rect 70 8182 136 8216
rect 86 8108 120 8124
rect 86 8058 120 8074
rect 4094 8003 4122 8037
rect 4094 7763 4122 7797
rect 86 7726 120 7742
rect 86 7676 120 7692
rect 70 7584 136 7618
rect 70 7392 136 7426
rect 86 7318 120 7334
rect 86 7268 120 7284
rect 4094 7213 4122 7247
rect 4094 6973 4122 7007
rect 86 6936 120 6952
rect 86 6886 120 6902
rect 70 6794 136 6828
rect 70 6602 136 6636
rect 86 6528 120 6544
rect 86 6478 120 6494
rect 4094 6423 4122 6457
rect 4094 6183 4122 6217
rect 86 6146 120 6162
rect 86 6096 120 6112
rect 70 6004 136 6038
rect 70 5812 136 5846
rect 86 5738 120 5754
rect 86 5688 120 5704
rect 4094 5633 4122 5667
rect 4094 5393 4122 5427
rect 86 5356 120 5372
rect 86 5306 120 5322
rect 70 5214 136 5248
rect 70 5022 136 5056
rect 86 4948 120 4964
rect 86 4898 120 4914
rect 4094 4843 4122 4877
rect 4094 4603 4122 4637
rect 86 4566 120 4582
rect 86 4516 120 4532
rect 70 4424 136 4458
rect 70 4232 136 4266
rect 86 4158 120 4174
rect 86 4108 120 4124
rect 4094 4053 4122 4087
rect 4094 3813 4122 3847
rect 86 3776 120 3792
rect 86 3726 120 3742
rect 70 3634 136 3668
rect 70 3442 136 3476
rect 86 3368 120 3384
rect 86 3318 120 3334
rect 4094 3263 4122 3297
rect 4094 3023 4122 3057
rect 86 2986 120 3002
rect 86 2936 120 2952
rect 70 2844 136 2878
rect 70 2652 136 2686
rect 86 2578 120 2594
rect 86 2528 120 2544
rect 4094 2473 4122 2507
rect 4094 2233 4122 2267
rect 86 2196 120 2212
rect 86 2146 120 2162
rect 70 2054 136 2088
rect 70 1862 136 1896
rect 86 1788 120 1804
rect 86 1738 120 1754
rect 4094 1683 4122 1717
rect 4094 1443 4122 1477
rect 86 1406 120 1422
rect 86 1356 120 1372
rect 70 1264 136 1298
rect 70 1072 136 1106
rect 86 998 120 1014
rect 86 948 120 964
rect 4094 893 4122 927
rect 4094 653 4122 687
rect 86 616 120 632
rect 86 566 120 582
rect 70 474 136 508
rect 70 282 136 316
rect 86 208 120 224
rect 86 158 120 174
rect 4094 103 4122 137
<< viali >>
rect 86 50352 120 50386
rect 86 49944 120 49978
rect 86 49562 120 49596
rect 86 49154 120 49188
rect 86 48772 120 48806
rect 86 48364 120 48398
rect 86 47982 120 48016
rect 86 47574 120 47608
rect 86 47192 120 47226
rect 86 46784 120 46818
rect 86 46402 120 46436
rect 86 45994 120 46028
rect 86 45612 120 45646
rect 86 45204 120 45238
rect 86 44822 120 44856
rect 86 44414 120 44448
rect 86 44032 120 44066
rect 86 43624 120 43658
rect 86 43242 120 43276
rect 86 42834 120 42868
rect 86 42452 120 42486
rect 86 42044 120 42078
rect 86 41662 120 41696
rect 86 41254 120 41288
rect 86 40872 120 40906
rect 86 40464 120 40498
rect 86 40082 120 40116
rect 86 39674 120 39708
rect 86 39292 120 39326
rect 86 38884 120 38918
rect 86 38502 120 38536
rect 86 38094 120 38128
rect 86 37712 120 37746
rect 86 37304 120 37338
rect 86 36922 120 36956
rect 86 36514 120 36548
rect 86 36132 120 36166
rect 86 35724 120 35758
rect 86 35342 120 35376
rect 86 34934 120 34968
rect 86 34552 120 34586
rect 86 34144 120 34178
rect 86 33762 120 33796
rect 86 33354 120 33388
rect 86 32972 120 33006
rect 86 32564 120 32598
rect 86 32182 120 32216
rect 86 31774 120 31808
rect 86 31392 120 31426
rect 86 30984 120 31018
rect 86 30602 120 30636
rect 86 30194 120 30228
rect 86 29812 120 29846
rect 86 29404 120 29438
rect 86 29022 120 29056
rect 86 28614 120 28648
rect 86 28232 120 28266
rect 86 27824 120 27858
rect 86 27442 120 27476
rect 86 27034 120 27068
rect 86 26652 120 26686
rect 86 26244 120 26278
rect 86 25862 120 25896
rect 86 25454 120 25488
rect 86 25072 120 25106
rect 86 24664 120 24698
rect 86 24282 120 24316
rect 86 23874 120 23908
rect 86 23492 120 23526
rect 86 23084 120 23118
rect 86 22702 120 22736
rect 86 22294 120 22328
rect 86 21912 120 21946
rect 86 21504 120 21538
rect 86 21122 120 21156
rect 86 20714 120 20748
rect 86 20332 120 20366
rect 86 19924 120 19958
rect 86 19542 120 19576
rect 86 19134 120 19168
rect 86 18752 120 18786
rect 86 18344 120 18378
rect 86 17962 120 17996
rect 86 17554 120 17588
rect 86 17172 120 17206
rect 86 16764 120 16798
rect 86 16382 120 16416
rect 86 15974 120 16008
rect 86 15592 120 15626
rect 86 15184 120 15218
rect 86 14802 120 14836
rect 86 14394 120 14428
rect 86 14012 120 14046
rect 86 13604 120 13638
rect 86 13222 120 13256
rect 86 12814 120 12848
rect 86 12432 120 12466
rect 86 12024 120 12058
rect 86 11642 120 11676
rect 86 11234 120 11268
rect 86 10852 120 10886
rect 86 10444 120 10478
rect 86 10062 120 10096
rect 86 9654 120 9688
rect 86 9272 120 9306
rect 86 8864 120 8898
rect 86 8482 120 8516
rect 86 8074 120 8108
rect 86 7692 120 7726
rect 86 7284 120 7318
rect 86 6902 120 6936
rect 86 6494 120 6528
rect 86 6112 120 6146
rect 86 5704 120 5738
rect 86 5322 120 5356
rect 86 4914 120 4948
rect 86 4532 120 4566
rect 86 4124 120 4158
rect 86 3742 120 3776
rect 86 3334 120 3368
rect 86 2952 120 2986
rect 86 2544 120 2578
rect 86 2162 120 2196
rect 86 1754 120 1788
rect 86 1372 120 1406
rect 86 964 120 998
rect 86 582 120 616
rect 86 174 120 208
<< metal1 >>
rect 71 50343 77 50395
rect 129 50343 135 50395
rect 71 49935 77 49987
rect 129 49935 135 49987
rect 71 49553 77 49605
rect 129 49553 135 49605
rect 71 49145 77 49197
rect 129 49145 135 49197
rect 71 48763 77 48815
rect 129 48763 135 48815
rect 71 48355 77 48407
rect 129 48355 135 48407
rect 71 47973 77 48025
rect 129 47973 135 48025
rect 71 47565 77 47617
rect 129 47565 135 47617
rect 71 47183 77 47235
rect 129 47183 135 47235
rect 71 46775 77 46827
rect 129 46775 135 46827
rect 71 46393 77 46445
rect 129 46393 135 46445
rect 71 45985 77 46037
rect 129 45985 135 46037
rect 71 45603 77 45655
rect 129 45603 135 45655
rect 71 45195 77 45247
rect 129 45195 135 45247
rect 71 44813 77 44865
rect 129 44813 135 44865
rect 71 44405 77 44457
rect 129 44405 135 44457
rect 71 44023 77 44075
rect 129 44023 135 44075
rect 71 43615 77 43667
rect 129 43615 135 43667
rect 71 43233 77 43285
rect 129 43233 135 43285
rect 71 42825 77 42877
rect 129 42825 135 42877
rect 71 42443 77 42495
rect 129 42443 135 42495
rect 71 42035 77 42087
rect 129 42035 135 42087
rect 71 41653 77 41705
rect 129 41653 135 41705
rect 71 41245 77 41297
rect 129 41245 135 41297
rect 71 40863 77 40915
rect 129 40863 135 40915
rect 71 40455 77 40507
rect 129 40455 135 40507
rect 71 40073 77 40125
rect 129 40073 135 40125
rect 71 39665 77 39717
rect 129 39665 135 39717
rect 71 39283 77 39335
rect 129 39283 135 39335
rect 71 38875 77 38927
rect 129 38875 135 38927
rect 71 38493 77 38545
rect 129 38493 135 38545
rect 71 38085 77 38137
rect 129 38085 135 38137
rect 71 37703 77 37755
rect 129 37703 135 37755
rect 71 37295 77 37347
rect 129 37295 135 37347
rect 71 36913 77 36965
rect 129 36913 135 36965
rect 71 36505 77 36557
rect 129 36505 135 36557
rect 71 36123 77 36175
rect 129 36123 135 36175
rect 71 35715 77 35767
rect 129 35715 135 35767
rect 71 35333 77 35385
rect 129 35333 135 35385
rect 71 34925 77 34977
rect 129 34925 135 34977
rect 71 34543 77 34595
rect 129 34543 135 34595
rect 71 34135 77 34187
rect 129 34135 135 34187
rect 71 33753 77 33805
rect 129 33753 135 33805
rect 71 33345 77 33397
rect 129 33345 135 33397
rect 71 32963 77 33015
rect 129 32963 135 33015
rect 71 32555 77 32607
rect 129 32555 135 32607
rect 71 32173 77 32225
rect 129 32173 135 32225
rect 71 31765 77 31817
rect 129 31765 135 31817
rect 71 31383 77 31435
rect 129 31383 135 31435
rect 71 30975 77 31027
rect 129 30975 135 31027
rect 71 30593 77 30645
rect 129 30593 135 30645
rect 71 30185 77 30237
rect 129 30185 135 30237
rect 71 29803 77 29855
rect 129 29803 135 29855
rect 71 29395 77 29447
rect 129 29395 135 29447
rect 71 29013 77 29065
rect 129 29013 135 29065
rect 71 28605 77 28657
rect 129 28605 135 28657
rect 71 28223 77 28275
rect 129 28223 135 28275
rect 71 27815 77 27867
rect 129 27815 135 27867
rect 71 27433 77 27485
rect 129 27433 135 27485
rect 71 27025 77 27077
rect 129 27025 135 27077
rect 71 26643 77 26695
rect 129 26643 135 26695
rect 71 26235 77 26287
rect 129 26235 135 26287
rect 71 25853 77 25905
rect 129 25853 135 25905
rect 71 25445 77 25497
rect 129 25445 135 25497
rect 71 25063 77 25115
rect 129 25063 135 25115
rect 71 24655 77 24707
rect 129 24655 135 24707
rect 71 24273 77 24325
rect 129 24273 135 24325
rect 71 23865 77 23917
rect 129 23865 135 23917
rect 71 23483 77 23535
rect 129 23483 135 23535
rect 71 23075 77 23127
rect 129 23075 135 23127
rect 71 22693 77 22745
rect 129 22693 135 22745
rect 71 22285 77 22337
rect 129 22285 135 22337
rect 71 21903 77 21955
rect 129 21903 135 21955
rect 71 21495 77 21547
rect 129 21495 135 21547
rect 71 21113 77 21165
rect 129 21113 135 21165
rect 71 20705 77 20757
rect 129 20705 135 20757
rect 71 20323 77 20375
rect 129 20323 135 20375
rect 71 19915 77 19967
rect 129 19915 135 19967
rect 71 19533 77 19585
rect 129 19533 135 19585
rect 71 19125 77 19177
rect 129 19125 135 19177
rect 71 18743 77 18795
rect 129 18743 135 18795
rect 71 18335 77 18387
rect 129 18335 135 18387
rect 71 17953 77 18005
rect 129 17953 135 18005
rect 71 17545 77 17597
rect 129 17545 135 17597
rect 71 17163 77 17215
rect 129 17163 135 17215
rect 71 16755 77 16807
rect 129 16755 135 16807
rect 71 16373 77 16425
rect 129 16373 135 16425
rect 71 15965 77 16017
rect 129 15965 135 16017
rect 71 15583 77 15635
rect 129 15583 135 15635
rect 71 15175 77 15227
rect 129 15175 135 15227
rect 71 14793 77 14845
rect 129 14793 135 14845
rect 71 14385 77 14437
rect 129 14385 135 14437
rect 71 14003 77 14055
rect 129 14003 135 14055
rect 71 13595 77 13647
rect 129 13595 135 13647
rect 71 13213 77 13265
rect 129 13213 135 13265
rect 71 12805 77 12857
rect 129 12805 135 12857
rect 71 12423 77 12475
rect 129 12423 135 12475
rect 71 12015 77 12067
rect 129 12015 135 12067
rect 71 11633 77 11685
rect 129 11633 135 11685
rect 71 11225 77 11277
rect 129 11225 135 11277
rect 71 10843 77 10895
rect 129 10843 135 10895
rect 71 10435 77 10487
rect 129 10435 135 10487
rect 71 10053 77 10105
rect 129 10053 135 10105
rect 71 9645 77 9697
rect 129 9645 135 9697
rect 71 9263 77 9315
rect 129 9263 135 9315
rect 71 8855 77 8907
rect 129 8855 135 8907
rect 71 8473 77 8525
rect 129 8473 135 8525
rect 71 8065 77 8117
rect 129 8065 135 8117
rect 71 7683 77 7735
rect 129 7683 135 7735
rect 71 7275 77 7327
rect 129 7275 135 7327
rect 71 6893 77 6945
rect 129 6893 135 6945
rect 71 6485 77 6537
rect 129 6485 135 6537
rect 71 6103 77 6155
rect 129 6103 135 6155
rect 71 5695 77 5747
rect 129 5695 135 5747
rect 71 5313 77 5365
rect 129 5313 135 5365
rect 71 4905 77 4957
rect 129 4905 135 4957
rect 71 4523 77 4575
rect 129 4523 135 4575
rect 71 4115 77 4167
rect 129 4115 135 4167
rect 71 3733 77 3785
rect 129 3733 135 3785
rect 71 3325 77 3377
rect 129 3325 135 3377
rect 71 2943 77 2995
rect 129 2943 135 2995
rect 71 2535 77 2587
rect 129 2535 135 2587
rect 71 2153 77 2205
rect 129 2153 135 2205
rect 71 1745 77 1797
rect 129 1745 135 1797
rect 71 1363 77 1415
rect 129 1363 135 1415
rect 71 955 77 1007
rect 129 955 135 1007
rect 71 573 77 625
rect 129 573 135 625
rect 71 165 77 217
rect 129 165 135 217
rect 256 -30 284 50560
rect 681 -32 709 50560
rect 1724 0 1752 50560
rect 3372 0 3400 50560
<< via1 >>
rect 77 50386 129 50395
rect 77 50352 86 50386
rect 86 50352 120 50386
rect 120 50352 129 50386
rect 77 50343 129 50352
rect 77 49978 129 49987
rect 77 49944 86 49978
rect 86 49944 120 49978
rect 120 49944 129 49978
rect 77 49935 129 49944
rect 77 49596 129 49605
rect 77 49562 86 49596
rect 86 49562 120 49596
rect 120 49562 129 49596
rect 77 49553 129 49562
rect 77 49188 129 49197
rect 77 49154 86 49188
rect 86 49154 120 49188
rect 120 49154 129 49188
rect 77 49145 129 49154
rect 77 48806 129 48815
rect 77 48772 86 48806
rect 86 48772 120 48806
rect 120 48772 129 48806
rect 77 48763 129 48772
rect 77 48398 129 48407
rect 77 48364 86 48398
rect 86 48364 120 48398
rect 120 48364 129 48398
rect 77 48355 129 48364
rect 77 48016 129 48025
rect 77 47982 86 48016
rect 86 47982 120 48016
rect 120 47982 129 48016
rect 77 47973 129 47982
rect 77 47608 129 47617
rect 77 47574 86 47608
rect 86 47574 120 47608
rect 120 47574 129 47608
rect 77 47565 129 47574
rect 77 47226 129 47235
rect 77 47192 86 47226
rect 86 47192 120 47226
rect 120 47192 129 47226
rect 77 47183 129 47192
rect 77 46818 129 46827
rect 77 46784 86 46818
rect 86 46784 120 46818
rect 120 46784 129 46818
rect 77 46775 129 46784
rect 77 46436 129 46445
rect 77 46402 86 46436
rect 86 46402 120 46436
rect 120 46402 129 46436
rect 77 46393 129 46402
rect 77 46028 129 46037
rect 77 45994 86 46028
rect 86 45994 120 46028
rect 120 45994 129 46028
rect 77 45985 129 45994
rect 77 45646 129 45655
rect 77 45612 86 45646
rect 86 45612 120 45646
rect 120 45612 129 45646
rect 77 45603 129 45612
rect 77 45238 129 45247
rect 77 45204 86 45238
rect 86 45204 120 45238
rect 120 45204 129 45238
rect 77 45195 129 45204
rect 77 44856 129 44865
rect 77 44822 86 44856
rect 86 44822 120 44856
rect 120 44822 129 44856
rect 77 44813 129 44822
rect 77 44448 129 44457
rect 77 44414 86 44448
rect 86 44414 120 44448
rect 120 44414 129 44448
rect 77 44405 129 44414
rect 77 44066 129 44075
rect 77 44032 86 44066
rect 86 44032 120 44066
rect 120 44032 129 44066
rect 77 44023 129 44032
rect 77 43658 129 43667
rect 77 43624 86 43658
rect 86 43624 120 43658
rect 120 43624 129 43658
rect 77 43615 129 43624
rect 77 43276 129 43285
rect 77 43242 86 43276
rect 86 43242 120 43276
rect 120 43242 129 43276
rect 77 43233 129 43242
rect 77 42868 129 42877
rect 77 42834 86 42868
rect 86 42834 120 42868
rect 120 42834 129 42868
rect 77 42825 129 42834
rect 77 42486 129 42495
rect 77 42452 86 42486
rect 86 42452 120 42486
rect 120 42452 129 42486
rect 77 42443 129 42452
rect 77 42078 129 42087
rect 77 42044 86 42078
rect 86 42044 120 42078
rect 120 42044 129 42078
rect 77 42035 129 42044
rect 77 41696 129 41705
rect 77 41662 86 41696
rect 86 41662 120 41696
rect 120 41662 129 41696
rect 77 41653 129 41662
rect 77 41288 129 41297
rect 77 41254 86 41288
rect 86 41254 120 41288
rect 120 41254 129 41288
rect 77 41245 129 41254
rect 77 40906 129 40915
rect 77 40872 86 40906
rect 86 40872 120 40906
rect 120 40872 129 40906
rect 77 40863 129 40872
rect 77 40498 129 40507
rect 77 40464 86 40498
rect 86 40464 120 40498
rect 120 40464 129 40498
rect 77 40455 129 40464
rect 77 40116 129 40125
rect 77 40082 86 40116
rect 86 40082 120 40116
rect 120 40082 129 40116
rect 77 40073 129 40082
rect 77 39708 129 39717
rect 77 39674 86 39708
rect 86 39674 120 39708
rect 120 39674 129 39708
rect 77 39665 129 39674
rect 77 39326 129 39335
rect 77 39292 86 39326
rect 86 39292 120 39326
rect 120 39292 129 39326
rect 77 39283 129 39292
rect 77 38918 129 38927
rect 77 38884 86 38918
rect 86 38884 120 38918
rect 120 38884 129 38918
rect 77 38875 129 38884
rect 77 38536 129 38545
rect 77 38502 86 38536
rect 86 38502 120 38536
rect 120 38502 129 38536
rect 77 38493 129 38502
rect 77 38128 129 38137
rect 77 38094 86 38128
rect 86 38094 120 38128
rect 120 38094 129 38128
rect 77 38085 129 38094
rect 77 37746 129 37755
rect 77 37712 86 37746
rect 86 37712 120 37746
rect 120 37712 129 37746
rect 77 37703 129 37712
rect 77 37338 129 37347
rect 77 37304 86 37338
rect 86 37304 120 37338
rect 120 37304 129 37338
rect 77 37295 129 37304
rect 77 36956 129 36965
rect 77 36922 86 36956
rect 86 36922 120 36956
rect 120 36922 129 36956
rect 77 36913 129 36922
rect 77 36548 129 36557
rect 77 36514 86 36548
rect 86 36514 120 36548
rect 120 36514 129 36548
rect 77 36505 129 36514
rect 77 36166 129 36175
rect 77 36132 86 36166
rect 86 36132 120 36166
rect 120 36132 129 36166
rect 77 36123 129 36132
rect 77 35758 129 35767
rect 77 35724 86 35758
rect 86 35724 120 35758
rect 120 35724 129 35758
rect 77 35715 129 35724
rect 77 35376 129 35385
rect 77 35342 86 35376
rect 86 35342 120 35376
rect 120 35342 129 35376
rect 77 35333 129 35342
rect 77 34968 129 34977
rect 77 34934 86 34968
rect 86 34934 120 34968
rect 120 34934 129 34968
rect 77 34925 129 34934
rect 77 34586 129 34595
rect 77 34552 86 34586
rect 86 34552 120 34586
rect 120 34552 129 34586
rect 77 34543 129 34552
rect 77 34178 129 34187
rect 77 34144 86 34178
rect 86 34144 120 34178
rect 120 34144 129 34178
rect 77 34135 129 34144
rect 77 33796 129 33805
rect 77 33762 86 33796
rect 86 33762 120 33796
rect 120 33762 129 33796
rect 77 33753 129 33762
rect 77 33388 129 33397
rect 77 33354 86 33388
rect 86 33354 120 33388
rect 120 33354 129 33388
rect 77 33345 129 33354
rect 77 33006 129 33015
rect 77 32972 86 33006
rect 86 32972 120 33006
rect 120 32972 129 33006
rect 77 32963 129 32972
rect 77 32598 129 32607
rect 77 32564 86 32598
rect 86 32564 120 32598
rect 120 32564 129 32598
rect 77 32555 129 32564
rect 77 32216 129 32225
rect 77 32182 86 32216
rect 86 32182 120 32216
rect 120 32182 129 32216
rect 77 32173 129 32182
rect 77 31808 129 31817
rect 77 31774 86 31808
rect 86 31774 120 31808
rect 120 31774 129 31808
rect 77 31765 129 31774
rect 77 31426 129 31435
rect 77 31392 86 31426
rect 86 31392 120 31426
rect 120 31392 129 31426
rect 77 31383 129 31392
rect 77 31018 129 31027
rect 77 30984 86 31018
rect 86 30984 120 31018
rect 120 30984 129 31018
rect 77 30975 129 30984
rect 77 30636 129 30645
rect 77 30602 86 30636
rect 86 30602 120 30636
rect 120 30602 129 30636
rect 77 30593 129 30602
rect 77 30228 129 30237
rect 77 30194 86 30228
rect 86 30194 120 30228
rect 120 30194 129 30228
rect 77 30185 129 30194
rect 77 29846 129 29855
rect 77 29812 86 29846
rect 86 29812 120 29846
rect 120 29812 129 29846
rect 77 29803 129 29812
rect 77 29438 129 29447
rect 77 29404 86 29438
rect 86 29404 120 29438
rect 120 29404 129 29438
rect 77 29395 129 29404
rect 77 29056 129 29065
rect 77 29022 86 29056
rect 86 29022 120 29056
rect 120 29022 129 29056
rect 77 29013 129 29022
rect 77 28648 129 28657
rect 77 28614 86 28648
rect 86 28614 120 28648
rect 120 28614 129 28648
rect 77 28605 129 28614
rect 77 28266 129 28275
rect 77 28232 86 28266
rect 86 28232 120 28266
rect 120 28232 129 28266
rect 77 28223 129 28232
rect 77 27858 129 27867
rect 77 27824 86 27858
rect 86 27824 120 27858
rect 120 27824 129 27858
rect 77 27815 129 27824
rect 77 27476 129 27485
rect 77 27442 86 27476
rect 86 27442 120 27476
rect 120 27442 129 27476
rect 77 27433 129 27442
rect 77 27068 129 27077
rect 77 27034 86 27068
rect 86 27034 120 27068
rect 120 27034 129 27068
rect 77 27025 129 27034
rect 77 26686 129 26695
rect 77 26652 86 26686
rect 86 26652 120 26686
rect 120 26652 129 26686
rect 77 26643 129 26652
rect 77 26278 129 26287
rect 77 26244 86 26278
rect 86 26244 120 26278
rect 120 26244 129 26278
rect 77 26235 129 26244
rect 77 25896 129 25905
rect 77 25862 86 25896
rect 86 25862 120 25896
rect 120 25862 129 25896
rect 77 25853 129 25862
rect 77 25488 129 25497
rect 77 25454 86 25488
rect 86 25454 120 25488
rect 120 25454 129 25488
rect 77 25445 129 25454
rect 77 25106 129 25115
rect 77 25072 86 25106
rect 86 25072 120 25106
rect 120 25072 129 25106
rect 77 25063 129 25072
rect 77 24698 129 24707
rect 77 24664 86 24698
rect 86 24664 120 24698
rect 120 24664 129 24698
rect 77 24655 129 24664
rect 77 24316 129 24325
rect 77 24282 86 24316
rect 86 24282 120 24316
rect 120 24282 129 24316
rect 77 24273 129 24282
rect 77 23908 129 23917
rect 77 23874 86 23908
rect 86 23874 120 23908
rect 120 23874 129 23908
rect 77 23865 129 23874
rect 77 23526 129 23535
rect 77 23492 86 23526
rect 86 23492 120 23526
rect 120 23492 129 23526
rect 77 23483 129 23492
rect 77 23118 129 23127
rect 77 23084 86 23118
rect 86 23084 120 23118
rect 120 23084 129 23118
rect 77 23075 129 23084
rect 77 22736 129 22745
rect 77 22702 86 22736
rect 86 22702 120 22736
rect 120 22702 129 22736
rect 77 22693 129 22702
rect 77 22328 129 22337
rect 77 22294 86 22328
rect 86 22294 120 22328
rect 120 22294 129 22328
rect 77 22285 129 22294
rect 77 21946 129 21955
rect 77 21912 86 21946
rect 86 21912 120 21946
rect 120 21912 129 21946
rect 77 21903 129 21912
rect 77 21538 129 21547
rect 77 21504 86 21538
rect 86 21504 120 21538
rect 120 21504 129 21538
rect 77 21495 129 21504
rect 77 21156 129 21165
rect 77 21122 86 21156
rect 86 21122 120 21156
rect 120 21122 129 21156
rect 77 21113 129 21122
rect 77 20748 129 20757
rect 77 20714 86 20748
rect 86 20714 120 20748
rect 120 20714 129 20748
rect 77 20705 129 20714
rect 77 20366 129 20375
rect 77 20332 86 20366
rect 86 20332 120 20366
rect 120 20332 129 20366
rect 77 20323 129 20332
rect 77 19958 129 19967
rect 77 19924 86 19958
rect 86 19924 120 19958
rect 120 19924 129 19958
rect 77 19915 129 19924
rect 77 19576 129 19585
rect 77 19542 86 19576
rect 86 19542 120 19576
rect 120 19542 129 19576
rect 77 19533 129 19542
rect 77 19168 129 19177
rect 77 19134 86 19168
rect 86 19134 120 19168
rect 120 19134 129 19168
rect 77 19125 129 19134
rect 77 18786 129 18795
rect 77 18752 86 18786
rect 86 18752 120 18786
rect 120 18752 129 18786
rect 77 18743 129 18752
rect 77 18378 129 18387
rect 77 18344 86 18378
rect 86 18344 120 18378
rect 120 18344 129 18378
rect 77 18335 129 18344
rect 77 17996 129 18005
rect 77 17962 86 17996
rect 86 17962 120 17996
rect 120 17962 129 17996
rect 77 17953 129 17962
rect 77 17588 129 17597
rect 77 17554 86 17588
rect 86 17554 120 17588
rect 120 17554 129 17588
rect 77 17545 129 17554
rect 77 17206 129 17215
rect 77 17172 86 17206
rect 86 17172 120 17206
rect 120 17172 129 17206
rect 77 17163 129 17172
rect 77 16798 129 16807
rect 77 16764 86 16798
rect 86 16764 120 16798
rect 120 16764 129 16798
rect 77 16755 129 16764
rect 77 16416 129 16425
rect 77 16382 86 16416
rect 86 16382 120 16416
rect 120 16382 129 16416
rect 77 16373 129 16382
rect 77 16008 129 16017
rect 77 15974 86 16008
rect 86 15974 120 16008
rect 120 15974 129 16008
rect 77 15965 129 15974
rect 77 15626 129 15635
rect 77 15592 86 15626
rect 86 15592 120 15626
rect 120 15592 129 15626
rect 77 15583 129 15592
rect 77 15218 129 15227
rect 77 15184 86 15218
rect 86 15184 120 15218
rect 120 15184 129 15218
rect 77 15175 129 15184
rect 77 14836 129 14845
rect 77 14802 86 14836
rect 86 14802 120 14836
rect 120 14802 129 14836
rect 77 14793 129 14802
rect 77 14428 129 14437
rect 77 14394 86 14428
rect 86 14394 120 14428
rect 120 14394 129 14428
rect 77 14385 129 14394
rect 77 14046 129 14055
rect 77 14012 86 14046
rect 86 14012 120 14046
rect 120 14012 129 14046
rect 77 14003 129 14012
rect 77 13638 129 13647
rect 77 13604 86 13638
rect 86 13604 120 13638
rect 120 13604 129 13638
rect 77 13595 129 13604
rect 77 13256 129 13265
rect 77 13222 86 13256
rect 86 13222 120 13256
rect 120 13222 129 13256
rect 77 13213 129 13222
rect 77 12848 129 12857
rect 77 12814 86 12848
rect 86 12814 120 12848
rect 120 12814 129 12848
rect 77 12805 129 12814
rect 77 12466 129 12475
rect 77 12432 86 12466
rect 86 12432 120 12466
rect 120 12432 129 12466
rect 77 12423 129 12432
rect 77 12058 129 12067
rect 77 12024 86 12058
rect 86 12024 120 12058
rect 120 12024 129 12058
rect 77 12015 129 12024
rect 77 11676 129 11685
rect 77 11642 86 11676
rect 86 11642 120 11676
rect 120 11642 129 11676
rect 77 11633 129 11642
rect 77 11268 129 11277
rect 77 11234 86 11268
rect 86 11234 120 11268
rect 120 11234 129 11268
rect 77 11225 129 11234
rect 77 10886 129 10895
rect 77 10852 86 10886
rect 86 10852 120 10886
rect 120 10852 129 10886
rect 77 10843 129 10852
rect 77 10478 129 10487
rect 77 10444 86 10478
rect 86 10444 120 10478
rect 120 10444 129 10478
rect 77 10435 129 10444
rect 77 10096 129 10105
rect 77 10062 86 10096
rect 86 10062 120 10096
rect 120 10062 129 10096
rect 77 10053 129 10062
rect 77 9688 129 9697
rect 77 9654 86 9688
rect 86 9654 120 9688
rect 120 9654 129 9688
rect 77 9645 129 9654
rect 77 9306 129 9315
rect 77 9272 86 9306
rect 86 9272 120 9306
rect 120 9272 129 9306
rect 77 9263 129 9272
rect 77 8898 129 8907
rect 77 8864 86 8898
rect 86 8864 120 8898
rect 120 8864 129 8898
rect 77 8855 129 8864
rect 77 8516 129 8525
rect 77 8482 86 8516
rect 86 8482 120 8516
rect 120 8482 129 8516
rect 77 8473 129 8482
rect 77 8108 129 8117
rect 77 8074 86 8108
rect 86 8074 120 8108
rect 120 8074 129 8108
rect 77 8065 129 8074
rect 77 7726 129 7735
rect 77 7692 86 7726
rect 86 7692 120 7726
rect 120 7692 129 7726
rect 77 7683 129 7692
rect 77 7318 129 7327
rect 77 7284 86 7318
rect 86 7284 120 7318
rect 120 7284 129 7318
rect 77 7275 129 7284
rect 77 6936 129 6945
rect 77 6902 86 6936
rect 86 6902 120 6936
rect 120 6902 129 6936
rect 77 6893 129 6902
rect 77 6528 129 6537
rect 77 6494 86 6528
rect 86 6494 120 6528
rect 120 6494 129 6528
rect 77 6485 129 6494
rect 77 6146 129 6155
rect 77 6112 86 6146
rect 86 6112 120 6146
rect 120 6112 129 6146
rect 77 6103 129 6112
rect 77 5738 129 5747
rect 77 5704 86 5738
rect 86 5704 120 5738
rect 120 5704 129 5738
rect 77 5695 129 5704
rect 77 5356 129 5365
rect 77 5322 86 5356
rect 86 5322 120 5356
rect 120 5322 129 5356
rect 77 5313 129 5322
rect 77 4948 129 4957
rect 77 4914 86 4948
rect 86 4914 120 4948
rect 120 4914 129 4948
rect 77 4905 129 4914
rect 77 4566 129 4575
rect 77 4532 86 4566
rect 86 4532 120 4566
rect 120 4532 129 4566
rect 77 4523 129 4532
rect 77 4158 129 4167
rect 77 4124 86 4158
rect 86 4124 120 4158
rect 120 4124 129 4158
rect 77 4115 129 4124
rect 77 3776 129 3785
rect 77 3742 86 3776
rect 86 3742 120 3776
rect 120 3742 129 3776
rect 77 3733 129 3742
rect 77 3368 129 3377
rect 77 3334 86 3368
rect 86 3334 120 3368
rect 120 3334 129 3368
rect 77 3325 129 3334
rect 77 2986 129 2995
rect 77 2952 86 2986
rect 86 2952 120 2986
rect 120 2952 129 2986
rect 77 2943 129 2952
rect 77 2578 129 2587
rect 77 2544 86 2578
rect 86 2544 120 2578
rect 120 2544 129 2578
rect 77 2535 129 2544
rect 77 2196 129 2205
rect 77 2162 86 2196
rect 86 2162 120 2196
rect 120 2162 129 2196
rect 77 2153 129 2162
rect 77 1788 129 1797
rect 77 1754 86 1788
rect 86 1754 120 1788
rect 120 1754 129 1788
rect 77 1745 129 1754
rect 77 1406 129 1415
rect 77 1372 86 1406
rect 86 1372 120 1406
rect 120 1372 129 1406
rect 77 1363 129 1372
rect 77 998 129 1007
rect 77 964 86 998
rect 86 964 120 998
rect 120 964 129 998
rect 77 955 129 964
rect 77 616 129 625
rect 77 582 86 616
rect 86 582 120 616
rect 120 582 129 616
rect 77 573 129 582
rect 77 208 129 217
rect 77 174 86 208
rect 86 174 120 208
rect 120 174 129 208
rect 77 165 129 174
<< metal2 >>
rect 70 50401 98 50560
rect 70 50395 129 50401
rect 70 50343 77 50395
rect 70 50337 129 50343
rect 70 49993 98 50337
rect 70 49987 129 49993
rect 70 49935 77 49987
rect 70 49929 129 49935
rect 70 49611 98 49929
rect 70 49605 129 49611
rect 70 49553 77 49605
rect 70 49547 129 49553
rect 70 49203 98 49547
rect 70 49197 129 49203
rect 70 49145 77 49197
rect 70 49139 129 49145
rect 70 48821 98 49139
rect 70 48815 129 48821
rect 70 48763 77 48815
rect 70 48757 129 48763
rect 70 48413 98 48757
rect 70 48407 129 48413
rect 70 48355 77 48407
rect 70 48349 129 48355
rect 70 48031 98 48349
rect 70 48025 129 48031
rect 70 47973 77 48025
rect 70 47967 129 47973
rect 70 47623 98 47967
rect 70 47617 129 47623
rect 70 47565 77 47617
rect 70 47559 129 47565
rect 70 47241 98 47559
rect 70 47235 129 47241
rect 70 47183 77 47235
rect 70 47177 129 47183
rect 70 46833 98 47177
rect 70 46827 129 46833
rect 70 46775 77 46827
rect 70 46769 129 46775
rect 70 46451 98 46769
rect 70 46445 129 46451
rect 70 46393 77 46445
rect 70 46387 129 46393
rect 70 46043 98 46387
rect 70 46037 129 46043
rect 70 45985 77 46037
rect 70 45979 129 45985
rect 70 45661 98 45979
rect 70 45655 129 45661
rect 70 45603 77 45655
rect 70 45597 129 45603
rect 70 45253 98 45597
rect 70 45247 129 45253
rect 70 45195 77 45247
rect 70 45189 129 45195
rect 70 44871 98 45189
rect 70 44865 129 44871
rect 70 44813 77 44865
rect 70 44807 129 44813
rect 70 44463 98 44807
rect 70 44457 129 44463
rect 70 44405 77 44457
rect 70 44399 129 44405
rect 70 44081 98 44399
rect 70 44075 129 44081
rect 70 44023 77 44075
rect 70 44017 129 44023
rect 70 43673 98 44017
rect 70 43667 129 43673
rect 70 43615 77 43667
rect 70 43609 129 43615
rect 70 43291 98 43609
rect 70 43285 129 43291
rect 70 43233 77 43285
rect 70 43227 129 43233
rect 70 42883 98 43227
rect 70 42877 129 42883
rect 70 42825 77 42877
rect 70 42819 129 42825
rect 70 42501 98 42819
rect 70 42495 129 42501
rect 70 42443 77 42495
rect 70 42437 129 42443
rect 70 42093 98 42437
rect 70 42087 129 42093
rect 70 42035 77 42087
rect 70 42029 129 42035
rect 70 41711 98 42029
rect 70 41705 129 41711
rect 70 41653 77 41705
rect 70 41647 129 41653
rect 70 41303 98 41647
rect 70 41297 129 41303
rect 70 41245 77 41297
rect 70 41239 129 41245
rect 70 40921 98 41239
rect 70 40915 129 40921
rect 70 40863 77 40915
rect 70 40857 129 40863
rect 70 40513 98 40857
rect 70 40507 129 40513
rect 70 40455 77 40507
rect 70 40449 129 40455
rect 70 40131 98 40449
rect 70 40125 129 40131
rect 70 40073 77 40125
rect 70 40067 129 40073
rect 70 39723 98 40067
rect 70 39717 129 39723
rect 70 39665 77 39717
rect 70 39659 129 39665
rect 70 39341 98 39659
rect 70 39335 129 39341
rect 70 39283 77 39335
rect 70 39277 129 39283
rect 70 38933 98 39277
rect 70 38927 129 38933
rect 70 38875 77 38927
rect 70 38869 129 38875
rect 70 38551 98 38869
rect 70 38545 129 38551
rect 70 38493 77 38545
rect 70 38487 129 38493
rect 70 38143 98 38487
rect 70 38137 129 38143
rect 70 38085 77 38137
rect 70 38079 129 38085
rect 70 37761 98 38079
rect 70 37755 129 37761
rect 70 37703 77 37755
rect 70 37697 129 37703
rect 70 37353 98 37697
rect 70 37347 129 37353
rect 70 37295 77 37347
rect 70 37289 129 37295
rect 70 36971 98 37289
rect 70 36965 129 36971
rect 70 36913 77 36965
rect 70 36907 129 36913
rect 70 36563 98 36907
rect 70 36557 129 36563
rect 70 36505 77 36557
rect 70 36499 129 36505
rect 70 36181 98 36499
rect 70 36175 129 36181
rect 70 36123 77 36175
rect 70 36117 129 36123
rect 70 35773 98 36117
rect 70 35767 129 35773
rect 70 35715 77 35767
rect 70 35709 129 35715
rect 70 35391 98 35709
rect 70 35385 129 35391
rect 70 35333 77 35385
rect 70 35327 129 35333
rect 70 34983 98 35327
rect 70 34977 129 34983
rect 70 34925 77 34977
rect 70 34919 129 34925
rect 70 34601 98 34919
rect 70 34595 129 34601
rect 70 34543 77 34595
rect 70 34537 129 34543
rect 70 34193 98 34537
rect 70 34187 129 34193
rect 70 34135 77 34187
rect 70 34129 129 34135
rect 70 33811 98 34129
rect 70 33805 129 33811
rect 70 33753 77 33805
rect 70 33747 129 33753
rect 70 33403 98 33747
rect 70 33397 129 33403
rect 70 33345 77 33397
rect 70 33339 129 33345
rect 70 33021 98 33339
rect 70 33015 129 33021
rect 70 32963 77 33015
rect 70 32957 129 32963
rect 70 32613 98 32957
rect 70 32607 129 32613
rect 70 32555 77 32607
rect 70 32549 129 32555
rect 70 32231 98 32549
rect 70 32225 129 32231
rect 70 32173 77 32225
rect 70 32167 129 32173
rect 70 31823 98 32167
rect 70 31817 129 31823
rect 70 31765 77 31817
rect 70 31759 129 31765
rect 70 31441 98 31759
rect 70 31435 129 31441
rect 70 31383 77 31435
rect 70 31377 129 31383
rect 70 31033 98 31377
rect 70 31027 129 31033
rect 70 30975 77 31027
rect 70 30969 129 30975
rect 70 30651 98 30969
rect 70 30645 129 30651
rect 70 30593 77 30645
rect 70 30587 129 30593
rect 70 30243 98 30587
rect 70 30237 129 30243
rect 70 30185 77 30237
rect 70 30179 129 30185
rect 70 29861 98 30179
rect 70 29855 129 29861
rect 70 29803 77 29855
rect 70 29797 129 29803
rect 70 29453 98 29797
rect 70 29447 129 29453
rect 70 29395 77 29447
rect 70 29389 129 29395
rect 70 29071 98 29389
rect 70 29065 129 29071
rect 70 29013 77 29065
rect 70 29007 129 29013
rect 70 28663 98 29007
rect 70 28657 129 28663
rect 70 28605 77 28657
rect 70 28599 129 28605
rect 70 28281 98 28599
rect 70 28275 129 28281
rect 70 28223 77 28275
rect 70 28217 129 28223
rect 70 27873 98 28217
rect 70 27867 129 27873
rect 70 27815 77 27867
rect 70 27809 129 27815
rect 70 27491 98 27809
rect 70 27485 129 27491
rect 70 27433 77 27485
rect 70 27427 129 27433
rect 70 27083 98 27427
rect 70 27077 129 27083
rect 70 27025 77 27077
rect 70 27019 129 27025
rect 70 26701 98 27019
rect 70 26695 129 26701
rect 70 26643 77 26695
rect 70 26637 129 26643
rect 70 26293 98 26637
rect 70 26287 129 26293
rect 70 26235 77 26287
rect 70 26229 129 26235
rect 70 25911 98 26229
rect 70 25905 129 25911
rect 70 25853 77 25905
rect 70 25847 129 25853
rect 70 25503 98 25847
rect 70 25497 129 25503
rect 70 25445 77 25497
rect 70 25439 129 25445
rect 70 25121 98 25439
rect 70 25115 129 25121
rect 70 25063 77 25115
rect 70 25057 129 25063
rect 70 24713 98 25057
rect 70 24707 129 24713
rect 70 24655 77 24707
rect 70 24649 129 24655
rect 70 24331 98 24649
rect 70 24325 129 24331
rect 70 24273 77 24325
rect 70 24267 129 24273
rect 70 23923 98 24267
rect 70 23917 129 23923
rect 70 23865 77 23917
rect 70 23859 129 23865
rect 70 23541 98 23859
rect 70 23535 129 23541
rect 70 23483 77 23535
rect 70 23477 129 23483
rect 70 23133 98 23477
rect 70 23127 129 23133
rect 70 23075 77 23127
rect 70 23069 129 23075
rect 70 22751 98 23069
rect 70 22745 129 22751
rect 70 22693 77 22745
rect 70 22687 129 22693
rect 70 22343 98 22687
rect 70 22337 129 22343
rect 70 22285 77 22337
rect 70 22279 129 22285
rect 70 21961 98 22279
rect 70 21955 129 21961
rect 70 21903 77 21955
rect 70 21897 129 21903
rect 70 21553 98 21897
rect 70 21547 129 21553
rect 70 21495 77 21547
rect 70 21489 129 21495
rect 70 21171 98 21489
rect 70 21165 129 21171
rect 70 21113 77 21165
rect 70 21107 129 21113
rect 70 20763 98 21107
rect 70 20757 129 20763
rect 70 20705 77 20757
rect 70 20699 129 20705
rect 70 20381 98 20699
rect 70 20375 129 20381
rect 70 20323 77 20375
rect 70 20317 129 20323
rect 70 19973 98 20317
rect 70 19967 129 19973
rect 70 19915 77 19967
rect 70 19909 129 19915
rect 70 19591 98 19909
rect 70 19585 129 19591
rect 70 19533 77 19585
rect 70 19527 129 19533
rect 70 19183 98 19527
rect 70 19177 129 19183
rect 70 19125 77 19177
rect 70 19119 129 19125
rect 70 18801 98 19119
rect 70 18795 129 18801
rect 70 18743 77 18795
rect 70 18737 129 18743
rect 70 18393 98 18737
rect 70 18387 129 18393
rect 70 18335 77 18387
rect 70 18329 129 18335
rect 70 18011 98 18329
rect 70 18005 129 18011
rect 70 17953 77 18005
rect 70 17947 129 17953
rect 70 17603 98 17947
rect 70 17597 129 17603
rect 70 17545 77 17597
rect 70 17539 129 17545
rect 70 17221 98 17539
rect 70 17215 129 17221
rect 70 17163 77 17215
rect 70 17157 129 17163
rect 70 16813 98 17157
rect 70 16807 129 16813
rect 70 16755 77 16807
rect 70 16749 129 16755
rect 70 16431 98 16749
rect 70 16425 129 16431
rect 70 16373 77 16425
rect 70 16367 129 16373
rect 70 16023 98 16367
rect 70 16017 129 16023
rect 70 15965 77 16017
rect 70 15959 129 15965
rect 70 15641 98 15959
rect 70 15635 129 15641
rect 70 15583 77 15635
rect 70 15577 129 15583
rect 70 15233 98 15577
rect 70 15227 129 15233
rect 70 15175 77 15227
rect 70 15169 129 15175
rect 70 14851 98 15169
rect 70 14845 129 14851
rect 70 14793 77 14845
rect 70 14787 129 14793
rect 70 14443 98 14787
rect 70 14437 129 14443
rect 70 14385 77 14437
rect 70 14379 129 14385
rect 70 14061 98 14379
rect 70 14055 129 14061
rect 70 14003 77 14055
rect 70 13997 129 14003
rect 70 13653 98 13997
rect 70 13647 129 13653
rect 70 13595 77 13647
rect 70 13589 129 13595
rect 70 13271 98 13589
rect 70 13265 129 13271
rect 70 13213 77 13265
rect 70 13207 129 13213
rect 70 12863 98 13207
rect 70 12857 129 12863
rect 70 12805 77 12857
rect 70 12799 129 12805
rect 70 12481 98 12799
rect 70 12475 129 12481
rect 70 12423 77 12475
rect 70 12417 129 12423
rect 70 12073 98 12417
rect 70 12067 129 12073
rect 70 12015 77 12067
rect 70 12009 129 12015
rect 70 11691 98 12009
rect 70 11685 129 11691
rect 70 11633 77 11685
rect 70 11627 129 11633
rect 70 11283 98 11627
rect 70 11277 129 11283
rect 70 11225 77 11277
rect 70 11219 129 11225
rect 70 10901 98 11219
rect 70 10895 129 10901
rect 70 10843 77 10895
rect 70 10837 129 10843
rect 70 10493 98 10837
rect 70 10487 129 10493
rect 70 10435 77 10487
rect 70 10429 129 10435
rect 70 10111 98 10429
rect 70 10105 129 10111
rect 70 10053 77 10105
rect 70 10047 129 10053
rect 70 9703 98 10047
rect 70 9697 129 9703
rect 70 9645 77 9697
rect 70 9639 129 9645
rect 70 9321 98 9639
rect 70 9315 129 9321
rect 70 9263 77 9315
rect 70 9257 129 9263
rect 70 8913 98 9257
rect 70 8907 129 8913
rect 70 8855 77 8907
rect 70 8849 129 8855
rect 70 8531 98 8849
rect 70 8525 129 8531
rect 70 8473 77 8525
rect 70 8467 129 8473
rect 70 8123 98 8467
rect 70 8117 129 8123
rect 70 8065 77 8117
rect 70 8059 129 8065
rect 70 7741 98 8059
rect 70 7735 129 7741
rect 70 7683 77 7735
rect 70 7677 129 7683
rect 70 7333 98 7677
rect 70 7327 129 7333
rect 70 7275 77 7327
rect 70 7269 129 7275
rect 70 6951 98 7269
rect 70 6945 129 6951
rect 70 6893 77 6945
rect 70 6887 129 6893
rect 70 6543 98 6887
rect 70 6537 129 6543
rect 70 6485 77 6537
rect 70 6479 129 6485
rect 70 6161 98 6479
rect 70 6155 129 6161
rect 70 6103 77 6155
rect 70 6097 129 6103
rect 70 5753 98 6097
rect 70 5747 129 5753
rect 70 5695 77 5747
rect 70 5689 129 5695
rect 70 5371 98 5689
rect 70 5365 129 5371
rect 70 5313 77 5365
rect 70 5307 129 5313
rect 70 4963 98 5307
rect 70 4957 129 4963
rect 70 4905 77 4957
rect 70 4899 129 4905
rect 70 4581 98 4899
rect 70 4575 129 4581
rect 70 4523 77 4575
rect 70 4517 129 4523
rect 70 4173 98 4517
rect 70 4167 129 4173
rect 70 4115 77 4167
rect 70 4109 129 4115
rect 70 3791 98 4109
rect 70 3785 129 3791
rect 70 3733 77 3785
rect 70 3727 129 3733
rect 70 3383 98 3727
rect 70 3377 129 3383
rect 70 3325 77 3377
rect 70 3319 129 3325
rect 70 3001 98 3319
rect 70 2995 129 3001
rect 70 2943 77 2995
rect 70 2937 129 2943
rect 70 2593 98 2937
rect 70 2587 129 2593
rect 70 2535 77 2587
rect 70 2529 129 2535
rect 70 2211 98 2529
rect 70 2205 129 2211
rect 70 2153 77 2205
rect 70 2147 129 2153
rect 70 1803 98 2147
rect 70 1797 129 1803
rect 70 1745 77 1797
rect 70 1739 129 1745
rect 70 1421 98 1739
rect 70 1415 129 1421
rect 70 1363 77 1415
rect 70 1357 129 1363
rect 70 1013 98 1357
rect 70 1007 129 1013
rect 70 955 77 1007
rect 70 949 129 955
rect 70 631 98 949
rect 70 625 129 631
rect 70 573 77 625
rect 70 567 129 573
rect 70 223 98 567
rect 70 217 129 223
rect 70 165 77 217
rect 70 159 129 165
rect 70 0 98 159
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_0
timestamp 1644511149
transform 1 0 74 0 1 12416
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_1
timestamp 1644511149
transform 1 0 74 0 1 12008
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_2
timestamp 1644511149
transform 1 0 74 0 1 11626
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_3
timestamp 1644511149
transform 1 0 74 0 1 11218
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_4
timestamp 1644511149
transform 1 0 74 0 1 10836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_5
timestamp 1644511149
transform 1 0 74 0 1 10428
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_6
timestamp 1644511149
transform 1 0 74 0 1 10046
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_7
timestamp 1644511149
transform 1 0 74 0 1 9638
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_8
timestamp 1644511149
transform 1 0 74 0 1 9256
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_9
timestamp 1644511149
transform 1 0 74 0 1 8848
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_10
timestamp 1644511149
transform 1 0 74 0 1 8466
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_11
timestamp 1644511149
transform 1 0 74 0 1 8058
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_12
timestamp 1644511149
transform 1 0 74 0 1 7676
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_13
timestamp 1644511149
transform 1 0 74 0 1 7268
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_14
timestamp 1644511149
transform 1 0 74 0 1 6886
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_15
timestamp 1644511149
transform 1 0 74 0 1 6478
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_16
timestamp 1644511149
transform 1 0 74 0 1 6096
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_17
timestamp 1644511149
transform 1 0 74 0 1 5688
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_18
timestamp 1644511149
transform 1 0 74 0 1 5306
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_19
timestamp 1644511149
transform 1 0 74 0 1 4898
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_20
timestamp 1644511149
transform 1 0 74 0 1 4516
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_21
timestamp 1644511149
transform 1 0 74 0 1 4108
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_22
timestamp 1644511149
transform 1 0 74 0 1 3726
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_23
timestamp 1644511149
transform 1 0 74 0 1 3318
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_24
timestamp 1644511149
transform 1 0 74 0 1 2936
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_25
timestamp 1644511149
transform 1 0 74 0 1 2528
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_26
timestamp 1644511149
transform 1 0 74 0 1 2146
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_27
timestamp 1644511149
transform 1 0 74 0 1 1738
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_28
timestamp 1644511149
transform 1 0 74 0 1 1356
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_29
timestamp 1644511149
transform 1 0 74 0 1 948
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_30
timestamp 1644511149
transform 1 0 74 0 1 566
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_31
timestamp 1644511149
transform 1 0 74 0 1 158
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_32
timestamp 1644511149
transform 1 0 74 0 1 12798
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_33
timestamp 1644511149
transform 1 0 74 0 1 13206
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_34
timestamp 1644511149
transform 1 0 74 0 1 25056
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_35
timestamp 1644511149
transform 1 0 74 0 1 24648
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_36
timestamp 1644511149
transform 1 0 74 0 1 24266
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_37
timestamp 1644511149
transform 1 0 74 0 1 23858
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_38
timestamp 1644511149
transform 1 0 74 0 1 23476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_39
timestamp 1644511149
transform 1 0 74 0 1 23068
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_40
timestamp 1644511149
transform 1 0 74 0 1 22686
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_41
timestamp 1644511149
transform 1 0 74 0 1 22278
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_42
timestamp 1644511149
transform 1 0 74 0 1 21896
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_43
timestamp 1644511149
transform 1 0 74 0 1 21488
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_44
timestamp 1644511149
transform 1 0 74 0 1 21106
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_45
timestamp 1644511149
transform 1 0 74 0 1 20698
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_46
timestamp 1644511149
transform 1 0 74 0 1 20316
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_47
timestamp 1644511149
transform 1 0 74 0 1 19908
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_48
timestamp 1644511149
transform 1 0 74 0 1 19526
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_49
timestamp 1644511149
transform 1 0 74 0 1 19118
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_50
timestamp 1644511149
transform 1 0 74 0 1 18736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_51
timestamp 1644511149
transform 1 0 74 0 1 18328
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_52
timestamp 1644511149
transform 1 0 74 0 1 17946
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_53
timestamp 1644511149
transform 1 0 74 0 1 17538
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_54
timestamp 1644511149
transform 1 0 74 0 1 17156
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_55
timestamp 1644511149
transform 1 0 74 0 1 16748
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_56
timestamp 1644511149
transform 1 0 74 0 1 16366
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_57
timestamp 1644511149
transform 1 0 74 0 1 15958
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_58
timestamp 1644511149
transform 1 0 74 0 1 15576
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_59
timestamp 1644511149
transform 1 0 74 0 1 15168
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_60
timestamp 1644511149
transform 1 0 74 0 1 14786
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_61
timestamp 1644511149
transform 1 0 74 0 1 14378
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_62
timestamp 1644511149
transform 1 0 74 0 1 13996
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_63
timestamp 1644511149
transform 1 0 74 0 1 13588
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_64
timestamp 1644511149
transform 1 0 74 0 1 31758
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_65
timestamp 1644511149
transform 1 0 74 0 1 31376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_66
timestamp 1644511149
transform 1 0 74 0 1 30968
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_67
timestamp 1644511149
transform 1 0 74 0 1 30586
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_68
timestamp 1644511149
transform 1 0 74 0 1 30178
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_69
timestamp 1644511149
transform 1 0 74 0 1 29796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_70
timestamp 1644511149
transform 1 0 74 0 1 29388
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_71
timestamp 1644511149
transform 1 0 74 0 1 29006
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_72
timestamp 1644511149
transform 1 0 74 0 1 28598
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_73
timestamp 1644511149
transform 1 0 74 0 1 28216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_74
timestamp 1644511149
transform 1 0 74 0 1 27808
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_75
timestamp 1644511149
transform 1 0 74 0 1 27426
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_76
timestamp 1644511149
transform 1 0 74 0 1 27018
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_77
timestamp 1644511149
transform 1 0 74 0 1 26636
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_78
timestamp 1644511149
transform 1 0 74 0 1 26228
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_79
timestamp 1644511149
transform 1 0 74 0 1 25846
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_80
timestamp 1644511149
transform 1 0 74 0 1 25438
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_81
timestamp 1644511149
transform 1 0 74 0 1 37696
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_82
timestamp 1644511149
transform 1 0 74 0 1 37288
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_83
timestamp 1644511149
transform 1 0 74 0 1 36906
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_84
timestamp 1644511149
transform 1 0 74 0 1 36498
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_85
timestamp 1644511149
transform 1 0 74 0 1 36116
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_86
timestamp 1644511149
transform 1 0 74 0 1 35708
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_87
timestamp 1644511149
transform 1 0 74 0 1 35326
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_88
timestamp 1644511149
transform 1 0 74 0 1 34918
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_89
timestamp 1644511149
transform 1 0 74 0 1 34536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_90
timestamp 1644511149
transform 1 0 74 0 1 34128
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_91
timestamp 1644511149
transform 1 0 74 0 1 33746
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_92
timestamp 1644511149
transform 1 0 74 0 1 33338
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_93
timestamp 1644511149
transform 1 0 74 0 1 32956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_94
timestamp 1644511149
transform 1 0 74 0 1 32548
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_95
timestamp 1644511149
transform 1 0 74 0 1 32166
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_96
timestamp 1644511149
transform 1 0 74 0 1 50336
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_97
timestamp 1644511149
transform 1 0 74 0 1 49928
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_98
timestamp 1644511149
transform 1 0 74 0 1 49546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_99
timestamp 1644511149
transform 1 0 74 0 1 49138
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_100
timestamp 1644511149
transform 1 0 74 0 1 48756
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_101
timestamp 1644511149
transform 1 0 74 0 1 48348
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_102
timestamp 1644511149
transform 1 0 74 0 1 47966
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_103
timestamp 1644511149
transform 1 0 74 0 1 47558
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_104
timestamp 1644511149
transform 1 0 74 0 1 47176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_105
timestamp 1644511149
transform 1 0 74 0 1 46768
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_106
timestamp 1644511149
transform 1 0 74 0 1 46386
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_107
timestamp 1644511149
transform 1 0 74 0 1 45978
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_108
timestamp 1644511149
transform 1 0 74 0 1 45596
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_109
timestamp 1644511149
transform 1 0 74 0 1 45188
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_110
timestamp 1644511149
transform 1 0 74 0 1 44806
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_111
timestamp 1644511149
transform 1 0 74 0 1 44398
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_112
timestamp 1644511149
transform 1 0 74 0 1 44016
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_113
timestamp 1644511149
transform 1 0 74 0 1 43608
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_114
timestamp 1644511149
transform 1 0 74 0 1 43226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_115
timestamp 1644511149
transform 1 0 74 0 1 42818
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_116
timestamp 1644511149
transform 1 0 74 0 1 42436
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_117
timestamp 1644511149
transform 1 0 74 0 1 42028
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_118
timestamp 1644511149
transform 1 0 74 0 1 41646
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_119
timestamp 1644511149
transform 1 0 74 0 1 41238
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_120
timestamp 1644511149
transform 1 0 74 0 1 40856
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_121
timestamp 1644511149
transform 1 0 74 0 1 40448
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_122
timestamp 1644511149
transform 1 0 74 0 1 40066
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_123
timestamp 1644511149
transform 1 0 74 0 1 39658
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_124
timestamp 1644511149
transform 1 0 74 0 1 39276
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_125
timestamp 1644511149
transform 1 0 74 0 1 38868
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_126
timestamp 1644511149
transform 1 0 74 0 1 38486
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_14  sky130_sram_1kbyte_1rw1r_32x256_8_contact_14_127
timestamp 1644511149
transform 1 0 74 0 1 38078
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_0
timestamp 1644511149
transform 1 0 71 0 1 12417
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_1
timestamp 1644511149
transform 1 0 71 0 1 12009
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_2
timestamp 1644511149
transform 1 0 71 0 1 11627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_3
timestamp 1644511149
transform 1 0 71 0 1 11219
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_4
timestamp 1644511149
transform 1 0 71 0 1 10837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_5
timestamp 1644511149
transform 1 0 71 0 1 10429
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_6
timestamp 1644511149
transform 1 0 71 0 1 10047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_7
timestamp 1644511149
transform 1 0 71 0 1 9639
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_8
timestamp 1644511149
transform 1 0 71 0 1 9257
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_9
timestamp 1644511149
transform 1 0 71 0 1 8849
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_10
timestamp 1644511149
transform 1 0 71 0 1 8467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_11
timestamp 1644511149
transform 1 0 71 0 1 8059
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_12
timestamp 1644511149
transform 1 0 71 0 1 7677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_13
timestamp 1644511149
transform 1 0 71 0 1 7269
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_14
timestamp 1644511149
transform 1 0 71 0 1 6887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_15
timestamp 1644511149
transform 1 0 71 0 1 6479
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_16
timestamp 1644511149
transform 1 0 71 0 1 6097
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_17
timestamp 1644511149
transform 1 0 71 0 1 5689
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_18
timestamp 1644511149
transform 1 0 71 0 1 5307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_19
timestamp 1644511149
transform 1 0 71 0 1 4899
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_20
timestamp 1644511149
transform 1 0 71 0 1 4517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_21
timestamp 1644511149
transform 1 0 71 0 1 4109
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_22
timestamp 1644511149
transform 1 0 71 0 1 3727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_23
timestamp 1644511149
transform 1 0 71 0 1 3319
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_24
timestamp 1644511149
transform 1 0 71 0 1 2937
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_25
timestamp 1644511149
transform 1 0 71 0 1 2529
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_26
timestamp 1644511149
transform 1 0 71 0 1 2147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_27
timestamp 1644511149
transform 1 0 71 0 1 1739
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_28
timestamp 1644511149
transform 1 0 71 0 1 1357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_29
timestamp 1644511149
transform 1 0 71 0 1 949
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_30
timestamp 1644511149
transform 1 0 71 0 1 567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_31
timestamp 1644511149
transform 1 0 71 0 1 159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_32
timestamp 1644511149
transform 1 0 71 0 1 12799
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_33
timestamp 1644511149
transform 1 0 71 0 1 25057
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_34
timestamp 1644511149
transform 1 0 71 0 1 24649
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_35
timestamp 1644511149
transform 1 0 71 0 1 24267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_36
timestamp 1644511149
transform 1 0 71 0 1 23859
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_37
timestamp 1644511149
transform 1 0 71 0 1 23477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_38
timestamp 1644511149
transform 1 0 71 0 1 23069
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_39
timestamp 1644511149
transform 1 0 71 0 1 22687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_40
timestamp 1644511149
transform 1 0 71 0 1 22279
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_41
timestamp 1644511149
transform 1 0 71 0 1 21897
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_42
timestamp 1644511149
transform 1 0 71 0 1 21489
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_43
timestamp 1644511149
transform 1 0 71 0 1 21107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_44
timestamp 1644511149
transform 1 0 71 0 1 20699
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_45
timestamp 1644511149
transform 1 0 71 0 1 20317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_46
timestamp 1644511149
transform 1 0 71 0 1 19909
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_47
timestamp 1644511149
transform 1 0 71 0 1 19527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_48
timestamp 1644511149
transform 1 0 71 0 1 19119
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_49
timestamp 1644511149
transform 1 0 71 0 1 18737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_50
timestamp 1644511149
transform 1 0 71 0 1 18329
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_51
timestamp 1644511149
transform 1 0 71 0 1 17947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_52
timestamp 1644511149
transform 1 0 71 0 1 17539
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_53
timestamp 1644511149
transform 1 0 71 0 1 17157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_54
timestamp 1644511149
transform 1 0 71 0 1 16749
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_55
timestamp 1644511149
transform 1 0 71 0 1 16367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_56
timestamp 1644511149
transform 1 0 71 0 1 15959
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_57
timestamp 1644511149
transform 1 0 71 0 1 15577
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_58
timestamp 1644511149
transform 1 0 71 0 1 15169
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_59
timestamp 1644511149
transform 1 0 71 0 1 14787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_60
timestamp 1644511149
transform 1 0 71 0 1 14379
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_61
timestamp 1644511149
transform 1 0 71 0 1 13997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_62
timestamp 1644511149
transform 1 0 71 0 1 13589
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_63
timestamp 1644511149
transform 1 0 71 0 1 13207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_64
timestamp 1644511149
transform 1 0 71 0 1 31759
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_65
timestamp 1644511149
transform 1 0 71 0 1 31377
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_66
timestamp 1644511149
transform 1 0 71 0 1 30969
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_67
timestamp 1644511149
transform 1 0 71 0 1 30587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_68
timestamp 1644511149
transform 1 0 71 0 1 30179
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_69
timestamp 1644511149
transform 1 0 71 0 1 29797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_70
timestamp 1644511149
transform 1 0 71 0 1 29389
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_71
timestamp 1644511149
transform 1 0 71 0 1 29007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_72
timestamp 1644511149
transform 1 0 71 0 1 28599
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_73
timestamp 1644511149
transform 1 0 71 0 1 28217
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_74
timestamp 1644511149
transform 1 0 71 0 1 27809
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_75
timestamp 1644511149
transform 1 0 71 0 1 27427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_76
timestamp 1644511149
transform 1 0 71 0 1 27019
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_77
timestamp 1644511149
transform 1 0 71 0 1 26637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_78
timestamp 1644511149
transform 1 0 71 0 1 26229
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_79
timestamp 1644511149
transform 1 0 71 0 1 25847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_80
timestamp 1644511149
transform 1 0 71 0 1 25439
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_81
timestamp 1644511149
transform 1 0 71 0 1 37697
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_82
timestamp 1644511149
transform 1 0 71 0 1 37289
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_83
timestamp 1644511149
transform 1 0 71 0 1 36907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_84
timestamp 1644511149
transform 1 0 71 0 1 36499
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_85
timestamp 1644511149
transform 1 0 71 0 1 36117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_86
timestamp 1644511149
transform 1 0 71 0 1 35709
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_87
timestamp 1644511149
transform 1 0 71 0 1 35327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_88
timestamp 1644511149
transform 1 0 71 0 1 34919
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_89
timestamp 1644511149
transform 1 0 71 0 1 34537
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_90
timestamp 1644511149
transform 1 0 71 0 1 34129
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_91
timestamp 1644511149
transform 1 0 71 0 1 33747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_92
timestamp 1644511149
transform 1 0 71 0 1 33339
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_93
timestamp 1644511149
transform 1 0 71 0 1 32957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_94
timestamp 1644511149
transform 1 0 71 0 1 32549
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_95
timestamp 1644511149
transform 1 0 71 0 1 32167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_96
timestamp 1644511149
transform 1 0 71 0 1 50337
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_97
timestamp 1644511149
transform 1 0 71 0 1 49929
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_98
timestamp 1644511149
transform 1 0 71 0 1 49547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_99
timestamp 1644511149
transform 1 0 71 0 1 49139
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_100
timestamp 1644511149
transform 1 0 71 0 1 48757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_101
timestamp 1644511149
transform 1 0 71 0 1 48349
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_102
timestamp 1644511149
transform 1 0 71 0 1 47967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_103
timestamp 1644511149
transform 1 0 71 0 1 47559
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_104
timestamp 1644511149
transform 1 0 71 0 1 47177
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_105
timestamp 1644511149
transform 1 0 71 0 1 46769
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_106
timestamp 1644511149
transform 1 0 71 0 1 46387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_107
timestamp 1644511149
transform 1 0 71 0 1 45979
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_108
timestamp 1644511149
transform 1 0 71 0 1 45597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_109
timestamp 1644511149
transform 1 0 71 0 1 45189
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_110
timestamp 1644511149
transform 1 0 71 0 1 44807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_111
timestamp 1644511149
transform 1 0 71 0 1 44399
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_112
timestamp 1644511149
transform 1 0 71 0 1 44017
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_113
timestamp 1644511149
transform 1 0 71 0 1 43609
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_114
timestamp 1644511149
transform 1 0 71 0 1 43227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_115
timestamp 1644511149
transform 1 0 71 0 1 42819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_116
timestamp 1644511149
transform 1 0 71 0 1 42437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_117
timestamp 1644511149
transform 1 0 71 0 1 42029
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_118
timestamp 1644511149
transform 1 0 71 0 1 41647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_119
timestamp 1644511149
transform 1 0 71 0 1 41239
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_120
timestamp 1644511149
transform 1 0 71 0 1 40857
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_121
timestamp 1644511149
transform 1 0 71 0 1 40449
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_122
timestamp 1644511149
transform 1 0 71 0 1 40067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_123
timestamp 1644511149
transform 1 0 71 0 1 39659
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_124
timestamp 1644511149
transform 1 0 71 0 1 39277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_125
timestamp 1644511149
transform 1 0 71 0 1 38869
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_126
timestamp 1644511149
transform 1 0 71 0 1 38487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_contact_19  sky130_sram_1kbyte_1rw1r_32x256_8_contact_19_127
timestamp 1644511149
transform 1 0 71 0 1 38079
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_0
timestamp 1644511149
transform 1 0 0 0 -1 2370
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_1
timestamp 1644511149
transform 1 0 0 0 -1 790
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_2
timestamp 1644511149
transform 1 0 0 0 1 0
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_3
timestamp 1644511149
transform 1 0 0 0 1 1580
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_4
timestamp 1644511149
transform 1 0 0 0 -1 1580
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_5
timestamp 1644511149
transform 1 0 0 0 1 790
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_6
timestamp 1644511149
transform 1 0 0 0 1 11850
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_7
timestamp 1644511149
transform 1 0 0 0 -1 11850
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_8
timestamp 1644511149
transform 1 0 0 0 1 11060
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_9
timestamp 1644511149
transform 1 0 0 0 -1 11060
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_10
timestamp 1644511149
transform 1 0 0 0 1 10270
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_11
timestamp 1644511149
transform 1 0 0 0 -1 10270
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_12
timestamp 1644511149
transform 1 0 0 0 1 9480
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_13
timestamp 1644511149
transform 1 0 0 0 -1 9480
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_14
timestamp 1644511149
transform 1 0 0 0 1 8690
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_15
timestamp 1644511149
transform 1 0 0 0 -1 8690
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_16
timestamp 1644511149
transform 1 0 0 0 1 7900
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_17
timestamp 1644511149
transform 1 0 0 0 -1 7900
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_18
timestamp 1644511149
transform 1 0 0 0 1 7110
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_19
timestamp 1644511149
transform 1 0 0 0 -1 7110
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_20
timestamp 1644511149
transform 1 0 0 0 1 6320
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_21
timestamp 1644511149
transform 1 0 0 0 -1 6320
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_22
timestamp 1644511149
transform 1 0 0 0 1 5530
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_23
timestamp 1644511149
transform 1 0 0 0 -1 5530
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_24
timestamp 1644511149
transform 1 0 0 0 1 4740
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_25
timestamp 1644511149
transform 1 0 0 0 -1 4740
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_26
timestamp 1644511149
transform 1 0 0 0 1 3950
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_27
timestamp 1644511149
transform 1 0 0 0 -1 3950
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_28
timestamp 1644511149
transform 1 0 0 0 1 3160
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_29
timestamp 1644511149
transform 1 0 0 0 -1 3160
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_30
timestamp 1644511149
transform 1 0 0 0 1 2370
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_31
timestamp 1644511149
transform 1 0 0 0 1 24490
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_32
timestamp 1644511149
transform 1 0 0 0 -1 24490
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_33
timestamp 1644511149
transform 1 0 0 0 1 23700
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_34
timestamp 1644511149
transform 1 0 0 0 -1 23700
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_35
timestamp 1644511149
transform 1 0 0 0 1 22910
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_36
timestamp 1644511149
transform 1 0 0 0 -1 22910
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_37
timestamp 1644511149
transform 1 0 0 0 1 22120
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_38
timestamp 1644511149
transform 1 0 0 0 -1 22120
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_39
timestamp 1644511149
transform 1 0 0 0 1 21330
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_40
timestamp 1644511149
transform 1 0 0 0 -1 21330
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_41
timestamp 1644511149
transform 1 0 0 0 1 20540
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_42
timestamp 1644511149
transform 1 0 0 0 -1 20540
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_43
timestamp 1644511149
transform 1 0 0 0 1 19750
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_44
timestamp 1644511149
transform 1 0 0 0 -1 19750
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_45
timestamp 1644511149
transform 1 0 0 0 1 18960
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_46
timestamp 1644511149
transform 1 0 0 0 -1 18960
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_47
timestamp 1644511149
transform 1 0 0 0 1 18170
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_48
timestamp 1644511149
transform 1 0 0 0 -1 18170
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_49
timestamp 1644511149
transform 1 0 0 0 1 17380
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_50
timestamp 1644511149
transform 1 0 0 0 -1 17380
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_51
timestamp 1644511149
transform 1 0 0 0 1 16590
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_52
timestamp 1644511149
transform 1 0 0 0 -1 16590
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_53
timestamp 1644511149
transform 1 0 0 0 1 15800
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_54
timestamp 1644511149
transform 1 0 0 0 -1 15800
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_55
timestamp 1644511149
transform 1 0 0 0 1 15010
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_56
timestamp 1644511149
transform 1 0 0 0 -1 15010
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_57
timestamp 1644511149
transform 1 0 0 0 1 14220
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_58
timestamp 1644511149
transform 1 0 0 0 -1 14220
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_59
timestamp 1644511149
transform 1 0 0 0 1 13430
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_60
timestamp 1644511149
transform 1 0 0 0 -1 13430
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_61
timestamp 1644511149
transform 1 0 0 0 1 12640
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_62
timestamp 1644511149
transform 1 0 0 0 -1 12640
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_63
timestamp 1644511149
transform 1 0 0 0 -1 26860
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_64
timestamp 1644511149
transform 1 0 0 0 1 26070
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_65
timestamp 1644511149
transform 1 0 0 0 -1 26070
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_66
timestamp 1644511149
transform 1 0 0 0 1 37130
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_67
timestamp 1644511149
transform 1 0 0 0 -1 37130
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_68
timestamp 1644511149
transform 1 0 0 0 1 36340
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_69
timestamp 1644511149
transform 1 0 0 0 -1 36340
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_70
timestamp 1644511149
transform 1 0 0 0 1 35550
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_71
timestamp 1644511149
transform 1 0 0 0 -1 35550
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_72
timestamp 1644511149
transform 1 0 0 0 1 34760
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_73
timestamp 1644511149
transform 1 0 0 0 -1 34760
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_74
timestamp 1644511149
transform 1 0 0 0 1 33970
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_75
timestamp 1644511149
transform 1 0 0 0 -1 33970
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_76
timestamp 1644511149
transform 1 0 0 0 1 33180
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_77
timestamp 1644511149
transform 1 0 0 0 -1 33180
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_78
timestamp 1644511149
transform 1 0 0 0 1 32390
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_79
timestamp 1644511149
transform 1 0 0 0 -1 32390
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_80
timestamp 1644511149
transform 1 0 0 0 1 31600
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_81
timestamp 1644511149
transform 1 0 0 0 -1 31600
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_82
timestamp 1644511149
transform 1 0 0 0 1 30810
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_83
timestamp 1644511149
transform 1 0 0 0 -1 30810
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_84
timestamp 1644511149
transform 1 0 0 0 1 30020
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_85
timestamp 1644511149
transform 1 0 0 0 -1 30020
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_86
timestamp 1644511149
transform 1 0 0 0 1 29230
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_87
timestamp 1644511149
transform 1 0 0 0 -1 29230
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_88
timestamp 1644511149
transform 1 0 0 0 1 28440
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_89
timestamp 1644511149
transform 1 0 0 0 -1 28440
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_90
timestamp 1644511149
transform 1 0 0 0 1 27650
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_91
timestamp 1644511149
transform 1 0 0 0 -1 27650
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_92
timestamp 1644511149
transform 1 0 0 0 1 26860
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_93
timestamp 1644511149
transform 1 0 0 0 -1 50560
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_94
timestamp 1644511149
transform 1 0 0 0 1 49770
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_95
timestamp 1644511149
transform 1 0 0 0 -1 49770
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_96
timestamp 1644511149
transform 1 0 0 0 1 48980
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_97
timestamp 1644511149
transform 1 0 0 0 -1 48980
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_98
timestamp 1644511149
transform 1 0 0 0 1 48190
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_99
timestamp 1644511149
transform 1 0 0 0 -1 48190
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_100
timestamp 1644511149
transform 1 0 0 0 1 47400
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_101
timestamp 1644511149
transform 1 0 0 0 -1 47400
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_102
timestamp 1644511149
transform 1 0 0 0 1 46610
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_103
timestamp 1644511149
transform 1 0 0 0 -1 46610
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_104
timestamp 1644511149
transform 1 0 0 0 1 45820
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_105
timestamp 1644511149
transform 1 0 0 0 -1 45820
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_106
timestamp 1644511149
transform 1 0 0 0 1 45030
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_107
timestamp 1644511149
transform 1 0 0 0 -1 45030
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_108
timestamp 1644511149
transform 1 0 0 0 1 44240
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_109
timestamp 1644511149
transform 1 0 0 0 -1 44240
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_110
timestamp 1644511149
transform 1 0 0 0 1 43450
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_111
timestamp 1644511149
transform 1 0 0 0 -1 43450
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_112
timestamp 1644511149
transform 1 0 0 0 1 42660
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_113
timestamp 1644511149
transform 1 0 0 0 -1 42660
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_114
timestamp 1644511149
transform 1 0 0 0 1 41870
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_115
timestamp 1644511149
transform 1 0 0 0 -1 41870
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_116
timestamp 1644511149
transform 1 0 0 0 1 41080
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_117
timestamp 1644511149
transform 1 0 0 0 -1 41080
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_118
timestamp 1644511149
transform 1 0 0 0 1 40290
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_119
timestamp 1644511149
transform 1 0 0 0 -1 40290
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_120
timestamp 1644511149
transform 1 0 0 0 1 39500
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_121
timestamp 1644511149
transform 1 0 0 0 -1 39500
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_122
timestamp 1644511149
transform 1 0 0 0 1 38710
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_123
timestamp 1644511149
transform 1 0 0 0 -1 38710
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_124
timestamp 1644511149
transform 1 0 0 0 1 37920
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_125
timestamp 1644511149
transform 1 0 0 0 -1 37920
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_126
timestamp 1644511149
transform 1 0 0 0 1 25280
box 70 -56 4140 490
use sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver  sky130_sram_1kbyte_1rw1r_32x256_8_wordline_driver_127
timestamp 1644511149
transform 1 0 0 0 -1 25280
box 70 -56 4140 490
<< labels >>
rlabel metal2 s 70 0 98 50560 4 en
port 1 nsew
rlabel metal1 s 681 -32 709 50560 4 vdd
port 2 nsew
rlabel metal1 s 3372 0 3400 50560 4 vdd
port 2 nsew
rlabel metal1 s 256 -30 284 50560 4 gnd
port 3 nsew
rlabel metal1 s 1724 0 1752 50560 4 gnd
port 3 nsew
rlabel locali s 4108 25400 4108 25400 4 wl_64
port 4 nsew
rlabel locali s 4108 25950 4108 25950 4 wl_65
port 5 nsew
rlabel locali s 4108 26190 4108 26190 4 wl_66
port 6 nsew
rlabel locali s 4108 26740 4108 26740 4 wl_67
port 7 nsew
rlabel locali s 4108 26980 4108 26980 4 wl_68
port 8 nsew
rlabel locali s 4108 27530 4108 27530 4 wl_69
port 9 nsew
rlabel locali s 4108 27770 4108 27770 4 wl_70
port 10 nsew
rlabel locali s 4108 28320 4108 28320 4 wl_71
port 11 nsew
rlabel locali s 4108 28560 4108 28560 4 wl_72
port 12 nsew
rlabel locali s 4108 29110 4108 29110 4 wl_73
port 13 nsew
rlabel locali s 4108 29350 4108 29350 4 wl_74
port 14 nsew
rlabel locali s 4108 29900 4108 29900 4 wl_75
port 15 nsew
rlabel locali s 4108 30140 4108 30140 4 wl_76
port 16 nsew
rlabel locali s 4108 30690 4108 30690 4 wl_77
port 17 nsew
rlabel locali s 4108 30930 4108 30930 4 wl_78
port 18 nsew
rlabel locali s 4108 31480 4108 31480 4 wl_79
port 19 nsew
rlabel locali s 4108 31720 4108 31720 4 wl_80
port 20 nsew
rlabel locali s 4108 32270 4108 32270 4 wl_81
port 21 nsew
rlabel locali s 4108 32510 4108 32510 4 wl_82
port 22 nsew
rlabel locali s 4108 33060 4108 33060 4 wl_83
port 23 nsew
rlabel locali s 4108 33300 4108 33300 4 wl_84
port 24 nsew
rlabel locali s 4108 33850 4108 33850 4 wl_85
port 25 nsew
rlabel locali s 4108 34090 4108 34090 4 wl_86
port 26 nsew
rlabel locali s 4108 34640 4108 34640 4 wl_87
port 27 nsew
rlabel locali s 4108 34880 4108 34880 4 wl_88
port 28 nsew
rlabel locali s 4108 35430 4108 35430 4 wl_89
port 29 nsew
rlabel locali s 4108 35670 4108 35670 4 wl_90
port 30 nsew
rlabel locali s 4108 36220 4108 36220 4 wl_91
port 31 nsew
rlabel locali s 4108 36460 4108 36460 4 wl_92
port 32 nsew
rlabel locali s 4108 37010 4108 37010 4 wl_93
port 33 nsew
rlabel locali s 4108 37250 4108 37250 4 wl_94
port 34 nsew
rlabel locali s 4108 37800 4108 37800 4 wl_95
port 35 nsew
rlabel locali s 4108 38040 4108 38040 4 wl_96
port 36 nsew
rlabel locali s 4108 38590 4108 38590 4 wl_97
port 37 nsew
rlabel locali s 4108 38830 4108 38830 4 wl_98
port 38 nsew
rlabel locali s 4108 39380 4108 39380 4 wl_99
port 39 nsew
rlabel locali s 4108 39620 4108 39620 4 wl_100
port 40 nsew
rlabel locali s 4108 40170 4108 40170 4 wl_101
port 41 nsew
rlabel locali s 4108 40410 4108 40410 4 wl_102
port 42 nsew
rlabel locali s 4108 40960 4108 40960 4 wl_103
port 43 nsew
rlabel locali s 4108 41200 4108 41200 4 wl_104
port 44 nsew
rlabel locali s 4108 41750 4108 41750 4 wl_105
port 45 nsew
rlabel locali s 4108 41990 4108 41990 4 wl_106
port 46 nsew
rlabel locali s 4108 42540 4108 42540 4 wl_107
port 47 nsew
rlabel locali s 4108 42780 4108 42780 4 wl_108
port 48 nsew
rlabel locali s 4108 43330 4108 43330 4 wl_109
port 49 nsew
rlabel locali s 4108 43570 4108 43570 4 wl_110
port 50 nsew
rlabel locali s 4108 44120 4108 44120 4 wl_111
port 51 nsew
rlabel locali s 4108 44360 4108 44360 4 wl_112
port 52 nsew
rlabel locali s 4108 44910 4108 44910 4 wl_113
port 53 nsew
rlabel locali s 4108 45150 4108 45150 4 wl_114
port 54 nsew
rlabel locali s 4108 45700 4108 45700 4 wl_115
port 55 nsew
rlabel locali s 4108 45940 4108 45940 4 wl_116
port 56 nsew
rlabel locali s 4108 46490 4108 46490 4 wl_117
port 57 nsew
rlabel locali s 4108 46730 4108 46730 4 wl_118
port 58 nsew
rlabel locali s 4108 47280 4108 47280 4 wl_119
port 59 nsew
rlabel locali s 4108 47520 4108 47520 4 wl_120
port 60 nsew
rlabel locali s 4108 48070 4108 48070 4 wl_121
port 61 nsew
rlabel locali s 4108 48310 4108 48310 4 wl_122
port 62 nsew
rlabel locali s 4108 48860 4108 48860 4 wl_123
port 63 nsew
rlabel locali s 4108 49100 4108 49100 4 wl_124
port 64 nsew
rlabel locali s 4108 49650 4108 49650 4 wl_125
port 65 nsew
rlabel locali s 4108 49890 4108 49890 4 wl_126
port 66 nsew
rlabel locali s 4108 50440 4108 50440 4 wl_127
port 67 nsew
rlabel locali s 103 38219 103 38219 4 in_96
port 68 nsew
rlabel locali s 103 31899 103 31899 4 in_80
port 69 nsew
rlabel locali s 103 38411 103 38411 4 in_97
port 70 nsew
rlabel locali s 103 28739 103 28739 4 in_72
port 71 nsew
rlabel locali s 103 39009 103 39009 4 in_98
port 72 nsew
rlabel locali s 103 32091 103 32091 4 in_81
port 73 nsew
rlabel locali s 103 39201 103 39201 4 in_99
port 74 nsew
rlabel locali s 103 27159 103 27159 4 in_68
port 75 nsew
rlabel locali s 103 39799 103 39799 4 in_100
port 76 nsew
rlabel locali s 103 32689 103 32689 4 in_82
port 77 nsew
rlabel locali s 103 39991 103 39991 4 in_101
port 78 nsew
rlabel locali s 103 28931 103 28931 4 in_73
port 79 nsew
rlabel locali s 103 40589 103 40589 4 in_102
port 80 nsew
rlabel locali s 103 32881 103 32881 4 in_83
port 81 nsew
rlabel locali s 103 40781 103 40781 4 in_103
port 82 nsew
rlabel locali s 103 26369 103 26369 4 in_66
port 83 nsew
rlabel locali s 103 41379 103 41379 4 in_104
port 84 nsew
rlabel locali s 103 33479 103 33479 4 in_84
port 85 nsew
rlabel locali s 103 41571 103 41571 4 in_105
port 86 nsew
rlabel locali s 103 29529 103 29529 4 in_74
port 87 nsew
rlabel locali s 103 42169 103 42169 4 in_106
port 88 nsew
rlabel locali s 103 33671 103 33671 4 in_85
port 89 nsew
rlabel locali s 103 42361 103 42361 4 in_107
port 90 nsew
rlabel locali s 103 27351 103 27351 4 in_69
port 91 nsew
rlabel locali s 103 42959 103 42959 4 in_108
port 92 nsew
rlabel locali s 103 34269 103 34269 4 in_86
port 93 nsew
rlabel locali s 103 43151 103 43151 4 in_109
port 94 nsew
rlabel locali s 103 29721 103 29721 4 in_75
port 95 nsew
rlabel locali s 103 43749 103 43749 4 in_110
port 96 nsew
rlabel locali s 103 34461 103 34461 4 in_87
port 97 nsew
rlabel locali s 103 43941 103 43941 4 in_111
port 98 nsew
rlabel locali s 103 25771 103 25771 4 in_65
port 99 nsew
rlabel locali s 103 44539 103 44539 4 in_112
port 100 nsew
rlabel locali s 103 35059 103 35059 4 in_88
port 101 nsew
rlabel locali s 103 44731 103 44731 4 in_113
port 102 nsew
rlabel locali s 103 30319 103 30319 4 in_76
port 103 nsew
rlabel locali s 103 45329 103 45329 4 in_114
port 104 nsew
rlabel locali s 103 35251 103 35251 4 in_89
port 105 nsew
rlabel locali s 103 45521 103 45521 4 in_115
port 106 nsew
rlabel locali s 103 27949 103 27949 4 in_70
port 107 nsew
rlabel locali s 103 46119 103 46119 4 in_116
port 108 nsew
rlabel locali s 103 35849 103 35849 4 in_90
port 109 nsew
rlabel locali s 103 46311 103 46311 4 in_117
port 110 nsew
rlabel locali s 103 30511 103 30511 4 in_77
port 111 nsew
rlabel locali s 103 46909 103 46909 4 in_118
port 112 nsew
rlabel locali s 103 36041 103 36041 4 in_91
port 113 nsew
rlabel locali s 103 47101 103 47101 4 in_119
port 114 nsew
rlabel locali s 103 26561 103 26561 4 in_67
port 115 nsew
rlabel locali s 103 47699 103 47699 4 in_120
port 116 nsew
rlabel locali s 103 36639 103 36639 4 in_92
port 117 nsew
rlabel locali s 103 47891 103 47891 4 in_121
port 118 nsew
rlabel locali s 103 31109 103 31109 4 in_78
port 119 nsew
rlabel locali s 103 48489 103 48489 4 in_122
port 120 nsew
rlabel locali s 103 36831 103 36831 4 in_93
port 121 nsew
rlabel locali s 103 48681 103 48681 4 in_123
port 122 nsew
rlabel locali s 103 28141 103 28141 4 in_71
port 123 nsew
rlabel locali s 103 49279 103 49279 4 in_124
port 124 nsew
rlabel locali s 103 37429 103 37429 4 in_94
port 125 nsew
rlabel locali s 103 49471 103 49471 4 in_125
port 126 nsew
rlabel locali s 103 31301 103 31301 4 in_79
port 127 nsew
rlabel locali s 103 50069 103 50069 4 in_126
port 128 nsew
rlabel locali s 103 37621 103 37621 4 in_95
port 129 nsew
rlabel locali s 103 50261 103 50261 4 in_127
port 130 nsew
rlabel locali s 103 25579 103 25579 4 in_64
port 131 nsew
rlabel locali s 103 299 103 299 4 in_0
port 132 nsew
rlabel locali s 103 491 103 491 4 in_1
port 133 nsew
rlabel locali s 103 1089 103 1089 4 in_2
port 134 nsew
rlabel locali s 103 1281 103 1281 4 in_3
port 135 nsew
rlabel locali s 103 1879 103 1879 4 in_4
port 136 nsew
rlabel locali s 103 2071 103 2071 4 in_5
port 137 nsew
rlabel locali s 103 2669 103 2669 4 in_6
port 138 nsew
rlabel locali s 103 2861 103 2861 4 in_7
port 139 nsew
rlabel locali s 103 3459 103 3459 4 in_8
port 140 nsew
rlabel locali s 103 3651 103 3651 4 in_9
port 141 nsew
rlabel locali s 103 4249 103 4249 4 in_10
port 142 nsew
rlabel locali s 103 4441 103 4441 4 in_11
port 143 nsew
rlabel locali s 103 5039 103 5039 4 in_12
port 144 nsew
rlabel locali s 103 5231 103 5231 4 in_13
port 145 nsew
rlabel locali s 103 5829 103 5829 4 in_14
port 146 nsew
rlabel locali s 103 6021 103 6021 4 in_15
port 147 nsew
rlabel locali s 103 6619 103 6619 4 in_16
port 148 nsew
rlabel locali s 103 6811 103 6811 4 in_17
port 149 nsew
rlabel locali s 103 7409 103 7409 4 in_18
port 150 nsew
rlabel locali s 103 7601 103 7601 4 in_19
port 151 nsew
rlabel locali s 103 8199 103 8199 4 in_20
port 152 nsew
rlabel locali s 103 8391 103 8391 4 in_21
port 153 nsew
rlabel locali s 103 8989 103 8989 4 in_22
port 154 nsew
rlabel locali s 103 9181 103 9181 4 in_23
port 155 nsew
rlabel locali s 103 9779 103 9779 4 in_24
port 156 nsew
rlabel locali s 103 9971 103 9971 4 in_25
port 157 nsew
rlabel locali s 103 10569 103 10569 4 in_26
port 158 nsew
rlabel locali s 103 10761 103 10761 4 in_27
port 159 nsew
rlabel locali s 103 11359 103 11359 4 in_28
port 160 nsew
rlabel locali s 103 11551 103 11551 4 in_29
port 161 nsew
rlabel locali s 103 12149 103 12149 4 in_30
port 162 nsew
rlabel locali s 103 12341 103 12341 4 in_31
port 163 nsew
rlabel locali s 103 12939 103 12939 4 in_32
port 164 nsew
rlabel locali s 103 13131 103 13131 4 in_33
port 165 nsew
rlabel locali s 103 13729 103 13729 4 in_34
port 166 nsew
rlabel locali s 103 13921 103 13921 4 in_35
port 167 nsew
rlabel locali s 103 14519 103 14519 4 in_36
port 168 nsew
rlabel locali s 103 14711 103 14711 4 in_37
port 169 nsew
rlabel locali s 103 15309 103 15309 4 in_38
port 170 nsew
rlabel locali s 103 15501 103 15501 4 in_39
port 171 nsew
rlabel locali s 103 16099 103 16099 4 in_40
port 172 nsew
rlabel locali s 103 16291 103 16291 4 in_41
port 173 nsew
rlabel locali s 103 16889 103 16889 4 in_42
port 174 nsew
rlabel locali s 103 17081 103 17081 4 in_43
port 175 nsew
rlabel locali s 103 17679 103 17679 4 in_44
port 176 nsew
rlabel locali s 103 17871 103 17871 4 in_45
port 177 nsew
rlabel locali s 103 18469 103 18469 4 in_46
port 178 nsew
rlabel locali s 103 18661 103 18661 4 in_47
port 179 nsew
rlabel locali s 103 19259 103 19259 4 in_48
port 180 nsew
rlabel locali s 103 19451 103 19451 4 in_49
port 181 nsew
rlabel locali s 103 20049 103 20049 4 in_50
port 182 nsew
rlabel locali s 103 20241 103 20241 4 in_51
port 183 nsew
rlabel locali s 103 20839 103 20839 4 in_52
port 184 nsew
rlabel locali s 103 21031 103 21031 4 in_53
port 185 nsew
rlabel locali s 103 21629 103 21629 4 in_54
port 186 nsew
rlabel locali s 103 21821 103 21821 4 in_55
port 187 nsew
rlabel locali s 103 22419 103 22419 4 in_56
port 188 nsew
rlabel locali s 103 22611 103 22611 4 in_57
port 189 nsew
rlabel locali s 103 23209 103 23209 4 in_58
port 190 nsew
rlabel locali s 103 23401 103 23401 4 in_59
port 191 nsew
rlabel locali s 103 23999 103 23999 4 in_60
port 192 nsew
rlabel locali s 103 24191 103 24191 4 in_61
port 193 nsew
rlabel locali s 103 24789 103 24789 4 in_62
port 194 nsew
rlabel locali s 103 24981 103 24981 4 in_63
port 195 nsew
rlabel locali s 4108 120 4108 120 4 wl_0
port 196 nsew
rlabel locali s 4108 12760 4108 12760 4 wl_32
port 197 nsew
rlabel locali s 4108 6440 4108 6440 4 wl_16
port 198 nsew
rlabel locali s 4108 13310 4108 13310 4 wl_33
port 199 nsew
rlabel locali s 4108 3280 4108 3280 4 wl_8
port 200 nsew
rlabel locali s 4108 13550 4108 13550 4 wl_34
port 201 nsew
rlabel locali s 4108 6990 4108 6990 4 wl_17
port 202 nsew
rlabel locali s 4108 14100 4108 14100 4 wl_35
port 203 nsew
rlabel locali s 4108 1700 4108 1700 4 wl_4
port 204 nsew
rlabel locali s 4108 14340 4108 14340 4 wl_36
port 205 nsew
rlabel locali s 4108 7230 4108 7230 4 wl_18
port 206 nsew
rlabel locali s 4108 14890 4108 14890 4 wl_37
port 207 nsew
rlabel locali s 4108 3830 4108 3830 4 wl_9
port 208 nsew
rlabel locali s 4108 15130 4108 15130 4 wl_38
port 209 nsew
rlabel locali s 4108 7780 4108 7780 4 wl_19
port 210 nsew
rlabel locali s 4108 15680 4108 15680 4 wl_39
port 211 nsew
rlabel locali s 4108 910 4108 910 4 wl_2
port 212 nsew
rlabel locali s 4108 15920 4108 15920 4 wl_40
port 213 nsew
rlabel locali s 4108 8020 4108 8020 4 wl_20
port 214 nsew
rlabel locali s 4108 16470 4108 16470 4 wl_41
port 215 nsew
rlabel locali s 4108 4070 4108 4070 4 wl_10
port 216 nsew
rlabel locali s 4108 16710 4108 16710 4 wl_42
port 217 nsew
rlabel locali s 4108 8570 4108 8570 4 wl_21
port 218 nsew
rlabel locali s 4108 17260 4108 17260 4 wl_43
port 219 nsew
rlabel locali s 4108 2250 4108 2250 4 wl_5
port 220 nsew
rlabel locali s 4108 17500 4108 17500 4 wl_44
port 221 nsew
rlabel locali s 4108 8810 4108 8810 4 wl_22
port 222 nsew
rlabel locali s 4108 18050 4108 18050 4 wl_45
port 223 nsew
rlabel locali s 4108 4620 4108 4620 4 wl_11
port 224 nsew
rlabel locali s 4108 18290 4108 18290 4 wl_46
port 225 nsew
rlabel locali s 4108 9360 4108 9360 4 wl_23
port 226 nsew
rlabel locali s 4108 18840 4108 18840 4 wl_47
port 227 nsew
rlabel locali s 4108 670 4108 670 4 wl_1
port 228 nsew
rlabel locali s 4108 19080 4108 19080 4 wl_48
port 229 nsew
rlabel locali s 4108 9600 4108 9600 4 wl_24
port 230 nsew
rlabel locali s 4108 19630 4108 19630 4 wl_49
port 231 nsew
rlabel locali s 4108 4860 4108 4860 4 wl_12
port 232 nsew
rlabel locali s 4108 19870 4108 19870 4 wl_50
port 233 nsew
rlabel locali s 4108 10150 4108 10150 4 wl_25
port 234 nsew
rlabel locali s 4108 20420 4108 20420 4 wl_51
port 235 nsew
rlabel locali s 4108 2490 4108 2490 4 wl_6
port 236 nsew
rlabel locali s 4108 20660 4108 20660 4 wl_52
port 237 nsew
rlabel locali s 4108 10390 4108 10390 4 wl_26
port 238 nsew
rlabel locali s 4108 21210 4108 21210 4 wl_53
port 239 nsew
rlabel locali s 4108 5410 4108 5410 4 wl_13
port 240 nsew
rlabel locali s 4108 21450 4108 21450 4 wl_54
port 241 nsew
rlabel locali s 4108 10940 4108 10940 4 wl_27
port 242 nsew
rlabel locali s 4108 22000 4108 22000 4 wl_55
port 243 nsew
rlabel locali s 4108 1460 4108 1460 4 wl_3
port 244 nsew
rlabel locali s 4108 22240 4108 22240 4 wl_56
port 245 nsew
rlabel locali s 4108 11180 4108 11180 4 wl_28
port 246 nsew
rlabel locali s 4108 22790 4108 22790 4 wl_57
port 247 nsew
rlabel locali s 4108 5650 4108 5650 4 wl_14
port 248 nsew
rlabel locali s 4108 23030 4108 23030 4 wl_58
port 249 nsew
rlabel locali s 4108 11730 4108 11730 4 wl_29
port 250 nsew
rlabel locali s 4108 23580 4108 23580 4 wl_59
port 251 nsew
rlabel locali s 4108 3040 4108 3040 4 wl_7
port 252 nsew
rlabel locali s 4108 23820 4108 23820 4 wl_60
port 253 nsew
rlabel locali s 4108 11970 4108 11970 4 wl_30
port 254 nsew
rlabel locali s 4108 24370 4108 24370 4 wl_61
port 255 nsew
rlabel locali s 4108 6200 4108 6200 4 wl_15
port 256 nsew
rlabel locali s 4108 24610 4108 24610 4 wl_62
port 257 nsew
rlabel locali s 4108 12520 4108 12520 4 wl_31
port 258 nsew
rlabel locali s 4108 25160 4108 25160 4 wl_63
port 259 nsew
<< properties >>
string FIXED_BBOX 0 0 4158 50560
string GDS_END 462238
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_32x256_8.gds
string GDS_START 395230
<< end >>
