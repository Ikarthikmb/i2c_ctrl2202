magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 808 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 437 47 467 177
rect 521 47 551 177
rect 605 47 635 177
rect 689 47 719 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 437 297 467 497
rect 521 297 551 497
rect 605 297 635 497
rect 689 297 719 497
<< ndiff >>
rect 27 165 79 177
rect 27 131 35 165
rect 69 131 79 165
rect 27 97 79 131
rect 27 63 35 97
rect 69 63 79 97
rect 27 47 79 63
rect 109 95 163 177
rect 109 61 119 95
rect 153 61 163 95
rect 109 47 163 61
rect 193 165 247 177
rect 193 131 203 165
rect 237 131 247 165
rect 193 97 247 131
rect 193 63 203 97
rect 237 63 247 97
rect 193 47 247 63
rect 277 95 437 177
rect 277 61 287 95
rect 321 61 393 95
rect 427 61 437 95
rect 277 47 437 61
rect 467 163 521 177
rect 467 129 477 163
rect 511 129 521 163
rect 467 95 521 129
rect 467 61 477 95
rect 511 61 521 95
rect 467 47 521 61
rect 551 95 605 177
rect 551 61 561 95
rect 595 61 605 95
rect 551 47 605 61
rect 635 163 689 177
rect 635 129 645 163
rect 679 129 689 163
rect 635 95 689 129
rect 635 61 645 95
rect 679 61 689 95
rect 635 47 689 61
rect 719 95 782 177
rect 719 61 729 95
rect 763 61 782 95
rect 719 47 782 61
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 297 163 497
rect 193 297 247 497
rect 277 485 437 497
rect 277 451 300 485
rect 334 451 393 485
rect 427 451 437 485
rect 277 417 437 451
rect 277 383 300 417
rect 334 383 393 417
rect 427 383 437 417
rect 277 297 437 383
rect 467 477 521 497
rect 467 443 477 477
rect 511 443 521 477
rect 467 409 521 443
rect 467 375 477 409
rect 511 375 521 409
rect 467 341 521 375
rect 467 307 477 341
rect 511 307 521 341
rect 467 297 521 307
rect 551 477 605 497
rect 551 443 561 477
rect 595 443 605 477
rect 551 409 605 443
rect 551 375 561 409
rect 595 375 605 409
rect 551 297 605 375
rect 635 477 689 497
rect 635 443 645 477
rect 679 443 689 477
rect 635 409 689 443
rect 635 375 645 409
rect 679 375 689 409
rect 635 341 689 375
rect 635 307 645 341
rect 679 307 689 341
rect 635 297 689 307
rect 719 477 791 497
rect 719 443 729 477
rect 763 443 791 477
rect 719 409 791 443
rect 719 375 729 409
rect 763 375 791 409
rect 719 297 791 375
<< ndiffc >>
rect 35 131 69 165
rect 35 63 69 97
rect 119 61 153 95
rect 203 131 237 165
rect 203 63 237 97
rect 287 61 321 95
rect 393 61 427 95
rect 477 129 511 163
rect 477 61 511 95
rect 561 61 595 95
rect 645 129 679 163
rect 645 61 679 95
rect 729 61 763 95
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 300 451 334 485
rect 393 451 427 485
rect 300 383 334 417
rect 393 383 427 417
rect 477 443 511 477
rect 477 375 511 409
rect 477 307 511 341
rect 561 443 595 477
rect 561 375 595 409
rect 645 443 679 477
rect 645 375 679 409
rect 645 307 679 341
rect 729 443 763 477
rect 729 375 763 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 437 497 467 523
rect 521 497 551 523
rect 605 497 635 523
rect 689 497 719 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 437 265 467 297
rect 521 265 551 297
rect 605 265 635 297
rect 689 265 719 297
rect 25 249 109 265
rect 25 215 35 249
rect 69 215 109 249
rect 25 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 249 305 265
rect 247 215 261 249
rect 295 215 305 249
rect 247 199 305 215
rect 380 249 719 265
rect 380 215 396 249
rect 430 215 464 249
rect 498 215 532 249
rect 566 215 600 249
rect 634 215 668 249
rect 702 215 719 249
rect 380 199 719 215
rect 79 177 109 199
rect 163 177 193 199
rect 247 177 277 199
rect 437 177 467 199
rect 521 177 551 199
rect 605 177 635 199
rect 689 177 719 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 437 21 467 47
rect 521 21 551 47
rect 605 21 635 47
rect 689 21 719 47
<< polycont >>
rect 35 215 69 249
rect 161 215 195 249
rect 261 215 295 249
rect 396 215 430 249
rect 464 215 498 249
rect 532 215 566 249
rect 600 215 634 249
rect 668 215 702 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 485 253 493
rect 17 451 35 485
rect 69 459 253 485
rect 69 451 85 459
rect 17 417 85 451
rect 17 383 35 417
rect 69 383 85 417
rect 17 349 85 383
rect 17 315 35 349
rect 69 315 85 349
rect 17 299 85 315
rect 119 265 166 410
rect 200 333 253 459
rect 287 485 427 527
rect 287 451 300 485
rect 334 451 393 485
rect 287 417 427 451
rect 287 383 300 417
rect 334 383 393 417
rect 287 367 427 383
rect 469 477 519 493
rect 469 443 477 477
rect 511 443 519 477
rect 469 409 519 443
rect 469 375 477 409
rect 511 375 519 409
rect 469 341 519 375
rect 553 477 603 527
rect 553 443 561 477
rect 595 443 603 477
rect 553 409 603 443
rect 553 375 561 409
rect 595 375 603 409
rect 553 359 603 375
rect 637 477 687 493
rect 637 443 645 477
rect 679 443 687 477
rect 637 409 687 443
rect 637 375 645 409
rect 679 375 687 409
rect 200 299 418 333
rect 17 249 85 265
rect 17 215 35 249
rect 69 215 85 249
rect 119 249 211 265
rect 119 215 161 249
rect 195 215 211 249
rect 245 249 340 265
rect 245 215 261 249
rect 295 215 340 249
rect 374 249 418 299
rect 469 307 477 341
rect 511 325 519 341
rect 637 341 687 375
rect 721 477 771 527
rect 721 443 729 477
rect 763 443 771 477
rect 721 409 771 443
rect 721 375 729 409
rect 763 375 771 409
rect 721 359 771 375
rect 637 325 645 341
rect 511 307 645 325
rect 679 325 687 341
rect 679 307 811 325
rect 469 291 811 307
rect 374 215 396 249
rect 430 215 464 249
rect 498 215 532 249
rect 566 215 600 249
rect 634 215 668 249
rect 702 215 719 249
rect 374 181 418 215
rect 753 181 811 291
rect 17 165 418 181
rect 17 131 35 165
rect 69 145 203 165
rect 69 131 85 145
rect 17 97 85 131
rect 187 131 203 145
rect 237 145 418 165
rect 461 163 811 181
rect 237 131 253 145
rect 17 63 35 97
rect 69 63 85 97
rect 17 51 85 63
rect 119 95 153 111
rect 119 17 153 61
rect 187 97 253 131
rect 461 129 477 163
rect 511 147 645 163
rect 511 129 527 147
rect 187 63 203 97
rect 237 63 253 97
rect 187 51 253 63
rect 287 95 427 111
rect 321 61 393 95
rect 287 17 427 61
rect 461 95 527 129
rect 629 129 645 147
rect 679 147 811 163
rect 679 129 695 147
rect 461 61 477 95
rect 511 61 527 95
rect 461 53 527 61
rect 561 95 595 111
rect 561 17 595 61
rect 629 95 695 129
rect 629 61 645 95
rect 679 61 695 95
rect 629 53 695 61
rect 729 95 763 111
rect 729 17 763 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 306 221 340 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 766 153 800 187 0 FreeSans 200 0 0 0 X
port 8 nsew signal output
flabel locali s 122 357 156 391 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 C
port 3 nsew signal input
flabel locali s 122 289 156 323 0 FreeSans 400 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
rlabel comment s 0 0 0 0 4 or3_4
rlabel metal1 s 0 -48 828 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 1038760
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1031702
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.140 0.000 
<< end >>
