magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -36 679 620 1471
<< pwell >>
rect 448 25 550 159
<< psubdiff >>
rect 474 109 524 133
rect 474 75 482 109
rect 516 75 524 109
rect 474 51 524 75
<< nsubdiff >>
rect 474 1339 524 1363
rect 474 1305 482 1339
rect 516 1305 524 1339
rect 474 1281 524 1305
<< psubdiffcont >>
rect 482 75 516 109
<< nsubdiffcont >>
rect 482 1305 516 1339
<< poly >>
rect 114 740 144 907
rect 48 724 144 740
rect 48 690 64 724
rect 98 690 144 724
rect 48 674 144 690
rect 114 507 144 674
<< polycont >>
rect 64 690 98 724
<< locali >>
rect 0 1397 584 1431
rect 62 1130 96 1397
rect 274 1130 308 1397
rect 482 1339 516 1397
rect 482 1289 516 1305
rect 64 724 98 740
rect 64 674 98 690
rect 272 724 306 1096
rect 272 690 323 724
rect 272 318 306 690
rect 62 17 96 218
rect 274 17 308 218
rect 482 109 516 125
rect 482 17 516 75
rect 0 -17 584 17
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_16  sky130_sram_2kbyte_1rw1r_32x512_8_contact_16_0
timestamp 1644511149
transform 1 0 48 0 1 674
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_28  sky130_sram_2kbyte_1rw1r_32x512_8_contact_28_0
timestamp 1644511149
transform 1 0 474 0 1 1281
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_contact_29  sky130_sram_2kbyte_1rw1r_32x512_8_contact_29_0
timestamp 1644511149
transform 1 0 474 0 1 51
box 0 0 1 1
use sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m3_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_nmos_m3_w2_000_sli_dli_da_p_0
timestamp 1644511149
transform 1 0 54 0 1 51
box -26 -26 392 456
use sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m3_w2_000_sli_dli_da_p  sky130_sram_2kbyte_1rw1r_32x512_8_pmos_m3_w2_000_sli_dli_da_p_0
timestamp 1644511149
transform 1 0 54 0 1 963
box -59 -56 425 454
<< labels >>
rlabel locali s 81 707 81 707 4 A
port 1 nsew
rlabel locali s 306 707 306 707 4 Z
port 2 nsew
rlabel locali s 292 0 292 0 4 gnd
port 3 nsew
rlabel locali s 292 1414 292 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 584 1414
string GDS_END 377690
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_2kbyte_1rw1r_32x512_8.gds
string GDS_START 375692
<< end >>
