magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -8 676 1176 1467
<< pwell >>
rect 2 76 1166 328
rect 2 -43 1088 76
<< scnmos >>
rect 81 102 111 302
rect 167 102 197 302
rect 239 102 269 302
rect 359 102 389 302
rect 431 102 461 302
rect 517 102 547 302
rect 589 102 619 302
rect 709 102 739 302
rect 781 102 811 302
rect 867 102 897 302
rect 1057 102 1087 302
<< scpmos >>
rect 81 712 111 1312
rect 167 712 197 1312
rect 239 712 269 1312
rect 359 712 389 1312
rect 431 712 461 1312
rect 517 712 547 1312
rect 589 712 619 1312
rect 709 712 739 1312
rect 781 712 811 1312
rect 867 712 897 1312
rect 1057 712 1087 1312
<< ndiff >>
rect 28 237 81 302
rect 28 203 36 237
rect 70 203 81 237
rect 28 169 81 203
rect 28 135 36 169
rect 70 135 81 169
rect 28 102 81 135
rect 111 237 167 302
rect 111 203 122 237
rect 156 203 167 237
rect 111 169 167 203
rect 111 135 122 169
rect 156 135 167 169
rect 111 102 167 135
rect 197 102 239 302
rect 269 237 359 302
rect 269 203 297 237
rect 331 203 359 237
rect 269 169 359 203
rect 269 135 297 169
rect 331 135 359 169
rect 269 102 359 135
rect 389 102 431 302
rect 461 237 517 302
rect 461 203 472 237
rect 506 203 517 237
rect 461 169 517 203
rect 461 135 472 169
rect 506 135 517 169
rect 461 102 517 135
rect 547 102 589 302
rect 619 237 709 302
rect 619 203 647 237
rect 681 203 709 237
rect 619 169 709 203
rect 619 135 647 169
rect 681 135 709 169
rect 619 102 709 135
rect 739 102 781 302
rect 811 237 867 302
rect 811 203 822 237
rect 856 203 867 237
rect 811 169 867 203
rect 811 135 822 169
rect 856 135 867 169
rect 811 102 867 135
rect 897 237 950 302
rect 897 203 908 237
rect 942 203 950 237
rect 897 169 950 203
rect 897 135 908 169
rect 942 135 950 169
rect 897 102 950 135
rect 1004 237 1057 302
rect 1004 203 1012 237
rect 1046 203 1057 237
rect 1004 169 1057 203
rect 1004 135 1012 169
rect 1046 135 1057 169
rect 1004 102 1057 135
rect 1087 237 1140 302
rect 1087 203 1098 237
rect 1132 203 1140 237
rect 1087 169 1140 203
rect 1087 135 1098 169
rect 1132 135 1140 169
rect 1087 102 1140 135
<< pdiff >>
rect 28 1279 81 1312
rect 28 1245 36 1279
rect 70 1245 81 1279
rect 28 1211 81 1245
rect 28 1177 36 1211
rect 70 1177 81 1211
rect 28 1143 81 1177
rect 28 1109 36 1143
rect 70 1109 81 1143
rect 28 1075 81 1109
rect 28 1041 36 1075
rect 70 1041 81 1075
rect 28 1007 81 1041
rect 28 973 36 1007
rect 70 973 81 1007
rect 28 939 81 973
rect 28 905 36 939
rect 70 905 81 939
rect 28 871 81 905
rect 28 837 36 871
rect 70 837 81 871
rect 28 712 81 837
rect 111 1279 167 1312
rect 111 1245 122 1279
rect 156 1245 167 1279
rect 111 1211 167 1245
rect 111 1177 122 1211
rect 156 1177 167 1211
rect 111 1143 167 1177
rect 111 1109 122 1143
rect 156 1109 167 1143
rect 111 1075 167 1109
rect 111 1041 122 1075
rect 156 1041 167 1075
rect 111 1007 167 1041
rect 111 973 122 1007
rect 156 973 167 1007
rect 111 939 167 973
rect 111 905 122 939
rect 156 905 167 939
rect 111 871 167 905
rect 111 837 122 871
rect 156 837 167 871
rect 111 712 167 837
rect 197 712 239 1312
rect 269 1279 359 1312
rect 269 1245 297 1279
rect 331 1245 359 1279
rect 269 1211 359 1245
rect 269 1177 297 1211
rect 331 1177 359 1211
rect 269 1143 359 1177
rect 269 1109 297 1143
rect 331 1109 359 1143
rect 269 1075 359 1109
rect 269 1041 297 1075
rect 331 1041 359 1075
rect 269 1007 359 1041
rect 269 973 297 1007
rect 331 973 359 1007
rect 269 939 359 973
rect 269 905 297 939
rect 331 905 359 939
rect 269 871 359 905
rect 269 837 297 871
rect 331 837 359 871
rect 269 712 359 837
rect 389 712 431 1312
rect 461 1279 517 1312
rect 461 1245 472 1279
rect 506 1245 517 1279
rect 461 1211 517 1245
rect 461 1177 472 1211
rect 506 1177 517 1211
rect 461 1143 517 1177
rect 461 1109 472 1143
rect 506 1109 517 1143
rect 461 1075 517 1109
rect 461 1041 472 1075
rect 506 1041 517 1075
rect 461 1007 517 1041
rect 461 973 472 1007
rect 506 973 517 1007
rect 461 939 517 973
rect 461 905 472 939
rect 506 905 517 939
rect 461 871 517 905
rect 461 837 472 871
rect 506 837 517 871
rect 461 712 517 837
rect 547 712 589 1312
rect 619 1279 709 1312
rect 619 1245 647 1279
rect 681 1245 709 1279
rect 619 1211 709 1245
rect 619 1177 647 1211
rect 681 1177 709 1211
rect 619 1143 709 1177
rect 619 1109 647 1143
rect 681 1109 709 1143
rect 619 1075 709 1109
rect 619 1041 647 1075
rect 681 1041 709 1075
rect 619 1007 709 1041
rect 619 973 647 1007
rect 681 973 709 1007
rect 619 939 709 973
rect 619 905 647 939
rect 681 905 709 939
rect 619 871 709 905
rect 619 837 647 871
rect 681 837 709 871
rect 619 712 709 837
rect 739 712 781 1312
rect 811 1279 867 1312
rect 811 1245 822 1279
rect 856 1245 867 1279
rect 811 1211 867 1245
rect 811 1177 822 1211
rect 856 1177 867 1211
rect 811 1143 867 1177
rect 811 1109 822 1143
rect 856 1109 867 1143
rect 811 1075 867 1109
rect 811 1041 822 1075
rect 856 1041 867 1075
rect 811 1007 867 1041
rect 811 973 822 1007
rect 856 973 867 1007
rect 811 939 867 973
rect 811 905 822 939
rect 856 905 867 939
rect 811 871 867 905
rect 811 837 822 871
rect 856 837 867 871
rect 811 712 867 837
rect 897 1279 950 1312
rect 897 1245 908 1279
rect 942 1245 950 1279
rect 897 1211 950 1245
rect 897 1177 908 1211
rect 942 1177 950 1211
rect 897 1143 950 1177
rect 897 1109 908 1143
rect 942 1109 950 1143
rect 897 1075 950 1109
rect 897 1041 908 1075
rect 942 1041 950 1075
rect 897 1007 950 1041
rect 897 973 908 1007
rect 942 973 950 1007
rect 897 939 950 973
rect 897 905 908 939
rect 942 905 950 939
rect 897 871 950 905
rect 897 837 908 871
rect 942 837 950 871
rect 897 712 950 837
rect 1004 1279 1057 1312
rect 1004 1245 1012 1279
rect 1046 1245 1057 1279
rect 1004 1211 1057 1245
rect 1004 1177 1012 1211
rect 1046 1177 1057 1211
rect 1004 1143 1057 1177
rect 1004 1109 1012 1143
rect 1046 1109 1057 1143
rect 1004 1075 1057 1109
rect 1004 1041 1012 1075
rect 1046 1041 1057 1075
rect 1004 1007 1057 1041
rect 1004 973 1012 1007
rect 1046 973 1057 1007
rect 1004 939 1057 973
rect 1004 905 1012 939
rect 1046 905 1057 939
rect 1004 871 1057 905
rect 1004 837 1012 871
rect 1046 837 1057 871
rect 1004 712 1057 837
rect 1087 1279 1140 1312
rect 1087 1245 1098 1279
rect 1132 1245 1140 1279
rect 1087 1211 1140 1245
rect 1087 1177 1098 1211
rect 1132 1177 1140 1211
rect 1087 1143 1140 1177
rect 1087 1109 1098 1143
rect 1132 1109 1140 1143
rect 1087 1075 1140 1109
rect 1087 1041 1098 1075
rect 1132 1041 1140 1075
rect 1087 1007 1140 1041
rect 1087 973 1098 1007
rect 1132 973 1140 1007
rect 1087 939 1140 973
rect 1087 905 1098 939
rect 1132 905 1140 939
rect 1087 871 1140 905
rect 1087 837 1098 871
rect 1132 837 1140 871
rect 1087 712 1140 837
<< ndiffc >>
rect 36 203 70 237
rect 36 135 70 169
rect 122 203 156 237
rect 122 135 156 169
rect 297 203 331 237
rect 297 135 331 169
rect 472 203 506 237
rect 472 135 506 169
rect 647 203 681 237
rect 647 135 681 169
rect 822 203 856 237
rect 822 135 856 169
rect 908 203 942 237
rect 908 135 942 169
rect 1012 203 1046 237
rect 1012 135 1046 169
rect 1098 203 1132 237
rect 1098 135 1132 169
<< pdiffc >>
rect 36 1245 70 1279
rect 36 1177 70 1211
rect 36 1109 70 1143
rect 36 1041 70 1075
rect 36 973 70 1007
rect 36 905 70 939
rect 36 837 70 871
rect 122 1245 156 1279
rect 122 1177 156 1211
rect 122 1109 156 1143
rect 122 1041 156 1075
rect 122 973 156 1007
rect 122 905 156 939
rect 122 837 156 871
rect 297 1245 331 1279
rect 297 1177 331 1211
rect 297 1109 331 1143
rect 297 1041 331 1075
rect 297 973 331 1007
rect 297 905 331 939
rect 297 837 331 871
rect 472 1245 506 1279
rect 472 1177 506 1211
rect 472 1109 506 1143
rect 472 1041 506 1075
rect 472 973 506 1007
rect 472 905 506 939
rect 472 837 506 871
rect 647 1245 681 1279
rect 647 1177 681 1211
rect 647 1109 681 1143
rect 647 1041 681 1075
rect 647 973 681 1007
rect 647 905 681 939
rect 647 837 681 871
rect 822 1245 856 1279
rect 822 1177 856 1211
rect 822 1109 856 1143
rect 822 1041 856 1075
rect 822 973 856 1007
rect 822 905 856 939
rect 822 837 856 871
rect 908 1245 942 1279
rect 908 1177 942 1211
rect 908 1109 942 1143
rect 908 1041 942 1075
rect 908 973 942 1007
rect 908 905 942 939
rect 908 837 942 871
rect 1012 1245 1046 1279
rect 1012 1177 1046 1211
rect 1012 1109 1046 1143
rect 1012 1041 1046 1075
rect 1012 973 1046 1007
rect 1012 905 1046 939
rect 1012 837 1046 871
rect 1098 1245 1132 1279
rect 1098 1177 1132 1211
rect 1098 1109 1132 1143
rect 1098 1041 1132 1075
rect 1098 973 1132 1007
rect 1098 905 1132 939
rect 1098 837 1132 871
<< psubdiff >>
rect 28 -17 52 17
rect 86 -17 110 17
rect 164 -17 188 17
rect 222 -17 246 17
rect 300 -17 324 17
rect 358 -17 382 17
rect 436 -17 460 17
rect 494 -17 518 17
rect 572 -17 596 17
rect 630 -17 654 17
rect 708 -17 732 17
rect 766 -17 790 17
rect 844 -17 868 17
rect 902 -17 926 17
rect 980 -17 1004 17
rect 1038 -17 1062 17
<< nsubdiff >>
rect 28 1397 52 1431
rect 86 1397 110 1431
rect 164 1397 188 1431
rect 222 1397 246 1431
rect 300 1397 324 1431
rect 358 1397 382 1431
rect 436 1397 460 1431
rect 494 1397 518 1431
rect 572 1397 596 1431
rect 630 1397 654 1431
rect 708 1397 732 1431
rect 766 1397 790 1431
rect 844 1397 868 1431
rect 902 1397 926 1431
rect 980 1397 1004 1431
rect 1038 1397 1062 1431
<< psubdiffcont >>
rect 52 -17 86 17
rect 188 -17 222 17
rect 324 -17 358 17
rect 460 -17 494 17
rect 596 -17 630 17
rect 732 -17 766 17
rect 868 -17 902 17
rect 1004 -17 1038 17
<< nsubdiffcont >>
rect 52 1397 86 1431
rect 188 1397 222 1431
rect 324 1397 358 1431
rect 460 1397 494 1431
rect 596 1397 630 1431
rect 732 1397 766 1431
rect 868 1397 902 1431
rect 1004 1397 1038 1431
<< poly >>
rect 81 1312 111 1338
rect 167 1312 197 1338
rect 239 1312 269 1338
rect 359 1312 389 1338
rect 431 1312 461 1338
rect 517 1312 547 1338
rect 589 1312 619 1338
rect 709 1312 739 1338
rect 781 1312 811 1338
rect 867 1312 897 1338
rect 1057 1312 1087 1338
rect 81 697 111 712
rect 70 677 111 697
rect 47 667 111 677
rect 47 661 101 667
rect 47 627 57 661
rect 91 627 101 661
rect 47 611 101 627
rect 71 447 101 611
rect 167 597 197 712
rect 239 672 269 712
rect 239 656 293 672
rect 239 622 249 656
rect 283 622 293 656
rect 239 606 293 622
rect 143 581 197 597
rect 143 547 153 581
rect 187 547 197 581
rect 143 531 197 547
rect 359 531 389 712
rect 431 667 461 712
rect 517 667 547 712
rect 431 657 547 667
rect 431 623 472 657
rect 506 623 547 657
rect 431 613 547 623
rect 589 531 619 712
rect 709 672 739 712
rect 685 656 739 672
rect 685 622 695 656
rect 729 622 739 656
rect 685 606 739 622
rect 781 597 811 712
rect 867 677 897 712
rect 867 661 938 677
rect 867 647 894 661
rect 878 627 894 647
rect 928 627 938 661
rect 878 611 938 627
rect 781 581 835 597
rect 781 547 791 581
rect 825 547 835 581
rect 781 531 835 547
rect 71 417 111 447
rect 81 302 111 417
rect 167 302 197 531
rect 239 501 739 531
rect 239 302 269 501
rect 685 467 695 501
rect 729 467 739 501
rect 685 451 739 467
rect 335 421 389 437
rect 335 387 345 421
rect 379 387 389 421
rect 335 371 389 387
rect 359 302 389 371
rect 431 421 547 431
rect 431 387 472 421
rect 506 387 547 421
rect 431 377 547 387
rect 431 302 461 377
rect 517 302 547 377
rect 589 421 643 437
rect 589 387 599 421
rect 633 387 643 421
rect 589 371 643 387
rect 589 302 619 371
rect 709 302 739 451
rect 781 302 811 531
rect 878 481 908 611
rect 1057 517 1087 712
rect 867 371 908 481
rect 1033 501 1087 517
rect 1033 467 1043 501
rect 1077 467 1087 501
rect 1033 451 1087 467
rect 867 302 897 371
rect 1057 302 1087 451
rect 81 76 111 102
rect 167 76 197 102
rect 239 76 269 102
rect 359 76 389 102
rect 431 76 461 102
rect 517 76 547 102
rect 589 76 619 102
rect 709 76 739 102
rect 781 76 811 102
rect 867 76 897 102
rect 1057 76 1087 102
<< polycont >>
rect 57 627 91 661
rect 249 622 283 656
rect 153 547 187 581
rect 472 623 506 657
rect 695 622 729 656
rect 894 627 928 661
rect 791 547 825 581
rect 695 467 729 501
rect 345 387 379 421
rect 472 387 506 421
rect 599 387 633 421
rect 1043 467 1077 501
<< locali >>
rect 0 1431 1168 1432
rect 0 1397 52 1431
rect 86 1397 188 1431
rect 222 1397 324 1431
rect 358 1397 460 1431
rect 494 1397 596 1431
rect 630 1397 732 1431
rect 766 1397 868 1431
rect 902 1397 1004 1431
rect 1038 1397 1168 1431
rect 0 1396 1168 1397
rect 36 1279 70 1312
rect 36 1211 70 1245
rect 36 1143 70 1177
rect 36 1075 70 1109
rect 36 1007 70 1041
rect 36 939 70 973
rect 36 871 70 905
rect 36 821 70 837
rect 122 1279 156 1396
rect 122 1211 156 1245
rect 122 1143 156 1177
rect 122 1075 156 1109
rect 122 1007 156 1041
rect 122 939 156 973
rect 122 871 156 905
rect 122 804 156 837
rect 280 1279 348 1312
rect 280 1245 297 1279
rect 331 1245 348 1279
rect 280 1211 348 1245
rect 280 1177 297 1211
rect 331 1177 348 1211
rect 280 1143 348 1177
rect 280 1109 297 1143
rect 331 1109 348 1143
rect 280 1075 348 1109
rect 280 1041 297 1075
rect 331 1041 348 1075
rect 280 1007 348 1041
rect 280 973 297 1007
rect 331 973 348 1007
rect 280 939 348 973
rect 280 905 297 939
rect 331 905 348 939
rect 280 871 348 905
rect 280 837 297 871
rect 331 837 348 871
rect 280 821 348 837
rect 280 804 297 821
rect 331 804 348 821
rect 472 1279 506 1396
rect 472 1211 506 1245
rect 472 1143 506 1177
rect 472 1075 506 1109
rect 472 1007 506 1041
rect 472 939 506 973
rect 472 871 506 905
rect 472 804 506 837
rect 630 1279 698 1312
rect 630 1245 647 1279
rect 681 1245 698 1279
rect 630 1211 698 1245
rect 630 1177 647 1211
rect 681 1177 698 1211
rect 630 1143 698 1177
rect 630 1109 647 1143
rect 681 1109 698 1143
rect 630 1075 698 1109
rect 630 1041 647 1075
rect 681 1041 698 1075
rect 630 1007 698 1041
rect 630 973 647 1007
rect 681 973 698 1007
rect 630 939 698 973
rect 630 905 647 939
rect 681 905 698 939
rect 630 871 698 905
rect 630 837 647 871
rect 681 837 698 871
rect 630 821 698 837
rect 630 804 647 821
rect 681 804 698 821
rect 822 1279 856 1396
rect 822 1211 856 1245
rect 822 1143 856 1177
rect 822 1075 856 1109
rect 822 1007 856 1041
rect 822 939 856 973
rect 822 871 856 905
rect 822 804 856 837
rect 908 1279 942 1312
rect 908 1211 942 1245
rect 908 1143 942 1177
rect 908 1075 942 1109
rect 908 1007 942 1041
rect 908 939 942 973
rect 908 871 942 905
rect 908 821 942 837
rect 1012 1279 1046 1396
rect 1012 1211 1046 1245
rect 1012 1143 1046 1177
rect 1012 1075 1046 1109
rect 1012 1007 1046 1041
rect 1012 939 1046 973
rect 1012 871 1046 905
rect 1012 804 1046 837
rect 1098 1279 1132 1312
rect 1098 1211 1132 1245
rect 1098 1143 1132 1177
rect 1098 1075 1132 1109
rect 1098 1007 1132 1041
rect 1098 939 1132 973
rect 1098 871 1132 905
rect 1098 821 1132 837
rect 41 707 379 741
rect 413 707 1132 741
rect 41 627 57 661
rect 91 627 113 661
rect 249 656 283 707
rect 456 623 472 657
rect 506 623 522 657
rect 249 606 283 622
rect 137 547 153 581
rect 187 547 203 581
rect 472 566 506 623
rect 239 532 506 566
rect 239 501 273 532
rect 70 467 273 501
rect 472 421 506 532
rect 599 421 633 707
rect 695 656 729 707
rect 894 661 928 707
rect 878 627 894 661
rect 928 627 944 661
rect 695 606 729 622
rect 1098 581 1132 618
rect 775 547 791 581
rect 825 547 1132 581
rect 679 467 695 501
rect 729 467 908 501
rect 1012 467 1020 501
rect 1077 467 1093 501
rect 328 387 345 421
rect 456 387 472 421
rect 506 387 522 421
rect 583 387 599 421
rect 633 387 649 421
rect 1012 341 1046 467
rect 647 307 1046 341
rect 647 270 681 307
rect 36 261 70 270
rect 36 169 70 203
rect 36 102 70 135
rect 122 237 156 270
rect 122 169 156 203
rect 122 20 156 135
rect 280 261 348 270
rect 280 203 297 261
rect 331 203 348 261
rect 280 169 348 203
rect 280 135 297 169
rect 331 135 348 169
rect 280 102 348 135
rect 472 237 506 270
rect 472 169 506 203
rect 472 20 506 135
rect 630 261 698 270
rect 630 203 647 261
rect 681 203 698 261
rect 630 169 698 203
rect 630 135 647 169
rect 681 135 698 169
rect 630 102 698 135
rect 822 237 856 270
rect 822 169 856 203
rect 822 20 856 135
rect 908 261 942 271
rect 908 169 942 203
rect 908 102 942 135
rect 1012 237 1046 270
rect 1012 169 1046 203
rect 1012 20 1046 135
rect 1098 261 1132 271
rect 1098 169 1132 203
rect 1098 102 1132 135
rect 0 17 1168 20
rect 0 -17 52 17
rect 86 -17 188 17
rect 222 -17 324 17
rect 358 -17 460 17
rect 494 -17 596 17
rect 630 -17 732 17
rect 766 -17 868 17
rect 902 -17 1004 17
rect 1038 -17 1168 17
rect 0 -20 1168 -17
<< viali >>
rect 36 787 70 821
rect 297 787 331 821
rect 647 787 681 821
rect 908 787 942 821
rect 1098 787 1132 821
rect 379 707 413 741
rect 113 627 147 661
rect 153 547 187 581
rect 36 467 70 501
rect 1098 618 1132 652
rect 908 467 942 501
rect 1020 467 1043 501
rect 1043 467 1054 501
rect 379 387 413 421
rect 36 237 70 261
rect 36 227 70 237
rect 297 237 331 261
rect 297 227 331 237
rect 647 237 681 261
rect 647 227 681 237
rect 908 237 942 261
rect 908 227 942 237
rect 1098 237 1132 261
rect 1098 227 1132 237
<< metal1 >>
rect 24 821 82 827
rect 24 787 36 821
rect 70 787 82 821
rect 24 781 82 787
rect 285 821 343 827
rect 285 787 297 821
rect 331 787 343 821
rect 285 781 343 787
rect 635 821 693 827
rect 635 787 647 821
rect 681 787 693 821
rect 635 781 693 787
rect 896 821 954 827
rect 896 787 908 821
rect 942 787 954 821
rect 896 781 954 787
rect 1086 821 1144 827
rect 1086 787 1098 821
rect 1132 787 1144 821
rect 1086 781 1144 787
rect 36 507 70 781
rect 101 661 159 667
rect 297 661 331 781
rect 369 750 423 756
rect 369 747 370 750
rect 367 701 370 747
rect 422 747 423 750
rect 369 698 370 701
rect 422 701 425 747
rect 422 698 423 701
rect 369 692 423 698
rect 101 627 113 661
rect 147 627 331 661
rect 101 621 159 627
rect 137 538 144 590
rect 196 538 203 590
rect 24 501 82 507
rect 24 467 36 501
rect 70 467 82 501
rect 24 461 82 467
rect 36 267 70 461
rect 297 267 331 627
rect 379 436 413 692
rect 369 427 423 436
rect 367 421 425 427
rect 367 387 379 421
rect 413 387 425 421
rect 367 381 425 387
rect 369 372 423 381
rect 647 267 681 781
rect 908 507 942 781
rect 1098 661 1132 781
rect 1082 609 1089 661
rect 1141 609 1148 661
rect 896 501 954 507
rect 896 467 908 501
rect 942 467 954 501
rect 896 461 954 467
rect 908 267 942 461
rect 1004 458 1011 510
rect 1063 458 1070 510
rect 1098 267 1132 609
rect 24 261 82 267
rect 24 227 36 261
rect 70 227 82 261
rect 24 221 82 227
rect 285 261 343 267
rect 285 227 297 261
rect 331 227 343 261
rect 285 221 343 227
rect 635 261 693 267
rect 635 227 647 261
rect 681 227 693 261
rect 635 221 693 227
rect 896 261 954 267
rect 896 227 908 261
rect 942 227 954 261
rect 896 221 954 227
rect 1086 261 1144 267
rect 1086 227 1098 261
rect 1132 227 1144 261
rect 1086 221 1144 227
<< via1 >>
rect 370 741 422 750
rect 370 707 379 741
rect 379 707 413 741
rect 413 707 422 741
rect 370 698 422 707
rect 144 581 196 590
rect 144 547 153 581
rect 153 547 187 581
rect 187 547 196 581
rect 144 538 196 547
rect 1089 652 1141 661
rect 1089 618 1098 652
rect 1098 618 1132 652
rect 1132 618 1141 652
rect 1089 609 1141 618
rect 1011 501 1063 510
rect 1011 467 1020 501
rect 1020 467 1054 501
rect 1054 467 1063 501
rect 1011 458 1063 467
<< metal2 >>
rect 369 750 423 756
rect 369 698 370 750
rect 422 698 423 750
rect 369 692 423 698
rect 1082 609 1089 661
rect 1141 609 1148 661
rect 137 538 144 590
rect 196 538 203 590
rect 1004 458 1011 510
rect 1063 458 1070 510
<< labels >>
rlabel locali s 544 0 544 0 4 gnd
rlabel locali s 548 1416 548 1416 4 vdd
rlabel locali s 584 1414 584 1414 4 vdd
port 4 nsew
rlabel locali s 584 0 584 0 4 gnd
port 5 nsew
rlabel metal2 s 1146 659 1146 659 4 Q
port 2 nsew
rlabel metal2 s 419 753 419 753 4 clk
port 3 nsew
rlabel metal2 s 1007 504 1007 504 4 ON
port 5 nsew
rlabel metal2 s 139 586 139 586 4 D
port 1 nsew
rlabel metal2 s 170 564 170 564 4 D
port 1 nsew
rlabel metal2 s 1115 635 1115 635 4 Q
port 2 nsew
rlabel metal2 s 396 724 396 724 4 clk
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1168 1414
string GDS_END 96512
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 75892
<< end >>
