magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect 56 1081 1082 1486
rect 56 931 550 1081
<< pwell >>
rect 183 591 973 843
rect 1143 732 2189 1314
rect 657 96 2090 389
rect 146 10 2090 96
<< mvnmos >>
rect 736 163 836 363
rect 892 163 992 363
rect 1048 163 1148 363
rect 1204 163 1304 363
rect 1476 163 1576 363
rect 1632 163 1732 363
rect 1911 163 2011 363
<< mvpmos >>
rect 175 997 275 1297
rect 331 997 431 1297
rect 597 1147 697 1297
rect 863 1147 963 1297
<< mvnnmos >>
rect 1222 1088 1402 1288
rect 1458 1088 1638 1288
rect 1694 1088 1874 1288
rect 1930 1088 2110 1288
rect 1222 758 1402 958
rect 1458 758 1638 958
rect 1694 758 1874 958
rect 1930 758 2110 958
<< nmoslvt >>
rect 262 617 292 817
rect 348 617 378 817
rect 434 617 464 817
rect 520 617 550 817
rect 606 617 636 817
rect 692 617 722 817
rect 778 617 808 817
rect 864 617 894 817
<< ndiff >>
rect 209 805 262 817
rect 209 771 217 805
rect 251 771 262 805
rect 209 737 262 771
rect 209 703 217 737
rect 251 703 262 737
rect 209 669 262 703
rect 209 635 217 669
rect 251 635 262 669
rect 209 617 262 635
rect 292 805 348 817
rect 292 771 303 805
rect 337 771 348 805
rect 292 737 348 771
rect 292 703 303 737
rect 337 703 348 737
rect 292 669 348 703
rect 292 635 303 669
rect 337 635 348 669
rect 292 617 348 635
rect 378 805 434 817
rect 378 771 389 805
rect 423 771 434 805
rect 378 737 434 771
rect 378 703 389 737
rect 423 703 434 737
rect 378 669 434 703
rect 378 635 389 669
rect 423 635 434 669
rect 378 617 434 635
rect 464 805 520 817
rect 464 771 475 805
rect 509 771 520 805
rect 464 737 520 771
rect 464 703 475 737
rect 509 703 520 737
rect 464 669 520 703
rect 464 635 475 669
rect 509 635 520 669
rect 464 617 520 635
rect 550 805 606 817
rect 550 771 561 805
rect 595 771 606 805
rect 550 737 606 771
rect 550 703 561 737
rect 595 703 606 737
rect 550 669 606 703
rect 550 635 561 669
rect 595 635 606 669
rect 550 617 606 635
rect 636 805 692 817
rect 636 771 647 805
rect 681 771 692 805
rect 636 737 692 771
rect 636 703 647 737
rect 681 703 692 737
rect 636 669 692 703
rect 636 635 647 669
rect 681 635 692 669
rect 636 617 692 635
rect 722 805 778 817
rect 722 771 733 805
rect 767 771 778 805
rect 722 737 778 771
rect 722 703 733 737
rect 767 703 778 737
rect 722 669 778 703
rect 722 635 733 669
rect 767 635 778 669
rect 722 617 778 635
rect 808 805 864 817
rect 808 771 819 805
rect 853 771 864 805
rect 808 737 864 771
rect 808 703 819 737
rect 853 703 864 737
rect 808 669 864 703
rect 808 635 819 669
rect 853 635 864 669
rect 808 617 864 635
rect 894 805 947 817
rect 894 771 905 805
rect 939 771 947 805
rect 894 737 947 771
rect 894 703 905 737
rect 939 703 947 737
rect 894 669 947 703
rect 894 635 905 669
rect 939 635 947 669
rect 894 617 947 635
<< mvndiff >>
rect 1169 1276 1222 1288
rect 1169 1242 1177 1276
rect 1211 1242 1222 1276
rect 1169 1208 1222 1242
rect 1169 1174 1177 1208
rect 1211 1174 1222 1208
rect 1169 1140 1222 1174
rect 1169 1106 1177 1140
rect 1211 1106 1222 1140
rect 1169 1088 1222 1106
rect 1402 1276 1458 1288
rect 1402 1242 1413 1276
rect 1447 1242 1458 1276
rect 1402 1208 1458 1242
rect 1402 1174 1413 1208
rect 1447 1174 1458 1208
rect 1402 1140 1458 1174
rect 1402 1106 1413 1140
rect 1447 1106 1458 1140
rect 1402 1088 1458 1106
rect 1638 1276 1694 1288
rect 1638 1242 1649 1276
rect 1683 1242 1694 1276
rect 1638 1208 1694 1242
rect 1638 1174 1649 1208
rect 1683 1174 1694 1208
rect 1638 1140 1694 1174
rect 1638 1106 1649 1140
rect 1683 1106 1694 1140
rect 1638 1088 1694 1106
rect 1874 1276 1930 1288
rect 1874 1242 1885 1276
rect 1919 1242 1930 1276
rect 1874 1208 1930 1242
rect 1874 1174 1885 1208
rect 1919 1174 1930 1208
rect 1874 1140 1930 1174
rect 1874 1106 1885 1140
rect 1919 1106 1930 1140
rect 1874 1088 1930 1106
rect 2110 1276 2163 1288
rect 2110 1242 2121 1276
rect 2155 1242 2163 1276
rect 2110 1208 2163 1242
rect 2110 1174 2121 1208
rect 2155 1174 2163 1208
rect 2110 1140 2163 1174
rect 2110 1106 2121 1140
rect 2155 1106 2163 1140
rect 2110 1088 2163 1106
rect 1169 940 1222 958
rect 1169 906 1177 940
rect 1211 906 1222 940
rect 1169 872 1222 906
rect 1169 838 1177 872
rect 1211 838 1222 872
rect 1169 804 1222 838
rect 1169 770 1177 804
rect 1211 770 1222 804
rect 1169 758 1222 770
rect 1402 940 1458 958
rect 1402 906 1413 940
rect 1447 906 1458 940
rect 1402 872 1458 906
rect 1402 838 1413 872
rect 1447 838 1458 872
rect 1402 804 1458 838
rect 1402 770 1413 804
rect 1447 770 1458 804
rect 1402 758 1458 770
rect 1638 940 1694 958
rect 1638 906 1649 940
rect 1683 906 1694 940
rect 1638 872 1694 906
rect 1638 838 1649 872
rect 1683 838 1694 872
rect 1638 804 1694 838
rect 1638 770 1649 804
rect 1683 770 1694 804
rect 1638 758 1694 770
rect 1874 940 1930 958
rect 1874 906 1885 940
rect 1919 906 1930 940
rect 1874 872 1930 906
rect 1874 838 1885 872
rect 1919 838 1930 872
rect 1874 804 1930 838
rect 1874 770 1885 804
rect 1919 770 1930 804
rect 1874 758 1930 770
rect 2110 940 2163 958
rect 2110 906 2121 940
rect 2155 906 2163 940
rect 2110 872 2163 906
rect 2110 838 2121 872
rect 2155 838 2163 872
rect 2110 804 2163 838
rect 2110 770 2121 804
rect 2155 770 2163 804
rect 2110 758 2163 770
rect 683 345 736 363
rect 683 311 691 345
rect 725 311 736 345
rect 683 277 736 311
rect 683 243 691 277
rect 725 243 736 277
rect 683 209 736 243
rect 683 175 691 209
rect 725 175 736 209
rect 683 163 736 175
rect 836 345 892 363
rect 836 311 847 345
rect 881 311 892 345
rect 836 277 892 311
rect 836 243 847 277
rect 881 243 892 277
rect 836 209 892 243
rect 836 175 847 209
rect 881 175 892 209
rect 836 163 892 175
rect 992 345 1048 363
rect 992 311 1003 345
rect 1037 311 1048 345
rect 992 277 1048 311
rect 992 243 1003 277
rect 1037 243 1048 277
rect 992 209 1048 243
rect 992 175 1003 209
rect 1037 175 1048 209
rect 992 163 1048 175
rect 1148 345 1204 363
rect 1148 311 1159 345
rect 1193 311 1204 345
rect 1148 277 1204 311
rect 1148 243 1159 277
rect 1193 243 1204 277
rect 1148 209 1204 243
rect 1148 175 1159 209
rect 1193 175 1204 209
rect 1148 163 1204 175
rect 1304 345 1357 363
rect 1304 311 1315 345
rect 1349 311 1357 345
rect 1304 277 1357 311
rect 1304 243 1315 277
rect 1349 243 1357 277
rect 1304 209 1357 243
rect 1304 175 1315 209
rect 1349 175 1357 209
rect 1304 163 1357 175
rect 1423 351 1476 363
rect 1423 317 1431 351
rect 1465 317 1476 351
rect 1423 283 1476 317
rect 1423 249 1431 283
rect 1465 249 1476 283
rect 1423 215 1476 249
rect 1423 181 1431 215
rect 1465 181 1476 215
rect 1423 163 1476 181
rect 1576 351 1632 363
rect 1576 317 1587 351
rect 1621 317 1632 351
rect 1576 283 1632 317
rect 1576 249 1587 283
rect 1621 249 1632 283
rect 1576 215 1632 249
rect 1576 181 1587 215
rect 1621 181 1632 215
rect 1576 163 1632 181
rect 1732 351 1785 363
rect 1732 317 1743 351
rect 1777 317 1785 351
rect 1732 283 1785 317
rect 1732 249 1743 283
rect 1777 249 1785 283
rect 1732 215 1785 249
rect 1732 181 1743 215
rect 1777 181 1785 215
rect 1732 163 1785 181
rect 1858 351 1911 363
rect 1858 317 1866 351
rect 1900 317 1911 351
rect 1858 283 1911 317
rect 1858 249 1866 283
rect 1900 249 1911 283
rect 1858 215 1911 249
rect 1858 181 1866 215
rect 1900 181 1911 215
rect 1858 163 1911 181
rect 2011 351 2064 363
rect 2011 317 2022 351
rect 2056 317 2064 351
rect 2011 283 2064 317
rect 2011 249 2022 283
rect 2056 249 2064 283
rect 2011 215 2064 249
rect 2011 181 2022 215
rect 2056 181 2064 215
rect 2011 163 2064 181
<< mvpdiff >>
rect 122 1285 175 1297
rect 122 1251 130 1285
rect 164 1251 175 1285
rect 122 1217 175 1251
rect 122 1183 130 1217
rect 164 1183 175 1217
rect 122 1149 175 1183
rect 122 1115 130 1149
rect 164 1115 175 1149
rect 122 1081 175 1115
rect 122 1047 130 1081
rect 164 1047 175 1081
rect 122 997 175 1047
rect 275 1285 331 1297
rect 275 1251 286 1285
rect 320 1251 331 1285
rect 275 1217 331 1251
rect 275 1183 286 1217
rect 320 1183 331 1217
rect 275 1149 331 1183
rect 275 1115 286 1149
rect 320 1115 331 1149
rect 275 1081 331 1115
rect 275 1047 286 1081
rect 320 1047 331 1081
rect 275 997 331 1047
rect 431 1285 484 1297
rect 431 1251 442 1285
rect 476 1251 484 1285
rect 431 1217 484 1251
rect 431 1183 442 1217
rect 476 1183 484 1217
rect 431 1149 484 1183
rect 431 1115 442 1149
rect 476 1115 484 1149
rect 544 1285 597 1297
rect 544 1251 552 1285
rect 586 1251 597 1285
rect 544 1217 597 1251
rect 544 1183 552 1217
rect 586 1183 597 1217
rect 544 1147 597 1183
rect 697 1285 750 1297
rect 697 1251 708 1285
rect 742 1251 750 1285
rect 697 1217 750 1251
rect 697 1183 708 1217
rect 742 1183 750 1217
rect 697 1147 750 1183
rect 810 1285 863 1297
rect 810 1251 818 1285
rect 852 1251 863 1285
rect 810 1217 863 1251
rect 810 1183 818 1217
rect 852 1183 863 1217
rect 810 1147 863 1183
rect 963 1285 1016 1297
rect 963 1251 974 1285
rect 1008 1251 1016 1285
rect 963 1217 1016 1251
rect 963 1183 974 1217
rect 1008 1183 1016 1217
rect 963 1147 1016 1183
rect 431 1081 484 1115
rect 431 1047 442 1081
rect 476 1047 484 1081
rect 431 997 484 1047
<< ndiffc >>
rect 217 771 251 805
rect 217 703 251 737
rect 217 635 251 669
rect 303 771 337 805
rect 303 703 337 737
rect 303 635 337 669
rect 389 771 423 805
rect 389 703 423 737
rect 389 635 423 669
rect 475 771 509 805
rect 475 703 509 737
rect 475 635 509 669
rect 561 771 595 805
rect 561 703 595 737
rect 561 635 595 669
rect 647 771 681 805
rect 647 703 681 737
rect 647 635 681 669
rect 733 771 767 805
rect 733 703 767 737
rect 733 635 767 669
rect 819 771 853 805
rect 819 703 853 737
rect 819 635 853 669
rect 905 771 939 805
rect 905 703 939 737
rect 905 635 939 669
<< mvndiffc >>
rect 1177 1242 1211 1276
rect 1177 1174 1211 1208
rect 1177 1106 1211 1140
rect 1413 1242 1447 1276
rect 1413 1174 1447 1208
rect 1413 1106 1447 1140
rect 1649 1242 1683 1276
rect 1649 1174 1683 1208
rect 1649 1106 1683 1140
rect 1885 1242 1919 1276
rect 1885 1174 1919 1208
rect 1885 1106 1919 1140
rect 2121 1242 2155 1276
rect 2121 1174 2155 1208
rect 2121 1106 2155 1140
rect 1177 906 1211 940
rect 1177 838 1211 872
rect 1177 770 1211 804
rect 1413 906 1447 940
rect 1413 838 1447 872
rect 1413 770 1447 804
rect 1649 906 1683 940
rect 1649 838 1683 872
rect 1649 770 1683 804
rect 1885 906 1919 940
rect 1885 838 1919 872
rect 1885 770 1919 804
rect 2121 906 2155 940
rect 2121 838 2155 872
rect 2121 770 2155 804
rect 691 311 725 345
rect 691 243 725 277
rect 691 175 725 209
rect 847 311 881 345
rect 847 243 881 277
rect 847 175 881 209
rect 1003 311 1037 345
rect 1003 243 1037 277
rect 1003 175 1037 209
rect 1159 311 1193 345
rect 1159 243 1193 277
rect 1159 175 1193 209
rect 1315 311 1349 345
rect 1315 243 1349 277
rect 1315 175 1349 209
rect 1431 317 1465 351
rect 1431 249 1465 283
rect 1431 181 1465 215
rect 1587 317 1621 351
rect 1587 249 1621 283
rect 1587 181 1621 215
rect 1743 317 1777 351
rect 1743 249 1777 283
rect 1743 181 1777 215
rect 1866 317 1900 351
rect 1866 249 1900 283
rect 1866 181 1900 215
rect 2022 317 2056 351
rect 2022 249 2056 283
rect 2022 181 2056 215
<< mvpdiffc >>
rect 130 1251 164 1285
rect 130 1183 164 1217
rect 130 1115 164 1149
rect 130 1047 164 1081
rect 286 1251 320 1285
rect 286 1183 320 1217
rect 286 1115 320 1149
rect 286 1047 320 1081
rect 442 1251 476 1285
rect 442 1183 476 1217
rect 442 1115 476 1149
rect 552 1251 586 1285
rect 552 1183 586 1217
rect 708 1251 742 1285
rect 708 1183 742 1217
rect 818 1251 852 1285
rect 818 1183 852 1217
rect 974 1251 1008 1285
rect 974 1183 1008 1217
rect 442 1047 476 1081
<< mvpsubdiff >>
rect 172 36 196 70
rect 230 36 266 70
rect 300 36 336 70
rect 370 36 406 70
rect 440 36 476 70
rect 510 36 546 70
rect 580 36 616 70
rect 650 36 686 70
rect 720 36 756 70
rect 790 36 826 70
rect 860 36 896 70
rect 930 36 966 70
rect 1000 36 1036 70
rect 1070 36 1106 70
rect 1140 36 1176 70
rect 1210 36 1246 70
rect 1280 36 1316 70
rect 1350 36 1385 70
rect 1419 36 1454 70
rect 1488 36 1523 70
rect 1557 36 1592 70
rect 1626 36 1661 70
rect 1695 36 1730 70
rect 1764 36 1799 70
rect 1833 36 1868 70
rect 1902 36 1937 70
rect 1971 36 2006 70
rect 2040 36 2064 70
<< mvnsubdiff >>
rect 122 1386 146 1420
rect 180 1386 220 1420
rect 254 1386 294 1420
rect 328 1386 368 1420
rect 402 1386 442 1420
rect 476 1386 516 1420
rect 550 1386 590 1420
rect 624 1386 664 1420
rect 698 1386 738 1420
rect 772 1386 812 1420
rect 846 1386 885 1420
rect 919 1386 958 1420
rect 992 1386 1016 1420
<< mvpsubdiffcont >>
rect 196 36 230 70
rect 266 36 300 70
rect 336 36 370 70
rect 406 36 440 70
rect 476 36 510 70
rect 546 36 580 70
rect 616 36 650 70
rect 686 36 720 70
rect 756 36 790 70
rect 826 36 860 70
rect 896 36 930 70
rect 966 36 1000 70
rect 1036 36 1070 70
rect 1106 36 1140 70
rect 1176 36 1210 70
rect 1246 36 1280 70
rect 1316 36 1350 70
rect 1385 36 1419 70
rect 1454 36 1488 70
rect 1523 36 1557 70
rect 1592 36 1626 70
rect 1661 36 1695 70
rect 1730 36 1764 70
rect 1799 36 1833 70
rect 1868 36 1902 70
rect 1937 36 1971 70
rect 2006 36 2040 70
<< mvnsubdiffcont >>
rect 146 1386 180 1420
rect 220 1386 254 1420
rect 294 1386 328 1420
rect 368 1386 402 1420
rect 442 1386 476 1420
rect 516 1386 550 1420
rect 590 1386 624 1420
rect 664 1386 698 1420
rect 738 1386 772 1420
rect 812 1386 846 1420
rect 885 1386 919 1420
rect 958 1386 992 1420
<< poly >>
rect 175 1297 275 1329
rect 331 1297 431 1329
rect 597 1297 697 1329
rect 863 1297 963 1329
rect 1222 1288 1402 1320
rect 1458 1288 1638 1320
rect 1694 1288 1874 1320
rect 1930 1288 2110 1320
rect 597 1089 697 1147
rect 863 1115 963 1147
rect 862 1111 963 1115
rect 597 1055 631 1089
rect 665 1055 697 1089
rect 597 1021 697 1055
rect 812 1095 963 1111
rect 812 1061 828 1095
rect 862 1061 896 1095
rect 930 1061 963 1095
rect 812 1045 963 1061
rect 1222 1056 1402 1088
rect 1458 1056 1638 1088
rect 1694 1056 1874 1088
rect 1930 1056 2110 1088
rect 175 965 275 997
rect 141 949 275 965
rect 141 915 157 949
rect 191 915 225 949
rect 259 915 275 949
rect 141 899 275 915
rect 331 965 431 997
rect 597 987 631 1021
rect 665 987 697 1021
rect 597 971 697 987
rect 1222 1040 2110 1056
rect 1222 1006 1238 1040
rect 1272 1006 1306 1040
rect 1340 1006 1374 1040
rect 1408 1006 1442 1040
rect 1476 1006 1510 1040
rect 1544 1006 1578 1040
rect 1612 1006 1646 1040
rect 1680 1006 1715 1040
rect 1749 1006 1784 1040
rect 1818 1006 1853 1040
rect 1887 1006 1922 1040
rect 1956 1006 1991 1040
rect 2025 1006 2060 1040
rect 2094 1006 2110 1040
rect 1222 990 2110 1006
rect 331 949 465 965
rect 1222 958 1402 990
rect 1458 958 1638 990
rect 1694 958 1874 990
rect 1930 958 2110 990
rect 331 915 347 949
rect 381 915 415 949
rect 449 915 465 949
rect 331 899 465 915
rect 262 817 292 849
rect 348 817 378 849
rect 434 817 464 849
rect 520 817 550 849
rect 606 817 636 849
rect 692 817 722 849
rect 778 817 808 849
rect 864 817 894 849
rect 1222 726 1402 758
rect 1458 726 1638 758
rect 1694 726 1874 758
rect 1930 726 2110 758
rect 262 585 292 617
rect 348 585 378 617
rect 434 585 464 617
rect 520 585 550 617
rect 262 569 550 585
rect 262 535 278 569
rect 312 535 352 569
rect 386 535 426 569
rect 460 535 500 569
rect 534 535 550 569
rect 262 519 550 535
rect 606 585 636 617
rect 692 585 722 617
rect 778 585 808 617
rect 864 585 894 617
rect 606 569 894 585
rect 606 535 622 569
rect 656 535 696 569
rect 730 535 770 569
rect 804 535 844 569
rect 878 535 894 569
rect 606 519 894 535
rect 1476 517 1576 537
rect 1476 483 1506 517
rect 1540 483 1576 517
rect 736 439 1304 455
rect 736 405 752 439
rect 786 405 823 439
rect 857 405 894 439
rect 928 405 966 439
rect 1000 405 1038 439
rect 1072 405 1110 439
rect 1144 405 1182 439
rect 1216 405 1254 439
rect 1288 405 1304 439
rect 736 389 1304 405
rect 736 363 836 389
rect 892 363 992 389
rect 1048 363 1148 389
rect 1204 363 1304 389
rect 1476 449 1576 483
rect 1476 415 1506 449
rect 1540 415 1576 449
rect 1476 363 1576 415
rect 1632 517 1732 533
rect 1632 483 1669 517
rect 1703 483 1732 517
rect 1632 449 1732 483
rect 1632 415 1669 449
rect 1703 415 1732 449
rect 1632 363 1732 415
rect 1911 517 2011 533
rect 1911 483 1947 517
rect 1981 483 2011 517
rect 1911 449 2011 483
rect 1911 415 1947 449
rect 1981 415 2011 449
rect 1911 363 2011 415
rect 736 137 836 163
rect 892 137 992 163
rect 1048 137 1148 163
rect 1204 137 1304 163
rect 1476 131 1576 163
rect 1632 131 1732 163
rect 1911 131 2011 163
<< polycont >>
rect 631 1055 665 1089
rect 828 1061 862 1095
rect 896 1061 930 1095
rect 157 915 191 949
rect 225 915 259 949
rect 631 987 665 1021
rect 1238 1006 1272 1040
rect 1306 1006 1340 1040
rect 1374 1006 1408 1040
rect 1442 1006 1476 1040
rect 1510 1006 1544 1040
rect 1578 1006 1612 1040
rect 1646 1006 1680 1040
rect 1715 1006 1749 1040
rect 1784 1006 1818 1040
rect 1853 1006 1887 1040
rect 1922 1006 1956 1040
rect 1991 1006 2025 1040
rect 2060 1006 2094 1040
rect 347 915 381 949
rect 415 915 449 949
rect 278 535 312 569
rect 352 535 386 569
rect 426 535 460 569
rect 500 535 534 569
rect 622 535 656 569
rect 696 535 730 569
rect 770 535 804 569
rect 844 535 878 569
rect 1506 483 1540 517
rect 752 405 786 439
rect 823 405 857 439
rect 894 405 928 439
rect 966 405 1000 439
rect 1038 405 1072 439
rect 1110 405 1144 439
rect 1182 405 1216 439
rect 1254 405 1288 439
rect 1506 415 1540 449
rect 1669 483 1703 517
rect 1669 415 1703 449
rect 1947 483 1981 517
rect 1947 415 1981 449
<< locali >>
rect 122 1386 144 1420
rect 180 1386 220 1420
rect 254 1386 294 1420
rect 330 1386 368 1420
rect 406 1386 442 1420
rect 482 1386 516 1420
rect 558 1386 590 1420
rect 634 1386 664 1420
rect 710 1386 738 1420
rect 787 1386 812 1420
rect 864 1386 885 1420
rect 941 1386 958 1420
rect 130 1285 164 1301
rect 130 1217 164 1251
rect 286 1285 320 1314
rect 553 1301 587 1314
rect 286 1217 320 1242
rect 164 1183 178 1196
rect 140 1162 178 1183
rect 130 1149 164 1162
rect 130 1081 164 1115
rect 130 1031 164 1047
rect 286 1149 320 1183
rect 442 1285 476 1301
rect 442 1217 476 1251
rect 442 1149 476 1183
rect 552 1285 587 1301
rect 586 1276 587 1285
rect 552 1242 553 1251
rect 708 1285 784 1301
rect 742 1251 784 1285
rect 552 1217 586 1242
rect 552 1167 586 1183
rect 708 1217 784 1251
rect 742 1183 784 1217
rect 708 1167 784 1183
rect 818 1285 852 1314
rect 818 1217 852 1242
rect 818 1167 852 1183
rect 974 1285 1105 1301
rect 1008 1251 1105 1285
rect 974 1217 1105 1251
rect 1008 1183 1105 1217
rect 974 1167 1105 1183
rect 286 1081 320 1115
rect 406 1115 442 1120
rect 406 1086 444 1115
rect 629 1094 667 1128
rect 605 1089 701 1094
rect 286 1031 320 1047
rect 442 1081 476 1086
rect 442 1031 476 1047
rect 605 1055 631 1089
rect 665 1055 701 1089
rect 605 1021 701 1055
rect 605 997 631 1021
rect 331 987 631 997
rect 665 987 701 1021
rect 735 1095 784 1167
rect 980 1128 1105 1167
rect 735 1061 828 1095
rect 862 1061 896 1095
rect 930 1061 946 1095
rect 735 1037 946 1061
rect 735 1003 755 1037
rect 789 1003 829 1037
rect 863 1003 903 1037
rect 937 1003 946 1037
rect 980 1094 995 1128
rect 1029 1094 1071 1128
rect 331 969 701 987
rect 980 969 1105 1094
rect 1177 1276 1211 1292
rect 1177 1208 1211 1242
rect 1413 1276 1447 1292
rect 1413 1212 1447 1242
rect 1649 1276 1683 1292
rect 1412 1208 1450 1212
rect 1412 1178 1413 1208
rect 1177 1140 1211 1174
rect 1447 1178 1450 1208
rect 1649 1208 1683 1242
rect 1885 1276 1919 1292
rect 1885 1212 1919 1242
rect 2121 1276 2155 1292
rect 1413 1140 1447 1174
rect 1211 1096 1249 1130
rect 1883 1208 1921 1212
rect 1883 1178 1885 1208
rect 1649 1140 1683 1174
rect 1177 1090 1211 1096
rect 1413 1090 1447 1106
rect 1648 1106 1649 1130
rect 1919 1178 1921 1208
rect 2121 1208 2155 1242
rect 1885 1140 1919 1174
rect 1683 1106 1686 1130
rect 1648 1096 1686 1106
rect 2121 1140 2155 1174
rect 1649 1090 1683 1096
rect 1885 1090 1919 1106
rect 2083 1096 2121 1130
rect 2121 1090 2155 1096
rect 1399 1040 1439 1041
rect 1473 1040 1513 1041
rect 1547 1040 1587 1041
rect 1621 1040 1660 1041
rect 1694 1040 1733 1041
rect 1767 1040 1806 1041
rect 1840 1040 1879 1041
rect 1913 1040 1952 1041
rect 1222 1006 1238 1040
rect 1272 1006 1306 1040
rect 1340 1007 1365 1040
rect 1408 1007 1439 1040
rect 1340 1006 1374 1007
rect 1408 1006 1442 1007
rect 1476 1006 1510 1040
rect 1547 1007 1578 1040
rect 1621 1007 1646 1040
rect 1694 1007 1715 1040
rect 1767 1007 1784 1040
rect 1840 1007 1853 1040
rect 1913 1007 1922 1040
rect 1986 1007 1991 1040
rect 1544 1006 1578 1007
rect 1612 1006 1646 1007
rect 1680 1006 1715 1007
rect 1749 1006 1784 1007
rect 1818 1006 1853 1007
rect 1887 1006 1922 1007
rect 1956 1006 1991 1007
rect 2025 1006 2060 1040
rect 2094 1006 2110 1040
rect 191 949 229 963
rect 331 949 1105 969
rect 141 915 157 949
rect 191 915 225 949
rect 263 929 275 949
rect 259 915 275 929
rect 331 915 347 949
rect 381 915 415 949
rect 449 915 1105 949
rect 217 805 251 821
rect 217 737 251 771
rect 217 669 251 689
rect 303 809 337 847
rect 303 737 337 771
rect 303 669 337 703
rect 303 619 337 635
rect 389 805 423 821
rect 389 737 423 771
rect 389 669 423 689
rect 475 809 509 847
rect 475 737 509 771
rect 475 669 509 703
rect 475 619 509 635
rect 561 805 595 821
rect 561 737 595 771
rect 561 669 595 689
rect 647 809 681 847
rect 647 737 681 771
rect 647 669 681 703
rect 647 619 681 635
rect 733 805 767 821
rect 733 737 767 771
rect 733 669 767 689
rect 819 809 853 847
rect 819 737 853 771
rect 819 669 853 703
rect 819 619 853 635
rect 905 805 939 821
rect 905 737 939 771
rect 905 669 939 689
rect 973 570 1105 915
rect 1177 940 1211 956
rect 1413 940 1447 956
rect 1649 940 1683 956
rect 1885 946 1919 956
rect 1885 940 2006 946
rect 1412 906 1413 940
rect 1447 906 1450 940
rect 1883 906 1885 940
rect 1919 906 1921 940
rect 1955 906 2006 940
rect 1177 872 1211 906
rect 1177 804 1211 838
rect 1173 770 1177 795
rect 1413 872 1447 906
rect 1413 804 1447 838
rect 1173 761 1211 770
rect 1649 872 1683 906
rect 1649 804 1683 838
rect 1177 754 1211 761
rect 1413 754 1447 770
rect 1648 770 1649 795
rect 1885 872 2006 906
rect 1919 838 2006 872
rect 1885 804 2006 838
rect 1683 770 1686 795
rect 1648 761 1686 770
rect 1919 770 2006 804
rect 2121 940 2155 956
rect 2121 872 2155 906
rect 2121 804 2155 838
rect 1649 754 1683 761
rect 1885 754 2006 770
rect 2080 761 2118 795
rect 2152 761 2155 770
rect 2121 754 2155 761
rect 262 535 278 569
rect 324 535 352 569
rect 386 535 397 569
rect 460 535 500 569
rect 538 535 550 569
rect 606 535 622 569
rect 656 535 696 569
rect 762 535 770 569
rect 804 535 834 569
rect 878 535 894 569
rect 973 536 984 570
rect 1018 536 1056 570
rect 1090 536 1105 570
rect 1894 535 2006 754
rect 1506 517 1540 530
rect 1506 449 1540 458
rect 838 439 882 444
rect 916 439 960 444
rect 994 439 1038 444
rect 1072 439 1116 444
rect 1150 439 1194 444
rect 736 405 752 439
rect 786 410 804 439
rect 857 410 882 439
rect 928 410 960 439
rect 786 405 823 410
rect 857 405 894 410
rect 928 405 966 410
rect 1000 405 1038 439
rect 1072 405 1110 439
rect 1150 410 1182 439
rect 1228 410 1254 439
rect 1144 405 1182 410
rect 1216 405 1254 410
rect 1288 405 1304 439
rect 1506 399 1540 415
rect 1669 525 1703 533
rect 1669 453 1703 483
rect 1669 399 1703 415
rect 1894 501 1942 535
rect 1976 517 2006 535
rect 1894 483 1947 501
rect 1981 483 2006 517
rect 1894 463 2006 483
rect 1894 429 1942 463
rect 1976 449 2006 463
rect 1894 415 1947 429
rect 1981 415 2006 449
rect 1894 401 2006 415
rect 1947 399 1981 401
rect 1388 373 1472 385
rect 691 345 725 361
rect 862 345 900 370
rect 881 336 900 345
rect 1003 345 1037 361
rect 691 277 725 311
rect 691 214 725 243
rect 691 142 725 175
rect 847 277 881 311
rect 847 209 881 243
rect 847 159 881 175
rect 1161 345 1199 370
rect 1193 336 1199 345
rect 1315 345 1349 361
rect 1003 277 1037 311
rect 1003 214 1037 243
rect 1003 142 1037 175
rect 1159 277 1193 311
rect 1159 209 1193 243
rect 1159 159 1193 175
rect 1315 277 1349 311
rect 1315 214 1349 243
rect 1315 142 1349 175
rect 1388 317 1431 373
rect 1465 317 1472 373
rect 1388 301 1472 317
rect 1388 249 1431 301
rect 1465 249 1472 301
rect 1388 215 1472 249
rect 1388 181 1431 215
rect 1465 181 1472 215
rect 1388 159 1472 181
rect 1587 351 1621 367
rect 1743 351 1777 367
rect 1866 351 1900 367
rect 1587 283 1621 317
rect 1777 317 1788 339
rect 1750 305 1788 317
rect 1587 215 1621 249
rect 1587 142 1621 180
rect 1743 283 1777 305
rect 1743 215 1777 249
rect 1743 165 1777 181
rect 1866 283 1900 317
rect 1866 215 1900 249
rect 1866 142 1900 180
rect 2022 351 2056 367
rect 2022 294 2056 317
rect 2056 260 2094 294
rect 2022 215 2056 249
rect 2022 165 2056 181
rect 172 36 194 70
rect 230 36 266 70
rect 300 36 336 70
rect 372 36 406 70
rect 444 36 476 70
rect 516 36 546 70
rect 588 36 616 70
rect 660 36 686 70
rect 732 36 756 70
rect 804 36 826 70
rect 876 36 896 70
rect 948 36 966 70
rect 1020 36 1036 70
rect 1092 36 1106 70
rect 1165 36 1176 70
rect 1238 36 1246 70
rect 1311 36 1316 70
rect 1384 36 1385 70
rect 1419 36 1423 70
rect 1488 36 1496 70
rect 1557 36 1569 70
rect 1626 36 1642 70
rect 1695 36 1715 70
rect 1764 36 1788 70
rect 1833 36 1861 70
rect 1902 36 1934 70
rect 1971 36 2006 70
rect 2041 36 2080 70
<< viali >>
rect 144 1386 146 1420
rect 146 1386 178 1420
rect 220 1386 254 1420
rect 296 1386 328 1420
rect 328 1386 330 1420
rect 372 1386 402 1420
rect 402 1386 406 1420
rect 448 1386 476 1420
rect 476 1386 482 1420
rect 524 1386 550 1420
rect 550 1386 558 1420
rect 600 1386 624 1420
rect 624 1386 634 1420
rect 676 1386 698 1420
rect 698 1386 710 1420
rect 753 1386 772 1420
rect 772 1386 787 1420
rect 830 1386 846 1420
rect 846 1386 864 1420
rect 907 1386 919 1420
rect 919 1386 941 1420
rect 984 1386 992 1420
rect 992 1386 1018 1420
rect 286 1314 320 1348
rect 553 1314 587 1348
rect 818 1314 852 1348
rect 286 1251 320 1276
rect 286 1242 320 1251
rect 106 1183 130 1196
rect 130 1183 140 1196
rect 106 1162 140 1183
rect 178 1162 212 1196
rect 553 1251 586 1276
rect 586 1251 587 1276
rect 553 1242 587 1251
rect 818 1251 852 1276
rect 818 1242 852 1251
rect 372 1086 406 1120
rect 444 1115 476 1120
rect 476 1115 478 1120
rect 444 1086 478 1115
rect 595 1094 629 1128
rect 667 1094 701 1128
rect 755 1003 789 1037
rect 829 1003 863 1037
rect 903 1003 937 1037
rect 995 1094 1029 1128
rect 1071 1094 1105 1128
rect 1378 1178 1412 1212
rect 1450 1178 1484 1212
rect 1177 1106 1211 1130
rect 1177 1096 1211 1106
rect 1249 1096 1283 1130
rect 1849 1178 1883 1212
rect 1614 1096 1648 1130
rect 1921 1178 1955 1212
rect 1686 1096 1720 1130
rect 2049 1096 2083 1130
rect 2121 1106 2155 1130
rect 2121 1096 2155 1106
rect 1365 1040 1399 1041
rect 1439 1040 1473 1041
rect 1513 1040 1547 1041
rect 1587 1040 1621 1041
rect 1660 1040 1694 1041
rect 1733 1040 1767 1041
rect 1806 1040 1840 1041
rect 1879 1040 1913 1041
rect 1952 1040 1986 1041
rect 1365 1007 1374 1040
rect 1374 1007 1399 1040
rect 1439 1007 1442 1040
rect 1442 1007 1473 1040
rect 1513 1007 1544 1040
rect 1544 1007 1547 1040
rect 1587 1007 1612 1040
rect 1612 1007 1621 1040
rect 1660 1007 1680 1040
rect 1680 1007 1694 1040
rect 1733 1007 1749 1040
rect 1749 1007 1767 1040
rect 1806 1007 1818 1040
rect 1818 1007 1840 1040
rect 1879 1007 1887 1040
rect 1887 1007 1913 1040
rect 1952 1007 1956 1040
rect 1956 1007 1986 1040
rect 157 949 191 963
rect 229 949 263 963
rect 157 929 191 949
rect 229 929 259 949
rect 259 929 263 949
rect 303 847 337 881
rect 217 703 251 723
rect 217 689 251 703
rect 217 635 251 651
rect 217 617 251 635
rect 475 847 509 881
rect 303 805 337 809
rect 303 775 337 805
rect 389 703 423 723
rect 389 689 423 703
rect 389 635 423 651
rect 389 617 423 635
rect 647 847 681 881
rect 475 805 509 809
rect 475 775 509 805
rect 561 703 595 723
rect 561 689 595 703
rect 561 635 595 651
rect 561 617 595 635
rect 819 847 853 881
rect 647 805 681 809
rect 647 775 681 805
rect 733 703 767 723
rect 733 689 767 703
rect 733 635 767 651
rect 733 617 767 635
rect 819 805 853 809
rect 819 775 853 805
rect 905 703 939 723
rect 905 689 939 703
rect 905 635 939 651
rect 905 617 939 635
rect 1378 906 1412 940
rect 1450 906 1484 940
rect 1849 906 1883 940
rect 1921 906 1955 940
rect 1139 761 1173 795
rect 1211 761 1245 795
rect 1614 761 1648 795
rect 1686 761 1720 795
rect 2046 761 2080 795
rect 2118 770 2121 795
rect 2121 770 2152 795
rect 2118 761 2152 770
rect 290 535 312 569
rect 312 535 324 569
rect 397 535 426 569
rect 426 535 431 569
rect 504 535 534 569
rect 534 535 538 569
rect 622 535 656 569
rect 728 535 730 569
rect 730 535 762 569
rect 834 535 844 569
rect 844 535 868 569
rect 984 536 1018 570
rect 1056 536 1090 570
rect 1506 530 1540 564
rect 1506 483 1540 492
rect 1506 458 1540 483
rect 804 439 838 444
rect 882 439 916 444
rect 960 439 994 444
rect 1038 439 1072 444
rect 1116 439 1150 444
rect 1194 439 1228 444
rect 804 410 823 439
rect 823 410 838 439
rect 882 410 894 439
rect 894 410 916 439
rect 960 410 966 439
rect 966 410 994 439
rect 1038 410 1072 439
rect 1116 410 1144 439
rect 1144 410 1150 439
rect 1194 410 1216 439
rect 1216 410 1228 439
rect 1669 517 1703 525
rect 1669 491 1703 517
rect 1669 449 1703 453
rect 1669 419 1703 449
rect 1942 517 1976 535
rect 1942 501 1947 517
rect 1947 501 1976 517
rect 1942 449 1976 463
rect 1942 429 1947 449
rect 1947 429 1976 449
rect 828 345 862 370
rect 828 336 847 345
rect 847 336 862 345
rect 900 336 934 370
rect 691 209 725 214
rect 691 180 725 209
rect 1127 345 1161 370
rect 1127 336 1159 345
rect 1159 336 1161 345
rect 1199 336 1233 370
rect 1003 209 1037 214
rect 1003 180 1037 209
rect 691 108 725 142
rect 1315 209 1349 214
rect 1315 180 1349 209
rect 1003 108 1037 142
rect 1431 351 1465 373
rect 1431 339 1465 351
rect 1431 283 1465 301
rect 1431 267 1465 283
rect 1716 317 1743 339
rect 1743 317 1750 339
rect 1716 305 1750 317
rect 1788 305 1822 339
rect 1587 181 1621 214
rect 1587 180 1621 181
rect 1315 108 1349 142
rect 1866 181 1900 214
rect 1866 180 1900 181
rect 1587 108 1621 142
rect 2022 283 2056 294
rect 2022 260 2056 283
rect 2094 260 2128 294
rect 1866 108 1900 142
rect 194 36 196 70
rect 196 36 228 70
rect 266 36 300 70
rect 338 36 370 70
rect 370 36 372 70
rect 410 36 440 70
rect 440 36 444 70
rect 482 36 510 70
rect 510 36 516 70
rect 554 36 580 70
rect 580 36 588 70
rect 626 36 650 70
rect 650 36 660 70
rect 698 36 720 70
rect 720 36 732 70
rect 770 36 790 70
rect 790 36 804 70
rect 842 36 860 70
rect 860 36 876 70
rect 914 36 930 70
rect 930 36 948 70
rect 986 36 1000 70
rect 1000 36 1020 70
rect 1058 36 1070 70
rect 1070 36 1092 70
rect 1131 36 1140 70
rect 1140 36 1165 70
rect 1204 36 1210 70
rect 1210 36 1238 70
rect 1277 36 1280 70
rect 1280 36 1311 70
rect 1350 36 1384 70
rect 1423 36 1454 70
rect 1454 36 1457 70
rect 1496 36 1523 70
rect 1523 36 1530 70
rect 1569 36 1592 70
rect 1592 36 1603 70
rect 1642 36 1661 70
rect 1661 36 1676 70
rect 1715 36 1730 70
rect 1730 36 1749 70
rect 1788 36 1799 70
rect 1799 36 1822 70
rect 1861 36 1868 70
rect 1868 36 1895 70
rect 1934 36 1937 70
rect 1937 36 1968 70
rect 2007 36 2040 70
rect 2040 36 2041 70
rect 2080 36 2114 70
<< metal1 >>
rect 115 1420 1048 1426
rect 115 1386 144 1420
rect 178 1386 220 1420
rect 254 1386 296 1420
rect 330 1386 372 1420
rect 406 1386 448 1420
rect 482 1386 524 1420
rect 558 1386 600 1420
rect 634 1386 676 1420
rect 710 1386 753 1420
rect 787 1386 830 1420
rect 864 1386 907 1420
rect 941 1386 984 1420
rect 1018 1386 1048 1420
rect 115 1348 1048 1386
rect 115 1314 286 1348
rect 320 1314 553 1348
rect 587 1314 818 1348
rect 852 1333 1048 1348
rect 852 1314 1009 1333
rect 115 1294 1009 1314
tri 1009 1294 1048 1333 nw
rect 115 1276 951 1294
rect 115 1242 286 1276
rect 320 1242 553 1276
rect 587 1242 818 1276
rect 852 1242 951 1276
rect 115 1236 951 1242
tri 951 1236 1009 1294 nw
tri 1015 1236 1073 1294 se
rect 1073 1288 2113 1294
rect 1073 1254 2061 1288
tri 1073 1236 1091 1254 nw
tri 2028 1236 2046 1254 ne
rect 2046 1236 2061 1254
rect 115 1230 945 1236
tri 945 1230 951 1236 nw
tri 1009 1230 1015 1236 se
rect 1015 1230 1055 1236
tri 997 1218 1009 1230 se
rect 1009 1218 1055 1230
tri 1055 1218 1073 1236 nw
tri 2046 1221 2061 1236 ne
rect 2061 1224 2113 1236
tri 991 1212 997 1218 se
rect 997 1212 1049 1218
tri 1049 1212 1055 1218 nw
tri 1096 1212 1102 1218 se
rect 1102 1212 1967 1218
tri 981 1202 991 1212 se
rect 991 1202 1039 1212
tri 1039 1202 1049 1212 nw
tri 1086 1202 1096 1212 se
rect 1096 1202 1378 1212
rect 94 1196 1015 1202
rect 94 1162 106 1196
rect 140 1162 178 1196
rect 212 1178 1015 1196
tri 1015 1178 1039 1202 nw
tri 1062 1178 1086 1202 se
rect 1086 1178 1378 1202
rect 1412 1178 1450 1212
rect 1484 1178 1849 1212
rect 1883 1178 1921 1212
rect 1955 1178 1967 1212
rect 212 1172 1009 1178
tri 1009 1172 1015 1178 nw
tri 1056 1172 1062 1178 se
rect 1062 1172 1967 1178
rect 212 1162 999 1172
tri 999 1162 1009 1172 nw
tri 1046 1162 1056 1172 se
rect 1056 1166 1155 1172
tri 1155 1166 1161 1172 nw
rect 2061 1166 2113 1172
rect 1056 1162 1129 1166
rect 94 1156 258 1162
tri 258 1156 264 1162 nw
tri 1040 1156 1046 1162 se
rect 1046 1156 1129 1162
tri 1018 1134 1040 1156 se
rect 1040 1134 1129 1156
tri 1129 1140 1155 1166 nw
rect 583 1128 1129 1134
tri 74 1120 80 1126 se
rect 80 1120 490 1126
tri 53 1099 74 1120 se
rect 74 1099 372 1120
rect 53 1086 372 1099
rect 406 1086 444 1120
rect 478 1086 490 1120
rect 583 1094 595 1128
rect 629 1094 667 1128
rect 701 1094 995 1128
rect 1029 1094 1071 1128
rect 1105 1094 1129 1128
rect 583 1088 1129 1094
rect 1165 1130 2167 1136
rect 1165 1096 1177 1130
rect 1211 1096 1249 1130
rect 1283 1096 1614 1130
rect 1648 1096 1686 1130
rect 1720 1096 2049 1130
rect 2083 1096 2121 1130
rect 2155 1096 2167 1130
rect 1165 1090 2167 1096
tri 2045 1088 2047 1090 ne
rect 2047 1088 2125 1090
rect 53 1080 490 1086
tri 2047 1080 2055 1088 ne
rect 2055 1080 2125 1088
rect 53 1056 109 1080
tri 109 1056 133 1080 nw
tri 2055 1056 2079 1080 ne
rect 53 410 99 1056
tri 99 1046 109 1056 nw
tri 561 1041 563 1043 se
rect 563 1041 1019 1043
tri 1019 1041 1021 1043 sw
rect 1353 1041 1998 1047
tri 557 1037 561 1041 se
rect 561 1037 1021 1041
tri 532 1012 557 1037 se
rect 557 1012 755 1037
tri 523 1003 532 1012 se
rect 532 1003 755 1012
rect 789 1003 829 1037
rect 863 1003 903 1037
rect 937 1012 1021 1037
tri 1021 1012 1050 1041 sw
rect 937 1007 1050 1012
tri 1050 1007 1055 1012 sw
rect 1353 1007 1365 1041
rect 1399 1007 1439 1041
rect 1473 1007 1513 1041
rect 1547 1007 1587 1041
rect 1621 1007 1660 1041
rect 1694 1007 1733 1041
rect 1767 1007 1806 1041
rect 1840 1007 1879 1041
rect 1913 1007 1952 1041
rect 1986 1007 1998 1041
rect 937 1003 1055 1007
tri 497 977 523 1003 se
rect 523 997 1055 1003
rect 523 977 563 997
tri 563 977 583 997 nw
tri 999 977 1019 997 ne
rect 1019 977 1055 997
tri 489 969 497 977 se
rect 497 969 555 977
tri 555 969 563 977 nw
tri 1019 969 1027 977 ne
rect 1027 969 1055 977
rect 145 963 532 969
rect 145 929 157 963
rect 191 929 229 963
rect 263 946 532 963
tri 532 946 555 969 nw
tri 572 946 595 969 se
rect 595 946 972 969
tri 972 946 995 969 sw
tri 1027 946 1050 969 ne
rect 1050 946 1055 969
tri 1055 946 1116 1007 sw
rect 1353 1001 1998 1007
rect 263 943 529 946
tri 529 943 532 946 nw
tri 569 943 572 946 se
rect 572 943 995 946
rect 263 940 526 943
tri 526 940 529 943 nw
tri 566 940 569 943 se
rect 569 940 995 943
tri 995 940 1001 946 sw
tri 1050 940 1056 946 ne
rect 1056 940 1967 946
rect 263 929 509 940
rect 145 923 509 929
tri 509 923 526 940 nw
tri 564 938 566 940 se
rect 566 938 1001 940
tri 1001 938 1003 940 sw
tri 1056 938 1058 940 ne
rect 1058 938 1378 940
tri 549 923 564 938 se
rect 564 927 1003 938
tri 1003 927 1014 938 sw
tri 1058 927 1069 938 ne
rect 1069 927 1378 938
rect 564 923 1014 927
tri 1014 923 1018 927 sw
tri 1069 923 1073 927 ne
rect 1073 923 1378 927
tri 532 906 549 923 se
rect 549 906 598 923
tri 598 906 615 923 nw
tri 952 906 969 923 ne
rect 969 906 1018 923
tri 1018 906 1035 923 sw
tri 1073 906 1090 923 ne
rect 1090 906 1378 923
rect 1412 906 1450 940
rect 1484 906 1849 940
rect 1883 906 1921 940
rect 1955 906 1967 940
tri 529 903 532 906 se
rect 532 903 595 906
tri 595 903 598 906 nw
tri 969 903 972 906 ne
rect 972 903 1035 906
tri 519 893 529 903 se
rect 529 893 585 903
tri 585 893 595 903 nw
tri 972 893 982 903 ne
rect 982 900 1035 903
tri 1035 900 1041 906 sw
tri 1090 900 1096 906 ne
rect 1096 900 1967 906
tri 2068 900 2079 911 se
rect 2079 900 2125 1080
tri 2125 1056 2159 1090 nw
rect 982 893 1041 900
rect 297 881 573 893
tri 573 881 585 893 nw
rect 641 881 687 893
rect 297 847 303 881
rect 337 847 475 881
rect 509 872 564 881
tri 564 872 573 881 nw
rect 509 847 539 872
tri 539 847 564 872 nw
rect 641 847 647 881
rect 681 847 687 881
rect 297 809 515 847
tri 515 823 539 847 nw
rect 641 823 687 847
rect 813 881 859 893
rect 813 847 819 881
rect 853 847 859 881
tri 982 872 1003 893 ne
rect 1003 872 1041 893
tri 1041 872 1069 900 sw
tri 2040 872 2068 900 se
rect 2068 891 2125 900
rect 2068 872 2106 891
tri 2106 872 2125 891 nw
tri 687 823 709 845 sw
tri 791 823 813 845 se
rect 813 830 859 847
tri 1003 845 1030 872 ne
rect 1030 845 2064 872
tri 859 830 874 845 sw
tri 1030 830 1045 845 ne
rect 1045 830 2064 845
tri 2064 830 2106 872 nw
rect 813 823 874 830
tri 874 823 881 830 sw
rect 297 775 303 809
rect 337 775 475 809
rect 509 775 515 809
rect 297 763 515 775
rect 641 811 709 823
tri 709 811 721 823 sw
tri 779 811 791 823 se
rect 791 811 881 823
tri 881 811 893 823 sw
rect 641 809 1023 811
rect 641 775 647 809
rect 681 775 819 809
rect 853 801 1023 809
tri 1023 801 1033 811 sw
rect 853 795 2164 801
rect 853 775 1139 795
rect 641 763 1139 775
tri 1005 761 1007 763 ne
rect 1007 761 1139 763
rect 1173 761 1211 795
rect 1245 761 1614 795
rect 1648 761 1686 795
rect 1720 761 2046 795
rect 2080 761 2118 795
rect 2152 761 2164 795
tri 1007 755 1013 761 ne
rect 1013 755 2164 761
rect 150 723 945 735
rect 150 689 217 723
rect 251 689 389 723
rect 423 689 561 723
rect 595 689 733 723
rect 767 689 905 723
rect 939 689 945 723
rect 150 651 945 689
rect 150 617 217 651
rect 251 617 389 651
rect 423 617 561 651
rect 595 617 733 651
rect 767 617 905 651
rect 939 617 945 651
rect 150 605 945 617
rect 150 575 208 605
tri 208 575 238 605 nw
rect 150 570 203 575
tri 203 570 208 575 nw
rect 150 569 202 570
tri 202 569 203 570 nw
rect 267 569 550 575
rect 150 458 196 569
tri 196 563 202 569 nw
rect 267 535 290 569
rect 324 535 397 569
rect 431 535 504 569
rect 538 535 550 569
rect 267 529 550 535
rect 596 569 886 575
rect 596 535 622 569
rect 656 535 728 569
rect 762 535 834 569
rect 868 535 886 569
rect 596 529 886 535
rect 972 570 1546 576
rect 972 536 984 570
rect 1018 536 1056 570
rect 1090 564 1546 570
rect 1090 536 1506 564
rect 972 530 1506 536
rect 1540 530 1546 564
tri 1466 529 1467 530 ne
rect 1467 529 1546 530
tri 297 525 301 529 ne
rect 301 525 303 529
tri 1467 525 1471 529 ne
rect 1471 525 1546 529
tri 301 523 303 525 ne
tri 1471 523 1473 525 ne
rect 1473 523 1546 525
tri 1473 496 1500 523 ne
rect 1500 492 1546 523
tri 196 458 198 460 sw
rect 1500 458 1506 492
rect 1540 458 1546 492
rect 150 453 198 458
tri 198 453 203 458 sw
rect 150 444 203 453
tri 203 444 212 453 sw
rect 792 444 1240 450
rect 1500 446 1546 458
rect 1663 525 1709 537
rect 1663 491 1669 525
rect 1703 491 1709 525
rect 1663 453 1709 491
rect 150 440 212 444
tri 212 440 216 444 sw
tri 150 423 167 440 ne
rect 167 423 216 440
tri 99 410 112 423 sw
tri 167 410 180 423 ne
rect 180 410 216 423
tri 216 410 246 440 sw
rect 792 410 804 444
rect 838 410 882 444
rect 916 410 960 444
rect 994 410 1038 444
rect 1072 410 1116 444
rect 1150 410 1194 444
rect 1228 410 1240 444
rect 53 403 112 410
tri 53 373 83 403 ne
rect 83 374 112 403
tri 112 374 148 410 sw
tri 180 374 216 410 ne
rect 216 376 246 410
tri 246 376 280 410 sw
rect 792 404 1240 410
rect 1663 419 1669 453
rect 1703 419 1709 453
rect 1663 407 1709 419
rect 1936 535 1982 547
rect 1936 501 1942 535
rect 1976 501 1982 535
rect 1936 463 1982 501
rect 1936 429 1942 463
rect 1976 429 1982 463
tri 1416 376 1425 385 se
rect 1425 376 1471 385
rect 216 374 1245 376
rect 83 373 148 374
tri 148 373 149 374 sw
tri 216 373 217 374 ne
rect 217 373 1245 374
tri 1413 373 1416 376 se
rect 1416 373 1471 376
tri 83 370 86 373 ne
rect 86 370 149 373
tri 149 370 152 373 sw
tri 217 370 220 373 ne
rect 220 370 1245 373
tri 86 367 89 370 ne
rect 89 367 152 370
tri 152 367 155 370 sw
tri 220 367 223 370 ne
rect 223 367 828 370
tri 89 357 99 367 ne
rect 99 357 155 367
tri 99 336 120 357 ne
rect 120 336 155 357
tri 155 336 186 367 sw
tri 223 336 254 367 ne
rect 254 336 828 367
rect 862 336 900 370
rect 934 336 1127 370
rect 1161 336 1199 370
rect 1233 336 1245 370
tri 1379 339 1413 373 se
rect 1413 339 1431 373
rect 1465 339 1471 373
tri 1905 345 1936 376 se
rect 1936 356 1982 429
rect 1936 345 1971 356
tri 1971 345 1982 356 nw
rect 2061 376 2113 382
tri 120 305 151 336 ne
rect 151 330 186 336
tri 186 330 192 336 sw
tri 254 330 260 336 ne
rect 260 330 1245 336
tri 1370 330 1379 339 se
rect 1379 330 1471 339
rect 151 305 192 330
tri 192 305 217 330 sw
tri 1345 305 1370 330 se
rect 1370 305 1471 330
tri 151 301 155 305 ne
rect 155 301 217 305
tri 217 301 221 305 sw
tri 1341 301 1345 305 se
rect 1345 301 1471 305
tri 155 267 189 301 ne
rect 189 267 1431 301
rect 1465 267 1471 301
rect 1704 339 1956 345
rect 1704 305 1716 339
rect 1750 305 1788 339
rect 1822 330 1956 339
tri 1956 330 1971 345 nw
tri 2057 330 2061 334 se
rect 1822 305 1925 330
rect 1704 299 1925 305
tri 1925 299 1956 330 nw
tri 2054 327 2057 330 se
rect 2057 327 2061 330
tri 2027 300 2054 327 se
rect 2054 324 2061 327
rect 2054 312 2113 324
rect 2054 300 2061 312
tri 189 260 196 267 ne
rect 196 260 1471 267
tri 196 255 201 260 ne
rect 201 255 1471 260
rect 2010 294 2061 300
tri 2113 300 2140 327 sw
rect 2113 294 2140 300
rect 2010 260 2022 294
rect 2056 260 2061 294
rect 2128 260 2140 294
rect 2010 254 2140 260
rect 78 214 2203 226
rect 78 180 691 214
rect 725 180 1003 214
rect 1037 180 1315 214
rect 1349 180 1587 214
rect 1621 180 1866 214
rect 1900 180 2203 214
rect 78 142 2203 180
rect 78 108 691 142
rect 725 108 1003 142
rect 1037 108 1315 142
rect 1349 108 1587 142
rect 1621 108 1866 142
rect 1900 108 2203 142
rect 78 70 2203 108
rect 78 36 194 70
rect 228 36 266 70
rect 300 36 338 70
rect 372 36 410 70
rect 444 36 482 70
rect 516 36 554 70
rect 588 36 626 70
rect 660 36 698 70
rect 732 36 770 70
rect 804 36 842 70
rect 876 36 914 70
rect 948 36 986 70
rect 1020 36 1058 70
rect 1092 36 1131 70
rect 1165 36 1204 70
rect 1238 36 1277 70
rect 1311 36 1350 70
rect 1384 36 1423 70
rect 1457 36 1496 70
rect 1530 36 1569 70
rect 1603 36 1642 70
rect 1676 36 1715 70
rect 1749 36 1788 70
rect 1822 36 1861 70
rect 1895 36 1934 70
rect 1968 36 2007 70
rect 2041 36 2080 70
rect 2114 36 2203 70
rect 78 30 2203 36
<< via1 >>
rect 2061 1236 2113 1288
rect 2061 1172 2113 1224
rect 2061 324 2113 376
rect 2061 294 2113 312
rect 2061 260 2094 294
rect 2094 260 2113 294
<< metal2 >>
rect 2061 1288 2113 1294
rect 2061 1224 2113 1236
rect 2061 376 2113 1172
rect 2061 312 2113 324
rect 2061 254 2113 260
use sky130_fd_pr__nfet_01v8__example_55959141808463  sky130_fd_pr__nfet_01v8__example_55959141808463_0
timestamp 1644511149
transform 1 0 736 0 1 163
box -28 0 596 97
use sky130_fd_pr__nfet_01v8__example_55959141808464  sky130_fd_pr__nfet_01v8__example_55959141808464_0
timestamp 1644511149
transform -1 0 2110 0 -1 1288
box -28 0 916 97
use sky130_fd_pr__nfet_01v8__example_55959141808465  sky130_fd_pr__nfet_01v8__example_55959141808465_0
timestamp 1644511149
transform 1 0 1632 0 -1 363
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808465  sky130_fd_pr__nfet_01v8__example_55959141808465_1
timestamp 1644511149
transform -1 0 1576 0 -1 363
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808465  sky130_fd_pr__nfet_01v8__example_55959141808465_2
timestamp 1644511149
transform 1 0 1911 0 -1 363
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808466  sky130_fd_pr__nfet_01v8__example_55959141808466_0
timestamp 1644511149
transform -1 0 550 0 -1 817
box -28 0 316 97
use sky130_fd_pr__nfet_01v8__example_55959141808467  sky130_fd_pr__nfet_01v8__example_55959141808467_0
timestamp 1644511149
transform -1 0 894 0 -1 817
box -28 0 316 97
use sky130_fd_pr__nfet_01v8__example_55959141808468  sky130_fd_pr__nfet_01v8__example_55959141808468_0
timestamp 1644511149
transform -1 0 2110 0 1 758
box -28 0 916 97
use sky130_fd_pr__pfet_01v8__example_55959141808460  sky130_fd_pr__pfet_01v8__example_55959141808460_0
timestamp 1644511149
transform 1 0 863 0 -1 1297
box -28 0 128 63
use sky130_fd_pr__pfet_01v8__example_55959141808460  sky130_fd_pr__pfet_01v8__example_55959141808460_1
timestamp 1644511149
transform 1 0 597 0 -1 1297
box -28 0 128 63
use sky130_fd_pr__pfet_01v8__example_55959141808590  sky130_fd_pr__pfet_01v8__example_55959141808590_0
timestamp 1644511149
transform 1 0 331 0 -1 1297
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808590  sky130_fd_pr__pfet_01v8__example_55959141808590_1
timestamp 1644511149
transform -1 0 275 0 -1 1297
box -28 0 128 131
<< labels >>
flabel metal1 s 771 541 799 569 3 FreeSans 280 0 0 0 IN_B
port 1 nsew
flabel metal1 s 2070 263 2098 291 3 FreeSans 280 0 0 0 OUT_H_N
port 2 nsew
flabel metal1 s 1434 292 1462 320 3 FreeSans 280 0 0 0 OUT_H
port 3 nsew
flabel metal1 s 463 1341 491 1369 3 FreeSans 280 0 0 0 VPWR_HV
port 4 nsew
flabel metal1 s 1980 157 2008 185 3 FreeSans 280 0 0 0 VGND
port 5 nsew
flabel metal1 s 837 407 865 435 3 FreeSans 280 0 0 0 HLD_H_N
port 6 nsew
flabel metal1 s 1668 455 1696 483 3 FreeSans 280 0 0 0 RST_H
port 7 nsew
flabel metal1 s 422 540 450 568 3 FreeSans 280 0 0 0 IN
port 8 nsew
flabel metal1 s 1563 1010 1591 1038 3 FreeSans 280 0 0 0 VPWR_LV
port 9 nsew
<< properties >>
string GDS_END 8388348
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8358660
<< end >>
