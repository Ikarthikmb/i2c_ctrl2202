magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -66 377 1122 897
<< pwell >>
rect 772 283 1038 291
rect 4 43 1038 283
rect -26 -43 1082 43
<< mvnmos >>
rect 122 107 222 257
rect 264 107 364 257
rect 423 107 523 257
rect 581 107 681 257
rect 855 115 955 265
<< mvpmos >>
rect 122 443 222 743
rect 278 443 378 743
rect 439 443 539 743
rect 581 443 681 743
rect 850 443 950 743
<< mvndiff >>
rect 798 257 855 265
rect 30 245 122 257
rect 30 211 38 245
rect 72 211 122 245
rect 30 153 122 211
rect 30 119 38 153
rect 72 119 122 153
rect 30 107 122 119
rect 222 107 264 257
rect 364 179 423 257
rect 364 145 375 179
rect 409 145 423 179
rect 364 107 423 145
rect 523 249 581 257
rect 523 215 534 249
rect 568 215 581 249
rect 523 149 581 215
rect 523 115 534 149
rect 568 115 581 149
rect 523 107 581 115
rect 681 159 738 257
rect 681 125 692 159
rect 726 125 738 159
rect 681 107 738 125
rect 798 223 810 257
rect 844 223 855 257
rect 798 157 855 223
rect 798 123 810 157
rect 844 123 855 157
rect 798 115 855 123
rect 955 257 1012 265
rect 955 223 966 257
rect 1000 223 1012 257
rect 955 157 1012 223
rect 955 123 966 157
rect 1000 123 1012 157
rect 955 115 1012 123
<< mvpdiff >>
rect 65 735 122 743
rect 65 701 77 735
rect 111 701 122 735
rect 65 647 122 701
rect 65 613 77 647
rect 111 613 122 647
rect 65 560 122 613
rect 65 526 77 560
rect 111 526 122 560
rect 65 443 122 526
rect 222 735 278 743
rect 222 701 233 735
rect 267 701 278 735
rect 222 659 278 701
rect 222 625 233 659
rect 267 625 278 659
rect 222 582 278 625
rect 222 548 233 582
rect 267 548 278 582
rect 222 506 278 548
rect 222 472 233 506
rect 267 472 278 506
rect 222 443 278 472
rect 378 735 439 743
rect 378 701 389 735
rect 423 701 439 735
rect 378 655 439 701
rect 378 621 389 655
rect 423 621 439 655
rect 378 574 439 621
rect 378 540 389 574
rect 423 540 439 574
rect 378 494 439 540
rect 378 460 389 494
rect 423 460 439 494
rect 378 443 439 460
rect 539 443 581 743
rect 681 735 850 743
rect 681 701 805 735
rect 839 701 850 735
rect 681 652 850 701
rect 681 618 805 652
rect 839 618 850 652
rect 681 568 850 618
rect 681 534 805 568
rect 839 534 850 568
rect 681 485 850 534
rect 681 451 805 485
rect 839 451 850 485
rect 681 443 850 451
rect 950 735 1007 743
rect 950 701 961 735
rect 995 701 1007 735
rect 950 652 1007 701
rect 950 618 961 652
rect 995 618 1007 652
rect 950 568 1007 618
rect 950 534 961 568
rect 995 534 1007 568
rect 950 485 1007 534
rect 950 451 961 485
rect 995 451 1007 485
rect 950 443 1007 451
<< mvndiffc >>
rect 38 211 72 245
rect 38 119 72 153
rect 375 145 409 179
rect 534 215 568 249
rect 534 115 568 149
rect 692 125 726 159
rect 810 223 844 257
rect 810 123 844 157
rect 966 223 1000 257
rect 966 123 1000 157
<< mvpdiffc >>
rect 77 701 111 735
rect 77 613 111 647
rect 77 526 111 560
rect 233 701 267 735
rect 233 625 267 659
rect 233 548 267 582
rect 233 472 267 506
rect 389 701 423 735
rect 389 621 423 655
rect 389 540 423 574
rect 389 460 423 494
rect 805 701 839 735
rect 805 618 839 652
rect 805 534 839 568
rect 805 451 839 485
rect 961 701 995 735
rect 961 618 995 652
rect 961 534 995 568
rect 961 451 995 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
<< poly >>
rect 122 743 222 769
rect 278 743 378 769
rect 439 743 539 769
rect 581 743 681 769
rect 850 743 950 769
rect 122 417 222 443
rect 111 395 222 417
rect 111 361 131 395
rect 165 361 222 395
rect 278 383 378 443
rect 439 383 539 443
rect 111 283 222 361
rect 122 257 222 283
rect 264 350 539 383
rect 264 316 362 350
rect 396 316 539 350
rect 264 283 539 316
rect 581 395 681 443
rect 850 417 950 443
rect 581 361 601 395
rect 635 361 681 395
rect 264 257 364 283
rect 423 257 523 283
rect 581 257 681 361
rect 726 341 955 417
rect 726 307 746 341
rect 780 307 955 341
rect 726 287 955 307
rect 855 265 955 287
rect 122 81 222 107
rect 264 81 364 107
rect 423 81 523 107
rect 581 81 681 107
rect 855 89 955 115
<< polycont >>
rect 131 361 165 395
rect 362 316 396 350
rect 601 361 635 395
rect 746 307 780 341
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 18 735 197 751
rect 18 701 19 735
rect 53 701 77 735
rect 125 701 163 735
rect 18 647 197 701
rect 18 613 77 647
rect 111 613 197 647
rect 18 560 197 613
rect 18 526 77 560
rect 111 526 197 560
rect 233 735 267 751
rect 233 659 267 701
rect 233 582 267 625
rect 233 506 267 548
rect 22 472 233 490
rect 22 456 267 472
rect 303 735 769 751
rect 337 701 375 735
rect 423 701 447 735
rect 481 701 519 735
rect 553 701 591 735
rect 625 701 663 735
rect 697 701 735 735
rect 303 655 769 701
rect 303 621 389 655
rect 423 621 769 655
rect 303 574 769 621
rect 303 540 389 574
rect 423 540 769 574
rect 303 494 769 540
rect 303 460 389 494
rect 423 460 769 494
rect 805 735 855 751
rect 839 701 855 735
rect 805 652 855 701
rect 839 618 855 652
rect 805 568 855 618
rect 839 534 855 568
rect 805 485 855 534
rect 22 280 72 456
rect 839 451 855 485
rect 893 735 1011 751
rect 893 701 899 735
rect 933 701 961 735
rect 1005 701 1011 735
rect 893 652 1011 701
rect 893 618 961 652
rect 995 618 1011 652
rect 893 568 1011 618
rect 893 534 961 568
rect 995 534 1011 568
rect 893 485 1011 534
rect 893 451 961 485
rect 995 451 1011 485
rect 313 420 651 424
rect 115 395 651 420
rect 115 361 131 395
rect 165 386 601 395
rect 165 361 181 386
rect 585 361 601 386
rect 635 361 651 395
rect 805 415 855 451
rect 805 381 1031 415
rect 115 345 181 361
rect 217 316 362 350
rect 396 316 412 350
rect 730 341 796 345
rect 730 325 746 341
rect 448 307 746 325
rect 780 307 796 341
rect 889 309 1031 381
rect 448 291 796 307
rect 448 280 482 291
rect 22 246 482 280
rect 950 257 1031 309
rect 518 249 810 257
rect 22 245 88 246
rect 22 211 38 245
rect 72 211 88 245
rect 22 153 88 211
rect 518 215 534 249
rect 568 223 810 249
rect 844 223 860 257
rect 568 221 860 223
rect 568 215 584 221
rect 22 119 38 153
rect 72 119 88 153
rect 22 99 88 119
rect 122 179 482 210
rect 122 145 375 179
rect 409 145 482 179
rect 122 113 482 145
rect 122 79 160 113
rect 194 79 232 113
rect 266 79 304 113
rect 338 79 376 113
rect 410 79 448 113
rect 518 149 584 215
rect 518 115 534 149
rect 568 115 584 149
rect 518 99 584 115
rect 620 159 726 185
rect 620 125 692 159
rect 620 113 726 125
rect 122 73 482 79
rect 654 79 692 113
rect 794 157 860 221
rect 794 123 810 157
rect 844 123 860 157
rect 794 107 860 123
rect 950 223 966 257
rect 1000 223 1031 257
rect 950 157 1031 223
rect 950 123 966 157
rect 1000 123 1031 157
rect 950 107 1031 123
rect 620 73 726 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 19 701 53 735
rect 91 701 111 735
rect 111 701 125 735
rect 163 701 197 735
rect 303 701 337 735
rect 375 701 389 735
rect 389 701 409 735
rect 447 701 481 735
rect 519 701 553 735
rect 591 701 625 735
rect 663 701 697 735
rect 735 701 769 735
rect 899 701 933 735
rect 971 701 995 735
rect 995 701 1005 735
rect 160 79 194 113
rect 232 79 266 113
rect 304 79 338 113
rect 376 79 410 113
rect 448 79 482 113
rect 620 79 654 113
rect 692 79 726 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 831 1056 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 0 791 1056 797
rect 0 735 1056 763
rect 0 701 19 735
rect 53 701 91 735
rect 125 701 163 735
rect 197 701 303 735
rect 337 701 375 735
rect 409 701 447 735
rect 481 701 519 735
rect 553 701 591 735
rect 625 701 663 735
rect 697 701 735 735
rect 769 701 899 735
rect 933 701 971 735
rect 1005 701 1056 735
rect 0 689 1056 701
rect 0 113 1056 125
rect 0 79 160 113
rect 194 79 232 113
rect 266 79 304 113
rect 338 79 376 113
rect 410 79 448 113
rect 482 79 620 113
rect 654 79 692 113
rect 726 79 1056 113
rect 0 51 1056 79
rect 0 17 1056 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -23 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xnor2_1
flabel metal1 s 0 51 1056 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 1056 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 1056 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 1056 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 390 353 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
flabel locali s 895 316 929 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 991 316 1025 350 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
flabel locali s 991 242 1025 276 0 FreeSans 340 0 0 0 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1056 814
string GDS_END 731298
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 719110
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
