magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect 30 43 764 283
rect -26 -43 794 43
<< mvnmos >>
rect 113 107 213 257
rect 269 107 369 257
rect 425 107 525 257
rect 581 107 681 257
<< mvpmos >>
rect 113 443 213 743
rect 269 443 369 743
rect 425 443 525 743
rect 581 443 681 743
<< mvndiff >>
rect 56 249 113 257
rect 56 215 68 249
rect 102 215 113 249
rect 56 149 113 215
rect 56 115 68 149
rect 102 115 113 149
rect 56 107 113 115
rect 213 249 269 257
rect 213 215 224 249
rect 258 215 269 249
rect 213 149 269 215
rect 213 115 224 149
rect 258 115 269 149
rect 213 107 269 115
rect 369 179 425 257
rect 369 145 380 179
rect 414 145 425 179
rect 369 107 425 145
rect 525 249 581 257
rect 525 215 536 249
rect 570 215 581 249
rect 525 149 581 215
rect 525 115 536 149
rect 570 115 581 149
rect 525 107 581 115
rect 681 249 738 257
rect 681 215 692 249
rect 726 215 738 249
rect 681 149 738 215
rect 681 115 692 149
rect 726 115 738 149
rect 681 107 738 115
<< mvpdiff >>
rect 56 735 113 743
rect 56 701 68 735
rect 102 701 113 735
rect 56 652 113 701
rect 56 618 68 652
rect 102 618 113 652
rect 56 568 113 618
rect 56 534 68 568
rect 102 534 113 568
rect 56 485 113 534
rect 56 451 68 485
rect 102 451 113 485
rect 56 443 113 451
rect 213 735 269 743
rect 213 701 224 735
rect 258 701 269 735
rect 213 652 269 701
rect 213 618 224 652
rect 258 618 269 652
rect 213 568 269 618
rect 213 534 224 568
rect 258 534 269 568
rect 213 485 269 534
rect 213 451 224 485
rect 258 451 269 485
rect 213 443 269 451
rect 369 735 425 743
rect 369 701 380 735
rect 414 701 425 735
rect 369 654 425 701
rect 369 620 380 654
rect 414 620 425 654
rect 369 571 425 620
rect 369 537 380 571
rect 414 537 425 571
rect 369 490 425 537
rect 369 456 380 490
rect 414 456 425 490
rect 369 443 425 456
rect 525 735 581 743
rect 525 701 536 735
rect 570 701 581 735
rect 525 652 581 701
rect 525 618 536 652
rect 570 618 581 652
rect 525 568 581 618
rect 525 534 536 568
rect 570 534 581 568
rect 525 485 581 534
rect 525 451 536 485
rect 570 451 581 485
rect 525 443 581 451
rect 681 735 738 743
rect 681 701 692 735
rect 726 701 738 735
rect 681 654 738 701
rect 681 620 692 654
rect 726 620 738 654
rect 681 571 738 620
rect 681 537 692 571
rect 726 537 738 571
rect 681 490 738 537
rect 681 456 692 490
rect 726 456 738 490
rect 681 443 738 456
<< mvndiffc >>
rect 68 215 102 249
rect 68 115 102 149
rect 224 215 258 249
rect 224 115 258 149
rect 380 145 414 179
rect 536 215 570 249
rect 536 115 570 149
rect 692 215 726 249
rect 692 115 726 149
<< mvpdiffc >>
rect 68 701 102 735
rect 68 618 102 652
rect 68 534 102 568
rect 68 451 102 485
rect 224 701 258 735
rect 224 618 258 652
rect 224 534 258 568
rect 224 451 258 485
rect 380 701 414 735
rect 380 620 414 654
rect 380 537 414 571
rect 380 456 414 490
rect 536 701 570 735
rect 536 618 570 652
rect 536 534 570 568
rect 536 451 570 485
rect 692 701 726 735
rect 692 620 726 654
rect 692 537 726 571
rect 692 456 726 490
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
<< poly >>
rect 113 743 213 769
rect 269 743 369 769
rect 425 743 525 769
rect 581 743 681 769
rect 113 417 213 443
rect 269 417 369 443
rect 425 417 525 443
rect 581 417 681 443
rect 113 374 681 417
rect 21 350 681 374
rect 21 316 41 350
rect 75 316 109 350
rect 143 316 177 350
rect 211 316 245 350
rect 279 316 313 350
rect 347 316 381 350
rect 415 316 449 350
rect 483 316 517 350
rect 551 316 681 350
rect 21 283 681 316
rect 113 257 213 283
rect 269 257 369 283
rect 425 257 525 283
rect 581 257 681 283
rect 113 81 213 107
rect 269 81 369 107
rect 425 81 525 107
rect 581 81 681 107
<< polycont >>
rect 41 316 75 350
rect 109 316 143 350
rect 177 316 211 350
rect 245 316 279 350
rect 313 316 347 350
rect 381 316 415 350
rect 449 316 483 350
rect 517 316 551 350
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 18 735 136 751
rect 18 701 24 735
rect 58 701 68 735
rect 130 701 136 735
rect 18 652 136 701
rect 18 618 68 652
rect 102 618 136 652
rect 18 568 136 618
rect 18 534 68 568
rect 102 534 136 568
rect 18 485 136 534
rect 18 451 68 485
rect 102 451 136 485
rect 18 435 136 451
rect 208 735 274 751
rect 208 701 224 735
rect 258 701 274 735
rect 208 652 274 701
rect 208 618 224 652
rect 258 618 274 652
rect 208 568 274 618
rect 208 534 224 568
rect 258 534 274 568
rect 208 485 274 534
rect 208 451 224 485
rect 258 451 274 485
rect 310 735 500 751
rect 310 701 316 735
rect 350 701 380 735
rect 422 701 460 735
rect 494 701 500 735
rect 310 654 500 701
rect 310 620 380 654
rect 414 620 500 654
rect 310 571 500 620
rect 310 537 380 571
rect 414 537 500 571
rect 310 490 500 537
rect 310 456 380 490
rect 414 456 500 490
rect 536 735 586 751
rect 570 701 586 735
rect 536 652 586 701
rect 570 618 586 652
rect 536 568 586 618
rect 570 534 586 568
rect 536 485 586 534
rect 208 420 274 451
rect 570 451 586 485
rect 624 735 742 751
rect 624 701 630 735
rect 664 701 692 735
rect 736 701 742 735
rect 624 654 742 701
rect 624 620 692 654
rect 726 620 742 654
rect 624 571 742 620
rect 624 537 692 571
rect 726 537 742 571
rect 624 490 742 537
rect 624 456 692 490
rect 726 456 742 490
rect 536 420 586 451
rect 208 386 743 420
rect 25 316 41 350
rect 75 316 109 350
rect 143 316 177 350
rect 211 316 245 350
rect 279 316 313 350
rect 347 316 381 350
rect 415 316 449 350
rect 483 316 517 350
rect 551 316 567 350
rect 603 310 743 386
rect 603 280 637 310
rect 18 249 136 265
rect 18 215 68 249
rect 102 215 136 249
rect 18 149 136 215
rect 18 115 68 149
rect 102 115 136 149
rect 18 113 136 115
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 136 113
rect 208 249 637 280
rect 208 215 224 249
rect 258 246 536 249
rect 208 149 258 215
rect 520 215 536 246
rect 570 215 637 249
rect 208 115 224 149
rect 208 99 258 115
rect 294 179 484 210
rect 294 145 380 179
rect 414 145 484 179
rect 294 113 484 145
rect 18 73 136 79
rect 294 79 300 113
rect 334 79 372 113
rect 406 79 444 113
rect 478 79 484 113
rect 520 149 637 215
rect 520 115 536 149
rect 570 115 637 149
rect 520 99 637 115
rect 676 249 742 265
rect 676 215 692 249
rect 726 215 742 249
rect 676 149 742 215
rect 676 115 692 149
rect 726 115 742 149
rect 676 113 742 115
rect 294 73 484 79
rect 676 79 682 113
rect 716 79 742 113
rect 676 73 742 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 24 701 58 735
rect 96 701 102 735
rect 102 701 130 735
rect 316 701 350 735
rect 388 701 414 735
rect 414 701 422 735
rect 460 701 494 735
rect 630 701 664 735
rect 702 701 726 735
rect 726 701 736 735
rect 24 79 58 113
rect 96 79 130 113
rect 300 79 334 113
rect 372 79 406 113
rect 444 79 478 113
rect 682 79 716 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 735 768 763
rect 0 701 24 735
rect 58 701 96 735
rect 130 701 316 735
rect 350 701 388 735
rect 422 701 460 735
rect 494 701 630 735
rect 664 701 702 735
rect 736 701 768 735
rect 0 689 768 701
rect 0 113 768 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 300 113
rect 334 79 372 113
rect 406 79 444 113
rect 478 79 682 113
rect 716 79 768 113
rect 0 51 768 79
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel comment s 0 0 0 0 4 inv_4
flabel metal1 s 0 51 768 125 0 FreeSans 340 0 0 0 VGND
port 2 nsew ground bidirectional
flabel metal1 s 0 0 768 23 0 FreeSans 340 0 0 0 VNB
port 3 nsew ground bidirectional
flabel metal1 s 0 689 768 763 0 FreeSans 340 0 0 0 VPWR
port 5 nsew power bidirectional
flabel metal1 s 0 791 768 814 0 FreeSans 340 0 0 0 VPB
port 4 nsew power bidirectional
flabel locali s 607 316 641 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 Y
port 6 nsew signal output
flabel locali s 31 316 65 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 127 316 161 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 223 316 257 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 319 316 353 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 415 316 449 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 316 545 350 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 768 814
string GDS_END 69816
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 59660
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
