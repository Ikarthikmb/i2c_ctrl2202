magic
tech sky130A
timestamp 1644511149
<< properties >>
string GDS_END 30669790
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30669338
<< end >>
