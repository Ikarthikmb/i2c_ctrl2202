/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/rf_aura_blocking/sky130_fd_pr__rf_aura_blocking.spice