magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1423 203
rect 30 -17 64 21
<< locali >>
rect 291 333 357 493
rect 459 401 525 493
rect 627 401 693 493
rect 459 333 693 401
rect 795 333 861 493
rect 1067 333 1133 493
rect 1235 333 1301 493
rect 291 289 1301 333
rect 86 215 156 255
rect 559 215 620 289
rect 654 215 896 255
rect 958 215 1300 255
rect 559 181 593 215
rect 291 127 593 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 17 289 85 493
rect 119 289 257 527
rect 391 367 425 527
rect 559 435 593 527
rect 727 367 761 527
rect 895 367 1033 527
rect 1167 367 1201 527
rect 1335 289 1401 527
rect 17 181 52 289
rect 201 215 525 255
rect 201 181 257 215
rect 17 143 257 181
rect 17 51 85 143
rect 627 143 1301 181
rect 627 127 945 143
rect 119 17 169 109
rect 207 51 945 93
rect 983 17 1033 109
rect 1067 51 1133 143
rect 1167 17 1201 109
rect 1235 51 1301 143
rect 1335 17 1401 181
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
rlabel locali s 86 215 156 255 6 A_N
port 1 nsew signal input
rlabel locali s 654 215 896 255 6 B
port 2 nsew signal input
rlabel locali s 958 215 1300 255 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 1472 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1423 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1510 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1472 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 291 127 593 181 6 Y
port 8 nsew signal output
rlabel locali s 559 181 593 215 6 Y
port 8 nsew signal output
rlabel locali s 559 215 620 289 6 Y
port 8 nsew signal output
rlabel locali s 291 289 1301 333 6 Y
port 8 nsew signal output
rlabel locali s 1235 333 1301 493 6 Y
port 8 nsew signal output
rlabel locali s 1067 333 1133 493 6 Y
port 8 nsew signal output
rlabel locali s 795 333 861 493 6 Y
port 8 nsew signal output
rlabel locali s 459 333 693 401 6 Y
port 8 nsew signal output
rlabel locali s 627 401 693 493 6 Y
port 8 nsew signal output
rlabel locali s 459 401 525 493 6 Y
port 8 nsew signal output
rlabel locali s 291 333 357 493 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1472 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1876968
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1865182
<< end >>
