/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/res_generic_pd/sky130_fd_pr__res_generic_pd.model.spice