magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< dnwell >>
rect 80 80 2376 2305
<< nwell >>
rect 0 2099 2456 2385
rect 0 286 286 2099
rect 1381 1652 2456 2099
rect 1420 1144 2456 1652
rect 1738 286 2456 1144
rect 0 0 2456 286
<< pwell >>
rect 353 1706 439 1716
rect 353 1451 1119 1706
rect 353 1084 1342 1451
rect 353 402 1616 1084
rect 353 392 439 402
rect 1256 392 1342 402
<< mvnmos >>
rect 493 1527 1093 1627
rect 493 1261 1093 1361
rect 493 1105 1093 1205
rect 493 949 1093 1049
rect 1390 905 1590 1005
rect 493 793 1093 893
rect 493 637 1093 737
rect 493 481 1093 581
rect 1390 637 1590 737
rect 1390 481 1590 581
<< mvpmos >>
rect 1486 1263 1570 1463
rect 1929 1263 2013 1463
rect 1804 637 2104 737
rect 1804 481 2104 581
<< mvndiff >>
rect 493 1672 1093 1680
rect 493 1638 571 1672
rect 605 1638 639 1672
rect 673 1638 707 1672
rect 741 1638 775 1672
rect 809 1638 843 1672
rect 877 1638 911 1672
rect 945 1638 979 1672
rect 1013 1638 1047 1672
rect 1081 1638 1093 1672
rect 493 1627 1093 1638
rect 493 1516 1093 1527
rect 493 1482 571 1516
rect 605 1482 639 1516
rect 673 1482 707 1516
rect 741 1482 775 1516
rect 809 1482 843 1516
rect 877 1482 911 1516
rect 945 1482 979 1516
rect 1013 1482 1047 1516
rect 1081 1482 1093 1516
rect 493 1474 1093 1482
rect 493 1406 1093 1414
rect 493 1372 571 1406
rect 605 1372 639 1406
rect 673 1372 707 1406
rect 741 1372 775 1406
rect 809 1372 843 1406
rect 877 1372 911 1406
rect 945 1372 979 1406
rect 1013 1372 1047 1406
rect 1081 1372 1093 1406
rect 493 1361 1093 1372
rect 493 1250 1093 1261
rect 493 1216 571 1250
rect 605 1216 639 1250
rect 673 1216 707 1250
rect 741 1216 775 1250
rect 809 1216 843 1250
rect 877 1216 911 1250
rect 945 1216 979 1250
rect 1013 1216 1047 1250
rect 1081 1216 1093 1250
rect 493 1205 1093 1216
rect 493 1094 1093 1105
rect 493 1060 571 1094
rect 605 1060 639 1094
rect 673 1060 707 1094
rect 741 1060 775 1094
rect 809 1060 843 1094
rect 877 1060 911 1094
rect 945 1060 979 1094
rect 1013 1060 1047 1094
rect 1081 1060 1093 1094
rect 493 1049 1093 1060
rect 1390 1050 1590 1058
rect 1390 1016 1402 1050
rect 1436 1016 1470 1050
rect 1504 1016 1538 1050
rect 1572 1016 1590 1050
rect 1390 1005 1590 1016
rect 493 938 1093 949
rect 493 904 571 938
rect 605 904 639 938
rect 673 904 707 938
rect 741 904 775 938
rect 809 904 843 938
rect 877 904 911 938
rect 945 904 979 938
rect 1013 904 1047 938
rect 1081 904 1093 938
rect 493 893 1093 904
rect 493 782 1093 793
rect 493 748 571 782
rect 605 748 639 782
rect 673 748 707 782
rect 741 748 775 782
rect 809 748 843 782
rect 877 748 911 782
rect 945 748 979 782
rect 1013 748 1047 782
rect 1081 748 1093 782
rect 493 737 1093 748
rect 493 626 1093 637
rect 493 592 571 626
rect 605 592 639 626
rect 673 592 707 626
rect 741 592 775 626
rect 809 592 843 626
rect 877 592 911 626
rect 945 592 979 626
rect 1013 592 1047 626
rect 1081 592 1093 626
rect 493 581 1093 592
rect 1390 894 1590 905
rect 1390 860 1402 894
rect 1436 860 1470 894
rect 1504 860 1538 894
rect 1572 860 1590 894
rect 1390 852 1590 860
rect 1390 782 1590 790
rect 1390 748 1402 782
rect 1436 748 1470 782
rect 1504 748 1538 782
rect 1572 748 1590 782
rect 1390 737 1590 748
rect 1390 626 1590 637
rect 1390 592 1402 626
rect 1436 592 1470 626
rect 1504 592 1538 626
rect 1572 592 1590 626
rect 1390 581 1590 592
rect 493 470 1093 481
rect 493 436 571 470
rect 605 436 639 470
rect 673 436 707 470
rect 741 436 775 470
rect 809 436 843 470
rect 877 436 911 470
rect 945 436 979 470
rect 1013 436 1047 470
rect 1081 436 1093 470
rect 493 428 1093 436
rect 1390 470 1590 481
rect 1390 436 1402 470
rect 1436 436 1470 470
rect 1504 436 1538 470
rect 1572 436 1590 470
rect 1390 428 1590 436
<< mvpdiff >>
rect 1486 1508 1570 1516
rect 1486 1474 1498 1508
rect 1532 1474 1570 1508
rect 1486 1463 1570 1474
rect 1929 1508 2013 1516
rect 1929 1474 1967 1508
rect 2001 1474 2013 1508
rect 1929 1463 2013 1474
rect 1486 1252 1570 1263
rect 1486 1218 1498 1252
rect 1532 1218 1570 1252
rect 1486 1210 1570 1218
rect 1929 1252 2013 1263
rect 1929 1218 1967 1252
rect 2001 1218 2013 1252
rect 1929 1210 2013 1218
rect 1804 782 2104 790
rect 1804 748 1854 782
rect 1888 748 1922 782
rect 1956 748 1990 782
rect 2024 748 2058 782
rect 2092 748 2104 782
rect 1804 737 2104 748
rect 1804 626 2104 637
rect 1804 592 1854 626
rect 1888 592 1922 626
rect 1956 592 1990 626
rect 2024 592 2058 626
rect 2092 592 2104 626
rect 1804 581 2104 592
rect 1804 470 2104 481
rect 1804 436 1854 470
rect 1888 436 1922 470
rect 1956 436 1990 470
rect 2024 436 2058 470
rect 2092 436 2104 470
rect 1804 428 2104 436
<< mvndiffc >>
rect 571 1638 605 1672
rect 639 1638 673 1672
rect 707 1638 741 1672
rect 775 1638 809 1672
rect 843 1638 877 1672
rect 911 1638 945 1672
rect 979 1638 1013 1672
rect 1047 1638 1081 1672
rect 571 1482 605 1516
rect 639 1482 673 1516
rect 707 1482 741 1516
rect 775 1482 809 1516
rect 843 1482 877 1516
rect 911 1482 945 1516
rect 979 1482 1013 1516
rect 1047 1482 1081 1516
rect 571 1372 605 1406
rect 639 1372 673 1406
rect 707 1372 741 1406
rect 775 1372 809 1406
rect 843 1372 877 1406
rect 911 1372 945 1406
rect 979 1372 1013 1406
rect 1047 1372 1081 1406
rect 571 1216 605 1250
rect 639 1216 673 1250
rect 707 1216 741 1250
rect 775 1216 809 1250
rect 843 1216 877 1250
rect 911 1216 945 1250
rect 979 1216 1013 1250
rect 1047 1216 1081 1250
rect 571 1060 605 1094
rect 639 1060 673 1094
rect 707 1060 741 1094
rect 775 1060 809 1094
rect 843 1060 877 1094
rect 911 1060 945 1094
rect 979 1060 1013 1094
rect 1047 1060 1081 1094
rect 1402 1016 1436 1050
rect 1470 1016 1504 1050
rect 1538 1016 1572 1050
rect 571 904 605 938
rect 639 904 673 938
rect 707 904 741 938
rect 775 904 809 938
rect 843 904 877 938
rect 911 904 945 938
rect 979 904 1013 938
rect 1047 904 1081 938
rect 571 748 605 782
rect 639 748 673 782
rect 707 748 741 782
rect 775 748 809 782
rect 843 748 877 782
rect 911 748 945 782
rect 979 748 1013 782
rect 1047 748 1081 782
rect 571 592 605 626
rect 639 592 673 626
rect 707 592 741 626
rect 775 592 809 626
rect 843 592 877 626
rect 911 592 945 626
rect 979 592 1013 626
rect 1047 592 1081 626
rect 1402 860 1436 894
rect 1470 860 1504 894
rect 1538 860 1572 894
rect 1402 748 1436 782
rect 1470 748 1504 782
rect 1538 748 1572 782
rect 1402 592 1436 626
rect 1470 592 1504 626
rect 1538 592 1572 626
rect 571 436 605 470
rect 639 436 673 470
rect 707 436 741 470
rect 775 436 809 470
rect 843 436 877 470
rect 911 436 945 470
rect 979 436 1013 470
rect 1047 436 1081 470
rect 1402 436 1436 470
rect 1470 436 1504 470
rect 1538 436 1572 470
<< mvpdiffc >>
rect 1498 1474 1532 1508
rect 1967 1474 2001 1508
rect 1498 1218 1532 1252
rect 1967 1218 2001 1252
rect 1854 748 1888 782
rect 1922 748 1956 782
rect 1990 748 2024 782
rect 2058 748 2092 782
rect 1854 592 1888 626
rect 1922 592 1956 626
rect 1990 592 2024 626
rect 2058 592 2092 626
rect 1854 436 1888 470
rect 1922 436 1956 470
rect 1990 436 2024 470
rect 2058 436 2092 470
<< mvpsubdiff >>
rect 379 1666 413 1690
rect 379 1596 413 1632
rect 379 1526 413 1562
rect 379 1456 413 1492
rect 379 1386 413 1422
rect 1282 1401 1316 1425
rect 379 1316 413 1352
rect 379 1246 413 1282
rect 379 1176 413 1212
rect 379 1106 413 1142
rect 379 1036 413 1072
rect 379 966 413 1002
rect 1282 1329 1316 1367
rect 1282 1257 1316 1295
rect 1282 1186 1316 1223
rect 1282 1115 1316 1152
rect 1282 1044 1316 1081
rect 1282 973 1316 1010
rect 379 896 413 932
rect 1282 902 1316 939
rect 379 826 413 862
rect 379 756 413 792
rect 379 686 413 722
rect 379 616 413 652
rect 379 546 413 582
rect 379 476 413 512
rect 1282 831 1316 868
rect 1282 760 1316 797
rect 1282 689 1316 726
rect 1282 618 1316 655
rect 1282 547 1316 584
rect 379 418 413 442
rect 1282 476 1316 513
rect 1282 418 1316 442
<< mvnsubdiff >>
rect 126 2225 194 2259
rect 228 2225 262 2259
rect 296 2225 330 2259
rect 364 2225 398 2259
rect 432 2225 466 2259
rect 500 2225 534 2259
rect 568 2225 602 2259
rect 636 2225 670 2259
rect 704 2225 738 2259
rect 772 2225 806 2259
rect 840 2225 874 2259
rect 908 2225 942 2259
rect 976 2225 1010 2259
rect 1044 2225 1078 2259
rect 1112 2225 1146 2259
rect 1180 2225 1214 2259
rect 1248 2225 1282 2259
rect 1316 2225 1350 2259
rect 1384 2225 1418 2259
rect 1452 2225 1486 2259
rect 1520 2225 1554 2259
rect 1588 2225 1622 2259
rect 1656 2225 1690 2259
rect 1724 2225 1758 2259
rect 1792 2225 1826 2259
rect 1860 2225 1894 2259
rect 1928 2225 1962 2259
rect 1996 2225 2030 2259
rect 2064 2225 2098 2259
rect 2132 2225 2166 2259
rect 2200 2225 2330 2259
rect 126 2167 160 2225
rect 126 2064 160 2133
rect 126 1996 160 2030
rect 126 1928 160 1962
rect 126 1860 160 1894
rect 126 1792 160 1826
rect 126 1724 160 1758
rect 2296 2191 2330 2225
rect 2296 2123 2330 2157
rect 2296 2055 2330 2089
rect 2296 1987 2330 2021
rect 2296 1919 2330 1953
rect 2296 1851 2330 1885
rect 2296 1783 2330 1817
rect 2296 1715 2330 1749
rect 126 1656 160 1690
rect 126 1588 160 1622
rect 126 1520 160 1554
rect 126 1452 160 1486
rect 126 1384 160 1418
rect 126 1316 160 1350
rect 126 1248 160 1282
rect 126 1180 160 1214
rect 126 1112 160 1146
rect 126 1044 160 1078
rect 126 976 160 1010
rect 126 908 160 942
rect 126 840 160 874
rect 126 772 160 806
rect 126 704 160 738
rect 126 636 160 670
rect 126 568 160 602
rect 126 500 160 534
rect 126 432 160 466
rect 2296 1647 2330 1681
rect 2296 1579 2330 1613
rect 2296 1511 2330 1545
rect 2296 1443 2330 1477
rect 2296 1375 2330 1409
rect 2296 1307 2330 1341
rect 2296 1239 2330 1273
rect 2296 1171 2330 1205
rect 2296 1103 2330 1137
rect 2296 1035 2330 1069
rect 2296 967 2330 1001
rect 2296 899 2330 933
rect 2296 831 2330 865
rect 2296 763 2330 797
rect 2296 695 2330 729
rect 2296 627 2330 661
rect 2296 559 2330 593
rect 2296 491 2330 525
rect 2296 423 2330 457
rect 126 364 160 398
rect 126 296 160 330
rect 126 228 160 262
rect 126 160 160 194
rect 2296 355 2330 389
rect 2296 287 2330 321
rect 2296 160 2330 253
rect 126 126 256 160
rect 290 126 324 160
rect 358 126 392 160
rect 426 126 460 160
rect 494 126 528 160
rect 562 126 596 160
rect 630 126 664 160
rect 698 126 732 160
rect 766 126 800 160
rect 834 126 868 160
rect 902 126 936 160
rect 970 126 1004 160
rect 1038 126 1072 160
rect 1106 126 1140 160
rect 1174 126 1208 160
rect 1242 126 1276 160
rect 1310 126 1344 160
rect 1378 126 1412 160
rect 1446 126 1480 160
rect 1514 126 1548 160
rect 1582 126 1616 160
rect 1650 126 1684 160
rect 1718 126 1752 160
rect 1786 126 1820 160
rect 1854 126 1888 160
rect 1922 126 1956 160
rect 1990 126 2024 160
rect 2058 126 2092 160
rect 2126 126 2160 160
rect 2194 126 2228 160
rect 2262 126 2330 160
<< mvpsubdiffcont >>
rect 379 1632 413 1666
rect 379 1562 413 1596
rect 379 1492 413 1526
rect 379 1422 413 1456
rect 379 1352 413 1386
rect 1282 1367 1316 1401
rect 379 1282 413 1316
rect 379 1212 413 1246
rect 379 1142 413 1176
rect 379 1072 413 1106
rect 379 1002 413 1036
rect 379 932 413 966
rect 1282 1295 1316 1329
rect 1282 1223 1316 1257
rect 1282 1152 1316 1186
rect 1282 1081 1316 1115
rect 1282 1010 1316 1044
rect 379 862 413 896
rect 1282 939 1316 973
rect 379 792 413 826
rect 379 722 413 756
rect 379 652 413 686
rect 379 582 413 616
rect 379 512 413 546
rect 1282 868 1316 902
rect 1282 797 1316 831
rect 1282 726 1316 760
rect 1282 655 1316 689
rect 1282 584 1316 618
rect 1282 513 1316 547
rect 379 442 413 476
rect 1282 442 1316 476
<< mvnsubdiffcont >>
rect 194 2225 228 2259
rect 262 2225 296 2259
rect 330 2225 364 2259
rect 398 2225 432 2259
rect 466 2225 500 2259
rect 534 2225 568 2259
rect 602 2225 636 2259
rect 670 2225 704 2259
rect 738 2225 772 2259
rect 806 2225 840 2259
rect 874 2225 908 2259
rect 942 2225 976 2259
rect 1010 2225 1044 2259
rect 1078 2225 1112 2259
rect 1146 2225 1180 2259
rect 1214 2225 1248 2259
rect 1282 2225 1316 2259
rect 1350 2225 1384 2259
rect 1418 2225 1452 2259
rect 1486 2225 1520 2259
rect 1554 2225 1588 2259
rect 1622 2225 1656 2259
rect 1690 2225 1724 2259
rect 1758 2225 1792 2259
rect 1826 2225 1860 2259
rect 1894 2225 1928 2259
rect 1962 2225 1996 2259
rect 2030 2225 2064 2259
rect 2098 2225 2132 2259
rect 2166 2225 2200 2259
rect 126 2133 160 2167
rect 126 2030 160 2064
rect 126 1962 160 1996
rect 126 1894 160 1928
rect 126 1826 160 1860
rect 126 1758 160 1792
rect 126 1690 160 1724
rect 2296 2157 2330 2191
rect 2296 2089 2330 2123
rect 2296 2021 2330 2055
rect 2296 1953 2330 1987
rect 2296 1885 2330 1919
rect 2296 1817 2330 1851
rect 2296 1749 2330 1783
rect 126 1622 160 1656
rect 126 1554 160 1588
rect 126 1486 160 1520
rect 126 1418 160 1452
rect 126 1350 160 1384
rect 126 1282 160 1316
rect 126 1214 160 1248
rect 126 1146 160 1180
rect 126 1078 160 1112
rect 126 1010 160 1044
rect 126 942 160 976
rect 126 874 160 908
rect 126 806 160 840
rect 126 738 160 772
rect 126 670 160 704
rect 126 602 160 636
rect 126 534 160 568
rect 126 466 160 500
rect 126 398 160 432
rect 2296 1681 2330 1715
rect 2296 1613 2330 1647
rect 2296 1545 2330 1579
rect 2296 1477 2330 1511
rect 2296 1409 2330 1443
rect 2296 1341 2330 1375
rect 2296 1273 2330 1307
rect 2296 1205 2330 1239
rect 2296 1137 2330 1171
rect 2296 1069 2330 1103
rect 2296 1001 2330 1035
rect 2296 933 2330 967
rect 2296 865 2330 899
rect 2296 797 2330 831
rect 2296 729 2330 763
rect 2296 661 2330 695
rect 2296 593 2330 627
rect 2296 525 2330 559
rect 2296 457 2330 491
rect 126 330 160 364
rect 126 262 160 296
rect 126 194 160 228
rect 2296 389 2330 423
rect 2296 321 2330 355
rect 2296 253 2330 287
rect 256 126 290 160
rect 324 126 358 160
rect 392 126 426 160
rect 460 126 494 160
rect 528 126 562 160
rect 596 126 630 160
rect 664 126 698 160
rect 732 126 766 160
rect 800 126 834 160
rect 868 126 902 160
rect 936 126 970 160
rect 1004 126 1038 160
rect 1072 126 1106 160
rect 1140 126 1174 160
rect 1208 126 1242 160
rect 1276 126 1310 160
rect 1344 126 1378 160
rect 1412 126 1446 160
rect 1480 126 1514 160
rect 1548 126 1582 160
rect 1616 126 1650 160
rect 1684 126 1718 160
rect 1752 126 1786 160
rect 1820 126 1854 160
rect 1888 126 1922 160
rect 1956 126 1990 160
rect 2024 126 2058 160
rect 2092 126 2126 160
rect 2160 126 2194 160
rect 2228 126 2262 160
<< poly >>
rect 1125 1627 1191 1643
rect 461 1527 493 1627
rect 1093 1593 1141 1627
rect 1175 1593 1191 1627
rect 1093 1559 1191 1593
rect 1093 1527 1141 1559
rect 1125 1525 1141 1527
rect 1175 1525 1191 1559
rect 1125 1509 1191 1525
rect 461 1261 493 1361
rect 1093 1345 1191 1361
rect 1093 1311 1141 1345
rect 1175 1311 1191 1345
rect 1093 1276 1191 1311
rect 1093 1261 1141 1276
rect 1125 1242 1141 1261
rect 1175 1242 1191 1276
rect 1125 1207 1191 1242
rect 1125 1205 1141 1207
rect 461 1105 493 1205
rect 1093 1173 1141 1205
rect 1175 1173 1191 1207
rect 1093 1138 1191 1173
rect 1093 1105 1141 1138
rect 1125 1104 1141 1105
rect 1175 1104 1191 1138
rect 1125 1069 1191 1104
rect 1125 1049 1141 1069
rect 461 949 493 1049
rect 1093 1035 1141 1049
rect 1175 1035 1191 1069
rect 1093 999 1191 1035
rect 1093 965 1141 999
rect 1175 965 1191 999
rect 1093 949 1191 965
rect 1454 1263 1486 1463
rect 1570 1447 1668 1463
rect 1570 1413 1618 1447
rect 1652 1413 1668 1447
rect 1570 1313 1668 1413
rect 1570 1279 1618 1313
rect 1652 1279 1668 1313
rect 1570 1263 1668 1279
rect 1831 1447 1929 1463
rect 1831 1413 1847 1447
rect 1881 1413 1929 1447
rect 1831 1313 1929 1413
rect 1831 1279 1847 1313
rect 1881 1279 1929 1313
rect 1831 1263 1929 1279
rect 2013 1263 2045 1463
rect 1630 1023 1696 1039
rect 1630 1005 1646 1023
rect 1358 905 1390 1005
rect 1590 989 1646 1005
rect 1680 989 1696 1023
rect 1590 955 1696 989
rect 1590 921 1646 955
rect 1680 921 1696 955
rect 1590 905 1696 921
rect 461 793 493 893
rect 1093 877 1191 893
rect 1093 843 1141 877
rect 1175 843 1191 877
rect 1093 808 1191 843
rect 1093 793 1141 808
rect 1125 774 1141 793
rect 1175 774 1191 808
rect 1125 739 1191 774
rect 1125 737 1141 739
rect 461 637 493 737
rect 1093 705 1141 737
rect 1175 705 1191 739
rect 1093 670 1191 705
rect 1093 637 1141 670
rect 1125 636 1141 637
rect 1175 636 1191 670
rect 1125 601 1191 636
rect 1125 581 1141 601
rect 461 481 493 581
rect 1093 567 1141 581
rect 1175 567 1191 601
rect 1093 531 1191 567
rect 1093 497 1141 531
rect 1175 497 1191 531
rect 1093 481 1191 497
rect 1358 637 1390 737
rect 1590 705 1804 737
rect 1590 671 1654 705
rect 1688 671 1722 705
rect 1756 671 1804 705
rect 1590 637 1804 671
rect 2104 637 2136 737
rect 1358 481 1390 581
rect 1590 549 1804 581
rect 1590 515 1654 549
rect 1688 515 1722 549
rect 1756 515 1804 549
rect 1590 481 1804 515
rect 2104 481 2136 581
<< polycont >>
rect 1141 1593 1175 1627
rect 1141 1525 1175 1559
rect 1141 1311 1175 1345
rect 1141 1242 1175 1276
rect 1141 1173 1175 1207
rect 1141 1104 1175 1138
rect 1141 1035 1175 1069
rect 1141 965 1175 999
rect 1618 1413 1652 1447
rect 1618 1279 1652 1313
rect 1847 1413 1881 1447
rect 1847 1279 1881 1313
rect 1646 989 1680 1023
rect 1646 921 1680 955
rect 1141 843 1175 877
rect 1141 774 1175 808
rect 1141 705 1175 739
rect 1141 636 1175 670
rect 1141 567 1175 601
rect 1141 497 1175 531
rect 1654 671 1688 705
rect 1722 671 1756 705
rect 1654 515 1688 549
rect 1722 515 1756 549
<< locali >>
rect 126 2225 194 2259
rect 232 2225 262 2259
rect 305 2225 330 2259
rect 378 2225 398 2259
rect 451 2225 466 2259
rect 524 2225 534 2259
rect 597 2225 602 2259
rect 704 2225 709 2259
rect 772 2225 782 2259
rect 840 2225 855 2259
rect 908 2225 928 2259
rect 976 2225 1000 2259
rect 1044 2225 1072 2259
rect 1112 2225 1144 2259
rect 1180 2225 1214 2259
rect 1250 2225 1282 2259
rect 1322 2225 1350 2259
rect 1394 2225 1418 2259
rect 1466 2225 1486 2259
rect 1538 2225 1554 2259
rect 1610 2225 1622 2259
rect 1682 2225 1690 2259
rect 1754 2225 1758 2259
rect 1860 2225 1864 2259
rect 1928 2225 1936 2259
rect 1996 2225 2008 2259
rect 2064 2225 2080 2259
rect 2132 2225 2152 2259
rect 2200 2225 2224 2259
rect 2258 2225 2330 2259
rect 126 2187 160 2225
rect 126 2115 160 2133
rect 126 2064 160 2081
rect 126 1996 160 2009
rect 126 1928 160 1937
rect 126 1860 160 1865
rect 126 1792 160 1793
rect 126 1755 160 1758
rect 2296 2191 2330 2225
rect 2296 2123 2330 2153
rect 2296 2055 2330 2078
rect 2296 1987 2330 2003
rect 2296 1919 2330 1928
rect 2296 1851 2330 1853
rect 2296 1812 2330 1817
rect 2296 1737 2330 1749
rect 126 1683 160 1690
rect 126 1611 160 1622
rect 126 1539 160 1554
rect 126 1467 160 1486
rect 126 1395 160 1418
rect 126 1323 160 1350
rect 126 1251 160 1282
rect 126 1180 160 1214
rect 126 1112 160 1145
rect 126 1044 160 1073
rect 126 976 160 1001
rect 126 908 160 928
rect 126 840 160 855
rect 126 772 160 782
rect 126 704 160 709
rect 126 597 160 602
rect 126 524 160 534
rect 126 451 160 466
rect 379 1678 413 1690
rect 605 1638 635 1672
rect 673 1638 707 1672
rect 749 1638 775 1672
rect 829 1638 843 1672
rect 909 1638 911 1672
rect 945 1638 955 1672
rect 1013 1638 1035 1672
rect 1081 1638 1097 1672
rect 2296 1662 2330 1681
rect 379 1602 413 1632
rect 379 1526 413 1562
rect 1141 1627 1175 1643
rect 1141 1559 1175 1593
rect 379 1456 413 1492
rect 605 1482 630 1516
rect 673 1482 704 1516
rect 741 1482 775 1516
rect 812 1482 843 1516
rect 886 1482 911 1516
rect 960 1482 979 1516
rect 1013 1482 1047 1516
rect 1081 1482 1097 1516
rect 1141 1509 1175 1521
rect 2296 1587 2330 1613
rect 2296 1512 2330 1545
rect 1464 1474 1498 1508
rect 1536 1474 1548 1508
rect 1951 1474 1967 1508
rect 2001 1474 2013 1508
rect 2047 1474 2085 1508
rect 1618 1447 1652 1463
rect 379 1386 413 1416
rect 555 1372 571 1406
rect 605 1372 639 1406
rect 673 1372 676 1406
rect 741 1372 751 1406
rect 809 1372 825 1406
rect 877 1372 899 1406
rect 945 1372 973 1406
rect 1013 1372 1047 1406
rect 1081 1372 1097 1406
rect 1282 1401 1316 1425
rect 379 1316 413 1340
rect 379 1246 413 1264
rect 1141 1345 1175 1361
rect 1141 1276 1175 1311
rect 605 1216 630 1250
rect 673 1216 704 1250
rect 741 1216 775 1250
rect 812 1216 843 1250
rect 886 1216 911 1250
rect 960 1216 979 1250
rect 1013 1216 1047 1250
rect 1081 1216 1097 1250
rect 379 1176 413 1188
rect 379 1106 413 1112
rect 1141 1207 1175 1218
rect 1141 1148 1175 1173
rect 379 1070 413 1072
rect 555 1060 571 1094
rect 605 1060 639 1094
rect 673 1060 676 1094
rect 741 1060 751 1094
rect 809 1060 825 1094
rect 877 1060 899 1094
rect 945 1060 973 1094
rect 1013 1060 1047 1094
rect 1081 1060 1097 1094
rect 1141 1069 1175 1104
rect 379 994 413 1002
rect 1141 999 1175 1010
rect 1141 949 1175 965
rect 1282 1329 1316 1367
rect 1282 1282 1316 1295
rect 1618 1404 1652 1413
rect 1847 1447 1881 1463
rect 1618 1370 1619 1404
rect 1618 1332 1653 1370
rect 1847 1345 1881 1413
rect 1618 1313 1619 1332
rect 1880 1313 1881 1345
rect 1618 1263 1652 1279
rect 1846 1279 1847 1311
rect 2296 1443 2330 1477
rect 2296 1375 2330 1403
rect 2296 1307 2330 1329
rect 1846 1273 1881 1279
rect 1282 1207 1316 1223
rect 1532 1218 1548 1252
rect 1880 1263 1881 1273
rect 1934 1252 1968 1255
rect 1934 1218 1967 1252
rect 2001 1218 2035 1252
rect 2296 1239 2330 1255
rect 1934 1217 1968 1218
rect 1282 1132 1316 1152
rect 1282 1057 1316 1081
rect 2296 1171 2330 1181
rect 2296 1103 2330 1107
rect 2296 1067 2330 1069
rect 1436 1016 1458 1050
rect 1504 1016 1538 1050
rect 1572 1016 1588 1050
rect 1282 982 1316 1010
rect 379 918 413 932
rect 605 904 630 938
rect 673 904 704 938
rect 741 904 775 938
rect 812 904 843 938
rect 886 904 911 938
rect 960 904 979 938
rect 1013 904 1047 938
rect 1081 904 1097 938
rect 1282 908 1316 939
rect 1646 972 1680 989
rect 1646 905 1680 921
rect 2296 993 2330 1001
rect 2296 919 2330 933
rect 379 842 413 862
rect 379 766 413 792
rect 1141 881 1175 893
rect 1141 808 1175 843
rect 555 748 571 782
rect 605 748 639 782
rect 673 748 676 782
rect 741 748 751 782
rect 809 748 825 782
rect 877 748 899 782
rect 945 748 973 782
rect 1013 748 1047 782
rect 1081 748 1097 782
rect 379 690 413 722
rect 379 616 413 652
rect 1141 739 1175 770
rect 1141 670 1175 693
rect 605 592 630 626
rect 673 592 704 626
rect 741 592 775 626
rect 812 592 843 626
rect 886 592 911 626
rect 960 592 979 626
rect 1013 592 1047 626
rect 1081 592 1097 626
rect 1141 601 1175 615
rect 379 546 413 580
rect 379 476 413 505
rect 1141 531 1175 537
rect 1141 481 1175 497
rect 1282 834 1316 868
rect 1386 860 1402 894
rect 1436 860 1470 894
rect 1504 882 1538 894
rect 1572 882 1588 894
rect 1516 860 1538 882
rect 1516 848 1554 860
rect 1282 760 1316 797
rect 2296 845 2330 865
rect 1386 748 1402 782
rect 1436 748 1470 782
rect 1516 748 1538 782
rect 1838 748 1854 782
rect 1888 748 1922 782
rect 1960 748 1990 782
rect 2024 748 2058 782
rect 2092 748 2108 782
rect 2296 771 2330 797
rect 1282 689 1316 726
rect 1638 671 1645 705
rect 1688 671 1717 705
rect 1756 671 1772 705
rect 2296 697 2330 729
rect 1282 618 1316 652
rect 2296 627 2330 661
rect 1436 592 1458 626
rect 1504 592 1538 626
rect 1572 592 1588 626
rect 1838 592 1854 626
rect 1907 592 1922 626
rect 1956 592 1966 626
rect 2024 592 2058 626
rect 2092 592 2108 626
rect 1282 547 1316 578
rect 2296 559 2330 589
rect 1638 515 1645 549
rect 1688 515 1717 549
rect 1756 515 1772 549
rect 1282 476 1316 504
rect 555 436 571 470
rect 605 436 639 470
rect 673 436 676 470
rect 741 436 751 470
rect 809 436 825 470
rect 877 436 899 470
rect 945 436 973 470
rect 1013 436 1047 470
rect 1081 436 1097 470
rect 2296 491 2330 515
rect 379 418 413 430
rect 1386 436 1402 470
rect 1436 436 1470 470
rect 1516 436 1538 470
rect 1838 436 1854 470
rect 1888 436 1922 470
rect 1960 436 1990 470
rect 2024 436 2058 470
rect 2092 436 2108 470
rect 1282 418 1316 430
rect 2296 423 2330 441
rect 126 378 160 398
rect 126 305 160 330
rect 126 232 160 262
rect 126 160 160 194
rect 2296 355 2330 389
rect 2296 287 2330 321
rect 2296 160 2330 253
rect 126 126 198 160
rect 232 126 256 160
rect 304 126 324 160
rect 376 126 392 160
rect 448 126 460 160
rect 520 126 528 160
rect 592 126 596 160
rect 698 126 702 160
rect 766 126 774 160
rect 834 126 846 160
rect 902 126 918 160
rect 970 126 990 160
rect 1038 126 1062 160
rect 1106 126 1135 160
rect 1174 126 1208 160
rect 1242 126 1276 160
rect 1315 126 1344 160
rect 1378 126 1412 160
rect 1446 126 1480 160
rect 1514 126 1548 160
rect 1582 126 1616 160
rect 1650 126 1684 160
rect 1718 126 1752 160
rect 1786 126 1820 160
rect 1854 126 1888 160
rect 1922 126 1956 160
rect 1990 126 2024 160
rect 2058 126 2092 160
rect 2126 126 2160 160
rect 2194 126 2228 160
rect 2262 126 2330 160
<< viali >>
rect 198 2225 228 2259
rect 228 2225 232 2259
rect 271 2225 296 2259
rect 296 2225 305 2259
rect 344 2225 364 2259
rect 364 2225 378 2259
rect 417 2225 432 2259
rect 432 2225 451 2259
rect 490 2225 500 2259
rect 500 2225 524 2259
rect 563 2225 568 2259
rect 568 2225 597 2259
rect 636 2225 670 2259
rect 709 2225 738 2259
rect 738 2225 743 2259
rect 782 2225 806 2259
rect 806 2225 816 2259
rect 855 2225 874 2259
rect 874 2225 889 2259
rect 928 2225 942 2259
rect 942 2225 962 2259
rect 1000 2225 1010 2259
rect 1010 2225 1034 2259
rect 1072 2225 1078 2259
rect 1078 2225 1106 2259
rect 1144 2225 1146 2259
rect 1146 2225 1178 2259
rect 1216 2225 1248 2259
rect 1248 2225 1250 2259
rect 1288 2225 1316 2259
rect 1316 2225 1322 2259
rect 1360 2225 1384 2259
rect 1384 2225 1394 2259
rect 1432 2225 1452 2259
rect 1452 2225 1466 2259
rect 1504 2225 1520 2259
rect 1520 2225 1538 2259
rect 1576 2225 1588 2259
rect 1588 2225 1610 2259
rect 1648 2225 1656 2259
rect 1656 2225 1682 2259
rect 1720 2225 1724 2259
rect 1724 2225 1754 2259
rect 1792 2225 1826 2259
rect 1864 2225 1894 2259
rect 1894 2225 1898 2259
rect 1936 2225 1962 2259
rect 1962 2225 1970 2259
rect 2008 2225 2030 2259
rect 2030 2225 2042 2259
rect 2080 2225 2098 2259
rect 2098 2225 2114 2259
rect 2152 2225 2166 2259
rect 2166 2225 2186 2259
rect 2224 2225 2258 2259
rect 126 2167 160 2187
rect 126 2153 160 2167
rect 126 2081 160 2115
rect 126 2030 160 2043
rect 126 2009 160 2030
rect 126 1962 160 1971
rect 126 1937 160 1962
rect 126 1894 160 1899
rect 126 1865 160 1894
rect 126 1826 160 1827
rect 126 1793 160 1826
rect 126 1724 160 1755
rect 126 1721 160 1724
rect 2296 2157 2330 2187
rect 2296 2153 2330 2157
rect 2296 2089 2330 2112
rect 2296 2078 2330 2089
rect 2296 2021 2330 2037
rect 2296 2003 2330 2021
rect 2296 1953 2330 1962
rect 2296 1928 2330 1953
rect 2296 1885 2330 1887
rect 2296 1853 2330 1885
rect 2296 1783 2330 1812
rect 2296 1778 2330 1783
rect 2296 1715 2330 1737
rect 2296 1703 2330 1715
rect 126 1656 160 1683
rect 126 1649 160 1656
rect 126 1588 160 1611
rect 126 1577 160 1588
rect 126 1520 160 1539
rect 126 1505 160 1520
rect 126 1452 160 1467
rect 126 1433 160 1452
rect 126 1384 160 1395
rect 126 1361 160 1384
rect 126 1316 160 1323
rect 126 1289 160 1316
rect 126 1248 160 1251
rect 126 1217 160 1248
rect 126 1146 160 1179
rect 126 1145 160 1146
rect 126 1078 160 1107
rect 126 1073 160 1078
rect 126 1010 160 1035
rect 126 1001 160 1010
rect 126 942 160 962
rect 126 928 160 942
rect 126 874 160 889
rect 126 855 160 874
rect 126 806 160 816
rect 126 782 160 806
rect 126 738 160 743
rect 126 709 160 738
rect 126 636 160 670
rect 126 568 160 597
rect 126 563 160 568
rect 126 500 160 524
rect 126 490 160 500
rect 126 432 160 451
rect 126 417 160 432
rect 379 1666 413 1678
rect 379 1644 413 1666
rect 555 1638 571 1672
rect 571 1638 589 1672
rect 635 1638 639 1672
rect 639 1638 669 1672
rect 715 1638 741 1672
rect 741 1638 749 1672
rect 795 1638 809 1672
rect 809 1638 829 1672
rect 875 1638 877 1672
rect 877 1638 909 1672
rect 955 1638 979 1672
rect 979 1638 989 1672
rect 1035 1638 1047 1672
rect 1047 1638 1069 1672
rect 2296 1647 2330 1662
rect 379 1596 413 1602
rect 379 1568 413 1596
rect 379 1492 413 1526
rect 1141 1593 1175 1627
rect 1141 1525 1175 1555
rect 1141 1521 1175 1525
rect 555 1482 571 1516
rect 571 1482 589 1516
rect 630 1482 639 1516
rect 639 1482 664 1516
rect 704 1482 707 1516
rect 707 1482 738 1516
rect 778 1482 809 1516
rect 809 1482 812 1516
rect 852 1482 877 1516
rect 877 1482 886 1516
rect 926 1482 945 1516
rect 945 1482 960 1516
rect 2296 1628 2330 1647
rect 2296 1579 2330 1587
rect 2296 1553 2330 1579
rect 2296 1511 2330 1512
rect 1430 1474 1464 1508
rect 1502 1474 1532 1508
rect 1532 1474 1536 1508
rect 2013 1474 2047 1508
rect 2085 1474 2119 1508
rect 2296 1478 2330 1511
rect 379 1422 413 1450
rect 379 1416 413 1422
rect 379 1352 413 1374
rect 676 1372 707 1406
rect 707 1372 710 1406
rect 751 1372 775 1406
rect 775 1372 785 1406
rect 825 1372 843 1406
rect 843 1372 859 1406
rect 899 1372 911 1406
rect 911 1372 933 1406
rect 973 1372 979 1406
rect 979 1372 1007 1406
rect 1047 1372 1081 1406
rect 379 1340 413 1352
rect 379 1282 413 1298
rect 379 1264 413 1282
rect 379 1212 413 1222
rect 555 1216 571 1250
rect 571 1216 589 1250
rect 630 1216 639 1250
rect 639 1216 664 1250
rect 704 1216 707 1250
rect 707 1216 738 1250
rect 778 1216 809 1250
rect 809 1216 812 1250
rect 852 1216 877 1250
rect 877 1216 886 1250
rect 926 1216 945 1250
rect 945 1216 960 1250
rect 1141 1242 1175 1252
rect 1141 1218 1175 1242
rect 379 1188 413 1212
rect 379 1142 413 1146
rect 379 1112 413 1142
rect 1141 1138 1175 1148
rect 1141 1114 1175 1138
rect 379 1036 413 1070
rect 676 1060 707 1094
rect 707 1060 710 1094
rect 751 1060 775 1094
rect 775 1060 785 1094
rect 825 1060 843 1094
rect 843 1060 859 1094
rect 899 1060 911 1094
rect 911 1060 933 1094
rect 973 1060 979 1094
rect 979 1060 1007 1094
rect 1047 1060 1081 1094
rect 379 966 413 994
rect 379 960 413 966
rect 1141 1035 1175 1044
rect 1141 1010 1175 1035
rect 1282 1257 1316 1282
rect 1619 1370 1653 1404
rect 1619 1313 1653 1332
rect 1619 1298 1652 1313
rect 1652 1298 1653 1313
rect 1846 1313 1880 1345
rect 1846 1311 1847 1313
rect 1847 1311 1880 1313
rect 2296 1409 2330 1437
rect 2296 1403 2330 1409
rect 2296 1341 2330 1363
rect 2296 1329 2330 1341
rect 1282 1248 1316 1257
rect 1476 1218 1498 1252
rect 1498 1218 1510 1252
rect 1548 1218 1582 1252
rect 1846 1239 1880 1273
rect 1934 1255 1968 1289
rect 2296 1273 2330 1289
rect 2296 1255 2330 1273
rect 1282 1186 1316 1207
rect 1282 1173 1316 1186
rect 1934 1183 1968 1217
rect 2296 1205 2330 1215
rect 1282 1115 1316 1132
rect 1282 1098 1316 1115
rect 1282 1044 1316 1057
rect 2296 1181 2330 1205
rect 2296 1137 2330 1141
rect 2296 1107 2330 1137
rect 1282 1023 1316 1044
rect 1386 1016 1402 1050
rect 1402 1016 1420 1050
rect 1458 1016 1470 1050
rect 1470 1016 1492 1050
rect 1646 1023 1680 1044
rect 1282 973 1316 982
rect 1282 948 1316 973
rect 379 896 413 918
rect 555 904 571 938
rect 571 904 589 938
rect 630 904 639 938
rect 639 904 664 938
rect 704 904 707 938
rect 707 904 738 938
rect 778 904 809 938
rect 809 904 812 938
rect 852 904 877 938
rect 877 904 886 938
rect 926 904 945 938
rect 945 904 960 938
rect 379 884 413 896
rect 1282 902 1316 908
rect 1646 1010 1680 1023
rect 1646 955 1680 972
rect 1646 938 1680 955
rect 2296 1035 2330 1067
rect 2296 1033 2330 1035
rect 2296 967 2330 993
rect 2296 959 2330 967
rect 379 826 413 842
rect 379 808 413 826
rect 1141 877 1175 881
rect 1141 847 1175 877
rect 379 756 413 766
rect 379 732 413 756
rect 676 748 707 782
rect 707 748 710 782
rect 751 748 775 782
rect 775 748 785 782
rect 825 748 843 782
rect 843 748 859 782
rect 899 748 911 782
rect 911 748 933 782
rect 973 748 979 782
rect 979 748 1007 782
rect 1047 748 1081 782
rect 1141 774 1175 804
rect 1141 770 1175 774
rect 379 686 413 690
rect 379 656 413 686
rect 1141 705 1175 727
rect 1141 693 1175 705
rect 1141 636 1175 649
rect 379 582 413 614
rect 555 592 571 626
rect 571 592 589 626
rect 630 592 639 626
rect 639 592 664 626
rect 704 592 707 626
rect 707 592 738 626
rect 778 592 809 626
rect 809 592 812 626
rect 852 592 877 626
rect 877 592 886 626
rect 926 592 945 626
rect 945 592 960 626
rect 1141 615 1175 636
rect 379 580 413 582
rect 379 512 413 539
rect 379 505 413 512
rect 1141 567 1175 571
rect 1141 537 1175 567
rect 1282 874 1316 902
rect 2296 899 2330 919
rect 1482 860 1504 882
rect 1504 860 1516 882
rect 1554 860 1572 882
rect 1572 860 1588 882
rect 1482 848 1516 860
rect 1554 848 1588 860
rect 2296 885 2330 899
rect 1282 831 1316 834
rect 1282 800 1316 831
rect 2296 831 2330 845
rect 2296 811 2330 831
rect 1282 726 1316 760
rect 1482 748 1504 782
rect 1504 748 1516 782
rect 1554 748 1572 782
rect 1572 748 1588 782
rect 1854 748 1888 782
rect 1926 748 1956 782
rect 1956 748 1960 782
rect 2296 763 2330 771
rect 2296 737 2330 763
rect 1282 655 1316 686
rect 1645 671 1654 705
rect 1654 671 1679 705
rect 1717 671 1722 705
rect 1722 671 1751 705
rect 2296 695 2330 697
rect 1282 652 1316 655
rect 2296 663 2330 695
rect 1282 584 1316 612
rect 1386 592 1402 626
rect 1402 592 1420 626
rect 1458 592 1470 626
rect 1470 592 1492 626
rect 1873 592 1888 626
rect 1888 592 1907 626
rect 1966 592 1990 626
rect 1990 592 2000 626
rect 2058 592 2092 626
rect 2296 593 2330 623
rect 1282 578 1316 584
rect 2296 589 2330 593
rect 1282 513 1316 538
rect 1645 515 1654 549
rect 1654 515 1679 549
rect 1717 515 1722 549
rect 1722 515 1751 549
rect 2296 525 2330 549
rect 2296 515 2330 525
rect 1282 504 1316 513
rect 379 442 413 464
rect 379 430 413 442
rect 676 436 707 470
rect 707 436 710 470
rect 751 436 775 470
rect 775 436 785 470
rect 825 436 843 470
rect 843 436 859 470
rect 899 436 911 470
rect 911 436 933 470
rect 973 436 979 470
rect 979 436 1007 470
rect 1047 436 1081 470
rect 1282 442 1316 464
rect 1282 430 1316 442
rect 1482 436 1504 470
rect 1504 436 1516 470
rect 1554 436 1572 470
rect 1572 436 1588 470
rect 1854 436 1888 470
rect 1926 436 1956 470
rect 1956 436 1960 470
rect 2296 457 2330 475
rect 2296 441 2330 457
rect 126 364 160 378
rect 126 344 160 364
rect 126 296 160 305
rect 126 271 160 296
rect 126 228 160 232
rect 126 198 160 228
rect 198 126 232 160
rect 270 126 290 160
rect 290 126 304 160
rect 342 126 358 160
rect 358 126 376 160
rect 414 126 426 160
rect 426 126 448 160
rect 486 126 494 160
rect 494 126 520 160
rect 558 126 562 160
rect 562 126 592 160
rect 630 126 664 160
rect 702 126 732 160
rect 732 126 736 160
rect 774 126 800 160
rect 800 126 808 160
rect 846 126 868 160
rect 868 126 880 160
rect 918 126 936 160
rect 936 126 952 160
rect 990 126 1004 160
rect 1004 126 1024 160
rect 1062 126 1072 160
rect 1072 126 1096 160
rect 1135 126 1140 160
rect 1140 126 1169 160
rect 1208 126 1242 160
rect 1281 126 1310 160
rect 1310 126 1315 160
<< metal1 >>
rect 120 2259 2336 2265
rect 120 2225 198 2259
rect 232 2225 271 2259
rect 305 2225 344 2259
rect 378 2225 417 2259
rect 451 2225 490 2259
rect 524 2225 563 2259
rect 597 2225 636 2259
rect 670 2225 709 2259
rect 743 2225 782 2259
rect 816 2225 855 2259
rect 889 2225 928 2259
rect 962 2225 1000 2259
rect 1034 2225 1072 2259
rect 1106 2225 1144 2259
rect 1178 2225 1216 2259
rect 1250 2225 1288 2259
rect 1322 2225 1360 2259
rect 1394 2225 1432 2259
rect 1466 2225 1504 2259
rect 1538 2225 1576 2259
rect 1610 2225 1648 2259
rect 1682 2225 1720 2259
rect 1754 2225 1792 2259
rect 1826 2225 1864 2259
rect 1898 2225 1936 2259
rect 1970 2225 2008 2259
rect 2042 2225 2080 2259
rect 2114 2225 2152 2259
rect 2186 2225 2224 2259
rect 2258 2225 2336 2259
rect 120 2213 2336 2225
rect 120 2187 174 2213
tri 174 2187 200 2213 nw
tri 2256 2187 2282 2213 ne
rect 2282 2187 2336 2213
rect 120 2153 126 2187
rect 160 2153 166 2187
tri 166 2179 174 2187 nw
tri 2282 2179 2290 2187 ne
rect 120 2115 166 2153
rect 120 2081 126 2115
rect 160 2081 166 2115
rect 120 2043 166 2081
rect 120 2009 126 2043
rect 160 2009 166 2043
rect 120 1971 166 2009
rect 120 1937 126 1971
rect 160 1937 166 1971
rect 120 1899 166 1937
rect 120 1865 126 1899
rect 160 1865 166 1899
rect 120 1827 166 1865
rect 120 1793 126 1827
rect 160 1793 166 1827
rect 120 1755 166 1793
rect 120 1721 126 1755
rect 160 1721 166 1755
rect 120 1683 166 1721
rect 2290 2153 2296 2187
rect 2330 2153 2336 2187
rect 2290 2112 2336 2153
rect 2290 2078 2296 2112
rect 2330 2078 2336 2112
rect 2290 2037 2336 2078
rect 2290 2003 2296 2037
rect 2330 2003 2336 2037
rect 2290 1962 2336 2003
rect 2290 1928 2296 1962
rect 2330 1928 2336 1962
rect 2290 1887 2336 1928
rect 2290 1853 2296 1887
rect 2330 1853 2336 1887
rect 2290 1812 2336 1853
rect 2290 1778 2296 1812
rect 2330 1778 2336 1812
rect 2290 1737 2336 1778
rect 2290 1703 2296 1737
rect 2330 1703 2336 1737
rect 120 1649 126 1683
rect 160 1649 166 1683
rect 120 1611 166 1649
rect 120 1577 126 1611
rect 160 1577 166 1611
rect 120 1539 166 1577
rect 120 1505 126 1539
rect 160 1505 166 1539
rect 120 1467 166 1505
rect 120 1433 126 1467
rect 160 1433 166 1467
rect 120 1395 166 1433
rect 120 1361 126 1395
rect 160 1361 166 1395
rect 120 1323 166 1361
rect 120 1289 126 1323
rect 160 1289 166 1323
rect 120 1251 166 1289
rect 120 1217 126 1251
rect 160 1217 166 1251
rect 120 1179 166 1217
rect 120 1145 126 1179
rect 160 1145 166 1179
rect 120 1107 166 1145
rect 120 1073 126 1107
rect 160 1073 166 1107
rect 120 1035 166 1073
rect 120 1001 126 1035
rect 160 1001 166 1035
rect 120 962 166 1001
rect 120 928 126 962
rect 160 928 166 962
rect 120 889 166 928
rect 120 855 126 889
rect 160 855 166 889
rect 120 816 166 855
rect 120 782 126 816
rect 160 782 166 816
rect 120 743 166 782
rect 120 709 126 743
rect 160 709 166 743
rect 120 670 166 709
rect 120 636 126 670
rect 160 636 166 670
rect 120 597 166 636
rect 120 563 126 597
rect 160 563 166 597
rect 120 524 166 563
rect 120 490 126 524
rect 160 490 166 524
rect 120 451 166 490
rect 120 417 126 451
rect 160 417 166 451
rect 120 378 166 417
rect 120 344 126 378
rect 160 344 166 378
rect 120 305 166 344
rect 120 271 126 305
rect 160 271 166 305
rect 120 232 166 271
rect 219 1678 1081 1690
rect 219 1644 379 1678
rect 413 1672 1081 1678
rect 2290 1672 2336 1703
rect 413 1644 555 1672
rect 219 1638 555 1644
rect 589 1638 635 1672
rect 669 1638 715 1672
rect 749 1638 795 1672
rect 829 1638 875 1672
rect 909 1638 955 1672
rect 989 1638 1035 1672
rect 1069 1638 1081 1672
rect 2013 1662 2336 1672
rect 219 1632 1081 1638
rect 1135 1637 1181 1639
rect 219 1602 419 1632
rect 219 1568 379 1602
rect 413 1568 419 1602
rect 219 1526 419 1568
rect 219 1492 379 1526
rect 413 1492 419 1526
rect 1132 1631 1184 1637
rect 1132 1567 1184 1579
rect 219 1450 419 1492
rect 219 1416 379 1450
rect 413 1416 419 1450
rect 219 1374 419 1416
rect 219 1340 379 1374
rect 413 1340 419 1374
rect 219 1298 419 1340
rect 219 1264 379 1298
rect 413 1264 419 1298
rect 219 1222 419 1264
rect 219 1188 379 1222
rect 413 1188 419 1222
rect 219 1146 419 1188
rect 219 1112 379 1146
rect 413 1112 419 1146
rect 219 1070 419 1112
rect 219 1036 379 1070
rect 413 1036 419 1070
rect 219 994 419 1036
rect 219 960 379 994
rect 413 960 419 994
rect 219 918 419 960
rect 219 884 379 918
rect 413 884 419 918
rect 219 842 419 884
rect 219 808 379 842
rect 413 808 419 842
rect 219 766 419 808
rect 219 732 379 766
rect 413 732 419 766
rect 219 690 419 732
rect 219 656 379 690
rect 413 656 419 690
rect 219 614 419 656
rect 219 580 379 614
rect 413 580 419 614
rect 474 1516 972 1522
rect 474 1482 555 1516
rect 589 1482 630 1516
rect 664 1482 704 1516
rect 738 1482 778 1516
rect 812 1482 852 1516
rect 886 1482 926 1516
rect 960 1482 972 1516
rect 1132 1509 1184 1515
rect 2013 1628 2296 1662
rect 2330 1628 2336 1662
rect 2013 1587 2336 1628
rect 2013 1553 2296 1587
rect 2330 1553 2336 1587
rect 2013 1514 2336 1553
rect 1418 1512 2336 1514
rect 474 1476 972 1482
rect 1418 1508 2296 1512
rect 474 1256 574 1476
rect 1418 1474 1430 1508
rect 1464 1474 1502 1508
rect 1536 1474 2013 1508
rect 2047 1474 2085 1508
rect 2119 1478 2296 1508
rect 2330 1478 2336 1512
rect 2119 1474 2336 1478
rect 1418 1468 2336 1474
rect 2013 1437 2336 1468
rect 1613 1412 1774 1437
rect 664 1406 1774 1412
rect 664 1372 676 1406
rect 710 1372 751 1406
rect 785 1372 825 1406
rect 859 1372 899 1406
rect 933 1372 973 1406
rect 1007 1372 1047 1406
rect 1081 1404 1774 1406
rect 1081 1372 1619 1404
rect 664 1370 1619 1372
rect 1653 1385 1774 1404
rect 1826 1385 1838 1437
rect 1890 1385 1974 1437
rect 1653 1370 1659 1385
rect 664 1366 1659 1370
rect 1033 1332 1659 1366
rect 474 1250 972 1256
rect 474 1216 555 1250
rect 589 1216 630 1250
rect 664 1216 704 1250
rect 738 1216 778 1250
rect 812 1216 852 1250
rect 886 1216 926 1250
rect 960 1216 972 1250
rect 474 1210 972 1216
rect 474 944 574 1210
rect 1033 1100 1093 1332
rect 1613 1298 1619 1332
rect 1653 1298 1659 1332
rect 1276 1282 1322 1294
rect 1613 1286 1659 1298
rect 1840 1345 1886 1357
rect 1840 1311 1846 1345
rect 1880 1311 1886 1345
rect 1135 1252 1181 1264
rect 1135 1247 1141 1252
rect 1132 1241 1141 1247
rect 1175 1247 1181 1252
rect 1276 1248 1282 1282
rect 1316 1248 1322 1282
tri 1838 1273 1840 1275 se
rect 1840 1273 1886 1311
tri 1823 1258 1838 1273 se
rect 1838 1258 1846 1273
rect 1175 1241 1184 1247
rect 1132 1177 1184 1189
rect 1132 1119 1141 1125
rect 664 1094 1093 1100
rect 664 1060 676 1094
rect 710 1060 751 1094
rect 785 1060 825 1094
rect 859 1060 899 1094
rect 933 1060 973 1094
rect 1007 1060 1047 1094
rect 1081 1060 1093 1094
rect 664 1054 1093 1060
rect 1135 1114 1141 1119
rect 1175 1119 1184 1125
rect 1276 1207 1322 1248
rect 1276 1173 1282 1207
rect 1316 1173 1322 1207
rect 1464 1252 1846 1258
rect 1464 1218 1476 1252
rect 1510 1218 1548 1252
rect 1582 1218 1764 1252
rect 1464 1206 1764 1218
rect 1276 1132 1322 1173
rect 1175 1114 1181 1119
rect 1135 1044 1181 1114
rect 1135 1010 1141 1044
rect 1175 1010 1181 1044
rect 1135 998 1181 1010
rect 1276 1098 1282 1132
rect 1316 1098 1322 1132
rect 1816 1239 1846 1252
rect 1880 1239 1886 1273
rect 1816 1206 1886 1239
rect 1928 1289 1974 1385
rect 1928 1255 1934 1289
rect 1968 1255 1974 1289
rect 1928 1217 1974 1255
rect 1764 1188 1816 1200
rect 1928 1183 1934 1217
rect 1968 1183 1974 1217
rect 1928 1171 1974 1183
rect 2013 1403 2296 1437
rect 2330 1403 2336 1437
rect 2013 1363 2336 1403
rect 2013 1329 2296 1363
rect 2330 1329 2336 1363
rect 2013 1289 2336 1329
rect 2013 1255 2296 1289
rect 2330 1255 2336 1289
rect 2013 1215 2336 1255
rect 2013 1181 2296 1215
rect 2330 1181 2336 1215
rect 1764 1130 1816 1136
rect 2013 1141 2336 1181
rect 1276 1084 1322 1098
rect 2013 1107 2296 1141
rect 2330 1107 2336 1141
rect 1276 1057 1440 1084
rect 1276 1023 1282 1057
rect 1316 1056 1440 1057
rect 2013 1067 2336 1107
rect 1316 1050 1504 1056
rect 1640 1054 1686 1056
rect 1316 1023 1386 1050
rect 1276 1016 1386 1023
rect 1420 1016 1458 1050
rect 1492 1016 1504 1050
rect 1276 1010 1504 1016
rect 1637 1048 1689 1054
rect 1276 982 1440 1010
rect 1276 948 1282 982
rect 1316 948 1440 982
rect 474 938 972 944
rect 474 904 555 938
rect 589 904 630 938
rect 664 904 704 938
rect 738 904 778 938
rect 812 904 852 938
rect 886 904 926 938
rect 960 904 972 938
rect 474 898 972 904
rect 1276 908 1440 948
rect 1637 984 1689 996
rect 2013 1033 2296 1067
rect 2330 1033 2336 1067
rect 2013 993 2336 1033
rect 1637 926 1689 932
rect 1844 964 1896 970
rect 474 632 574 898
rect 1132 887 1184 893
rect 1132 823 1184 835
rect 664 782 1093 788
rect 664 748 676 782
rect 710 748 751 782
rect 785 748 825 782
rect 859 748 899 782
rect 933 748 973 782
rect 1007 748 1047 782
rect 1081 748 1093 782
rect 1132 770 1141 771
rect 1175 770 1184 771
rect 1132 765 1184 770
rect 1276 874 1282 908
rect 1316 874 1440 908
rect 1844 900 1896 912
rect 1276 834 1440 874
rect 1470 882 1844 888
rect 1470 848 1482 882
rect 1516 848 1554 882
rect 1588 848 1844 882
rect 1470 842 1896 848
rect 2013 959 2296 993
rect 2330 959 2336 993
rect 2013 919 2336 959
rect 2013 885 2296 919
rect 2330 885 2336 919
rect 2013 845 2336 885
rect 1276 800 1282 834
rect 1316 800 1440 834
rect 664 742 1093 748
rect 1033 708 1093 742
rect 1033 656 1041 708
rect 1033 644 1093 656
rect 474 626 972 632
rect 474 592 555 626
rect 589 592 630 626
rect 664 592 704 626
rect 738 592 778 626
rect 812 592 852 626
rect 886 592 926 626
rect 960 592 972 626
rect 474 586 972 592
rect 1033 592 1041 644
rect 219 539 419 580
rect 219 505 379 539
rect 413 505 419 539
rect 219 464 419 505
rect 1033 476 1093 592
rect 1135 727 1181 765
rect 1135 693 1141 727
rect 1175 693 1181 727
rect 1135 649 1181 693
rect 1135 615 1141 649
rect 1175 615 1181 649
rect 1135 571 1181 615
rect 1135 537 1141 571
rect 1175 537 1181 571
rect 1135 525 1181 537
rect 1276 760 1440 800
rect 2013 811 2296 845
rect 2330 811 2336 845
rect 1529 788 1535 794
rect 1276 726 1282 760
rect 1316 726 1440 760
rect 1470 782 1535 788
rect 1587 782 1599 794
rect 1470 748 1482 782
rect 1516 748 1535 782
rect 1588 748 1599 782
rect 1470 742 1535 748
rect 1587 742 1599 748
rect 1651 788 1657 794
rect 1651 782 1972 788
rect 1651 748 1854 782
rect 1888 748 1926 782
rect 1960 748 1972 782
rect 1651 742 1972 748
rect 2013 771 2336 811
rect 1276 686 1440 726
rect 2013 737 2296 771
rect 2330 737 2336 771
rect 1636 711 1642 714
rect 1276 652 1282 686
rect 1316 652 1440 686
rect 1633 665 1642 711
rect 1636 662 1642 665
rect 1694 662 1706 714
rect 1758 662 1764 714
rect 2013 697 2336 737
rect 2013 663 2296 697
rect 2330 663 2336 697
rect 1276 632 1440 652
rect 2013 632 2336 663
rect 1276 626 1504 632
rect 1276 612 1386 626
rect 1276 578 1282 612
rect 1316 592 1386 612
rect 1420 592 1458 626
rect 1492 592 1504 626
rect 1316 586 1504 592
rect 1861 626 2336 632
rect 1861 592 1873 626
rect 1907 592 1966 626
rect 2000 592 2058 626
rect 2092 623 2336 626
rect 2092 592 2296 623
rect 1861 589 2296 592
rect 2330 589 2336 623
rect 1861 586 2336 589
rect 1316 578 1440 586
rect 1276 538 1440 578
rect 1636 555 1642 558
rect 219 455 379 464
rect 219 403 225 455
rect 277 403 293 455
rect 345 403 361 455
rect 413 403 419 464
rect 664 470 1093 476
rect 664 436 676 470
rect 710 436 751 470
rect 785 436 825 470
rect 859 436 899 470
rect 933 436 973 470
rect 1007 436 1047 470
rect 1081 436 1093 470
rect 664 430 1093 436
rect 1276 504 1282 538
rect 1316 504 1440 538
rect 1633 509 1642 555
rect 1636 506 1642 509
rect 1694 506 1706 558
rect 1758 506 1764 558
rect 2013 549 2336 586
rect 2013 515 2296 549
rect 2330 515 2336 549
rect 1276 464 1440 504
rect 1276 449 1282 464
rect 1316 449 1440 464
rect 219 381 419 403
rect 219 329 225 381
rect 277 329 293 381
rect 345 329 361 381
rect 413 329 419 381
rect 219 307 419 329
rect 219 255 225 307
rect 277 255 293 307
rect 345 255 361 307
rect 413 255 419 307
rect 1328 397 1386 449
rect 1438 397 1440 449
rect 1470 470 1854 476
rect 1470 436 1482 470
rect 1516 436 1554 470
rect 1588 436 1854 470
rect 1470 430 1854 436
rect 1848 424 1854 430
rect 1906 424 1918 476
rect 1970 424 1976 476
rect 2013 475 2336 515
rect 2013 441 2296 475
rect 2330 441 2336 475
rect 2013 407 2336 441
rect 1276 381 1440 397
rect 1328 329 1386 381
rect 1438 329 1440 381
rect 1276 313 1440 329
rect 1328 261 1386 313
rect 1438 261 1440 313
rect 1276 255 1440 261
rect 120 198 126 232
rect 160 198 166 232
rect 120 166 166 198
tri 166 166 200 200 sw
rect 120 160 1327 166
rect 120 126 198 160
rect 232 126 270 160
rect 304 126 342 160
rect 376 126 414 160
rect 448 126 486 160
rect 520 126 558 160
rect 592 126 630 160
rect 664 126 702 160
rect 736 126 774 160
rect 808 126 846 160
rect 880 126 918 160
rect 952 126 990 160
rect 1024 126 1062 160
rect 1096 126 1135 160
rect 1169 126 1208 160
rect 1242 126 1281 160
rect 1315 126 1327 160
rect 120 120 1327 126
<< via1 >>
rect 1132 1627 1184 1631
rect 1132 1593 1141 1627
rect 1141 1593 1175 1627
rect 1175 1593 1184 1627
rect 1132 1579 1184 1593
rect 1132 1555 1184 1567
rect 1132 1521 1141 1555
rect 1141 1521 1175 1555
rect 1175 1521 1184 1555
rect 1132 1515 1184 1521
rect 1774 1385 1826 1437
rect 1838 1385 1890 1437
rect 1132 1218 1141 1241
rect 1141 1218 1175 1241
rect 1175 1218 1184 1241
rect 1132 1189 1184 1218
rect 1132 1148 1184 1177
rect 1132 1125 1141 1148
rect 1141 1125 1175 1148
rect 1175 1125 1184 1148
rect 1764 1200 1816 1252
rect 1764 1136 1816 1188
rect 1637 1044 1689 1048
rect 1637 1010 1646 1044
rect 1646 1010 1680 1044
rect 1680 1010 1689 1044
rect 1637 996 1689 1010
rect 1637 972 1689 984
rect 1637 938 1646 972
rect 1646 938 1680 972
rect 1680 938 1689 972
rect 1637 932 1689 938
rect 1132 881 1184 887
rect 1132 847 1141 881
rect 1141 847 1175 881
rect 1175 847 1184 881
rect 1132 835 1184 847
rect 1132 804 1184 823
rect 1132 771 1141 804
rect 1141 771 1175 804
rect 1175 771 1184 804
rect 1844 912 1896 964
rect 1844 848 1896 900
rect 1041 656 1093 708
rect 1041 592 1093 644
rect 1535 782 1587 794
rect 1535 748 1554 782
rect 1554 748 1587 782
rect 1535 742 1587 748
rect 1599 742 1651 794
rect 1642 705 1694 714
rect 1642 671 1645 705
rect 1645 671 1679 705
rect 1679 671 1694 705
rect 1642 662 1694 671
rect 1706 705 1758 714
rect 1706 671 1717 705
rect 1717 671 1751 705
rect 1751 671 1758 705
rect 1706 662 1758 671
rect 225 403 277 455
rect 293 403 345 455
rect 361 430 379 455
rect 379 430 413 455
rect 361 403 413 430
rect 1642 549 1694 558
rect 1642 515 1645 549
rect 1645 515 1679 549
rect 1679 515 1694 549
rect 1642 506 1694 515
rect 1706 549 1758 558
rect 1706 515 1717 549
rect 1717 515 1751 549
rect 1751 515 1758 549
rect 1706 506 1758 515
rect 1276 430 1282 449
rect 1282 430 1316 449
rect 1316 430 1328 449
rect 225 329 277 381
rect 293 329 345 381
rect 361 329 413 381
rect 225 255 277 307
rect 293 255 345 307
rect 361 255 413 307
rect 1276 397 1328 430
rect 1386 397 1438 449
rect 1854 470 1906 476
rect 1854 436 1888 470
rect 1888 436 1906 470
rect 1854 424 1906 436
rect 1918 470 1970 476
rect 1918 436 1926 470
rect 1926 436 1960 470
rect 1960 436 1970 470
rect 1918 424 1970 436
rect 1276 329 1328 381
rect 1386 329 1438 381
rect 1276 261 1328 313
rect 1386 261 1438 313
<< metal2 >>
rect 1132 1631 1184 2125
rect 1132 1567 1184 1579
rect 1132 1509 1184 1515
tri 1220 1441 1242 1463 se
rect 1242 1441 1294 2124
tri 1216 1437 1220 1441 se
rect 1220 1437 1290 1441
tri 1290 1437 1294 1441 nw
tri 1184 1405 1216 1437 se
rect 1216 1405 1258 1437
tri 1258 1405 1290 1437 nw
tri 1164 1385 1184 1405 se
rect 1184 1385 1238 1405
tri 1238 1385 1258 1405 nw
tri 1132 1353 1164 1385 se
rect 1164 1371 1224 1385
tri 1224 1371 1238 1385 nw
rect 1164 1353 1184 1371
rect 1132 1241 1184 1353
tri 1184 1331 1224 1371 nw
tri 1306 1331 1346 1371 se
rect 1346 1349 1398 2124
tri 1272 1297 1306 1331 se
rect 1306 1297 1346 1331
tri 1346 1297 1398 1349 nw
rect 1132 1177 1184 1189
rect 1132 1119 1184 1125
tri 1236 1261 1272 1297 se
rect 1272 1261 1310 1297
tri 1310 1261 1346 1297 nw
rect 1236 1252 1301 1261
tri 1301 1252 1310 1261 nw
tri 1220 932 1236 948 se
rect 1236 932 1288 1252
tri 1288 1239 1301 1252 nw
tri 1200 912 1220 932 se
rect 1220 926 1288 932
rect 1220 912 1274 926
tri 1274 912 1288 926 nw
tri 1188 900 1200 912 se
rect 1200 900 1262 912
tri 1262 900 1274 912 nw
tri 1181 893 1188 900 se
rect 1188 893 1253 900
rect 1132 891 1253 893
tri 1253 891 1262 900 nw
rect 1132 887 1231 891
rect 1184 835 1231 887
tri 1231 869 1253 891 nw
rect 1132 823 1231 835
rect 1184 771 1231 823
rect 1132 765 1231 771
rect 1529 794 1581 2128
rect 1637 1048 1689 2128
rect 1768 1385 1774 1437
rect 1826 1385 1838 1437
rect 1890 1385 1896 1437
rect 1637 984 1689 996
rect 1637 926 1689 932
rect 1764 1252 1816 1258
rect 1764 1188 1816 1200
rect 1529 742 1535 794
rect 1587 742 1599 794
rect 1651 742 1657 794
rect 1764 714 1816 1136
rect 1041 708 1642 714
rect 1093 662 1642 708
rect 1694 662 1706 714
rect 1758 662 1816 714
rect 1844 964 1896 1385
rect 1844 900 1896 912
rect 1041 644 1093 656
rect 1041 586 1093 592
rect 1844 558 1896 848
rect 1636 506 1642 558
rect 1694 506 1706 558
rect 1758 506 1896 558
rect 1924 476 1976 2120
rect 219 403 225 455
rect 277 403 293 455
rect 345 403 361 455
rect 413 449 1439 455
rect 413 403 1276 449
rect 219 397 1276 403
rect 1328 397 1386 449
rect 1438 397 1439 449
rect 1848 424 1854 476
rect 1906 424 1918 476
rect 1970 424 1976 476
rect 219 381 1439 397
rect 219 329 225 381
rect 277 329 293 381
rect 345 329 361 381
rect 413 329 1276 381
rect 1328 329 1386 381
rect 1438 329 1439 381
rect 219 313 1439 329
rect 219 307 1276 313
rect 219 255 225 307
rect 277 255 293 307
rect 345 255 361 307
rect 413 261 1276 307
rect 1328 261 1386 313
rect 1438 261 1439 313
rect 413 255 1439 261
use sky130_fd_pr__nfet_01v8__example_55959141808478  sky130_fd_pr__nfet_01v8__example_55959141808478_0
timestamp 1644511149
transform 0 1 1390 -1 0 581
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808478  sky130_fd_pr__nfet_01v8__example_55959141808478_1
timestamp 1644511149
transform 0 1 1390 1 0 637
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808478  sky130_fd_pr__nfet_01v8__example_55959141808478_2
timestamp 1644511149
transform 0 1 1390 1 0 905
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808479  sky130_fd_pr__nfet_01v8__example_55959141808479_0
timestamp 1644511149
transform 0 -1 1093 -1 0 1627
box -28 0 128 267
use sky130_fd_pr__nfet_01v8__example_55959141808480  sky130_fd_pr__nfet_01v8__example_55959141808480_0
timestamp 1644511149
transform 0 -1 1093 1 0 949
box -28 0 440 267
use sky130_fd_pr__nfet_01v8__example_55959141808480  sky130_fd_pr__nfet_01v8__example_55959141808480_1
timestamp 1644511149
transform 0 -1 1093 -1 0 893
box -28 0 440 267
use sky130_fd_pr__pfet_01v8__example_55959141808475  sky130_fd_pr__pfet_01v8__example_55959141808475_0
timestamp 1644511149
transform 0 -1 2104 -1 0 581
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808475  sky130_fd_pr__pfet_01v8__example_55959141808475_1
timestamp 1644511149
transform 0 -1 2104 1 0 637
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_0
timestamp 1644511149
transform 0 -1 2013 -1 0 1463
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_1
timestamp 1644511149
transform 0 1 1486 1 0 1263
box -28 0 228 29
<< labels >>
flabel metal1 s 2072 965 2299 1399 3 FreeSans 520 0 0 0 VPWR_HV
port 1 nsew
flabel metal1 s 235 1266 338 1612 3 FreeSans 520 0 0 0 VGND
port 2 nsew
flabel metal2 s 1646 2072 1681 2121 3 FreeSans 520 0 0 0 RST_H
port 3 nsew
flabel metal2 s 1536 2066 1566 2125 3 FreeSans 520 90 0 0 OUT_H
port 4 nsew
flabel metal2 s 1931 2074 1970 2114 3 FreeSans 520 0 0 0 OUT_H_N
port 5 nsew
flabel metal2 s 1352 2062 1390 2118 3 FreeSans 520 90 0 0 IN
port 6 nsew
flabel metal2 s 1250 2055 1284 2118 3 FreeSans 520 90 0 0 IN_B
port 7 nsew
flabel metal2 s 1137 2062 1179 2118 3 FreeSans 520 90 0 0 HLD_H
port 8 nsew
flabel comment s 329 1121 329 1121 0 FreeSans 440 270 0 0 CONDIODE
<< properties >>
string GDS_END 48764816
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48723036
<< end >>
