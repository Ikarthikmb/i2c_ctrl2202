magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< metal2 >>
rect -6231 23152 -1085 23500
rect -6231 22896 -6130 23152
rect -5874 22896 -5606 23152
rect -5350 22896 -5052 23152
rect -4796 22896 -4498 23152
rect -4242 22896 -3944 23152
rect -3688 22896 -3390 23152
rect -3134 22896 -2836 23152
rect -2580 22896 -2312 23152
rect -2056 22896 -1085 23152
rect -6231 22628 -1085 22896
rect -6231 22372 -6130 22628
rect -5874 22372 -5606 22628
rect -5350 22372 -5052 22628
rect -4796 22372 -4498 22628
rect -4242 22372 -3944 22628
rect -3688 22372 -3390 22628
rect -3134 22372 -2836 22628
rect -2580 22372 -2312 22628
rect -2056 22372 -1085 22628
rect -6231 22104 -1085 22372
rect -6231 21848 -6130 22104
rect -5874 21848 -5606 22104
rect -5350 21848 -5052 22104
rect -4796 21848 -4498 22104
rect -4242 21848 -3944 22104
rect -3688 21848 -3390 22104
rect -3134 21848 -2836 22104
rect -2580 21848 -2312 22104
rect -2056 21848 -1085 22104
rect -6231 21500 -1085 21848
tri -1085 21500 915 23500 sw
tri -1915 21330 -1745 21500 ne
rect -1745 21330 915 21500
tri 915 21330 1085 21500 sw
tri -1745 18500 1085 21330 ne
tri 1085 20500 1915 21330 sw
rect 1085 20151 6008 20500
rect 1085 19895 1833 20151
rect 2089 19895 2357 20151
rect 2613 19895 2911 20151
rect 3167 19895 3465 20151
rect 3721 19895 4019 20151
rect 4275 19895 4573 20151
rect 4829 19895 5127 20151
rect 5383 19895 5651 20151
rect 5907 19895 6008 20151
rect 1085 19627 6008 19895
rect 1085 19371 1833 19627
rect 2089 19371 2357 19627
rect 2613 19371 2911 19627
rect 3167 19371 3465 19627
rect 3721 19371 4019 19627
rect 4275 19371 4573 19627
rect 4829 19371 5127 19627
rect 5383 19371 5651 19627
rect 5907 19371 6008 19627
rect 1085 19103 6008 19371
rect 1085 18847 1833 19103
rect 2089 18847 2357 19103
rect 2613 18847 2911 19103
rect 3167 18847 3465 19103
rect 3721 18847 4019 19103
rect 4275 18847 4573 19103
rect 4829 18847 5127 19103
rect 5383 18847 5651 19103
rect 5907 18847 6008 19103
rect 1085 18500 6008 18847
rect -6231 17153 -1085 17500
rect -6231 16897 -6131 17153
rect -5875 16897 -5607 17153
rect -5351 16897 -5053 17153
rect -4797 16897 -4499 17153
rect -4243 16897 -3945 17153
rect -3689 16897 -3391 17153
rect -3135 16897 -2837 17153
rect -2581 16897 -2313 17153
rect -2057 16897 -1085 17153
rect -6231 16629 -1085 16897
rect -6231 16373 -6131 16629
rect -5875 16373 -5607 16629
rect -5351 16373 -5053 16629
rect -4797 16373 -4499 16629
rect -4243 16373 -3945 16629
rect -3689 16373 -3391 16629
rect -3135 16373 -2837 16629
rect -2581 16373 -2313 16629
rect -2057 16373 -1085 16629
rect -6231 16105 -1085 16373
rect -6231 15849 -6131 16105
rect -5875 15849 -5607 16105
rect -5351 15849 -5053 16105
rect -4797 15849 -4499 16105
rect -4243 15849 -3945 16105
rect -3689 15849 -3391 16105
rect -3135 15849 -2837 16105
rect -2581 15849 -2313 16105
rect -2057 15849 -1085 16105
rect -6231 15500 -1085 15849
tri -1085 15500 915 17500 sw
tri -1915 15330 -1745 15500 ne
rect -1745 15330 915 15500
tri 915 15330 1085 15500 sw
tri -1745 12500 1085 15330 ne
tri 1085 14500 1915 15330 sw
rect 1085 14153 6008 14500
rect 1085 13897 1833 14153
rect 2089 13897 2357 14153
rect 2613 13897 2911 14153
rect 3167 13897 3465 14153
rect 3721 13897 4019 14153
rect 4275 13897 4573 14153
rect 4829 13897 5127 14153
rect 5383 13897 5651 14153
rect 5907 13897 6008 14153
rect 1085 13629 6008 13897
rect 1085 13373 1833 13629
rect 2089 13373 2357 13629
rect 2613 13373 2911 13629
rect 3167 13373 3465 13629
rect 3721 13373 4019 13629
rect 4275 13373 4573 13629
rect 4829 13373 5127 13629
rect 5383 13373 5651 13629
rect 5907 13373 6008 13629
rect 1085 13105 6008 13373
rect 1085 12849 1833 13105
rect 2089 12849 2357 13105
rect 2613 12849 2911 13105
rect 3167 12849 3465 13105
rect 3721 12849 4019 13105
rect 4275 12849 4573 13105
rect 4829 12849 5127 13105
rect 5383 12849 5651 13105
rect 5907 12849 6008 13105
rect 1085 12500 6008 12849
rect 9908 652 27500 1000
rect 9908 396 10052 652
rect 10308 396 10576 652
rect 10832 396 11130 652
rect 11386 396 27500 652
rect 9908 128 27500 396
rect 9908 -128 10052 128
rect 10308 -128 10576 128
rect 10832 -128 11130 128
rect 11386 -128 27500 128
rect 9908 -396 27500 -128
rect 9908 -652 10052 -396
rect 10308 -652 10576 -396
rect 10832 -652 11130 -396
rect 11386 -652 27500 -396
rect 9908 -1000 27500 -652
tri -1745 -18330 1085 -15500 se
rect 1085 -15849 6008 -15500
rect 1085 -16105 1832 -15849
rect 2088 -16105 2356 -15849
rect 2612 -16105 2910 -15849
rect 3166 -16105 3464 -15849
rect 3720 -16105 4018 -15849
rect 4274 -16105 4572 -15849
rect 4828 -16105 5126 -15849
rect 5382 -16105 5650 -15849
rect 5906 -16105 6008 -15849
rect 1085 -16373 6008 -16105
rect 1085 -16629 1832 -16373
rect 2088 -16629 2356 -16373
rect 2612 -16629 2910 -16373
rect 3166 -16629 3464 -16373
rect 3720 -16629 4018 -16373
rect 4274 -16629 4572 -16373
rect 4828 -16629 5126 -16373
rect 5382 -16629 5650 -16373
rect 5906 -16629 6008 -16373
rect 1085 -16897 6008 -16629
rect 1085 -17153 1832 -16897
rect 2088 -17153 2356 -16897
rect 2612 -17153 2910 -16897
rect 3166 -17153 3464 -16897
rect 3720 -17153 4018 -16897
rect 4274 -17153 4572 -16897
rect 4828 -17153 5126 -16897
rect 5382 -17153 5650 -16897
rect 5906 -17153 6008 -16897
rect 1085 -17500 6008 -17153
tri 1085 -18330 1915 -17500 nw
tri -1915 -18500 -1745 -18330 se
rect -1745 -18500 915 -18330
tri 915 -18500 1085 -18330 nw
rect -6231 -18848 -1085 -18500
rect -6231 -19104 -6130 -18848
rect -5874 -19104 -5606 -18848
rect -5350 -19104 -5052 -18848
rect -4796 -19104 -4498 -18848
rect -4242 -19104 -3944 -18848
rect -3688 -19104 -3390 -18848
rect -3134 -19104 -2836 -18848
rect -2580 -19104 -2312 -18848
rect -2056 -19104 -1085 -18848
rect -6231 -19372 -1085 -19104
rect -6231 -19628 -6130 -19372
rect -5874 -19628 -5606 -19372
rect -5350 -19628 -5052 -19372
rect -4796 -19628 -4498 -19372
rect -4242 -19628 -3944 -19372
rect -3688 -19628 -3390 -19372
rect -3134 -19628 -2836 -19372
rect -2580 -19628 -2312 -19372
rect -2056 -19628 -1085 -19372
rect -6231 -19896 -1085 -19628
rect -6231 -20152 -6130 -19896
rect -5874 -20152 -5606 -19896
rect -5350 -20152 -5052 -19896
rect -4796 -20152 -4498 -19896
rect -4242 -20152 -3944 -19896
rect -3688 -20152 -3390 -19896
rect -3134 -20152 -2836 -19896
rect -2580 -20152 -2312 -19896
rect -2056 -20152 -1085 -19896
rect -6231 -20500 -1085 -20152
tri -1085 -20500 915 -18500 nw
tri -1745 -24330 1085 -21500 se
rect 1085 -21848 6008 -21500
rect 1085 -22104 1833 -21848
rect 2089 -22104 2357 -21848
rect 2613 -22104 2911 -21848
rect 3167 -22104 3465 -21848
rect 3721 -22104 4019 -21848
rect 4275 -22104 4573 -21848
rect 4829 -22104 5127 -21848
rect 5383 -22104 5651 -21848
rect 5907 -22104 6008 -21848
rect 1085 -22372 6008 -22104
rect 1085 -22628 1833 -22372
rect 2089 -22628 2357 -22372
rect 2613 -22628 2911 -22372
rect 3167 -22628 3465 -22372
rect 3721 -22628 4019 -22372
rect 4275 -22628 4573 -22372
rect 4829 -22628 5127 -22372
rect 5383 -22628 5651 -22372
rect 5907 -22628 6008 -22372
rect 1085 -22896 6008 -22628
rect 1085 -23152 1833 -22896
rect 2089 -23152 2357 -22896
rect 2613 -23152 2911 -22896
rect 3167 -23152 3465 -22896
rect 3721 -23152 4019 -22896
rect 4275 -23152 4573 -22896
rect 4829 -23152 5127 -22896
rect 5383 -23152 5651 -22896
rect 5907 -23152 6008 -22896
rect 1085 -23500 6008 -23152
tri 1085 -24330 1915 -23500 nw
tri -1915 -24500 -1745 -24330 se
rect -1745 -24500 915 -24330
tri 915 -24500 1085 -24330 nw
rect -6231 -24848 -1085 -24500
rect -6231 -25104 -6130 -24848
rect -5874 -25104 -5606 -24848
rect -5350 -25104 -5052 -24848
rect -4796 -25104 -4498 -24848
rect -4242 -25104 -3944 -24848
rect -3688 -25104 -3390 -24848
rect -3134 -25104 -2836 -24848
rect -2580 -25104 -2312 -24848
rect -2056 -25104 -1085 -24848
rect -6231 -25372 -1085 -25104
rect -6231 -25628 -6130 -25372
rect -5874 -25628 -5606 -25372
rect -5350 -25628 -5052 -25372
rect -4796 -25628 -4498 -25372
rect -4242 -25628 -3944 -25372
rect -3688 -25628 -3390 -25372
rect -3134 -25628 -2836 -25372
rect -2580 -25628 -2312 -25372
rect -2056 -25628 -1085 -25372
rect -6231 -25896 -1085 -25628
rect -6231 -26152 -6130 -25896
rect -5874 -26152 -5606 -25896
rect -5350 -26152 -5052 -25896
rect -4796 -26152 -4498 -25896
rect -4242 -26152 -3944 -25896
rect -3688 -26152 -3390 -25896
rect -3134 -26152 -2836 -25896
rect -2580 -26152 -2312 -25896
rect -2056 -26152 -1085 -25896
rect -6231 -26500 -1085 -26152
tri -1085 -26500 915 -24500 nw
<< via2 >>
rect -6130 22896 -5874 23152
rect -5606 22896 -5350 23152
rect -5052 22896 -4796 23152
rect -4498 22896 -4242 23152
rect -3944 22896 -3688 23152
rect -3390 22896 -3134 23152
rect -2836 22896 -2580 23152
rect -2312 22896 -2056 23152
rect -6130 22372 -5874 22628
rect -5606 22372 -5350 22628
rect -5052 22372 -4796 22628
rect -4498 22372 -4242 22628
rect -3944 22372 -3688 22628
rect -3390 22372 -3134 22628
rect -2836 22372 -2580 22628
rect -2312 22372 -2056 22628
rect -6130 21848 -5874 22104
rect -5606 21848 -5350 22104
rect -5052 21848 -4796 22104
rect -4498 21848 -4242 22104
rect -3944 21848 -3688 22104
rect -3390 21848 -3134 22104
rect -2836 21848 -2580 22104
rect -2312 21848 -2056 22104
rect 1833 19895 2089 20151
rect 2357 19895 2613 20151
rect 2911 19895 3167 20151
rect 3465 19895 3721 20151
rect 4019 19895 4275 20151
rect 4573 19895 4829 20151
rect 5127 19895 5383 20151
rect 5651 19895 5907 20151
rect 1833 19371 2089 19627
rect 2357 19371 2613 19627
rect 2911 19371 3167 19627
rect 3465 19371 3721 19627
rect 4019 19371 4275 19627
rect 4573 19371 4829 19627
rect 5127 19371 5383 19627
rect 5651 19371 5907 19627
rect 1833 18847 2089 19103
rect 2357 18847 2613 19103
rect 2911 18847 3167 19103
rect 3465 18847 3721 19103
rect 4019 18847 4275 19103
rect 4573 18847 4829 19103
rect 5127 18847 5383 19103
rect 5651 18847 5907 19103
rect -6131 16897 -5875 17153
rect -5607 16897 -5351 17153
rect -5053 16897 -4797 17153
rect -4499 16897 -4243 17153
rect -3945 16897 -3689 17153
rect -3391 16897 -3135 17153
rect -2837 16897 -2581 17153
rect -2313 16897 -2057 17153
rect -6131 16373 -5875 16629
rect -5607 16373 -5351 16629
rect -5053 16373 -4797 16629
rect -4499 16373 -4243 16629
rect -3945 16373 -3689 16629
rect -3391 16373 -3135 16629
rect -2837 16373 -2581 16629
rect -2313 16373 -2057 16629
rect -6131 15849 -5875 16105
rect -5607 15849 -5351 16105
rect -5053 15849 -4797 16105
rect -4499 15849 -4243 16105
rect -3945 15849 -3689 16105
rect -3391 15849 -3135 16105
rect -2837 15849 -2581 16105
rect -2313 15849 -2057 16105
rect 1833 13897 2089 14153
rect 2357 13897 2613 14153
rect 2911 13897 3167 14153
rect 3465 13897 3721 14153
rect 4019 13897 4275 14153
rect 4573 13897 4829 14153
rect 5127 13897 5383 14153
rect 5651 13897 5907 14153
rect 1833 13373 2089 13629
rect 2357 13373 2613 13629
rect 2911 13373 3167 13629
rect 3465 13373 3721 13629
rect 4019 13373 4275 13629
rect 4573 13373 4829 13629
rect 5127 13373 5383 13629
rect 5651 13373 5907 13629
rect 1833 12849 2089 13105
rect 2357 12849 2613 13105
rect 2911 12849 3167 13105
rect 3465 12849 3721 13105
rect 4019 12849 4275 13105
rect 4573 12849 4829 13105
rect 5127 12849 5383 13105
rect 5651 12849 5907 13105
rect 10052 396 10308 652
rect 10576 396 10832 652
rect 11130 396 11386 652
rect 10052 -128 10308 128
rect 10576 -128 10832 128
rect 11130 -128 11386 128
rect 10052 -652 10308 -396
rect 10576 -652 10832 -396
rect 11130 -652 11386 -396
rect 1832 -16105 2088 -15849
rect 2356 -16105 2612 -15849
rect 2910 -16105 3166 -15849
rect 3464 -16105 3720 -15849
rect 4018 -16105 4274 -15849
rect 4572 -16105 4828 -15849
rect 5126 -16105 5382 -15849
rect 5650 -16105 5906 -15849
rect 1832 -16629 2088 -16373
rect 2356 -16629 2612 -16373
rect 2910 -16629 3166 -16373
rect 3464 -16629 3720 -16373
rect 4018 -16629 4274 -16373
rect 4572 -16629 4828 -16373
rect 5126 -16629 5382 -16373
rect 5650 -16629 5906 -16373
rect 1832 -17153 2088 -16897
rect 2356 -17153 2612 -16897
rect 2910 -17153 3166 -16897
rect 3464 -17153 3720 -16897
rect 4018 -17153 4274 -16897
rect 4572 -17153 4828 -16897
rect 5126 -17153 5382 -16897
rect 5650 -17153 5906 -16897
rect -6130 -19104 -5874 -18848
rect -5606 -19104 -5350 -18848
rect -5052 -19104 -4796 -18848
rect -4498 -19104 -4242 -18848
rect -3944 -19104 -3688 -18848
rect -3390 -19104 -3134 -18848
rect -2836 -19104 -2580 -18848
rect -2312 -19104 -2056 -18848
rect -6130 -19628 -5874 -19372
rect -5606 -19628 -5350 -19372
rect -5052 -19628 -4796 -19372
rect -4498 -19628 -4242 -19372
rect -3944 -19628 -3688 -19372
rect -3390 -19628 -3134 -19372
rect -2836 -19628 -2580 -19372
rect -2312 -19628 -2056 -19372
rect -6130 -20152 -5874 -19896
rect -5606 -20152 -5350 -19896
rect -5052 -20152 -4796 -19896
rect -4498 -20152 -4242 -19896
rect -3944 -20152 -3688 -19896
rect -3390 -20152 -3134 -19896
rect -2836 -20152 -2580 -19896
rect -2312 -20152 -2056 -19896
rect 1833 -22104 2089 -21848
rect 2357 -22104 2613 -21848
rect 2911 -22104 3167 -21848
rect 3465 -22104 3721 -21848
rect 4019 -22104 4275 -21848
rect 4573 -22104 4829 -21848
rect 5127 -22104 5383 -21848
rect 5651 -22104 5907 -21848
rect 1833 -22628 2089 -22372
rect 2357 -22628 2613 -22372
rect 2911 -22628 3167 -22372
rect 3465 -22628 3721 -22372
rect 4019 -22628 4275 -22372
rect 4573 -22628 4829 -22372
rect 5127 -22628 5383 -22372
rect 5651 -22628 5907 -22372
rect 1833 -23152 2089 -22896
rect 2357 -23152 2613 -22896
rect 2911 -23152 3167 -22896
rect 3465 -23152 3721 -22896
rect 4019 -23152 4275 -22896
rect 4573 -23152 4829 -22896
rect 5127 -23152 5383 -22896
rect 5651 -23152 5907 -22896
rect -6130 -25104 -5874 -24848
rect -5606 -25104 -5350 -24848
rect -5052 -25104 -4796 -24848
rect -4498 -25104 -4242 -24848
rect -3944 -25104 -3688 -24848
rect -3390 -25104 -3134 -24848
rect -2836 -25104 -2580 -24848
rect -2312 -25104 -2056 -24848
rect -6130 -25628 -5874 -25372
rect -5606 -25628 -5350 -25372
rect -5052 -25628 -4796 -25372
rect -4498 -25628 -4242 -25372
rect -3944 -25628 -3688 -25372
rect -3390 -25628 -3134 -25372
rect -2836 -25628 -2580 -25372
rect -2312 -25628 -2056 -25372
rect -6130 -26152 -5874 -25896
rect -5606 -26152 -5350 -25896
rect -5052 -26152 -4796 -25896
rect -4498 -26152 -4242 -25896
rect -3944 -26152 -3688 -25896
rect -3390 -26152 -3134 -25896
rect -2836 -26152 -2580 -25896
rect -2312 -26152 -2056 -25896
<< metal3 >>
tri -12978 24500 -10978 26500 se
rect -10978 25118 10978 26500
tri 10978 25118 12360 26500 sw
rect -10978 24500 12360 25118
tri 12360 24500 12978 25118 sw
tri -13806 23672 -12978 24500 se
rect -12978 23672 -10978 24500
tri -10978 23672 -10150 24500 nw
tri 10150 23672 10978 24500 ne
rect 10978 23672 12978 24500
tri -14326 23152 -13806 23672 se
rect -13806 23500 -11150 23672
tri -11150 23500 -10978 23672 nw
tri 10978 23500 11150 23672 ne
rect 11150 23500 12978 23672
rect -13806 23152 -11498 23500
tri -11498 23152 -11150 23500 nw
tri -10084 23152 -9736 23500 se
rect -9736 23253 -2202 23500
tri -2202 23253 -1955 23500 sw
rect -9736 23152 -1955 23253
tri -14582 22896 -14326 23152 se
rect -14326 22896 -11754 23152
tri -11754 22896 -11498 23152 nw
tri -10340 22896 -10084 23152 se
rect -10084 22896 -6130 23152
rect -5874 22896 -5606 23152
rect -5350 22896 -5052 23152
rect -4796 22896 -4498 23152
rect -4242 22896 -3944 23152
rect -3688 22896 -3390 23152
rect -3134 22896 -2836 23152
rect -2580 22896 -2312 23152
rect -2056 22896 -1955 23152
tri -14850 22628 -14582 22896 se
rect -14582 22628 -12022 22896
tri -12022 22628 -11754 22896 nw
tri -10608 22628 -10340 22896 se
rect -10340 22628 -1955 22896
tri -15106 22372 -14850 22628 se
rect -14850 22372 -12278 22628
tri -12278 22372 -12022 22628 nw
tri -10864 22372 -10608 22628 se
rect -10608 22372 -6130 22628
rect -5874 22372 -5606 22628
rect -5350 22372 -5052 22628
rect -4796 22372 -4498 22628
rect -4242 22372 -3944 22628
rect -3688 22372 -3390 22628
rect -3134 22372 -2836 22628
rect -2580 22372 -2312 22628
rect -2056 22372 -1955 22628
tri -15188 22290 -15106 22372 se
rect -15106 22290 -12360 22372
tri -12360 22290 -12278 22372 nw
tri -10946 22290 -10864 22372 se
rect -10864 22290 -1955 22372
tri -125 22290 1085 23500 se
rect 1085 22462 9736 23500
tri 9736 22462 10774 23500 sw
tri 11150 22462 12188 23500 ne
rect 12188 22462 12978 23500
rect 1085 22290 10774 22462
tri 10774 22290 10946 22462 sw
tri 12188 22290 12360 22462 ne
rect 12360 22290 12978 22462
tri 12978 22290 15188 24500 sw
tri -15374 22104 -15188 22290 se
rect -15188 22104 -12546 22290
tri -12546 22104 -12360 22290 nw
tri -11132 22104 -10946 22290 se
rect -10946 22104 -1955 22290
tri -15630 21848 -15374 22104 se
rect -15374 22086 -12564 22104
tri -12564 22086 -12546 22104 nw
tri -11150 22086 -11132 22104 se
rect -11132 22086 -6130 22104
rect -15374 21848 -12802 22086
tri -12802 21848 -12564 22086 nw
tri -11388 21848 -11150 22086 se
rect -11150 21848 -6130 22086
rect -5874 21848 -5606 22104
rect -5350 21848 -5052 22104
rect -4796 21848 -4498 22104
rect -4242 21848 -3944 22104
rect -3688 21848 -3390 22104
rect -3134 21848 -2836 22104
rect -2580 21848 -2312 22104
rect -2056 21848 -1955 22104
tri -16634 20844 -15630 21848 se
rect -15630 20844 -13806 21848
tri -13806 20844 -12802 21848 nw
tri -12188 21048 -11388 21848 se
rect -11388 21747 -1955 21848
rect -11388 21500 -2202 21747
tri -2202 21500 -1955 21747 nw
tri -915 21500 -125 22290 se
rect -125 21500 10946 22290
rect -11388 21048 -9360 21500
tri -9360 21048 -8908 21500 nw
tri -1367 21048 -915 21500 se
rect -915 21048 1463 21500
tri 1463 21048 1915 21500 nw
tri 8908 21048 9360 21500 ne
rect 9360 21048 10946 21500
tri 10946 21048 12188 22290 sw
tri 12360 21048 13602 22290 ne
rect 13602 21048 15188 22290
tri -12392 20844 -12188 21048 se
rect -12188 20844 -9564 21048
tri -9564 20844 -9360 21048 nw
tri -1571 20844 -1367 21048 se
rect -1367 20844 1259 21048
tri 1259 20844 1463 21048 nw
tri 9360 20844 9564 21048 ne
rect 9564 20844 12188 21048
tri 12188 20844 12392 21048 sw
tri 13602 20844 13806 21048 ne
rect 13806 20844 15188 21048
tri -17327 20151 -16634 20844 se
rect -16634 20672 -13978 20844
tri -13978 20672 -13806 20844 nw
tri -12564 20672 -12392 20844 se
rect -12392 20672 -9736 20844
tri -9736 20672 -9564 20844 nw
tri -1743 20672 -1571 20844 se
rect -1571 20672 1087 20844
tri 1087 20672 1259 20844 nw
tri 9564 20672 9736 20844 ne
rect 9736 20672 12392 20844
rect -16634 20151 -14499 20672
tri -14499 20151 -13978 20672 nw
tri -13085 20151 -12564 20672 se
rect -12564 20500 -9908 20672
tri -9908 20500 -9736 20672 nw
tri -1745 20670 -1743 20672 se
rect -1743 20670 1085 20672
tri 1085 20670 1087 20672 nw
tri 9736 20670 9738 20672 ne
rect 9738 20670 12392 20672
tri -1915 20500 -1745 20670 se
rect -1745 20500 915 20670
tri 915 20500 1085 20670 nw
tri 9738 20500 9908 20670 ne
rect 9908 20500 12392 20670
rect -12564 20151 -10257 20500
tri -10257 20151 -9908 20500 nw
tri -8842 20151 -8493 20500 se
rect -8493 20151 566 20500
tri 566 20151 915 20500 nw
tri 1732 20253 1979 20500 se
rect 1979 20253 8493 20500
rect 1732 20151 8493 20253
tri -17583 19895 -17327 20151 se
rect -17327 19895 -14755 20151
tri -14755 19895 -14499 20151 nw
tri -13341 19895 -13085 20151 se
rect -13085 19895 -10513 20151
tri -10513 19895 -10257 20151 nw
tri -9098 19895 -8842 20151 se
rect -8842 19895 310 20151
tri 310 19895 566 20151 nw
rect 1732 19895 1833 20151
rect 2089 19895 2357 20151
rect 2613 19895 2911 20151
rect 3167 19895 3465 20151
rect 3721 19895 4019 20151
rect 4275 19895 4573 20151
rect 4829 19895 5127 20151
rect 5383 19895 5651 20151
rect 5907 19895 8493 20151
tri -17851 19627 -17583 19895 se
rect -17583 19627 -15023 19895
tri -15023 19627 -14755 19895 nw
tri -13609 19627 -13341 19895 se
rect -13341 19627 -10781 19895
tri -10781 19627 -10513 19895 nw
tri -9188 19805 -9098 19895 se
rect -9098 19805 220 19895
tri 220 19805 310 19895 nw
rect 1732 19805 8493 19895
tri 8493 19805 9188 20500 sw
tri 9908 19805 10603 20500 ne
rect 10603 19805 12392 20500
tri -9366 19627 -9188 19805 se
rect -9188 19627 42 19805
tri 42 19627 220 19805 nw
rect 1732 19627 9188 19805
tri -18016 19462 -17851 19627 se
rect -17851 19462 -15188 19627
tri -15188 19462 -15023 19627 nw
tri -13774 19462 -13609 19627 se
rect -13609 19462 -10946 19627
tri -10946 19462 -10781 19627 nw
tri -9531 19462 -9366 19627 se
rect -9366 19462 -123 19627
tri -123 19462 42 19627 nw
tri -18107 19371 -18016 19462 se
rect -18016 19371 -15279 19462
tri -15279 19371 -15188 19462 nw
tri -13865 19371 -13774 19462 se
rect -13774 19371 -11037 19462
tri -11037 19371 -10946 19462 nw
tri -9622 19371 -9531 19462 se
rect -9531 19371 -214 19462
tri -214 19371 -123 19462 nw
rect 1732 19371 1833 19627
rect 2089 19371 2357 19627
rect 2613 19371 2911 19627
rect 3167 19371 3465 19627
rect 3721 19371 4019 19627
rect 4275 19371 4573 19627
rect 4829 19371 5127 19627
rect 5383 19371 5651 19627
rect 5907 19462 9188 19627
tri 9188 19462 9531 19805 sw
tri 10603 19462 10946 19805 ne
rect 10946 19634 12392 19805
tri 12392 19634 13602 20844 sw
tri 13806 19634 15016 20844 ne
rect 15016 19634 15188 20844
rect 10946 19462 13602 19634
tri 13602 19462 13774 19634 sw
tri 15016 19462 15188 19634 ne
tri 15188 19462 18016 22290 sw
rect 5907 19371 9531 19462
tri -18375 19103 -18107 19371 se
rect -18107 19258 -15392 19371
tri -15392 19258 -15279 19371 nw
tri -13978 19258 -13865 19371 se
rect -13865 19258 -11305 19371
rect -18107 19103 -15547 19258
tri -15547 19103 -15392 19258 nw
tri -14133 19103 -13978 19258 se
rect -13978 19103 -11305 19258
tri -11305 19103 -11037 19371 nw
tri -9890 19103 -9622 19371 se
rect -9622 19103 -482 19371
tri -482 19103 -214 19371 nw
rect 1732 19103 9531 19371
tri -18631 18847 -18375 19103 se
rect -18375 18847 -15803 19103
tri -15803 18847 -15547 19103 nw
tri -14389 18847 -14133 19103 se
rect -14133 19087 -11321 19103
tri -11321 19087 -11305 19103 nw
tri -9906 19087 -9890 19103 se
rect -9890 19087 -738 19103
rect -14133 18847 -11561 19087
tri -11561 18847 -11321 19087 nw
tri -10146 18847 -9906 19087 se
rect -9906 18847 -738 19087
tri -738 18847 -482 19103 nw
rect 1732 18847 1833 19103
rect 2089 18847 2357 19103
rect 2613 18847 2911 19103
rect 3167 18847 3465 19103
rect 3721 18847 4019 19103
rect 4275 18847 4573 19103
rect 4829 18847 5127 19103
rect 5383 18847 5651 19103
rect 5907 18847 9531 19103
tri -19462 18016 -18631 18847 se
rect -18631 18016 -16634 18847
tri -16634 18016 -15803 18847 nw
tri -15016 18220 -14389 18847 se
rect -14389 18220 -12188 18847
tri -12188 18220 -11561 18847 nw
tri -10773 18220 -10146 18847 se
rect -10146 18500 -1085 18847
tri -1085 18500 -738 18847 nw
rect 1732 18747 9531 18847
tri 1732 18500 1979 18747 ne
rect 1979 18500 9531 18747
rect -10146 18220 -7945 18500
tri -7945 18220 -7665 18500 nw
tri 7665 18220 7945 18500 ne
rect 7945 18392 9531 18500
tri 9531 18392 10601 19462 sw
tri 10946 18392 12016 19462 ne
rect 12016 18392 13774 19462
rect 7945 18220 10601 18392
tri 10601 18220 10773 18392 sw
tri 12016 18220 12188 18392 ne
rect 12188 18220 13774 18392
tri 13774 18220 15016 19462 sw
tri 15188 18220 16430 19462 ne
rect 16430 18220 18016 19462
tri -15220 18016 -15016 18220 se
rect -15016 18016 -12392 18220
tri -12392 18016 -12188 18220 nw
tri -10977 18016 -10773 18220 se
rect -10773 18016 -8149 18220
tri -8149 18016 -7945 18220 nw
tri 7945 18016 8149 18220 ne
rect 8149 18016 10773 18220
tri 10773 18016 10977 18220 sw
tri 12188 18016 12392 18220 ne
rect 12392 18016 15016 18220
tri 15016 18016 15220 18220 sw
tri 16430 18016 16634 18220 ne
rect 16634 18016 18016 18220
tri -20325 17153 -19462 18016 se
rect -19462 17844 -16806 18016
tri -16806 17844 -16634 18016 nw
tri -15392 17844 -15220 18016 se
rect -15220 17844 -12564 18016
tri -12564 17844 -12392 18016 nw
tri -11149 17844 -10977 18016 se
rect -10977 17844 -8321 18016
tri -8321 17844 -8149 18016 nw
tri 8149 17844 8321 18016 ne
rect 8321 17844 10977 18016
tri 10977 17844 11149 18016 sw
tri 12392 17844 12564 18016 ne
rect 12564 17844 15220 18016
rect -19462 17153 -17497 17844
tri -17497 17153 -16806 17844 nw
tri -16083 17153 -15392 17844 se
rect -15392 17672 -12736 17844
tri -12736 17672 -12564 17844 nw
tri -11321 17672 -11149 17844 se
rect -11149 17672 -8493 17844
tri -8493 17672 -8321 17844 nw
tri 8321 17672 8493 17844 ne
rect 8493 17672 11149 17844
rect -15392 17153 -13255 17672
tri -13255 17153 -12736 17672 nw
tri -11840 17153 -11321 17672 se
rect -11321 17500 -8665 17672
tri -8665 17500 -8493 17672 nw
tri 8493 17500 8665 17672 ne
rect 8665 17500 11149 17672
rect -11321 17153 -9012 17500
tri -9012 17153 -8665 17500 nw
tri -7598 17153 -7251 17500 se
rect -7251 17253 -2202 17500
tri -2202 17253 -1955 17500 sw
rect -7251 17153 -1955 17253
tri -20581 16897 -20325 17153 se
rect -20325 16897 -17753 17153
tri -17753 16897 -17497 17153 nw
tri -16339 16897 -16083 17153 se
rect -16083 16897 -13511 17153
tri -13511 16897 -13255 17153 nw
tri -12016 16977 -11840 17153 se
rect -11840 16977 -9188 17153
tri -9188 16977 -9012 17153 nw
tri -7774 16977 -7598 17153 se
rect -7598 16977 -6131 17153
tri -12096 16897 -12016 16977 se
rect -12016 16897 -9268 16977
tri -9268 16897 -9188 16977 nw
tri -7854 16897 -7774 16977 se
rect -7774 16897 -6131 16977
rect -5875 16897 -5607 17153
rect -5351 16897 -5053 17153
rect -4797 16897 -4499 17153
rect -4243 16897 -3945 17153
rect -3689 16897 -3391 17153
rect -3135 16897 -2837 17153
rect -2581 16897 -2313 17153
rect -2057 16897 -1955 17153
tri 562 16977 1085 17500 se
rect 1085 17149 7251 17500
tri 7251 17149 7602 17500 sw
tri 8665 17149 9016 17500 ne
rect 9016 17149 11149 17500
rect 1085 16977 7602 17149
tri 7602 16977 7774 17149 sw
tri 9016 16977 9188 17149 ne
rect 9188 16977 11149 17149
tri 11149 16977 12016 17844 sw
tri 12564 16977 13431 17844 ne
rect 13431 16977 15220 17844
tri -20844 16634 -20581 16897 se
rect -20581 16634 -18016 16897
tri -18016 16634 -17753 16897 nw
tri -16602 16634 -16339 16897 se
rect -16339 16634 -13774 16897
tri -13774 16634 -13511 16897 nw
tri -12359 16634 -12096 16897 se
rect -12096 16634 -9531 16897
tri -9531 16634 -9268 16897 nw
tri -8117 16634 -7854 16897 se
rect -7854 16634 -1955 16897
tri 219 16634 562 16977 se
rect 562 16634 7774 16977
tri 7774 16634 8117 16977 sw
tri 9188 16634 9531 16977 ne
rect 9531 16634 12016 16977
tri 12016 16634 12359 16977 sw
tri 13431 16634 13774 16977 ne
rect 13774 16806 15220 16977
tri 15220 16806 16430 18016 sw
tri 16634 16806 17844 18016 ne
rect 17844 16806 18016 18016
rect 13774 16634 16430 16806
tri 16430 16634 16602 16806 sw
tri 17844 16634 18016 16806 ne
tri 18016 16634 20844 19462 sw
tri -20849 16629 -20844 16634 se
rect -20844 16629 -18021 16634
tri -18021 16629 -18016 16634 nw
tri -16607 16629 -16602 16634 se
rect -16602 16629 -13779 16634
tri -13779 16629 -13774 16634 nw
tri -12364 16629 -12359 16634 se
rect -12359 16629 -9536 16634
tri -9536 16629 -9531 16634 nw
tri -8122 16629 -8117 16634 se
rect -8117 16629 -1955 16634
tri -21105 16373 -20849 16629 se
rect -20849 16430 -18220 16629
tri -18220 16430 -18021 16629 nw
tri -16806 16430 -16607 16629 se
rect -16607 16430 -14035 16629
rect -20849 16373 -18277 16430
tri -18277 16373 -18220 16430 nw
tri -16863 16373 -16806 16430 se
rect -16806 16373 -14035 16430
tri -14035 16373 -13779 16629 nw
tri -12620 16373 -12364 16629 se
rect -12364 16373 -9792 16629
tri -9792 16373 -9536 16629 nw
tri -8378 16373 -8122 16629 se
rect -8122 16373 -6131 16629
rect -5875 16373 -5607 16629
rect -5351 16373 -5053 16629
rect -4797 16373 -4499 16629
rect -4243 16373 -3945 16629
rect -3689 16373 -3391 16629
rect -3135 16373 -2837 16629
rect -2581 16373 -2313 16629
rect -2057 16373 -1955 16629
tri -21373 16105 -21105 16373 se
rect -21105 16105 -18545 16373
tri -18545 16105 -18277 16373 nw
tri -17131 16105 -16863 16373 se
rect -16863 16259 -14149 16373
tri -14149 16259 -14035 16373 nw
tri -12734 16259 -12620 16373 se
rect -12620 16259 -10060 16373
rect -16863 16105 -14303 16259
tri -14303 16105 -14149 16259 nw
tri -12888 16105 -12734 16259 se
rect -12734 16105 -10060 16259
tri -10060 16105 -9792 16373 nw
tri -8646 16105 -8378 16373 se
rect -8378 16105 -1955 16373
tri -21629 15849 -21373 16105 se
rect -21373 15849 -18801 16105
tri -18801 15849 -18545 16105 nw
tri -17387 15849 -17131 16105 se
rect -17131 15849 -14559 16105
tri -14559 15849 -14303 16105 nw
tri -13144 15849 -12888 16105 se
rect -12888 16086 -10079 16105
tri -10079 16086 -10060 16105 nw
tri -8665 16086 -8646 16105 se
rect -8646 16086 -6131 16105
rect -12888 15849 -10316 16086
tri -10316 15849 -10079 16086 nw
tri -8902 15849 -8665 16086 se
rect -8665 15849 -6131 16086
rect -5875 15849 -5607 16105
rect -5351 15849 -5053 16105
rect -4797 15849 -4499 16105
rect -4243 15849 -3945 16105
rect -3689 15849 -3391 16105
rect -3135 15849 -2837 16105
rect -2581 15849 -2313 16105
rect -2057 15849 -1955 16105
tri -22290 15188 -21629 15849 se
rect -21629 15188 -19462 15849
tri -19462 15188 -18801 15849 nw
tri -17844 15392 -17387 15849 se
rect -17387 15392 -15016 15849
tri -15016 15392 -14559 15849 nw
tri -13601 15392 -13144 15849 se
rect -13144 15392 -10773 15849
tri -10773 15392 -10316 15849 nw
tri -9251 15500 -8902 15849 se
rect -8902 15747 -1955 15849
rect -8902 15735 -1967 15747
tri -1967 15735 -1955 15747 nw
tri -680 15735 219 16634 se
rect 219 15735 8117 16634
tri 8117 15735 9016 16634 sw
tri 9531 15735 10430 16634 ne
rect 10430 15735 12359 16634
rect -8902 15500 -2202 15735
tri -2202 15500 -1967 15735 nw
tri -915 15500 -680 15735 se
rect -680 15500 9016 15735
tri -9359 15392 -9251 15500 se
rect -9251 15392 -6531 15500
tri -6531 15392 -6423 15500 nw
tri -1023 15392 -915 15500 se
rect -915 15392 1807 15500
tri 1807 15392 1915 15500 nw
tri 6423 15392 6531 15500 ne
rect 6531 15392 9016 15500
tri 9016 15392 9359 15735 sw
tri 10430 15392 10773 15735 ne
rect 10773 15564 12359 15735
tri 12359 15564 13429 16634 sw
tri 13774 15564 14844 16634 ne
rect 14844 15564 16602 16634
rect 10773 15392 13429 15564
tri 13429 15392 13601 15564 sw
tri 14844 15392 15016 15564 ne
rect 15016 15392 16602 15564
tri 16602 15392 17844 16634 sw
tri 18016 15392 19258 16634 ne
rect 19258 15392 20844 16634
tri -18048 15188 -17844 15392 se
rect -17844 15188 -15220 15392
tri -15220 15188 -15016 15392 nw
tri -13805 15188 -13601 15392 se
rect -13601 15188 -10977 15392
tri -10977 15188 -10773 15392 nw
tri -9563 15188 -9359 15392 se
rect -9359 15188 -6735 15392
tri -6735 15188 -6531 15392 nw
tri -1227 15188 -1023 15392 se
rect -1023 15188 1603 15392
tri 1603 15188 1807 15392 nw
tri 6531 15188 6735 15392 ne
rect 6735 15188 9359 15392
tri 9359 15188 9563 15392 sw
tri 10773 15188 10977 15392 ne
rect 10977 15188 13601 15392
tri 13601 15188 13805 15392 sw
tri 15016 15188 15220 15392 ne
rect 15220 15188 17844 15392
tri 17844 15188 18048 15392 sw
tri 19258 15188 19462 15392 ne
rect 19462 15188 20844 15392
tri -23325 14153 -22290 15188 se
rect -22290 15016 -19634 15188
tri -19634 15016 -19462 15188 nw
tri -18220 15016 -18048 15188 se
rect -18048 15016 -15392 15188
tri -15392 15016 -15220 15188 nw
tri -13977 15016 -13805 15188 se
rect -13805 15016 -11149 15188
tri -11149 15016 -10977 15188 nw
tri -9735 15016 -9563 15188 se
rect -9563 15016 -6907 15188
tri -6907 15016 -6735 15188 nw
tri -1399 15016 -1227 15188 se
rect -1227 15016 1431 15188
tri 1431 15016 1603 15188 nw
tri 6735 15016 6907 15188 ne
rect 6907 15016 9563 15188
tri 9563 15016 9735 15188 sw
tri 10977 15016 11149 15188 ne
rect 11149 15016 13805 15188
tri 13805 15016 13977 15188 sw
tri 15220 15016 15392 15188 ne
rect 15392 15016 18048 15188
rect -22290 14153 -20497 15016
tri -20497 14153 -19634 15016 nw
tri -19083 14153 -18220 15016 se
rect -18220 14844 -15564 15016
tri -15564 14844 -15392 15016 nw
tri -14149 14844 -13977 15016 se
rect -13977 14844 -11321 15016
tri -11321 14844 -11149 15016 nw
tri -9907 14844 -9735 15016 se
rect -9735 14844 -7079 15016
tri -7079 14844 -6907 15016 nw
tri -1571 14844 -1399 15016 se
rect -1399 14844 1259 15016
tri 1259 14844 1431 15016 nw
tri 6907 14844 7079 15016 ne
rect 7079 14844 9735 15016
tri 9735 14844 9907 15016 sw
tri 11149 14844 11321 15016 ne
rect 11321 14844 13977 15016
rect -18220 14153 -16255 14844
tri -16255 14153 -15564 14844 nw
tri -14840 14153 -14149 14844 se
rect -14149 14672 -11493 14844
tri -11493 14672 -11321 14844 nw
tri -10079 14672 -9907 14844 se
rect -9907 14672 -7251 14844
tri -7251 14672 -7079 14844 nw
tri -1743 14672 -1571 14844 se
rect -1571 14672 1087 14844
tri 1087 14672 1259 14844 nw
tri 7079 14672 7251 14844 ne
rect 7251 14672 9907 14844
rect -14149 14153 -12012 14672
tri -12012 14153 -11493 14672 nw
tri -10598 14153 -10079 14672 se
rect -10079 14500 -7423 14672
tri -7423 14500 -7251 14672 nw
tri -1745 14670 -1743 14672 se
rect -1743 14670 1085 14672
tri 1085 14670 1087 14672 nw
tri 7251 14670 7253 14672 ne
rect 7253 14670 9907 14672
tri -1915 14500 -1745 14670 se
rect -1745 14500 915 14670
tri 915 14500 1085 14670 nw
tri 7253 14500 7423 14670 ne
rect 7423 14500 9907 14670
rect -10079 14153 -7770 14500
tri -7770 14153 -7423 14500 nw
tri -6355 14153 -6008 14500 se
rect -6008 14153 568 14500
tri 568 14153 915 14500 nw
tri 1732 14253 1979 14500 se
rect 1979 14492 6008 14500
tri 6008 14492 6016 14500 sw
tri 7423 14492 7431 14500 ne
rect 7431 14492 9907 14500
rect 1979 14253 6016 14492
rect 1732 14153 6016 14253
tri -23581 13897 -23325 14153 se
rect -23325 13897 -20753 14153
tri -20753 13897 -20497 14153 nw
tri -19339 13897 -19083 14153 se
rect -19083 13897 -16511 14153
tri -16511 13897 -16255 14153 nw
tri -14844 14149 -14840 14153 se
rect -14840 14149 -12016 14153
tri -12016 14149 -12012 14153 nw
tri -10602 14149 -10598 14153 se
rect -10598 14149 -7774 14153
tri -7774 14149 -7770 14153 nw
tri -6359 14149 -6355 14153 se
rect -6355 14149 312 14153
tri -15096 13897 -14844 14149 se
rect -14844 13897 -12268 14149
tri -12268 13897 -12016 14149 nw
tri -10854 13897 -10602 14149 se
rect -10602 13897 -8026 14149
tri -8026 13897 -7774 14149 nw
tri -6611 13897 -6359 14149 se
rect -6359 13897 312 14149
tri 312 13897 568 14153 nw
rect 1732 13897 1833 14153
rect 2089 13897 2357 14153
rect 2613 13897 2911 14153
rect 3167 13897 3465 14153
rect 3721 13897 4019 14153
rect 4275 13897 4573 14153
rect 4829 13897 5127 14153
rect 5383 13897 5651 14153
rect 5907 14149 6016 14153
tri 6016 14149 6359 14492 sw
tri 7431 14149 7774 14492 ne
rect 7774 14321 9907 14492
tri 9907 14321 10430 14844 sw
tri 11321 14321 11844 14844 ne
rect 11844 14321 13977 14844
rect 7774 14149 10430 14321
tri 10430 14149 10602 14321 sw
tri 11844 14149 12016 14321 ne
rect 12016 14149 13977 14321
tri 13977 14149 14844 15016 sw
tri 15392 14149 16259 15016 ne
rect 16259 14149 18048 15016
rect 5907 13897 6359 14149
tri -23672 13806 -23581 13897 se
rect -23581 13806 -20844 13897
tri -20844 13806 -20753 13897 nw
tri -19430 13806 -19339 13897 se
rect -19339 13806 -16602 13897
tri -16602 13806 -16511 13897 nw
tri -15187 13806 -15096 13897 se
rect -15096 13806 -12359 13897
tri -12359 13806 -12268 13897 nw
tri -10945 13806 -10854 13897 se
rect -10854 13806 -8117 13897
tri -8117 13806 -8026 13897 nw
tri -6702 13806 -6611 13897 se
rect -6611 13806 44 13897
tri -23849 13629 -23672 13806 se
rect -23672 13629 -21021 13806
tri -21021 13629 -20844 13806 nw
tri -19607 13629 -19430 13806 se
rect -19430 13629 -16779 13806
tri -16779 13629 -16602 13806 nw
tri -15364 13629 -15187 13806 se
rect -15187 13629 -12536 13806
tri -12536 13629 -12359 13806 nw
tri -11122 13629 -10945 13806 se
rect -10945 13629 -8294 13806
tri -8294 13629 -8117 13806 nw
tri -6879 13629 -6702 13806 se
rect -6702 13629 44 13806
tri 44 13629 312 13897 nw
rect 1732 13806 6359 13897
tri 6359 13806 6702 14149 sw
tri 7774 13806 8117 14149 ne
rect 8117 13806 10602 14149
tri 10602 13806 10945 14149 sw
tri 12016 13806 12359 14149 ne
rect 12359 13806 14844 14149
tri 14844 13806 15187 14149 sw
tri 16259 13806 16602 14149 ne
rect 16602 13978 18048 14149
tri 18048 13978 19258 15188 sw
tri 19462 13978 20672 15188 ne
rect 20672 13978 20844 15188
rect 16602 13806 19258 13978
tri 19258 13806 19430 13978 sw
tri 20672 13806 20844 13978 ne
tri 20844 13806 23672 16634 sw
rect 1732 13629 6702 13806
tri -24105 13373 -23849 13629 se
rect -23849 13602 -21048 13629
tri -21048 13602 -21021 13629 nw
tri -19634 13602 -19607 13629 se
rect -19607 13602 -16977 13629
rect -23849 13373 -21277 13602
tri -21277 13373 -21048 13602 nw
tri -19863 13373 -19634 13602 se
rect -19634 13431 -16977 13602
tri -16977 13431 -16779 13629 nw
tri -15562 13431 -15364 13629 se
rect -15364 13431 -12792 13629
rect -19634 13373 -17035 13431
tri -17035 13373 -16977 13431 nw
tri -15620 13373 -15562 13431 se
rect -15562 13373 -12792 13431
tri -12792 13373 -12536 13629 nw
tri -11378 13373 -11122 13629 se
rect -11122 13373 -8550 13629
tri -8550 13373 -8294 13629 nw
tri -7135 13373 -6879 13629 se
rect -6879 13373 -212 13629
tri -212 13373 44 13629 nw
rect 1732 13373 1833 13629
rect 2089 13373 2357 13629
rect 2613 13373 2911 13629
rect 3167 13373 3465 13629
rect 3721 13373 4019 13629
rect 4275 13373 4573 13629
rect 4829 13373 5127 13629
rect 5383 13373 5651 13629
rect 5907 13373 6702 13629
tri -24373 13105 -24105 13373 se
rect -24105 13105 -21545 13373
tri -21545 13105 -21277 13373 nw
tri -20131 13105 -19863 13373 se
rect -19863 13105 -17303 13373
tri -17303 13105 -17035 13373 nw
tri -15888 13105 -15620 13373 se
rect -15620 13258 -12907 13373
tri -12907 13258 -12792 13373 nw
tri -11493 13258 -11378 13373 se
rect -11378 13258 -8818 13373
rect -15620 13105 -13060 13258
tri -13060 13105 -12907 13258 nw
tri -11646 13105 -11493 13258 se
rect -11493 13105 -8818 13258
tri -8818 13105 -8550 13373 nw
tri -7403 13105 -7135 13373 se
rect -7135 13105 -480 13373
tri -480 13105 -212 13373 nw
rect 1732 13105 6702 13373
tri -24629 12849 -24373 13105 se
rect -24373 12849 -21801 13105
tri -21801 12849 -21545 13105 nw
tri -20387 12849 -20131 13105 se
rect -20131 12849 -17559 13105
tri -17559 12849 -17303 13105 nw
tri -16144 12849 -15888 13105 se
rect -15888 12849 -13316 13105
tri -13316 12849 -13060 13105 nw
tri -11844 12907 -11646 13105 se
rect -11646 13087 -8836 13105
tri -8836 13087 -8818 13105 nw
tri -7421 13087 -7403 13105 se
rect -7403 13087 -736 13105
rect -11646 12907 -9016 13087
tri -9016 12907 -8836 13087 nw
tri -7601 12907 -7421 13087 se
rect -7421 12907 -736 13087
tri -11902 12849 -11844 12907 se
rect -11844 12849 -9074 12907
tri -9074 12849 -9016 12907 nw
tri -7659 12849 -7601 12907 se
rect -7601 12849 -736 12907
tri -736 12849 -480 13105 nw
rect 1732 12849 1833 13105
rect 2089 12849 2357 13105
rect 2613 12849 2911 13105
rect 3167 12849 3465 13105
rect 3721 12849 4019 13105
rect 4275 12849 4573 13105
rect 4829 12849 5127 13105
rect 5383 12849 5651 13105
rect 5907 13079 6702 13105
tri 6702 13079 7429 13806 sw
tri 8117 13079 8844 13806 ne
rect 8844 13079 10945 13806
rect 5907 12907 7429 13079
tri 7429 12907 7601 13079 sw
tri 8844 12907 9016 13079 ne
rect 9016 12907 10945 13079
tri 10945 12907 11844 13806 sw
tri 12359 12907 13258 13806 ne
rect 13258 12907 15187 13806
rect 5907 12849 7601 12907
tri -25118 12360 -24629 12849 se
rect -24629 12360 -22290 12849
tri -22290 12360 -21801 12849 nw
tri -20672 12564 -20387 12849 se
rect -20387 12564 -17844 12849
tri -17844 12564 -17559 12849 nw
tri -16429 12564 -16144 12849 se
rect -16144 12564 -13601 12849
tri -13601 12564 -13316 12849 nw
tri -12187 12564 -11902 12849 se
rect -11902 12564 -9359 12849
tri -9359 12564 -9074 12849 nw
tri -7944 12564 -7659 12849 se
rect -7659 12564 -1021 12849
tri -1021 12564 -736 12849 nw
rect 1732 12747 7601 12849
tri 1732 12564 1915 12747 ne
rect 1915 12564 7601 12747
tri 7601 12564 7944 12907 sw
tri 9016 12564 9359 12907 ne
rect 9359 12564 11844 12907
tri 11844 12564 12187 12907 sw
tri 13258 12564 13601 12907 ne
rect 13601 12736 15187 12907
tri 15187 12736 16257 13806 sw
tri 16602 12736 17672 13806 ne
rect 17672 12736 19430 13806
rect 13601 12564 16257 12736
tri 16257 12564 16429 12736 sw
tri 17672 12564 17844 12736 ne
rect 17844 12564 19430 12736
tri 19430 12564 20672 13806 sw
tri 20844 12564 22086 13806 ne
rect 22086 12564 23672 13806
tri -20876 12360 -20672 12564 se
rect -20672 12360 -18048 12564
tri -18048 12360 -17844 12564 nw
tri -16633 12360 -16429 12564 se
rect -16429 12360 -13805 12564
tri -13805 12360 -13601 12564 nw
tri -12391 12360 -12187 12564 se
rect -12187 12360 -9563 12564
tri -9563 12360 -9359 12564 nw
tri -8008 12500 -7944 12564 se
rect -7944 12500 -1085 12564
tri -1085 12500 -1021 12564 nw
tri 1915 12500 1979 12564 ne
rect 1979 12500 7944 12564
tri 7944 12500 8008 12564 sw
tri 9359 12500 9423 12564 ne
rect 9423 12500 12187 12564
tri -8148 12360 -8008 12500 se
rect -8008 12360 -5320 12500
tri -5320 12360 -5180 12500 nw
tri 5180 12360 5320 12500 ne
rect 5320 12360 8008 12500
tri 8008 12360 8148 12500 sw
tri 9423 12360 9563 12500 ne
rect 9563 12360 12187 12500
tri 12187 12360 12391 12564 sw
tri 13601 12360 13805 12564 ne
rect 13805 12360 16429 12564
tri 16429 12360 16633 12564 sw
tri 17844 12360 18048 12564 ne
rect 18048 12360 20672 12564
tri 20672 12360 20876 12564 sw
tri 22086 12360 22290 12564 ne
rect 22290 12360 23672 12564
tri -26500 10978 -25118 12360 se
rect -25118 12188 -22462 12360
tri -22462 12188 -22290 12360 nw
tri -21048 12188 -20876 12360 se
rect -20876 12188 -18220 12360
tri -18220 12188 -18048 12360 nw
tri -16805 12188 -16633 12360 se
rect -16633 12188 -13977 12360
tri -13977 12188 -13805 12360 nw
tri -12563 12188 -12391 12360 se
rect -12391 12188 -9735 12360
tri -9735 12188 -9563 12360 nw
tri -8320 12188 -8148 12360 se
rect -8148 12188 -5492 12360
tri -5492 12188 -5320 12360 nw
tri 5320 12188 5492 12360 ne
rect 5492 12188 8148 12360
tri 8148 12188 8320 12360 sw
tri 9563 12188 9735 12360 ne
rect 9735 12188 12391 12360
tri 12391 12188 12563 12360 sw
tri 13805 12188 13977 12360 ne
rect 13977 12188 16633 12360
tri 16633 12188 16805 12360 sw
tri 18048 12188 18220 12360 ne
rect 18220 12188 20876 12360
rect -25118 11150 -23500 12188
tri -23500 11150 -22462 12188 nw
tri -22086 11150 -21048 12188 se
rect -21048 12016 -18392 12188
tri -18392 12016 -18220 12188 nw
tri -16977 12016 -16805 12188 se
rect -16805 12016 -14149 12188
tri -14149 12016 -13977 12188 nw
tri -12735 12016 -12563 12188 se
rect -12563 12016 -9907 12188
tri -9907 12016 -9735 12188 nw
tri -8492 12016 -8320 12188 se
rect -8320 12016 -5664 12188
tri -5664 12016 -5492 12188 nw
tri 5492 12016 5664 12188 ne
rect 5664 12016 8320 12188
tri 8320 12016 8492 12188 sw
tri 9735 12016 9907 12188 ne
rect 9907 12016 12563 12188
tri 12563 12016 12735 12188 sw
tri 13977 12016 14149 12188 ne
rect 14149 12016 16805 12188
rect -21048 11150 -19430 12016
rect -25118 10978 -23672 11150
tri -23672 10978 -23500 11150 nw
tri -22258 10978 -22086 11150 se
rect -22086 10978 -19430 11150
tri -19430 10978 -18392 12016 nw
tri -17672 11321 -16977 12016 se
rect -16977 11844 -14321 12016
tri -14321 11844 -14149 12016 nw
tri -12907 11844 -12735 12016 se
rect -12735 11844 -10079 12016
tri -10079 11844 -9907 12016 nw
tri -8664 11844 -8492 12016 se
rect -8492 11844 -5836 12016
tri -5836 11844 -5664 12016 nw
tri 5664 11844 5836 12016 ne
rect 5836 11844 8492 12016
tri 8492 11844 8664 12016 sw
tri 9907 11844 10079 12016 ne
rect 10079 11844 12735 12016
rect -16977 11321 -14844 11844
tri -14844 11321 -14321 11844 nw
tri -13430 11321 -12907 11844 se
rect -12907 11672 -10251 11844
tri -10251 11672 -10079 11844 nw
tri -8836 11672 -8664 11844 se
rect -8664 11672 -6008 11844
tri -6008 11672 -5836 11844 nw
tri 5836 11672 6008 11844 ne
rect 6008 11672 8664 11844
rect -12907 11321 -10602 11672
tri -10602 11321 -10251 11672 nw
tri -8844 11664 -8836 11672 se
rect -8836 11664 -6016 11672
tri -6016 11664 -6008 11672 nw
tri 6008 11664 6016 11672 ne
rect 6016 11664 8664 11672
tri 8664 11664 8844 11844 sw
tri 10079 11664 10259 11844 ne
rect 10259 11664 12735 11844
tri -9187 11321 -8844 11664 se
rect -8844 11321 -6359 11664
tri -6359 11321 -6016 11664 nw
tri 6016 11321 6359 11664 ne
rect 6359 11321 8844 11664
tri 8844 11321 9187 11664 sw
tri 10259 11321 10602 11664 ne
rect 10602 11493 12735 11664
tri 12735 11493 13258 12016 sw
tri 14149 11493 14672 12016 ne
rect 14672 11493 16805 12016
rect 10602 11321 13258 11493
tri 13258 11321 13430 11493 sw
tri 14672 11321 14844 11493 ne
rect 14844 11321 16805 11493
tri 16805 11321 17672 12188 sw
tri 18220 11321 19087 12188 ne
rect 19087 11321 20876 12188
tri -18015 10978 -17672 11321 se
rect -17672 10978 -15187 11321
tri -15187 10978 -14844 11321 nw
tri -13773 10978 -13430 11321 se
rect -13430 10978 -10945 11321
tri -10945 10978 -10602 11321 nw
tri -9530 10978 -9187 11321 se
rect -9187 10978 -6702 11321
tri -6702 10978 -6359 11321 nw
tri 6359 10978 6702 11321 ne
rect 6702 10978 9187 11321
tri 9187 10978 9530 11321 sw
tri 10602 10978 10945 11321 ne
rect 10945 10978 13430 11321
tri 13430 10978 13773 11321 sw
tri 14844 10978 15187 11321 ne
rect 15187 10978 17672 11321
tri 17672 10978 18015 11321 sw
tri 19087 10978 19430 11321 ne
rect 19430 11150 20876 11321
tri 20876 11150 22086 12360 sw
tri 22290 11150 23500 12360 ne
rect 23500 11150 23672 12360
rect 19430 10978 22086 11150
tri 22086 10978 22258 11150 sw
tri 23500 10978 23672 11150 ne
tri 23672 10978 26500 13806 sw
rect -26500 -10978 -24500 10978
tri -24500 10150 -23672 10978 nw
tri -23086 10150 -22258 10978 se
rect -22258 10603 -19805 10978
tri -19805 10603 -19430 10978 nw
tri -18390 10603 -18015 10978 se
rect -18015 10603 -15735 10978
rect -22258 10150 -20258 10603
tri -20258 10150 -19805 10603 nw
tri -18843 10150 -18390 10603 se
rect -18390 10430 -15735 10603
tri -15735 10430 -15187 10978 nw
tri -14321 10430 -13773 10978 se
rect -13773 10430 -11664 10978
rect -18390 10150 -16015 10430
tri -16015 10150 -15735 10430 nw
tri -14601 10150 -14321 10430 se
rect -14321 10259 -11664 10430
tri -11664 10259 -10945 10978 nw
tri -10249 10259 -9530 10978 se
rect -9530 10259 -7530 10978
rect -14321 10150 -11773 10259
tri -11773 10150 -11664 10259 nw
tri -10358 10150 -10249 10259 se
rect -10249 10150 -7530 10259
tri -7530 10150 -6702 10978 nw
tri 6702 10150 7530 10978 ne
rect 7530 10251 9530 10978
tri 9530 10251 10257 10978 sw
tri 10945 10251 11672 10978 ne
rect 11672 10251 13773 10978
rect 7530 10150 10257 10251
tri 10257 10150 10358 10251 sw
tri 11672 10150 11773 10251 ne
rect 11773 10150 13773 10251
tri 13773 10150 14601 10978 sw
tri 15187 10150 16015 10978 ne
rect 16015 10150 18015 10978
tri 18015 10150 18843 10978 sw
tri 19430 10150 20258 10978 ne
rect 20258 10150 22258 10978
tri 22258 10150 23086 10978 sw
tri 23672 10150 24500 10978 ne
tri -23500 9736 -23086 10150 se
rect -23086 9736 -20672 10150
tri -20672 9736 -20258 10150 nw
tri -19257 9736 -18843 10150 se
rect -18843 9736 -16429 10150
tri -16429 9736 -16015 10150 nw
tri -14672 10079 -14601 10150 se
rect -14601 10079 -11844 10150
tri -11844 10079 -11773 10150 nw
tri -10429 10079 -10358 10150 se
rect -10358 10079 -7601 10150
tri -7601 10079 -7530 10150 nw
tri 7530 10079 7601 10150 ne
rect 7601 10079 10358 10150
tri 10358 10079 10429 10150 sw
tri 11773 10079 11844 10150 ne
rect 11844 10079 14601 10150
tri 14601 10079 14672 10150 sw
tri 16015 10079 16086 10150 ne
rect 16086 10079 18843 10150
tri -15015 9736 -14672 10079 se
rect -14672 9736 -12187 10079
tri -12187 9736 -11844 10079 nw
tri -10772 9736 -10429 10079 se
rect -10429 9736 -7944 10079
tri -7944 9736 -7601 10079 nw
tri 7601 9736 7944 10079 ne
rect 7944 9736 10429 10079
tri 10429 9736 10772 10079 sw
tri 11844 9736 12187 10079 ne
rect 12187 9736 14672 10079
tri 14672 9736 15015 10079 sw
tri 16086 9736 16429 10079 ne
rect 16429 9908 18843 10079
tri 18843 9908 19085 10150 sw
tri 20258 9908 20500 10150 ne
rect 20500 9908 23086 10150
rect 16429 9736 19085 9908
tri 19085 9736 19257 9908 sw
tri 20500 9736 20672 9908 ne
rect 20672 9736 23086 9908
tri 23086 9736 23500 10150 sw
rect -23500 9564 -20844 9736
tri -20844 9564 -20672 9736 nw
tri -19429 9564 -19257 9736 se
rect -19257 9564 -16601 9736
tri -16601 9564 -16429 9736 nw
tri -15187 9564 -15015 9736 se
rect -15015 9564 -12359 9736
tri -12359 9564 -12187 9736 nw
tri -10944 9564 -10772 9736 se
rect -10772 9564 -8116 9736
tri -8116 9564 -7944 9736 nw
tri 7944 9564 8116 9736 ne
rect 8116 9564 10772 9736
tri 10772 9564 10944 9736 sw
tri 12187 9564 12359 9736 ne
rect 12359 9564 15015 9736
tri 15015 9564 15187 9736 sw
tri 16429 9564 16601 9736 ne
rect 16601 9564 19257 9736
tri 19257 9564 19429 9736 sw
tri 20672 9564 20844 9736 ne
rect 20844 9564 23500 9736
rect -23500 -9736 -21500 9564
tri -21500 8908 -20844 9564 nw
tri -19805 9188 -19429 9564 se
rect -19429 9188 -16977 9564
tri -16977 9188 -16601 9564 nw
tri -15563 9188 -15187 9564 se
rect -15187 9188 -12735 9564
tri -12735 9188 -12359 9564 nw
tri -11320 9188 -10944 9564 se
rect -10944 9188 -8492 9564
tri -8492 9188 -8116 9564 nw
tri 8116 9188 8492 9564 ne
rect 8492 9188 10944 9564
tri 10944 9188 11320 9564 sw
tri 12359 9188 12735 9564 ne
rect 12735 9188 15187 9564
tri 15187 9188 15563 9564 sw
tri 16601 9188 16977 9564 ne
rect 16977 9188 19429 9564
tri -20085 8908 -19805 9188 se
rect -19805 9016 -17149 9188
tri -17149 9016 -16977 9188 nw
tri -15735 9016 -15563 9188 se
rect -15563 9016 -12907 9188
tri -12907 9016 -12735 9188 nw
tri -11492 9016 -11320 9188 se
rect -11320 9016 -8664 9188
tri -8664 9016 -8492 9188 nw
tri 8492 9016 8664 9188 ne
rect 8664 9016 11320 9188
tri 11320 9016 11492 9188 sw
tri 12735 9016 12907 9188 ne
rect 12907 9016 15563 9188
rect -19805 8908 -17257 9016
tri -17257 8908 -17149 9016 nw
tri -15843 8908 -15735 9016 se
rect -15735 8908 -13015 9016
tri -13015 8908 -12907 9016 nw
tri -11600 8908 -11492 9016 se
rect -11492 8908 -8772 9016
tri -8772 8908 -8664 9016 nw
tri 8664 8908 8772 9016 ne
rect 8772 8908 11492 9016
tri 11492 8908 11600 9016 sw
tri 12907 8908 13015 9016 ne
rect 13015 8908 15563 9016
tri 15563 8908 15843 9188 sw
tri 16977 8908 17257 9188 ne
rect 17257 8908 19429 9188
tri 19429 8908 20085 9564 sw
tri 20844 8908 21500 9564 ne
tri -20500 8493 -20085 8908 se
rect -20085 8665 -17500 8908
tri -17500 8665 -17257 8908 nw
tri -16086 8665 -15843 8908 se
rect -15843 8844 -13079 8908
tri -13079 8844 -13015 8908 nw
tri -11664 8844 -11600 8908 se
rect -11600 8844 -8836 8908
tri -8836 8844 -8772 8908 nw
tri 8772 8844 8836 8908 ne
rect 8836 8844 11600 8908
rect -15843 8665 -13430 8844
rect -20085 8493 -17672 8665
tri -17672 8493 -17500 8665 nw
tri -16258 8493 -16086 8665 se
rect -16086 8493 -13430 8665
tri -13430 8493 -13079 8844 nw
tri -11672 8836 -11664 8844 se
rect -11664 8836 -8844 8844
tri -8844 8836 -8836 8844 nw
tri 8836 8836 8844 8844 ne
rect 8844 8836 11600 8844
tri 11600 8836 11672 8908 sw
tri 13015 8836 13087 8908 ne
rect 13087 8836 15843 8908
tri -12015 8493 -11672 8836 se
rect -11672 8493 -9187 8836
tri -9187 8493 -8844 8836 nw
tri 8844 8493 9187 8836 ne
rect 9187 8493 11672 8836
tri 11672 8493 12015 8836 sw
tri 13087 8493 13430 8836 ne
rect 13430 8665 15843 8836
tri 15843 8665 16086 8908 sw
tri 17257 8665 17500 8908 ne
rect 17500 8665 20085 8908
rect 13430 8493 16086 8665
tri 16086 8493 16258 8665 sw
tri 17500 8493 17672 8665 ne
rect 17672 8493 20085 8665
tri 20085 8493 20500 8908 sw
rect -20500 -8493 -18500 8493
tri -18500 7665 -17672 8493 nw
tri -17086 7665 -16258 8493 se
rect -16258 7665 -14258 8493
tri -14258 7665 -13430 8493 nw
tri -12843 7665 -12015 8493 se
rect -12015 7665 -10015 8493
tri -10015 7665 -9187 8493 nw
tri 9187 7665 10015 8493 ne
rect 10015 7665 12015 8493
tri 12015 7665 12843 8493 sw
tri 13430 7665 14258 8493 ne
rect 14258 7665 16258 8493
tri 16258 7665 17086 8493 sw
tri 17672 7665 18500 8493 ne
tri -17500 7251 -17086 7665 se
rect -17086 7431 -14492 7665
tri -14492 7431 -14258 7665 nw
tri -13077 7431 -12843 7665 se
rect -12843 7431 -10429 7665
rect -17086 7251 -14672 7431
tri -14672 7251 -14492 7431 nw
tri -13257 7251 -13077 7431 se
rect -13077 7251 -10429 7431
tri -10429 7251 -10015 7665 nw
tri 10015 7251 10429 7665 ne
rect 10429 7423 12843 7665
tri 12843 7423 13085 7665 sw
tri 14258 7423 14500 7665 ne
rect 14500 7423 17086 7665
rect 10429 7251 13085 7423
tri 13085 7251 13257 7423 sw
tri 14500 7251 14672 7423 ne
rect 14672 7251 17086 7423
tri 17086 7251 17500 7665 sw
rect -17500 -7251 -15500 7251
tri -15500 6423 -14672 7251 nw
tri -14085 6423 -13257 7251 se
rect -13257 6423 -11257 7251
tri -11257 6423 -10429 7251 nw
tri 10429 6423 11257 7251 ne
rect 11257 6423 13257 7251
tri 13257 6423 14085 7251 sw
tri 14672 6423 15500 7251 ne
tri -14492 6016 -14085 6423 se
rect -14085 6016 -11664 6423
tri -11664 6016 -11257 6423 nw
tri 11257 6016 11664 6423 ne
rect 11664 6016 14085 6423
tri -14500 6008 -14492 6016 se
rect -14492 6008 -11672 6016
tri -11672 6008 -11664 6016 nw
tri 11664 6008 11672 6016 ne
rect 11672 6008 14085 6016
tri 14085 6008 14500 6423 sw
rect -14500 1000 -12500 6008
tri -12500 5180 -11672 6008 nw
tri 11672 5180 12500 6008 ne
rect -14500 652 11500 1000
rect -14500 396 10052 652
rect 10308 396 10576 652
rect 10832 396 11130 652
rect 11386 396 11500 652
rect -14500 128 11500 396
rect -14500 -128 10052 128
rect 10308 -128 10576 128
rect 10832 -128 11130 128
rect 11386 -128 11500 128
rect -14500 -396 11500 -128
rect -14500 -652 10052 -396
rect 10308 -652 10576 -396
rect 10832 -652 11130 -396
rect 11386 -652 11500 -396
rect -14500 -1000 11500 -652
rect -14500 -6008 -12500 -1000
tri -12500 -6008 -11672 -5180 sw
tri 11672 -6008 12500 -5180 se
rect 12500 -6008 14500 6008
tri -14500 -6016 -14492 -6008 ne
rect -14492 -6016 -11672 -6008
tri -11672 -6016 -11664 -6008 sw
tri 11664 -6016 11672 -6008 se
rect 11672 -6016 14492 -6008
tri 14492 -6016 14500 -6008 nw
tri -14492 -6423 -14085 -6016 ne
rect -14085 -6423 -11664 -6016
tri -11664 -6423 -11257 -6016 sw
tri 11257 -6423 11664 -6016 se
rect 11664 -6423 14085 -6016
tri 14085 -6423 14492 -6016 nw
tri -15500 -7251 -14672 -6423 sw
tri -14085 -7251 -13257 -6423 ne
rect -13257 -7251 -11257 -6423
tri -11257 -7251 -10429 -6423 sw
tri 10429 -7251 11257 -6423 se
rect 11257 -7251 13257 -6423
tri 13257 -7251 14085 -6423 nw
tri 14672 -7251 15500 -6423 se
rect 15500 -7251 17500 7251
tri -17500 -7665 -17086 -7251 ne
rect -17086 -7423 -14672 -7251
tri -14672 -7423 -14500 -7251 sw
tri -13257 -7423 -13085 -7251 ne
rect -13085 -7423 -10429 -7251
rect -17086 -7665 -14500 -7423
tri -14500 -7665 -14258 -7423 sw
tri -13085 -7665 -12843 -7423 ne
rect -12843 -7665 -10429 -7423
tri -10429 -7665 -10015 -7251 sw
tri 10015 -7665 10429 -7251 se
rect 10429 -7431 13077 -7251
tri 13077 -7431 13257 -7251 nw
tri 14492 -7431 14672 -7251 se
rect 14672 -7431 17086 -7251
rect 10429 -7665 12843 -7431
tri 12843 -7665 13077 -7431 nw
tri 14258 -7665 14492 -7431 se
rect 14492 -7665 17086 -7431
tri 17086 -7665 17500 -7251 nw
tri -18500 -8493 -17672 -7665 sw
tri -17086 -8493 -16258 -7665 ne
rect -16258 -8493 -14258 -7665
tri -14258 -8493 -13430 -7665 sw
tri -12843 -8493 -12015 -7665 ne
rect -12015 -8493 -10015 -7665
tri -10015 -8493 -9187 -7665 sw
tri 9187 -8493 10015 -7665 se
rect 10015 -8493 12015 -7665
tri 12015 -8493 12843 -7665 nw
tri 13430 -8493 14258 -7665 se
rect 14258 -8493 16258 -7665
tri 16258 -8493 17086 -7665 nw
tri 17672 -8493 18500 -7665 se
rect 18500 -8493 20500 8493
tri -20500 -8908 -20085 -8493 ne
rect -20085 -8665 -17672 -8493
tri -17672 -8665 -17500 -8493 sw
tri -16258 -8665 -16086 -8493 ne
rect -16086 -8665 -13430 -8493
rect -20085 -8908 -17500 -8665
tri -17500 -8908 -17257 -8665 sw
tri -16086 -8908 -15843 -8665 ne
rect -15843 -8836 -13430 -8665
tri -13430 -8836 -13087 -8493 sw
tri -12015 -8836 -11672 -8493 ne
rect -11672 -8836 -9187 -8493
tri -9187 -8836 -8844 -8493 sw
tri 8844 -8836 9187 -8493 se
rect 9187 -8836 11664 -8493
rect -15843 -8908 -13087 -8836
tri -13087 -8908 -13015 -8836 sw
tri -11672 -8844 -11664 -8836 ne
rect -11664 -8844 -8844 -8836
tri -8844 -8844 -8836 -8836 sw
tri 8836 -8844 8844 -8836 se
rect 8844 -8844 11664 -8836
tri 11664 -8844 12015 -8493 nw
tri 13079 -8844 13430 -8493 se
rect 13430 -8665 16086 -8493
tri 16086 -8665 16258 -8493 nw
tri 17500 -8665 17672 -8493 se
rect 17672 -8665 20085 -8493
rect 13430 -8844 15843 -8665
tri -11664 -8908 -11600 -8844 ne
rect -11600 -8908 -8836 -8844
tri -8836 -8908 -8772 -8844 sw
tri 8772 -8908 8836 -8844 se
rect 8836 -8908 11600 -8844
tri 11600 -8908 11664 -8844 nw
tri 13015 -8908 13079 -8844 se
rect 13079 -8908 15843 -8844
tri 15843 -8908 16086 -8665 nw
tri 17257 -8908 17500 -8665 se
rect 17500 -8908 20085 -8665
tri 20085 -8908 20500 -8493 nw
tri -21500 -9736 -20672 -8908 sw
tri -20085 -9188 -19805 -8908 ne
rect -19805 -9188 -17257 -8908
tri -17257 -9188 -16977 -8908 sw
tri -15843 -9016 -15735 -8908 ne
rect -15735 -9016 -13015 -8908
tri -13015 -9016 -12907 -8908 sw
tri -11600 -9016 -11492 -8908 ne
rect -11492 -9016 -8772 -8908
tri -8772 -9016 -8664 -8908 sw
tri 8664 -9016 8772 -8908 se
rect 8772 -9016 11492 -8908
tri 11492 -9016 11600 -8908 nw
tri 12907 -9016 13015 -8908 se
rect 13015 -9016 15735 -8908
tri 15735 -9016 15843 -8908 nw
tri 17149 -9016 17257 -8908 se
rect 17257 -9016 19805 -8908
tri -15735 -9188 -15563 -9016 ne
rect -15563 -9188 -12907 -9016
tri -12907 -9188 -12735 -9016 sw
tri -11492 -9188 -11320 -9016 ne
rect -11320 -9188 -8664 -9016
tri -8664 -9188 -8492 -9016 sw
tri 8492 -9188 8664 -9016 se
rect 8664 -9188 11320 -9016
tri 11320 -9188 11492 -9016 nw
tri 12735 -9188 12907 -9016 se
rect 12907 -9188 15563 -9016
tri 15563 -9188 15735 -9016 nw
tri 16977 -9188 17149 -9016 se
rect 17149 -9188 19805 -9016
tri 19805 -9188 20085 -8908 nw
tri 21220 -9188 21500 -8908 se
rect 21500 -9188 23500 9564
rect 24500 5000 26500 10978
rect 24500 3000 27500 5000
tri -19805 -9736 -19257 -9188 ne
rect -19257 -9736 -16977 -9188
tri -16977 -9736 -16429 -9188 sw
tri -15563 -9736 -15015 -9188 ne
rect -15015 -9736 -12735 -9188
tri -12735 -9736 -12187 -9188 sw
tri -11320 -9736 -10772 -9188 ne
rect -10772 -9736 -8492 -9188
tri -8492 -9736 -7944 -9188 sw
tri 7944 -9736 8492 -9188 se
rect 8492 -9736 10772 -9188
tri 10772 -9736 11320 -9188 nw
tri 12187 -9736 12735 -9188 se
rect 12735 -9736 15015 -9188
tri 15015 -9736 15563 -9188 nw
tri 16429 -9736 16977 -9188 se
rect 16977 -9736 19257 -9188
tri 19257 -9736 19805 -9188 nw
tri 20672 -9736 21220 -9188 se
rect 21220 -9736 23500 -9188
tri -23500 -10150 -23086 -9736 ne
rect -23086 -9908 -20672 -9736
tri -20672 -9908 -20500 -9736 sw
tri -19257 -9908 -19085 -9736 ne
rect -19085 -9908 -16429 -9736
rect -23086 -10150 -20500 -9908
tri -20500 -10150 -20258 -9908 sw
tri -19085 -10150 -18843 -9908 ne
rect -18843 -10079 -16429 -9908
tri -16429 -10079 -16086 -9736 sw
tri -15015 -10079 -14672 -9736 ne
rect -14672 -10079 -12187 -9736
tri -12187 -10079 -11844 -9736 sw
tri -10772 -10079 -10429 -9736 ne
rect -10429 -10079 -7944 -9736
tri -7944 -10079 -7601 -9736 sw
tri 7601 -10079 7944 -9736 se
rect 7944 -10079 10429 -9736
tri 10429 -10079 10772 -9736 nw
tri 11844 -10079 12187 -9736 se
rect 12187 -10079 14601 -9736
rect -18843 -10150 -16086 -10079
tri -16086 -10150 -16015 -10079 sw
tri -14672 -10150 -14601 -10079 ne
rect -14601 -10150 -11844 -10079
tri -11844 -10150 -11773 -10079 sw
tri -10429 -10150 -10358 -10079 ne
rect -10358 -10150 -7601 -10079
tri -7601 -10150 -7530 -10079 sw
tri 7530 -10150 7601 -10079 se
rect 7601 -10150 10358 -10079
tri 10358 -10150 10429 -10079 nw
tri 11773 -10150 11844 -10079 se
rect 11844 -10150 14601 -10079
tri 14601 -10150 15015 -9736 nw
tri 16015 -10150 16429 -9736 se
rect 16429 -10150 18843 -9736
tri 18843 -10150 19257 -9736 nw
tri 20258 -10150 20672 -9736 se
rect 20672 -10150 23086 -9736
tri 23086 -10150 23500 -9736 nw
rect 24500 -5000 27500 -3000
tri -24500 -10978 -23672 -10150 sw
tri -23086 -10978 -22258 -10150 ne
rect -22258 -10978 -20258 -10150
tri -20258 -10978 -19430 -10150 sw
tri -18843 -10978 -18015 -10150 ne
rect -18015 -10978 -16015 -10150
tri -16015 -10978 -15187 -10150 sw
tri -14601 -10978 -13773 -10150 ne
rect -13773 -10251 -11773 -10150
tri -11773 -10251 -11672 -10150 sw
tri -10358 -10251 -10257 -10150 ne
rect -10257 -10251 -7530 -10150
rect -13773 -10978 -11672 -10251
tri -11672 -10978 -10945 -10251 sw
tri -10257 -10978 -9530 -10251 ne
rect -9530 -10978 -7530 -10251
tri -7530 -10978 -6702 -10150 sw
tri 6702 -10978 7530 -10150 se
rect 7530 -10259 10249 -10150
tri 10249 -10259 10358 -10150 nw
tri 11664 -10259 11773 -10150 se
rect 11773 -10259 14321 -10150
rect 7530 -10978 9530 -10259
tri 9530 -10978 10249 -10259 nw
tri 10945 -10978 11664 -10259 se
rect 11664 -10430 14321 -10259
tri 14321 -10430 14601 -10150 nw
tri 15735 -10430 16015 -10150 se
rect 16015 -10430 18390 -10150
rect 11664 -10978 13773 -10430
tri 13773 -10978 14321 -10430 nw
tri 15187 -10978 15735 -10430 se
rect 15735 -10603 18390 -10430
tri 18390 -10603 18843 -10150 nw
tri 19805 -10603 20258 -10150 se
rect 20258 -10603 22258 -10150
rect 15735 -10978 18015 -10603
tri 18015 -10978 18390 -10603 nw
tri 19430 -10978 19805 -10603 se
rect 19805 -10978 22258 -10603
tri 22258 -10978 23086 -10150 nw
tri 23672 -10978 24500 -10150 se
rect 24500 -10978 26500 -5000
tri -26500 -12360 -25118 -10978 ne
rect -25118 -11150 -23672 -10978
tri -23672 -11150 -23500 -10978 sw
tri -22258 -11150 -22086 -10978 ne
rect -22086 -11150 -19430 -10978
rect -25118 -12360 -23500 -11150
tri -23500 -12360 -22290 -11150 sw
tri -22086 -12188 -21048 -11150 ne
rect -21048 -11321 -19430 -11150
tri -19430 -11321 -19087 -10978 sw
tri -18015 -11321 -17672 -10978 ne
rect -17672 -11321 -15187 -10978
tri -15187 -11321 -14844 -10978 sw
tri -13773 -11321 -13430 -10978 ne
rect -13430 -11321 -10945 -10978
tri -10945 -11321 -10602 -10978 sw
tri -9530 -11321 -9187 -10978 ne
rect -9187 -11321 -6702 -10978
tri -6702 -11321 -6359 -10978 sw
tri 6359 -11321 6702 -10978 se
rect 6702 -11321 9187 -10978
tri 9187 -11321 9530 -10978 nw
tri 10602 -11321 10945 -10978 se
rect 10945 -11321 13430 -10978
tri 13430 -11321 13773 -10978 nw
tri 14844 -11321 15187 -10978 se
rect 15187 -11321 16977 -10978
rect -21048 -12188 -19087 -11321
tri -19087 -12188 -18220 -11321 sw
tri -17672 -12016 -16977 -11321 ne
rect -16977 -11493 -14844 -11321
tri -14844 -11493 -14672 -11321 sw
tri -13430 -11493 -13258 -11321 ne
rect -13258 -11493 -10602 -11321
rect -16977 -12016 -14672 -11493
tri -14672 -12016 -14149 -11493 sw
tri -13258 -11844 -12907 -11493 ne
rect -12907 -11664 -10602 -11493
tri -10602 -11664 -10259 -11321 sw
tri -9187 -11664 -8844 -11321 ne
rect -8844 -11664 -6359 -11321
tri -6359 -11664 -6016 -11321 sw
tri 6016 -11664 6359 -11321 se
rect 6359 -11664 8836 -11321
rect -12907 -11844 -10259 -11664
tri -10259 -11844 -10079 -11664 sw
tri -8844 -11672 -8836 -11664 ne
rect -8836 -11672 -6016 -11664
tri -6016 -11672 -6008 -11664 sw
tri 6008 -11672 6016 -11664 se
rect 6016 -11672 8836 -11664
tri 8836 -11672 9187 -11321 nw
tri 10251 -11672 10602 -11321 se
rect 10602 -11672 12907 -11321
tri -8836 -11844 -8664 -11672 ne
rect -8664 -11844 -6008 -11672
tri -6008 -11844 -5836 -11672 sw
tri 5836 -11844 6008 -11672 se
rect 6008 -11844 8664 -11672
tri 8664 -11844 8836 -11672 nw
tri 10079 -11844 10251 -11672 se
rect 10251 -11844 12907 -11672
tri 12907 -11844 13430 -11321 nw
tri 14321 -11844 14844 -11321 se
rect 14844 -11844 16977 -11321
tri -12907 -12016 -12735 -11844 ne
rect -12735 -12016 -10079 -11844
tri -10079 -12016 -9907 -11844 sw
tri -8664 -12016 -8492 -11844 ne
rect -8492 -12016 -5836 -11844
tri -5836 -12016 -5664 -11844 sw
tri 5664 -12016 5836 -11844 se
rect 5836 -12016 8492 -11844
tri 8492 -12016 8664 -11844 nw
tri 9907 -12016 10079 -11844 se
rect 10079 -12016 12735 -11844
tri 12735 -12016 12907 -11844 nw
tri 14149 -12016 14321 -11844 se
rect 14321 -12016 16977 -11844
tri 16977 -12016 18015 -10978 nw
tri 18392 -12016 19430 -10978 se
rect 19430 -11150 22086 -10978
tri 22086 -11150 22258 -10978 nw
tri 23500 -11150 23672 -10978 se
rect 23672 -11150 25118 -10978
rect 19430 -12016 21048 -11150
tri -16977 -12188 -16805 -12016 ne
rect -16805 -12188 -14149 -12016
tri -14149 -12188 -13977 -12016 sw
tri -12735 -12188 -12563 -12016 ne
rect -12563 -12188 -9907 -12016
tri -9907 -12188 -9735 -12016 sw
tri -8492 -12188 -8320 -12016 ne
rect -8320 -12188 -5664 -12016
tri -5664 -12188 -5492 -12016 sw
tri 5492 -12188 5664 -12016 se
rect 5664 -12188 8320 -12016
tri 8320 -12188 8492 -12016 nw
tri 9735 -12188 9907 -12016 se
rect 9907 -12188 12563 -12016
tri 12563 -12188 12735 -12016 nw
tri 13977 -12188 14149 -12016 se
rect 14149 -12188 16805 -12016
tri 16805 -12188 16977 -12016 nw
tri 18220 -12188 18392 -12016 se
rect 18392 -12188 21048 -12016
tri 21048 -12188 22086 -11150 nw
tri 22462 -12188 23500 -11150 se
rect 23500 -12188 25118 -11150
tri -21048 -12360 -20876 -12188 ne
rect -20876 -12360 -18220 -12188
tri -18220 -12360 -18048 -12188 sw
tri -16805 -12360 -16633 -12188 ne
rect -16633 -12360 -13977 -12188
tri -13977 -12360 -13805 -12188 sw
tri -12563 -12360 -12391 -12188 ne
rect -12391 -12360 -9735 -12188
tri -9735 -12360 -9563 -12188 sw
tri -8320 -12360 -8148 -12188 ne
rect -8148 -12360 -5492 -12188
tri -5492 -12360 -5320 -12188 sw
tri 5320 -12360 5492 -12188 se
rect 5492 -12360 8148 -12188
tri 8148 -12360 8320 -12188 nw
tri 9563 -12360 9735 -12188 se
rect 9735 -12360 12391 -12188
tri 12391 -12360 12563 -12188 nw
tri 13805 -12360 13977 -12188 se
rect 13977 -12360 16633 -12188
tri 16633 -12360 16805 -12188 nw
tri 18048 -12360 18220 -12188 se
rect 18220 -12360 20876 -12188
tri 20876 -12360 21048 -12188 nw
tri 22290 -12360 22462 -12188 se
rect 22462 -12360 25118 -12188
tri 25118 -12360 26500 -10978 nw
tri -25118 -13806 -23672 -12360 ne
rect -23672 -12564 -22290 -12360
tri -22290 -12564 -22086 -12360 sw
tri -20876 -12564 -20672 -12360 ne
rect -20672 -12564 -18048 -12360
tri -18048 -12564 -17844 -12360 sw
tri -16633 -12564 -16429 -12360 ne
rect -16429 -12564 -13805 -12360
tri -13805 -12564 -13601 -12360 sw
tri -12391 -12564 -12187 -12360 ne
rect -12187 -12564 -9563 -12360
tri -9563 -12564 -9359 -12360 sw
tri -8148 -12564 -7944 -12360 ne
rect -7944 -12500 -5320 -12360
tri -5320 -12500 -5180 -12360 sw
tri 5180 -12500 5320 -12360 se
rect 5320 -12500 7944 -12360
rect -7944 -12564 7944 -12500
tri 7944 -12564 8148 -12360 nw
tri 9359 -12564 9563 -12360 se
rect 9563 -12564 12187 -12360
tri 12187 -12564 12391 -12360 nw
tri 13601 -12564 13805 -12360 se
rect 13805 -12564 16429 -12360
tri 16429 -12564 16633 -12360 nw
tri 17844 -12564 18048 -12360 se
rect 18048 -12564 19634 -12360
rect -23672 -13806 -22086 -12564
tri -22086 -13806 -20844 -12564 sw
tri -20672 -13806 -19430 -12564 ne
rect -19430 -12736 -17844 -12564
tri -17844 -12736 -17672 -12564 sw
tri -16429 -12736 -16257 -12564 ne
rect -16257 -12736 -13601 -12564
rect -19430 -13806 -17672 -12736
tri -17672 -13806 -16602 -12736 sw
tri -16257 -13806 -15187 -12736 ne
rect -15187 -12907 -13601 -12736
tri -13601 -12907 -13258 -12564 sw
tri -12187 -12907 -11844 -12564 ne
rect -11844 -12907 -9359 -12564
tri -9359 -12907 -9016 -12564 sw
tri -7944 -12907 -7601 -12564 ne
rect -7601 -12907 7601 -12564
tri 7601 -12907 7944 -12564 nw
tri 9016 -12907 9359 -12564 se
rect 9359 -12907 11493 -12564
rect -15187 -13806 -13258 -12907
tri -13258 -13806 -12359 -12907 sw
tri -11844 -13806 -10945 -12907 ne
rect -10945 -13079 -9016 -12907
tri -9016 -13079 -8844 -12907 sw
tri -7601 -13079 -7429 -12907 ne
rect -7429 -13079 7421 -12907
rect -10945 -13806 -8844 -13079
tri -8844 -13806 -8117 -13079 sw
tri -7429 -13806 -6702 -13079 ne
rect -6702 -13087 7421 -13079
tri 7421 -13087 7601 -12907 nw
tri 8836 -13087 9016 -12907 se
rect 9016 -13087 11493 -12907
rect -6702 -13806 6702 -13087
tri 6702 -13806 7421 -13087 nw
tri 8117 -13806 8836 -13087 se
rect 8836 -13258 11493 -13087
tri 11493 -13258 12187 -12564 nw
tri 12907 -13258 13601 -12564 se
rect 13601 -13258 15562 -12564
rect 8836 -13806 10945 -13258
tri 10945 -13806 11493 -13258 nw
tri 12359 -13806 12907 -13258 se
rect 12907 -13431 15562 -13258
tri 15562 -13431 16429 -12564 nw
tri 16977 -13431 17844 -12564 se
rect 17844 -13431 19634 -12564
rect 12907 -13806 15187 -13431
tri 15187 -13806 15562 -13431 nw
tri 16602 -13806 16977 -13431 se
rect 16977 -13602 19634 -13431
tri 19634 -13602 20876 -12360 nw
tri 21048 -13602 22290 -12360 se
rect 16977 -13806 19430 -13602
tri 19430 -13806 19634 -13602 nw
tri 20844 -13806 21048 -13602 se
rect 21048 -13806 22290 -13602
tri -23672 -15188 -22290 -13806 ne
rect -22290 -13978 -20844 -13806
tri -20844 -13978 -20672 -13806 sw
tri -19430 -13978 -19258 -13806 ne
rect -19258 -13978 -16602 -13806
rect -22290 -15188 -20672 -13978
tri -20672 -15188 -19462 -13978 sw
tri -19258 -15016 -18220 -13978 ne
rect -18220 -14149 -16602 -13978
tri -16602 -14149 -16259 -13806 sw
tri -15187 -14149 -14844 -13806 ne
rect -14844 -14149 -12359 -13806
tri -12359 -14149 -12016 -13806 sw
tri -10945 -14149 -10602 -13806 ne
rect -10602 -14149 -8117 -13806
tri -8117 -14149 -7774 -13806 sw
tri -6702 -14149 -6359 -13806 ne
rect -6359 -14149 6359 -13806
tri 6359 -14149 6702 -13806 nw
tri 7774 -14149 8117 -13806 se
rect 8117 -14149 10602 -13806
tri 10602 -14149 10945 -13806 nw
tri 12016 -14149 12359 -13806 se
rect 12359 -14149 14149 -13806
rect -18220 -15016 -16259 -14149
tri -16259 -15016 -15392 -14149 sw
tri -14844 -14844 -14149 -14149 ne
rect -14149 -14321 -12016 -14149
tri -12016 -14321 -11844 -14149 sw
tri -10602 -14321 -10430 -14149 ne
rect -10430 -14321 -7774 -14149
rect -14149 -14844 -11844 -14321
tri -11844 -14844 -11321 -14321 sw
tri -10430 -14672 -10079 -14321 ne
rect -10079 -14492 -7774 -14321
tri -7774 -14492 -7431 -14149 sw
tri -6359 -14492 -6016 -14149 ne
rect -6016 -14492 6008 -14149
rect -10079 -14672 -7431 -14492
tri -7431 -14672 -7251 -14492 sw
tri -6016 -14500 -6008 -14492 ne
rect -6008 -14500 6008 -14492
tri 6008 -14500 6359 -14149 nw
tri 7423 -14500 7774 -14149 se
rect 7774 -14500 10079 -14149
tri 7251 -14672 7423 -14500 se
rect 7423 -14672 10079 -14500
tri 10079 -14672 10602 -14149 nw
tri 11493 -14672 12016 -14149 se
rect 12016 -14672 14149 -14149
tri -10079 -14844 -9907 -14672 ne
rect -9907 -14844 -7251 -14672
tri -7251 -14844 -7079 -14672 sw
tri 7079 -14844 7251 -14672 se
rect 7251 -14844 9907 -14672
tri 9907 -14844 10079 -14672 nw
tri 11321 -14844 11493 -14672 se
rect 11493 -14844 14149 -14672
tri 14149 -14844 15187 -13806 nw
tri 15564 -14844 16602 -13806 se
rect 16602 -14844 18220 -13806
tri -14149 -15016 -13977 -14844 ne
rect -13977 -15016 -11321 -14844
tri -11321 -15016 -11149 -14844 sw
tri -9907 -15016 -9735 -14844 ne
rect -9735 -15016 -7079 -14844
tri -7079 -15016 -6907 -14844 sw
tri 6907 -15016 7079 -14844 se
rect 7079 -15016 9735 -14844
tri 9735 -15016 9907 -14844 nw
tri 11149 -15016 11321 -14844 se
rect 11321 -15016 13977 -14844
tri 13977 -15016 14149 -14844 nw
tri 15392 -15016 15564 -14844 se
rect 15564 -15016 18220 -14844
tri 18220 -15016 19430 -13806 nw
tri 19634 -15016 20844 -13806 se
rect 20844 -15016 22290 -13806
tri -18220 -15188 -18048 -15016 ne
rect -18048 -15188 -15392 -15016
tri -15392 -15188 -15220 -15016 sw
tri -13977 -15188 -13805 -15016 ne
rect -13805 -15188 -11149 -15016
tri -11149 -15188 -10977 -15016 sw
tri -9735 -15188 -9563 -15016 ne
rect -9563 -15188 -6907 -15016
tri -6907 -15188 -6735 -15016 sw
tri 6735 -15188 6907 -15016 se
rect 6907 -15188 9563 -15016
tri 9563 -15188 9735 -15016 nw
tri 10977 -15188 11149 -15016 se
rect 11149 -15188 13805 -15016
tri 13805 -15188 13977 -15016 nw
tri 15220 -15188 15392 -15016 se
rect 15392 -15188 18048 -15016
tri 18048 -15188 18220 -15016 nw
tri 19462 -15188 19634 -15016 se
rect 19634 -15188 22290 -15016
tri 22290 -15188 25118 -12360 nw
tri -22290 -15849 -21629 -15188 ne
rect -21629 -15392 -19462 -15188
tri -19462 -15392 -19258 -15188 sw
tri -18048 -15392 -17844 -15188 ne
rect -17844 -15392 -15220 -15188
tri -15220 -15392 -15016 -15188 sw
tri -13805 -15392 -13601 -15188 ne
rect -13601 -15392 -10977 -15188
tri -10977 -15392 -10773 -15188 sw
tri -9563 -15392 -9359 -15188 ne
rect -9359 -15392 -6735 -15188
tri -6735 -15392 -6531 -15188 sw
tri 6531 -15392 6735 -15188 se
rect 6735 -15392 9359 -15188
tri 9359 -15392 9563 -15188 nw
tri 10773 -15392 10977 -15188 se
rect 10977 -15392 13601 -15188
tri 13601 -15392 13805 -15188 nw
tri 15016 -15392 15220 -15188 se
rect 15220 -15392 16806 -15188
rect -21629 -15849 -19258 -15392
tri -19258 -15849 -18801 -15392 sw
tri -17844 -15849 -17387 -15392 ne
rect -17387 -15564 -15016 -15392
tri -15016 -15564 -14844 -15392 sw
tri -13601 -15500 -13493 -15392 ne
rect -13493 -15500 -10773 -15392
tri -10773 -15500 -10665 -15392 sw
tri -9359 -15500 -9251 -15392 ne
rect -9251 -15500 -6531 -15392
tri -6531 -15500 -6423 -15392 sw
tri 6423 -15500 6531 -15392 se
rect 6531 -15500 9251 -15392
tri 9251 -15500 9359 -15392 nw
tri 10665 -15500 10773 -15392 se
rect 10773 -15500 13493 -15392
tri 13493 -15500 13601 -15392 nw
tri 14908 -15500 15016 -15392 se
rect 15016 -15500 16806 -15392
tri -13493 -15564 -13429 -15500 ne
rect -13429 -15564 -10665 -15500
rect -17387 -15849 -14844 -15564
tri -14844 -15849 -14559 -15564 sw
tri -13429 -15849 -13144 -15564 ne
rect -13144 -15735 -10665 -15564
tri -10665 -15735 -10430 -15500 sw
tri -9251 -15735 -9016 -15500 ne
rect -9016 -15735 -1085 -15500
rect -13144 -15849 -10430 -15735
tri -10430 -15849 -10316 -15735 sw
tri -9016 -15849 -8902 -15735 ne
rect -8902 -15849 -1085 -15735
tri -1085 -15849 -736 -15500 sw
tri 1732 -15747 1979 -15500 se
rect 1979 -15747 8665 -15500
rect 1732 -15849 8665 -15747
tri -21629 -16105 -21373 -15849 ne
rect -21373 -16105 -18801 -15849
tri -18801 -16105 -18545 -15849 sw
tri -17387 -16105 -17131 -15849 ne
rect -17131 -16105 -14559 -15849
tri -14559 -16105 -14303 -15849 sw
tri -13144 -16105 -12888 -15849 ne
rect -12888 -16105 -10316 -15849
tri -10316 -16105 -10060 -15849 sw
tri -8902 -16105 -8646 -15849 ne
rect -8646 -16105 -736 -15849
tri -736 -16105 -480 -15849 sw
rect 1732 -16105 1832 -15849
rect 2088 -16105 2356 -15849
rect 2612 -16105 2910 -15849
rect 3166 -16105 3464 -15849
rect 3720 -16105 4018 -15849
rect 4274 -16105 4572 -15849
rect 4828 -16105 5126 -15849
rect 5382 -16105 5650 -15849
rect 5906 -16086 8665 -15849
tri 8665 -16086 9251 -15500 nw
tri 10079 -16086 10665 -15500 se
rect 10665 -16086 12734 -15500
rect 5906 -16105 7251 -16086
tri -21373 -16373 -21105 -16105 ne
rect -21105 -16373 -18545 -16105
tri -18545 -16373 -18277 -16105 sw
tri -17131 -16373 -16863 -16105 ne
rect -16863 -16373 -14303 -16105
tri -14303 -16373 -14035 -16105 sw
tri -12888 -16373 -12620 -16105 ne
rect -12620 -16373 -10060 -16105
tri -10060 -16373 -9792 -16105 sw
tri -8646 -16373 -8378 -16105 ne
rect -8378 -16373 -480 -16105
tri -480 -16373 -212 -16105 sw
rect 1732 -16373 7251 -16105
tri -21105 -16629 -20849 -16373 ne
rect -20849 -16629 -18277 -16373
tri -18277 -16629 -18021 -16373 sw
tri -16863 -16629 -16607 -16373 ne
rect -16607 -16629 -14035 -16373
tri -14035 -16629 -13779 -16373 sw
tri -12620 -16629 -12364 -16373 ne
rect -12364 -16629 -9792 -16373
tri -9792 -16629 -9536 -16373 sw
tri -8378 -16629 -8122 -16373 ne
rect -8122 -16629 -212 -16373
tri -212 -16629 44 -16373 sw
rect 1732 -16629 1832 -16373
rect 2088 -16629 2356 -16373
rect 2612 -16629 2910 -16373
rect 3166 -16629 3464 -16373
rect 3720 -16629 4018 -16373
rect 4274 -16629 4572 -16373
rect 4828 -16629 5126 -16373
rect 5382 -16629 5650 -16373
rect 5906 -16629 7251 -16373
tri -20849 -16634 -20844 -16629 ne
rect -20844 -16634 -18021 -16629
tri -18021 -16634 -18016 -16629 sw
tri -16607 -16634 -16602 -16629 ne
rect -16602 -16634 -13779 -16629
tri -13779 -16634 -13774 -16629 sw
tri -12364 -16634 -12359 -16629 ne
rect -12359 -16634 -9536 -16629
tri -20844 -16897 -20581 -16634 ne
rect -20581 -16806 -18016 -16634
tri -18016 -16806 -17844 -16634 sw
tri -16602 -16806 -16430 -16634 ne
rect -16430 -16806 -13774 -16634
rect -20581 -16897 -17844 -16806
tri -17844 -16897 -17753 -16806 sw
tri -16430 -16897 -16339 -16806 ne
rect -16339 -16897 -13774 -16806
tri -13774 -16897 -13511 -16634 sw
tri -12359 -16897 -12096 -16634 ne
rect -12096 -16897 -9536 -16634
tri -9536 -16897 -9268 -16629 sw
tri -8122 -16897 -7854 -16629 ne
rect -7854 -16634 44 -16629
tri 44 -16634 49 -16629 sw
rect -7854 -16897 49 -16634
tri 49 -16897 312 -16634 sw
rect 1732 -16897 7251 -16629
tri -20581 -17153 -20325 -16897 ne
rect -20325 -17153 -17753 -16897
tri -17753 -17153 -17497 -16897 sw
tri -16339 -17153 -16083 -16897 ne
rect -16083 -16977 -13511 -16897
tri -13511 -16977 -13431 -16897 sw
tri -12096 -16977 -12016 -16897 ne
rect -12016 -16977 -9268 -16897
tri -9268 -16977 -9188 -16897 sw
tri -7854 -16977 -7774 -16897 ne
rect -7774 -16977 312 -16897
rect -16083 -17153 -13431 -16977
tri -13431 -17153 -13255 -16977 sw
tri -12016 -17153 -11840 -16977 ne
rect -11840 -17149 -9188 -16977
tri -9188 -17149 -9016 -16977 sw
tri -7774 -17149 -7602 -16977 ne
rect -7602 -17149 312 -16977
rect -11840 -17153 -9016 -17149
tri -9016 -17153 -9012 -17149 sw
tri -7602 -17153 -7598 -17149 ne
rect -7598 -17153 312 -17149
tri 312 -17153 568 -16897 sw
rect 1732 -17153 1832 -16897
rect 2088 -17153 2356 -16897
rect 2612 -17153 2910 -16897
rect 3166 -17153 3464 -16897
rect 3720 -17153 4018 -16897
rect 4274 -17153 4572 -16897
rect 4828 -17153 5126 -16897
rect 5382 -17153 5650 -16897
rect 5906 -17153 7251 -16897
tri -20325 -18016 -19462 -17153 ne
rect -19462 -18016 -17497 -17153
tri -17497 -18016 -16634 -17153 sw
tri -16083 -17844 -15392 -17153 ne
rect -15392 -17844 -13255 -17153
tri -13255 -17844 -12564 -17153 sw
tri -11840 -17500 -11493 -17153 ne
rect -11493 -17500 -9012 -17153
tri -9012 -17500 -8665 -17153 sw
tri -7598 -17500 -7251 -17153 ne
rect -7251 -17500 568 -17153
tri 568 -17500 915 -17153 sw
rect 1732 -17253 7251 -17153
tri 1732 -17500 1979 -17253 ne
rect 1979 -17500 7251 -17253
tri 7251 -17500 8665 -16086 nw
tri 8665 -17500 10079 -16086 se
rect 10079 -16259 12734 -16086
tri 12734 -16259 13493 -15500 nw
tri 14149 -16259 14908 -15500 se
rect 14908 -16259 16806 -15500
rect 10079 -16634 12359 -16259
tri 12359 -16634 12734 -16259 nw
tri 13774 -16634 14149 -16259 se
rect 14149 -16430 16806 -16259
tri 16806 -16430 18048 -15188 nw
tri 18220 -16430 19462 -15188 se
rect 14149 -16634 16602 -16430
tri 16602 -16634 16806 -16430 nw
tri 18016 -16634 18220 -16430 se
rect 18220 -16634 19462 -16430
rect 10079 -17500 11493 -16634
tri 11493 -17500 12359 -16634 nw
tri 12908 -17500 13774 -16634 se
rect 13774 -17500 15392 -16634
tri -11493 -17670 -11323 -17500 ne
rect -11323 -17670 -8665 -17500
tri -8665 -17670 -8495 -17500 sw
tri -1915 -17670 -1745 -17500 ne
rect -1745 -17670 915 -17500
tri 915 -17670 1085 -17500 sw
tri 8495 -17670 8665 -17500 se
rect 8665 -17670 11323 -17500
tri 11323 -17670 11493 -17500 nw
tri 12738 -17670 12908 -17500 se
rect 12908 -17670 15392 -17500
tri -11323 -17844 -11149 -17670 ne
rect -11149 -17844 -8495 -17670
tri -8495 -17844 -8321 -17670 sw
tri -1745 -17844 -1571 -17670 ne
rect -1571 -17844 1085 -17670
tri 1085 -17844 1259 -17670 sw
tri 8493 -17672 8495 -17670 se
rect 8495 -17672 11321 -17670
tri 11321 -17672 11323 -17670 nw
tri 12736 -17672 12738 -17670 se
rect 12738 -17672 15392 -17670
tri 8321 -17844 8493 -17672 se
rect 8493 -17844 11149 -17672
tri 11149 -17844 11321 -17672 nw
tri 12564 -17844 12736 -17672 se
rect 12736 -17844 15392 -17672
tri 15392 -17844 16602 -16634 nw
tri 16806 -17844 18016 -16634 se
rect 18016 -17844 19462 -16634
tri -15392 -18016 -15220 -17844 ne
rect -15220 -18016 -12564 -17844
tri -12564 -18016 -12392 -17844 sw
tri -11149 -18016 -10977 -17844 ne
rect -10977 -18016 -8321 -17844
tri -8321 -18016 -8149 -17844 sw
tri -1571 -18016 -1399 -17844 ne
rect -1399 -18016 1259 -17844
tri 1259 -18016 1431 -17844 sw
tri 8149 -18016 8321 -17844 se
rect 8321 -18016 10977 -17844
tri 10977 -18016 11149 -17844 nw
tri 12392 -18016 12564 -17844 se
rect 12564 -18016 15220 -17844
tri 15220 -18016 15392 -17844 nw
tri 16634 -18016 16806 -17844 se
rect 16806 -18016 19462 -17844
tri 19462 -18016 22290 -15188 nw
tri -19462 -18848 -18630 -18016 ne
rect -18630 -18220 -16634 -18016
tri -16634 -18220 -16430 -18016 sw
tri -15220 -18220 -15016 -18016 ne
rect -15016 -18220 -12392 -18016
tri -12392 -18220 -12188 -18016 sw
tri -10977 -18220 -10773 -18016 ne
rect -10773 -18220 -8149 -18016
tri -8149 -18220 -7945 -18016 sw
tri -1399 -18220 -1195 -18016 ne
rect -1195 -18220 1431 -18016
rect -18630 -18848 -16430 -18220
tri -16430 -18848 -15802 -18220 sw
tri -15016 -18848 -14388 -18220 ne
rect -14388 -18392 -12188 -18220
tri -12188 -18392 -12016 -18220 sw
tri -10773 -18392 -10601 -18220 ne
rect -10601 -18392 -7945 -18220
rect -14388 -18848 -12016 -18392
tri -12016 -18848 -11560 -18392 sw
tri -10601 -18848 -10145 -18392 ne
rect -10145 -18500 -7945 -18392
tri -7945 -18500 -7665 -18220 sw
tri -1195 -18500 -915 -18220 ne
rect -915 -18500 1431 -18220
tri 1431 -18500 1915 -18016 sw
tri 7665 -18500 8149 -18016 se
rect 8149 -18500 10493 -18016
tri 10493 -18500 10977 -18016 nw
tri 11908 -18500 12392 -18016 se
rect 12392 -18500 13978 -18016
rect -10145 -18747 -2202 -18500
tri -2202 -18747 -1955 -18500 sw
rect -10145 -18848 -1955 -18747
tri -18630 -19104 -18374 -18848 ne
rect -18374 -19104 -15802 -18848
tri -15802 -19104 -15546 -18848 sw
tri -14388 -19104 -14132 -18848 ne
rect -14132 -19104 -11560 -18848
tri -11560 -19104 -11304 -18848 sw
tri -10145 -19104 -9889 -18848 ne
rect -9889 -19104 -6130 -18848
rect -5874 -19104 -5606 -18848
rect -5350 -19104 -5052 -18848
rect -4796 -19104 -4498 -18848
rect -4242 -19104 -3944 -18848
rect -3688 -19104 -3390 -18848
rect -3134 -19104 -2836 -18848
rect -2580 -19104 -2312 -18848
rect -2056 -19104 -1955 -18848
tri -18374 -19372 -18106 -19104 ne
rect -18106 -19372 -15546 -19104
tri -15546 -19372 -15278 -19104 sw
tri -14132 -19372 -13864 -19104 ne
rect -13864 -19372 -11304 -19104
tri -11304 -19372 -11036 -19104 sw
tri -9889 -19372 -9621 -19104 ne
rect -9621 -19372 -1955 -19104
tri -18106 -19462 -18016 -19372 ne
rect -18016 -19462 -15278 -19372
tri -15278 -19462 -15188 -19372 sw
tri -13864 -19462 -13774 -19372 ne
rect -13774 -19462 -11036 -19372
tri -11036 -19462 -10946 -19372 sw
tri -9621 -19462 -9531 -19372 ne
rect -9531 -19462 -6130 -19372
tri -18016 -19628 -17850 -19462 ne
rect -17850 -19628 -15188 -19462
tri -15188 -19628 -15022 -19462 sw
tri -13774 -19628 -13608 -19462 ne
rect -13608 -19628 -10946 -19462
tri -10946 -19628 -10780 -19462 sw
tri -9531 -19628 -9365 -19462 ne
rect -9365 -19628 -6130 -19462
rect -5874 -19628 -5606 -19372
rect -5350 -19628 -5052 -19372
rect -4796 -19628 -4498 -19372
rect -4242 -19628 -3944 -19372
rect -3688 -19628 -3390 -19372
rect -3134 -19628 -2836 -19372
rect -2580 -19628 -2312 -19372
rect -2056 -19628 -1955 -19372
tri -915 -19462 47 -18500 ne
rect 47 -19087 9906 -18500
tri 9906 -19087 10493 -18500 nw
tri 11321 -19087 11908 -18500 se
rect 11908 -19087 13978 -18500
rect 47 -19462 9531 -19087
tri 9531 -19462 9906 -19087 nw
tri 10946 -19462 11321 -19087 se
rect 11321 -19258 13978 -19087
tri 13978 -19258 15220 -18016 nw
tri 15392 -19258 16634 -18016 se
rect 11321 -19462 13774 -19258
tri 13774 -19462 13978 -19258 nw
tri 15188 -19462 15392 -19258 se
rect 15392 -19462 16634 -19258
tri -17850 -19896 -17582 -19628 ne
rect -17582 -19634 -15022 -19628
tri -15022 -19634 -15016 -19628 sw
tri -13608 -19634 -13602 -19628 ne
rect -13602 -19634 -10780 -19628
rect -17582 -19896 -15016 -19634
tri -15016 -19896 -14754 -19634 sw
tri -13602 -19896 -13340 -19634 ne
rect -13340 -19805 -10780 -19634
tri -10780 -19805 -10603 -19628 sw
tri -9365 -19805 -9188 -19628 ne
rect -9188 -19805 -1955 -19628
rect -13340 -19896 -10603 -19805
tri -10603 -19896 -10512 -19805 sw
tri -9188 -19896 -9097 -19805 ne
rect -9097 -19896 -1955 -19805
tri -17582 -20152 -17326 -19896 ne
rect -17326 -20152 -14754 -19896
tri -14754 -20152 -14498 -19896 sw
tri -13340 -20152 -13084 -19896 ne
rect -13084 -20152 -10512 -19896
tri -10512 -20152 -10256 -19896 sw
tri -9097 -20152 -8841 -19896 ne
rect -8841 -20152 -6130 -19896
rect -5874 -20152 -5606 -19896
rect -5350 -20152 -5052 -19896
rect -4796 -20152 -4498 -19896
rect -4242 -20152 -3944 -19896
rect -3688 -20152 -3390 -19896
rect -3134 -20152 -2836 -19896
rect -2580 -20152 -2312 -19896
rect -2056 -20152 -1955 -19896
tri -17326 -20844 -16634 -20152 ne
rect -16634 -20844 -14498 -20152
tri -14498 -20844 -13806 -20152 sw
tri -13084 -20672 -12564 -20152 ne
rect -12564 -20672 -10256 -20152
tri -10256 -20672 -9736 -20152 sw
tri -8841 -20500 -8493 -20152 ne
rect -8493 -20253 -1955 -20152
rect -8493 -20500 -2202 -20253
tri -2202 -20500 -1955 -20253 nw
tri 47 -20500 1085 -19462 ne
rect 1085 -20500 8493 -19462
tri 8493 -20500 9531 -19462 nw
tri 9908 -20500 10946 -19462 se
rect 10946 -20500 12564 -19462
tri 9736 -20672 9908 -20500 se
rect 9908 -20672 12564 -20500
tri 12564 -20672 13774 -19462 nw
tri 13978 -20672 15188 -19462 se
rect 15188 -20672 16634 -19462
tri -12564 -20844 -12392 -20672 ne
rect -12392 -20844 -9736 -20672
tri -9736 -20844 -9564 -20672 sw
tri 9564 -20844 9736 -20672 se
rect 9736 -20844 12392 -20672
tri 12392 -20844 12564 -20672 nw
tri 13806 -20844 13978 -20672 se
rect 13978 -20844 16634 -20672
tri 16634 -20844 19462 -18016 nw
tri -16634 -21848 -15630 -20844 ne
rect -15630 -21048 -13806 -20844
tri -13806 -21048 -13602 -20844 sw
tri -12392 -21048 -12188 -20844 ne
rect -12188 -21048 -9564 -20844
tri -9564 -21048 -9360 -20844 sw
tri 9360 -21048 9564 -20844 se
rect 9564 -21048 11150 -20844
rect -15630 -21848 -13602 -21048
tri -13602 -21848 -12802 -21048 sw
tri -12188 -21848 -11388 -21048 ne
rect -11388 -21500 -9360 -21048
tri -9360 -21500 -8908 -21048 sw
tri 8908 -21500 9360 -21048 se
rect 9360 -21500 11150 -21048
rect -11388 -21848 -1085 -21500
tri -1085 -21848 -737 -21500 sw
tri 1732 -21747 1979 -21500 se
rect 1979 -21747 11150 -21500
rect 1732 -21848 11150 -21747
tri -15630 -22104 -15374 -21848 ne
rect -15374 -22104 -12802 -21848
tri -12802 -22104 -12546 -21848 sw
tri -11388 -22104 -11132 -21848 ne
rect -11132 -22104 -737 -21848
tri -737 -22104 -481 -21848 sw
rect 1732 -22104 1833 -21848
rect 2089 -22104 2357 -21848
rect 2613 -22104 2911 -21848
rect 3167 -22104 3465 -21848
rect 3721 -22104 4019 -21848
rect 4275 -22104 4573 -21848
rect 4829 -22104 5127 -21848
rect 5383 -22104 5651 -21848
rect 5907 -22086 11150 -21848
tri 11150 -22086 12392 -20844 nw
tri 12564 -22086 13806 -20844 se
rect 5907 -22104 10946 -22086
tri -15374 -22290 -15188 -22104 ne
rect -15188 -22290 -12546 -22104
tri -12546 -22290 -12360 -22104 sw
tri -11132 -22290 -10946 -22104 ne
rect -10946 -22290 -481 -22104
tri -481 -22290 -295 -22104 sw
rect 1732 -22290 10946 -22104
tri 10946 -22290 11150 -22086 nw
tri 12360 -22290 12564 -22086 se
rect 12564 -22290 13806 -22086
tri -15188 -22372 -15106 -22290 ne
rect -15106 -22372 -12360 -22290
tri -12360 -22372 -12278 -22290 sw
tri -10946 -22372 -10864 -22290 ne
rect -10864 -22372 -295 -22290
tri -295 -22372 -213 -22290 sw
rect 1732 -22372 9736 -22290
tri -15106 -22628 -14850 -22372 ne
rect -14850 -22462 -12278 -22372
tri -12278 -22462 -12188 -22372 sw
tri -10864 -22462 -10774 -22372 ne
rect -10774 -22462 -213 -22372
rect -14850 -22628 -12188 -22462
tri -12188 -22628 -12022 -22462 sw
tri -10774 -22628 -10608 -22462 ne
rect -10608 -22628 -213 -22462
tri -213 -22628 43 -22372 sw
rect 1732 -22628 1833 -22372
rect 2089 -22628 2357 -22372
rect 2613 -22628 2911 -22372
rect 3167 -22628 3465 -22372
rect 3721 -22628 4019 -22372
rect 4275 -22628 4573 -22372
rect 4829 -22628 5127 -22372
rect 5383 -22628 5651 -22372
rect 5907 -22628 9736 -22372
tri -14850 -22896 -14582 -22628 ne
rect -14582 -22896 -12022 -22628
tri -12022 -22896 -11754 -22628 sw
tri -10608 -22896 -10340 -22628 ne
rect -10340 -22896 43 -22628
tri 43 -22896 311 -22628 sw
rect 1732 -22896 9736 -22628
tri -14582 -23152 -14326 -22896 ne
rect -14326 -23152 -11754 -22896
tri -11754 -23152 -11498 -22896 sw
tri -10340 -23152 -10084 -22896 ne
rect -10084 -23152 311 -22896
tri 311 -23152 567 -22896 sw
rect 1732 -23152 1833 -22896
rect 2089 -23152 2357 -22896
rect 2613 -23152 2911 -22896
rect 3167 -23152 3465 -22896
rect 3721 -23152 4019 -22896
rect 4275 -23152 4573 -22896
rect 4829 -23152 5127 -22896
rect 5383 -23152 5651 -22896
rect 5907 -23152 9736 -22896
tri -14326 -23672 -13806 -23152 ne
rect -13806 -23500 -11498 -23152
tri -11498 -23500 -11150 -23152 sw
tri -10084 -23500 -9736 -23152 ne
rect -9736 -23500 567 -23152
tri 567 -23500 915 -23152 sw
rect 1732 -23253 9736 -23152
tri 1732 -23500 1979 -23253 ne
rect 1979 -23500 9736 -23253
tri 9736 -23500 10946 -22290 nw
tri 11150 -23500 12360 -22290 se
rect 12360 -23500 13806 -22290
rect -13806 -23672 -11150 -23500
tri -11150 -23672 -10978 -23500 sw
tri -1915 -23670 -1745 -23500 ne
rect -1745 -23670 915 -23500
tri 915 -23670 1085 -23500 sw
tri 10980 -23670 11150 -23500 se
rect 11150 -23670 13806 -23500
tri -1745 -23672 -1743 -23670 ne
rect -1743 -23672 1085 -23670
tri 1085 -23672 1087 -23670 sw
tri 10978 -23672 10980 -23670 se
rect 10980 -23672 13806 -23670
tri 13806 -23672 16634 -20844 nw
tri -13806 -24848 -12630 -23672 ne
rect -12630 -24500 -10978 -23672
tri -10978 -24500 -10150 -23672 sw
tri -1743 -24500 -915 -23672 ne
rect -915 -24500 1087 -23672
tri 1087 -24500 1915 -23672 sw
tri 10150 -24500 10978 -23672 se
rect -12630 -24747 -2202 -24500
tri -2202 -24747 -1955 -24500 sw
rect -12630 -24848 -1955 -24747
tri -12630 -25104 -12374 -24848 ne
rect -12374 -25104 -6130 -24848
rect -5874 -25104 -5606 -24848
rect -5350 -25104 -5052 -24848
rect -4796 -25104 -4498 -24848
rect -4242 -25104 -3944 -24848
rect -3688 -25104 -3390 -24848
rect -3134 -25104 -2836 -24848
rect -2580 -25104 -2312 -24848
rect -2056 -25104 -1955 -24848
tri -12374 -25118 -12360 -25104 ne
rect -12360 -25118 -1955 -25104
tri -915 -25118 -297 -24500 ne
rect -297 -25118 10978 -24500
tri -12360 -25372 -12106 -25118 ne
rect -12106 -25372 -1955 -25118
tri -12106 -25628 -11850 -25372 ne
rect -11850 -25628 -6130 -25372
rect -5874 -25628 -5606 -25372
rect -5350 -25628 -5052 -25372
rect -4796 -25628 -4498 -25372
rect -4242 -25628 -3944 -25372
rect -3688 -25628 -3390 -25372
rect -3134 -25628 -2836 -25372
rect -2580 -25628 -2312 -25372
rect -2056 -25628 -1955 -25372
tri -11850 -25896 -11582 -25628 ne
rect -11582 -25896 -1955 -25628
tri -11582 -26152 -11326 -25896 ne
rect -11326 -26152 -6130 -25896
rect -5874 -26152 -5606 -25896
rect -5350 -26152 -5052 -25896
rect -4796 -26152 -4498 -25896
rect -4242 -26152 -3944 -25896
rect -3688 -26152 -3390 -25896
rect -3134 -26152 -2836 -25896
rect -2580 -26152 -2312 -25896
rect -2056 -26152 -1955 -25896
tri -11326 -26500 -10978 -26152 ne
rect -10978 -26253 -1955 -26152
rect -10978 -26500 -2202 -26253
tri -2202 -26500 -1955 -26253 nw
tri -297 -26500 1085 -25118 ne
rect 1085 -26500 10978 -25118
tri 10978 -26500 13806 -23672 nw
<< comment >>
tri -10979 10979 -4548 26500 ne
rect -4548 10979 4548 26500
tri 4548 10979 10979 26500 nw
tri -26500 1884 -4548 10979 sw
tri -4548 1884 -781 10979 ne
rect -781 1884 781 10979
tri 781 1884 4548 10979 nw
tri 4548 1884 26500 10979 se
rect -26500 323 -4548 1884
tri -4548 323 -781 1884 sw
tri -781 323 -134 1884 ne
rect -134 323 134 1884
tri 134 323 781 1884 nw
tri 781 323 4548 1884 se
rect 4548 323 26500 1884
rect -26500 55 -780 323
tri -780 55 -134 323 sw
tri -134 55 -23 323 ne
rect -23 56 23 323
tri 23 56 134 323 nw
tri 134 56 781 323 se
rect 781 56 26500 323
rect -23 55 4 56
rect -26500 9 -134 55
tri -134 9 -23 55 sw
tri -23 9 -4 55 ne
rect -4 10 4 55
tri 4 10 23 56 nw
tri 23 10 134 56 se
rect 134 10 26500 56
rect -4 9 1 10
rect -26500 2 -23 9
tri -23 2 -4 9 sw
tri -4 2 -1 9 ne
rect -1 2 1 9
tri 1 2 4 10 nw
tri 4 2 23 10 se
rect 23 2 26500 10
rect -26500 -2 -4 2
tri -4 0 -1 2 sw
tri -1 0 0 2 ne
tri 0 0 1 2 nw
tri 1 0 4 2 se
rect 4 0 26500 2
tri -4 -2 -1 0 nw
tri -1 -2 0 0 se
tri 0 -1 1 0 ne
rect 1 -1 26500 0
rect -26500 -10 -23 -2
tri -23 -10 -4 -2 nw
tri -4 -10 -1 -2 se
rect -1 -3 0 -2
tri 0 -3 1 -1 sw
tri 1 -3 8 -1 ne
rect 8 -3 26500 -1
rect -1 -10 1 -3
tri 8 -4 9 -3 ne
rect 9 -4 26500 -3
rect -26500 -56 -134 -10
tri -134 -56 -23 -10 nw
tri -23 -56 -4 -10 se
rect -4 -23 1 -10
tri 1 -23 9 -4 sw
tri 9 -23 55 -4 ne
rect 55 -23 26500 -4
rect -4 -56 9 -23
rect -26500 -323 -781 -56
tri -781 -323 -134 -56 nw
tri -134 -323 -23 -56 se
rect -23 -134 9 -56
tri 9 -134 55 -23 sw
tri 55 -134 323 -23 ne
rect 323 -134 26500 -23
rect -23 -323 55 -134
rect -26500 -1884 -4548 -323
tri -4548 -1884 -781 -323 nw
tri -781 -1884 -134 -323 se
rect -134 -780 55 -323
tri 55 -780 323 -134 sw
tri 323 -780 1883 -134 ne
rect 1883 -780 26500 -134
rect -134 -1884 323 -780
tri 1883 -781 1884 -780 ne
rect 1884 -781 26500 -780
tri -26500 -10979 -4548 -1884 nw
tri -4548 -10979 -781 -1884 se
rect -781 -4548 323 -1884
tri 323 -4548 1884 -781 sw
tri 1884 -4548 10979 -781 ne
rect 10979 -4548 26500 -781
rect -781 -10978 1884 -4548
tri 1884 -10978 4548 -4548 sw
rect -781 -10979 4548 -10978
tri 10979 -10979 26500 -4548 ne
tri -10979 -26500 -4548 -10979 se
rect -4548 -26500 4548 -10979
tri 4548 -26500 10979 -10979 sw
<< properties >>
string GDS_END 10508074
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10489606
string gencell sky130_fd_pr__rf_test_coil2
string library sky130
string parameter m=1
string path 637.500 -274.450 637.500 -75.000 
<< end >>
