magic
tech sky130B
timestamp 1644511149
<< properties >>
string GDS_END 5606734
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 5603850
<< end >>
