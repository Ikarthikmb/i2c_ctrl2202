magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 29 -17 63 21
<< locali >>
rect 29 299 386 335
rect 29 207 129 299
rect 163 199 285 265
rect 321 249 386 299
rect 321 215 387 249
rect 463 157 523 423
rect 560 199 615 325
rect 191 123 523 157
rect 191 51 260 123
rect 459 51 523 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 22 421 74 493
rect 108 455 174 527
rect 210 421 244 493
rect 295 439 329 527
rect 363 457 618 493
rect 22 405 244 421
rect 363 405 429 457
rect 22 371 429 405
rect 20 17 79 173
rect 557 359 618 457
rect 352 17 418 89
rect 559 17 625 165
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 163 199 285 265 6 A1
port 1 nsew signal input
rlabel locali s 321 215 387 249 6 A2
port 2 nsew signal input
rlabel locali s 321 249 386 299 6 A2
port 2 nsew signal input
rlabel locali s 29 207 129 299 6 A2
port 2 nsew signal input
rlabel locali s 29 299 386 335 6 A2
port 2 nsew signal input
rlabel locali s 560 199 615 325 6 B1
port 3 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 643 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 459 51 523 123 6 Y
port 8 nsew signal output
rlabel locali s 191 51 260 123 6 Y
port 8 nsew signal output
rlabel locali s 191 123 523 157 6 Y
port 8 nsew signal output
rlabel locali s 463 157 523 423 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4034326
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4028462
<< end >>
