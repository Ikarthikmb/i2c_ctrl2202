magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 317 157 917 203
rect 1 139 917 157
rect 1 67 919 139
rect 1 21 315 67
rect 733 29 919 67
rect 733 21 917 29
rect 29 -17 63 21
<< locali >>
rect 85 325 155 391
rect 121 189 245 223
rect 121 153 163 189
rect 579 265 616 327
rect 670 265 709 327
rect 579 199 625 265
rect 670 199 721 265
rect 579 83 616 199
rect 670 84 709 199
rect 851 51 903 493
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 427 69 493
rect 131 451 197 527
rect 17 291 51 427
rect 245 417 283 493
rect 333 451 399 527
rect 441 417 475 493
rect 514 451 580 527
rect 632 417 666 493
rect 751 451 817 527
rect 245 383 393 417
rect 209 315 325 349
rect 209 291 243 315
rect 17 257 243 291
rect 359 281 393 383
rect 17 117 51 257
rect 279 247 393 281
rect 427 383 817 417
rect 279 151 313 247
rect 427 185 461 383
rect 17 51 69 117
rect 131 17 197 93
rect 233 85 313 151
rect 351 119 461 185
rect 495 85 529 265
rect 233 51 529 85
rect 783 199 817 383
rect 751 17 817 93
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 85 325 155 391 6 A_N
port 1 nsew signal input
rlabel locali s 121 153 163 189 6 B_N
port 2 nsew signal input
rlabel locali s 121 189 245 223 6 B_N
port 2 nsew signal input
rlabel locali s 579 83 616 199 6 C
port 3 nsew signal input
rlabel locali s 579 199 625 265 6 C
port 3 nsew signal input
rlabel locali s 579 265 616 327 6 C
port 3 nsew signal input
rlabel locali s 670 84 709 199 6 D
port 4 nsew signal input
rlabel locali s 670 199 721 265 6 D
port 4 nsew signal input
rlabel locali s 670 265 709 327 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 733 21 917 29 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 733 29 919 67 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 315 67 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 67 919 139 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 139 917 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 317 157 917 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 851 51 903 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 920 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3066900
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3058560
<< end >>
