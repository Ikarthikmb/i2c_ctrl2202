magic
tech sky130A
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdfl1sd2__example_55959141808306  sky130_fd_pr__hvdfl1sd2__example_55959141808306_0
timestamp 1644511149
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808306  sky130_fd_pr__hvdfl1sd2__example_55959141808306_1
timestamp 1644511149
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808306  sky130_fd_pr__hvdfl1sd2__example_55959141808306_2
timestamp 1644511149
transform 1 0 472 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808306  sky130_fd_pr__hvdfl1sd2__example_55959141808306_3
timestamp 1644511149
transform 1 0 648 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808306  sky130_fd_pr__hvdfl1sd2__example_55959141808306_4
timestamp 1644511149
transform 1 0 824 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808115  sky130_fd_pr__hvdfl1sd__example_55959141808115_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808115  sky130_fd_pr__hvdfl1sd__example_55959141808115_1
timestamp 1644511149
transform 1 0 1000 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 1028 267 1028 267 0 FreeSans 300 0 0 0 S
flabel comment s 852 267 852 267 0 FreeSans 300 0 0 0 D
flabel comment s 676 267 676 267 0 FreeSans 300 0 0 0 S
flabel comment s 500 267 500 267 0 FreeSans 300 0 0 0 D
flabel comment s 324 267 324 267 0 FreeSans 300 0 0 0 S
flabel comment s 148 267 148 267 0 FreeSans 300 0 0 0 D
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7013998
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7010482
<< end >>
