/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/cap_mim_m3/sky130_fd_pr__cap_mim_m3_2.model.spice