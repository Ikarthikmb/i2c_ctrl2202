magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< pwell >>
rect 15 163 615 1225
<< nmoslvt >>
rect 171 189 201 1199
rect 257 189 287 1199
rect 343 189 373 1199
rect 429 189 459 1199
<< ndiff >>
rect 111 1187 171 1199
rect 111 1153 126 1187
rect 160 1153 171 1187
rect 111 1119 171 1153
rect 111 1085 126 1119
rect 160 1085 171 1119
rect 111 1051 171 1085
rect 111 1017 126 1051
rect 160 1017 171 1051
rect 111 983 171 1017
rect 111 949 126 983
rect 160 949 171 983
rect 111 915 171 949
rect 111 881 126 915
rect 160 881 171 915
rect 111 847 171 881
rect 111 813 126 847
rect 160 813 171 847
rect 111 779 171 813
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 1187 257 1199
rect 201 889 212 1187
rect 246 889 257 1187
rect 201 843 257 889
rect 201 545 212 843
rect 246 545 257 843
rect 201 499 257 545
rect 201 201 212 499
rect 246 201 257 499
rect 201 189 257 201
rect 287 1187 343 1199
rect 287 889 298 1187
rect 332 889 343 1187
rect 287 843 343 889
rect 287 545 298 843
rect 332 545 343 843
rect 287 499 343 545
rect 287 201 298 499
rect 332 201 343 499
rect 287 189 343 201
rect 373 1187 429 1199
rect 373 889 384 1187
rect 418 889 429 1187
rect 373 843 429 889
rect 373 545 384 843
rect 418 545 429 843
rect 373 499 429 545
rect 373 201 384 499
rect 418 201 429 499
rect 373 189 429 201
rect 459 1187 519 1199
rect 459 1153 470 1187
rect 504 1153 519 1187
rect 459 1119 519 1153
rect 459 1085 470 1119
rect 504 1085 519 1119
rect 459 1051 519 1085
rect 459 1017 470 1051
rect 504 1017 519 1051
rect 459 983 519 1017
rect 459 949 470 983
rect 504 949 519 983
rect 459 915 519 949
rect 459 881 470 915
rect 504 881 519 915
rect 459 847 519 881
rect 459 813 470 847
rect 504 813 519 847
rect 459 779 519 813
rect 459 745 470 779
rect 504 745 519 779
rect 459 711 519 745
rect 459 677 470 711
rect 504 677 519 711
rect 459 643 519 677
rect 459 609 470 643
rect 504 609 519 643
rect 459 575 519 609
rect 459 541 470 575
rect 504 541 519 575
rect 459 507 519 541
rect 459 473 470 507
rect 504 473 519 507
rect 459 439 519 473
rect 459 405 470 439
rect 504 405 519 439
rect 459 371 519 405
rect 459 337 470 371
rect 504 337 519 371
rect 459 303 519 337
rect 459 269 470 303
rect 504 269 519 303
rect 459 235 519 269
rect 459 201 470 235
rect 504 201 519 235
rect 459 189 519 201
<< ndiffc >>
rect 126 1153 160 1187
rect 126 1085 160 1119
rect 126 1017 160 1051
rect 126 949 160 983
rect 126 881 160 915
rect 126 813 160 847
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 889 246 1187
rect 212 545 246 843
rect 212 201 246 499
rect 298 889 332 1187
rect 298 545 332 843
rect 298 201 332 499
rect 384 889 418 1187
rect 384 545 418 843
rect 384 201 418 499
rect 470 1153 504 1187
rect 470 1085 504 1119
rect 470 1017 504 1051
rect 470 949 504 983
rect 470 881 504 915
rect 470 813 504 847
rect 470 745 504 779
rect 470 677 504 711
rect 470 609 504 643
rect 470 541 504 575
rect 470 473 504 507
rect 470 405 504 439
rect 470 337 504 371
rect 470 269 504 303
rect 470 201 504 235
<< psubdiff >>
rect 41 1187 111 1199
rect 41 1153 58 1187
rect 92 1153 111 1187
rect 41 1119 111 1153
rect 41 1085 58 1119
rect 92 1085 111 1119
rect 41 1051 111 1085
rect 41 1017 58 1051
rect 92 1017 111 1051
rect 41 983 111 1017
rect 41 949 58 983
rect 92 949 111 983
rect 41 915 111 949
rect 41 881 58 915
rect 92 881 111 915
rect 41 847 111 881
rect 41 813 58 847
rect 92 813 111 847
rect 41 779 111 813
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 519 1187 589 1199
rect 519 1153 538 1187
rect 572 1153 589 1187
rect 519 1119 589 1153
rect 519 1085 538 1119
rect 572 1085 589 1119
rect 519 1051 589 1085
rect 519 1017 538 1051
rect 572 1017 589 1051
rect 519 983 589 1017
rect 519 949 538 983
rect 572 949 589 983
rect 519 915 589 949
rect 519 881 538 915
rect 572 881 589 915
rect 519 847 589 881
rect 519 813 538 847
rect 572 813 589 847
rect 519 779 589 813
rect 519 745 538 779
rect 572 745 589 779
rect 519 711 589 745
rect 519 677 538 711
rect 572 677 589 711
rect 519 643 589 677
rect 519 609 538 643
rect 572 609 589 643
rect 519 575 589 609
rect 519 541 538 575
rect 572 541 589 575
rect 519 507 589 541
rect 519 473 538 507
rect 572 473 589 507
rect 519 439 589 473
rect 519 405 538 439
rect 572 405 589 439
rect 519 371 589 405
rect 519 337 538 371
rect 572 337 589 371
rect 519 303 589 337
rect 519 269 538 303
rect 572 269 589 303
rect 519 235 589 269
rect 519 201 538 235
rect 572 201 589 235
rect 519 189 589 201
<< psubdiffcont >>
rect 58 1153 92 1187
rect 58 1085 92 1119
rect 58 1017 92 1051
rect 58 949 92 983
rect 58 881 92 915
rect 58 813 92 847
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 538 1153 572 1187
rect 538 1085 572 1119
rect 538 1017 572 1051
rect 538 949 572 983
rect 538 881 572 915
rect 538 813 572 847
rect 538 745 572 779
rect 538 677 572 711
rect 538 609 572 643
rect 538 541 572 575
rect 538 473 572 507
rect 538 405 572 439
rect 538 337 572 371
rect 538 269 572 303
rect 538 201 572 235
<< poly >>
rect 243 1299 387 1315
rect 120 1275 201 1291
rect 120 1241 136 1275
rect 170 1241 201 1275
rect 243 1265 264 1299
rect 366 1265 387 1299
rect 243 1249 387 1265
rect 429 1275 510 1291
rect 120 1225 201 1241
rect 171 1199 201 1225
rect 257 1199 287 1249
rect 343 1199 373 1249
rect 429 1241 460 1275
rect 494 1241 510 1275
rect 429 1225 510 1241
rect 429 1199 459 1225
rect 171 163 201 189
rect 120 147 201 163
rect 120 113 136 147
rect 170 113 201 147
rect 257 139 287 189
rect 343 139 373 189
rect 429 163 459 189
rect 429 147 510 163
rect 120 97 201 113
rect 243 123 387 139
rect 243 89 264 123
rect 366 89 387 123
rect 429 113 460 147
rect 494 113 510 147
rect 429 97 510 113
rect 243 73 387 89
<< polycont >>
rect 136 1241 170 1275
rect 264 1265 366 1299
rect 460 1241 494 1275
rect 136 113 170 147
rect 264 89 366 123
rect 460 113 494 147
<< locali >>
rect 248 1369 382 1388
rect 120 1275 186 1291
rect 120 1241 136 1275
rect 170 1241 186 1275
rect 248 1263 262 1369
rect 368 1263 382 1369
rect 248 1249 382 1263
rect 444 1275 510 1291
rect 120 1225 186 1241
rect 444 1241 460 1275
rect 494 1241 510 1275
rect 444 1225 510 1241
rect 120 1203 160 1225
rect 470 1203 510 1225
rect 41 1187 160 1203
rect 41 1153 58 1187
rect 92 1179 126 1187
rect 94 1153 126 1179
rect 41 1145 60 1153
rect 94 1145 160 1153
rect 41 1119 160 1145
rect 41 1085 58 1119
rect 92 1107 126 1119
rect 94 1085 126 1107
rect 41 1073 60 1085
rect 94 1073 160 1085
rect 41 1051 160 1073
rect 41 1017 58 1051
rect 92 1035 126 1051
rect 94 1017 126 1035
rect 41 1001 60 1017
rect 94 1001 160 1017
rect 41 983 160 1001
rect 41 949 58 983
rect 92 963 126 983
rect 94 949 126 963
rect 41 929 60 949
rect 94 929 160 949
rect 41 915 160 929
rect 41 881 58 915
rect 92 891 126 915
rect 94 881 126 891
rect 41 857 60 881
rect 94 857 160 881
rect 41 847 160 857
rect 41 813 58 847
rect 92 819 126 847
rect 94 813 126 819
rect 41 785 60 813
rect 94 785 160 813
rect 41 779 160 785
rect 41 745 58 779
rect 92 747 126 779
rect 94 745 126 747
rect 41 713 60 745
rect 94 713 160 745
rect 41 711 160 713
rect 41 677 58 711
rect 92 677 126 711
rect 41 675 160 677
rect 41 643 60 675
rect 94 643 160 675
rect 41 609 58 643
rect 94 641 126 643
rect 92 609 126 641
rect 41 603 160 609
rect 41 575 60 603
rect 94 575 160 603
rect 41 541 58 575
rect 94 569 126 575
rect 92 541 126 569
rect 41 531 160 541
rect 41 507 60 531
rect 94 507 160 531
rect 41 473 58 507
rect 94 497 126 507
rect 92 473 126 497
rect 41 459 160 473
rect 41 439 60 459
rect 94 439 160 459
rect 41 405 58 439
rect 94 425 126 439
rect 92 405 126 425
rect 41 387 160 405
rect 41 371 60 387
rect 94 371 160 387
rect 41 337 58 371
rect 94 353 126 371
rect 92 337 126 353
rect 41 315 160 337
rect 41 303 60 315
rect 94 303 160 315
rect 41 269 58 303
rect 94 281 126 303
rect 92 269 126 281
rect 41 243 160 269
rect 41 235 60 243
rect 94 235 160 243
rect 41 201 58 235
rect 94 209 126 235
rect 92 201 126 209
rect 41 185 160 201
rect 212 1187 246 1203
rect 212 843 246 857
rect 212 531 246 545
rect 212 185 246 201
rect 298 1187 332 1203
rect 298 843 332 857
rect 298 531 332 545
rect 298 185 332 201
rect 384 1187 418 1203
rect 384 843 418 857
rect 384 531 418 545
rect 384 185 418 201
rect 470 1187 589 1203
rect 504 1179 538 1187
rect 504 1153 536 1179
rect 572 1153 589 1187
rect 470 1145 536 1153
rect 570 1145 589 1153
rect 470 1119 589 1145
rect 504 1107 538 1119
rect 504 1085 536 1107
rect 572 1085 589 1119
rect 470 1073 536 1085
rect 570 1073 589 1085
rect 470 1051 589 1073
rect 504 1035 538 1051
rect 504 1017 536 1035
rect 572 1017 589 1051
rect 470 1001 536 1017
rect 570 1001 589 1017
rect 470 983 589 1001
rect 504 963 538 983
rect 504 949 536 963
rect 572 949 589 983
rect 470 929 536 949
rect 570 929 589 949
rect 470 915 589 929
rect 504 891 538 915
rect 504 881 536 891
rect 572 881 589 915
rect 470 857 536 881
rect 570 857 589 881
rect 470 847 589 857
rect 504 819 538 847
rect 504 813 536 819
rect 572 813 589 847
rect 470 785 536 813
rect 570 785 589 813
rect 470 779 589 785
rect 504 747 538 779
rect 504 745 536 747
rect 572 745 589 779
rect 470 713 536 745
rect 570 713 589 745
rect 470 711 589 713
rect 504 677 538 711
rect 572 677 589 711
rect 470 675 589 677
rect 470 643 536 675
rect 570 643 589 675
rect 504 641 536 643
rect 504 609 538 641
rect 572 609 589 643
rect 470 603 589 609
rect 470 575 536 603
rect 570 575 589 603
rect 504 569 536 575
rect 504 541 538 569
rect 572 541 589 575
rect 470 531 589 541
rect 470 507 536 531
rect 570 507 589 531
rect 504 497 536 507
rect 504 473 538 497
rect 572 473 589 507
rect 470 459 589 473
rect 470 439 536 459
rect 570 439 589 459
rect 504 425 536 439
rect 504 405 538 425
rect 572 405 589 439
rect 470 387 589 405
rect 470 371 536 387
rect 570 371 589 387
rect 504 353 536 371
rect 504 337 538 353
rect 572 337 589 371
rect 470 315 589 337
rect 470 303 536 315
rect 570 303 589 315
rect 504 281 536 303
rect 504 269 538 281
rect 572 269 589 303
rect 470 243 589 269
rect 470 235 536 243
rect 570 235 589 243
rect 504 209 536 235
rect 504 201 538 209
rect 572 201 589 235
rect 470 185 589 201
rect 120 163 160 185
rect 470 163 510 185
rect 120 147 186 163
rect 120 113 136 147
rect 170 113 186 147
rect 444 147 510 163
rect 120 97 186 113
rect 248 125 382 139
rect 248 19 262 125
rect 368 19 382 125
rect 444 113 460 147
rect 494 113 510 147
rect 444 97 510 113
rect 248 0 382 19
<< viali >>
rect 262 1299 368 1369
rect 262 1265 264 1299
rect 264 1265 366 1299
rect 366 1265 368 1299
rect 262 1263 368 1265
rect 60 1153 92 1179
rect 92 1153 94 1179
rect 60 1145 94 1153
rect 60 1085 92 1107
rect 92 1085 94 1107
rect 60 1073 94 1085
rect 60 1017 92 1035
rect 92 1017 94 1035
rect 60 1001 94 1017
rect 60 949 92 963
rect 92 949 94 963
rect 60 929 94 949
rect 60 881 92 891
rect 92 881 94 891
rect 60 857 94 881
rect 60 813 92 819
rect 92 813 94 819
rect 60 785 94 813
rect 60 745 92 747
rect 92 745 94 747
rect 60 713 94 745
rect 60 643 94 675
rect 60 641 92 643
rect 92 641 94 643
rect 60 575 94 603
rect 60 569 92 575
rect 92 569 94 575
rect 60 507 94 531
rect 60 497 92 507
rect 92 497 94 507
rect 60 439 94 459
rect 60 425 92 439
rect 92 425 94 439
rect 60 371 94 387
rect 60 353 92 371
rect 92 353 94 371
rect 60 303 94 315
rect 60 281 92 303
rect 92 281 94 303
rect 60 235 94 243
rect 60 209 92 235
rect 92 209 94 235
rect 212 1145 246 1179
rect 212 1073 246 1107
rect 212 1001 246 1035
rect 212 929 246 963
rect 212 889 246 891
rect 212 857 246 889
rect 212 785 246 819
rect 212 713 246 747
rect 212 641 246 675
rect 212 569 246 603
rect 212 499 246 531
rect 212 497 246 499
rect 212 425 246 459
rect 212 353 246 387
rect 212 281 246 315
rect 212 209 246 243
rect 298 1145 332 1179
rect 298 1073 332 1107
rect 298 1001 332 1035
rect 298 929 332 963
rect 298 889 332 891
rect 298 857 332 889
rect 298 785 332 819
rect 298 713 332 747
rect 298 641 332 675
rect 298 569 332 603
rect 298 499 332 531
rect 298 497 332 499
rect 298 425 332 459
rect 298 353 332 387
rect 298 281 332 315
rect 298 209 332 243
rect 384 1145 418 1179
rect 384 1073 418 1107
rect 384 1001 418 1035
rect 384 929 418 963
rect 384 889 418 891
rect 384 857 418 889
rect 384 785 418 819
rect 384 713 418 747
rect 384 641 418 675
rect 384 569 418 603
rect 384 499 418 531
rect 384 497 418 499
rect 384 425 418 459
rect 384 353 418 387
rect 384 281 418 315
rect 384 209 418 243
rect 536 1153 538 1179
rect 538 1153 570 1179
rect 536 1145 570 1153
rect 536 1085 538 1107
rect 538 1085 570 1107
rect 536 1073 570 1085
rect 536 1017 538 1035
rect 538 1017 570 1035
rect 536 1001 570 1017
rect 536 949 538 963
rect 538 949 570 963
rect 536 929 570 949
rect 536 881 538 891
rect 538 881 570 891
rect 536 857 570 881
rect 536 813 538 819
rect 538 813 570 819
rect 536 785 570 813
rect 536 745 538 747
rect 538 745 570 747
rect 536 713 570 745
rect 536 643 570 675
rect 536 641 538 643
rect 538 641 570 643
rect 536 575 570 603
rect 536 569 538 575
rect 538 569 570 575
rect 536 507 570 531
rect 536 497 538 507
rect 538 497 570 507
rect 536 439 570 459
rect 536 425 538 439
rect 538 425 570 439
rect 536 371 570 387
rect 536 353 538 371
rect 538 353 570 371
rect 536 303 570 315
rect 536 281 538 303
rect 538 281 570 303
rect 536 235 570 243
rect 536 209 538 235
rect 538 209 570 235
rect 262 123 368 125
rect 262 89 264 123
rect 264 89 366 123
rect 366 89 368 123
rect 262 19 368 89
<< metal1 >>
rect 250 1369 380 1388
rect 250 1263 262 1369
rect 368 1263 380 1369
rect 250 1251 380 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 203 1179 255 1191
rect 203 1145 212 1179
rect 246 1145 255 1179
rect 203 1107 255 1145
rect 203 1073 212 1107
rect 246 1073 255 1107
rect 203 1035 255 1073
rect 203 1001 212 1035
rect 246 1001 255 1035
rect 203 963 255 1001
rect 203 929 212 963
rect 246 929 255 963
rect 203 891 255 929
rect 203 857 212 891
rect 246 857 255 891
rect 203 819 255 857
rect 203 785 212 819
rect 246 785 255 819
rect 203 747 255 785
rect 203 713 212 747
rect 246 713 255 747
rect 203 675 255 713
rect 203 641 212 675
rect 246 641 255 675
rect 203 639 255 641
rect 203 575 212 587
rect 246 575 255 587
rect 203 511 212 523
rect 246 511 255 523
rect 203 447 212 459
rect 246 447 255 459
rect 203 387 255 395
rect 203 383 212 387
rect 246 383 255 387
rect 203 319 255 331
rect 203 255 255 267
rect 203 197 255 203
rect 289 1185 341 1191
rect 289 1121 341 1133
rect 289 1057 341 1069
rect 289 1001 298 1005
rect 332 1001 341 1005
rect 289 993 341 1001
rect 289 929 298 941
rect 332 929 341 941
rect 289 865 298 877
rect 332 865 341 877
rect 289 801 298 813
rect 332 801 341 813
rect 289 747 341 749
rect 289 713 298 747
rect 332 713 341 747
rect 289 675 341 713
rect 289 641 298 675
rect 332 641 341 675
rect 289 603 341 641
rect 289 569 298 603
rect 332 569 341 603
rect 289 531 341 569
rect 289 497 298 531
rect 332 497 341 531
rect 289 459 341 497
rect 289 425 298 459
rect 332 425 341 459
rect 289 387 341 425
rect 289 353 298 387
rect 332 353 341 387
rect 289 315 341 353
rect 289 281 298 315
rect 332 281 341 315
rect 289 243 341 281
rect 289 209 298 243
rect 332 209 341 243
rect 289 197 341 209
rect 375 1179 427 1191
rect 375 1145 384 1179
rect 418 1145 427 1179
rect 375 1107 427 1145
rect 375 1073 384 1107
rect 418 1073 427 1107
rect 375 1035 427 1073
rect 375 1001 384 1035
rect 418 1001 427 1035
rect 375 963 427 1001
rect 375 929 384 963
rect 418 929 427 963
rect 375 891 427 929
rect 375 857 384 891
rect 418 857 427 891
rect 375 819 427 857
rect 375 785 384 819
rect 418 785 427 819
rect 375 747 427 785
rect 375 713 384 747
rect 418 713 427 747
rect 375 675 427 713
rect 375 641 384 675
rect 418 641 427 675
rect 375 639 427 641
rect 375 575 384 587
rect 418 575 427 587
rect 375 511 384 523
rect 418 511 427 523
rect 375 447 384 459
rect 418 447 427 459
rect 375 387 427 395
rect 375 383 384 387
rect 418 383 427 387
rect 375 319 427 331
rect 375 255 427 267
rect 375 197 427 203
rect 530 1179 589 1191
rect 530 1145 536 1179
rect 570 1145 589 1179
rect 530 1107 589 1145
rect 530 1073 536 1107
rect 570 1073 589 1107
rect 530 1035 589 1073
rect 530 1001 536 1035
rect 570 1001 589 1035
rect 530 963 589 1001
rect 530 929 536 963
rect 570 929 589 963
rect 530 891 589 929
rect 530 857 536 891
rect 570 857 589 891
rect 530 819 589 857
rect 530 785 536 819
rect 570 785 589 819
rect 530 747 589 785
rect 530 713 536 747
rect 570 713 589 747
rect 530 675 589 713
rect 530 641 536 675
rect 570 641 589 675
rect 530 603 589 641
rect 530 569 536 603
rect 570 569 589 603
rect 530 531 589 569
rect 530 497 536 531
rect 570 497 589 531
rect 530 459 589 497
rect 530 425 536 459
rect 570 425 589 459
rect 530 387 589 425
rect 530 353 536 387
rect 570 353 589 387
rect 530 315 589 353
rect 530 281 536 315
rect 570 281 589 315
rect 530 243 589 281
rect 530 209 536 243
rect 570 209 589 243
rect 530 197 589 209
rect 250 125 380 137
rect 250 19 262 125
rect 368 19 380 125
rect 250 0 380 19
<< via1 >>
rect 203 603 255 639
rect 203 587 212 603
rect 212 587 246 603
rect 246 587 255 603
rect 203 569 212 575
rect 212 569 246 575
rect 246 569 255 575
rect 203 531 255 569
rect 203 523 212 531
rect 212 523 246 531
rect 246 523 255 531
rect 203 497 212 511
rect 212 497 246 511
rect 246 497 255 511
rect 203 459 255 497
rect 203 425 212 447
rect 212 425 246 447
rect 246 425 255 447
rect 203 395 255 425
rect 203 353 212 383
rect 212 353 246 383
rect 246 353 255 383
rect 203 331 255 353
rect 203 315 255 319
rect 203 281 212 315
rect 212 281 246 315
rect 246 281 255 315
rect 203 267 255 281
rect 203 243 255 255
rect 203 209 212 243
rect 212 209 246 243
rect 246 209 255 243
rect 203 203 255 209
rect 289 1179 341 1185
rect 289 1145 298 1179
rect 298 1145 332 1179
rect 332 1145 341 1179
rect 289 1133 341 1145
rect 289 1107 341 1121
rect 289 1073 298 1107
rect 298 1073 332 1107
rect 332 1073 341 1107
rect 289 1069 341 1073
rect 289 1035 341 1057
rect 289 1005 298 1035
rect 298 1005 332 1035
rect 332 1005 341 1035
rect 289 963 341 993
rect 289 941 298 963
rect 298 941 332 963
rect 332 941 341 963
rect 289 891 341 929
rect 289 877 298 891
rect 298 877 332 891
rect 332 877 341 891
rect 289 857 298 865
rect 298 857 332 865
rect 332 857 341 865
rect 289 819 341 857
rect 289 813 298 819
rect 298 813 332 819
rect 332 813 341 819
rect 289 785 298 801
rect 298 785 332 801
rect 332 785 341 801
rect 289 749 341 785
rect 375 603 427 639
rect 375 587 384 603
rect 384 587 418 603
rect 418 587 427 603
rect 375 569 384 575
rect 384 569 418 575
rect 418 569 427 575
rect 375 531 427 569
rect 375 523 384 531
rect 384 523 418 531
rect 418 523 427 531
rect 375 497 384 511
rect 384 497 418 511
rect 418 497 427 511
rect 375 459 427 497
rect 375 425 384 447
rect 384 425 418 447
rect 418 425 427 447
rect 375 395 427 425
rect 375 353 384 383
rect 384 353 418 383
rect 418 353 427 383
rect 375 331 427 353
rect 375 315 427 319
rect 375 281 384 315
rect 384 281 418 315
rect 418 281 427 315
rect 375 267 427 281
rect 375 243 427 255
rect 375 209 384 243
rect 384 209 418 243
rect 418 209 427 243
rect 375 203 427 209
<< metal2 >>
rect 14 1185 616 1191
rect 14 1133 289 1185
rect 341 1133 616 1185
rect 14 1121 616 1133
rect 14 1069 289 1121
rect 341 1069 616 1121
rect 14 1057 616 1069
rect 14 1005 289 1057
rect 341 1005 616 1057
rect 14 993 616 1005
rect 14 941 289 993
rect 341 941 616 993
rect 14 929 616 941
rect 14 877 289 929
rect 341 877 616 929
rect 14 865 616 877
rect 14 813 289 865
rect 341 813 616 865
rect 14 801 616 813
rect 14 749 289 801
rect 341 749 616 801
rect 14 719 616 749
rect 14 639 616 669
rect 14 587 203 639
rect 255 587 375 639
rect 427 587 616 639
rect 14 575 616 587
rect 14 523 203 575
rect 255 523 375 575
rect 427 523 616 575
rect 14 511 616 523
rect 14 459 203 511
rect 255 459 375 511
rect 427 459 616 511
rect 14 447 616 459
rect 14 395 203 447
rect 255 395 375 447
rect 427 395 616 447
rect 14 383 616 395
rect 14 331 203 383
rect 255 331 375 383
rect 427 331 616 383
rect 14 319 616 331
rect 14 267 203 319
rect 255 267 375 319
rect 427 267 616 319
rect 14 255 616 267
rect 14 203 203 255
rect 255 203 375 255
rect 427 203 616 255
rect 14 197 616 203
<< labels >>
flabel comment s 184 736 184 736 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 441 740 441 740 0 FreeSans 180 90 0 0 dummy_poly
flabel metal1 s 255 1288 374 1339 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 255 44 374 95 0 FreeSans 200 0 0 0 GATE
port 1 nsew
flabel metal1 s 530 683 589 713 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal1 s 41 675 100 705 0 FreeSans 200 90 0 0 SUBSTRATE
port 2 nsew
flabel metal2 s 14 384 35 512 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 908 35 1036 7 FreeSans 300 180 0 0 DRAIN
port 4 nsew
<< properties >>
string GDS_END 6673730
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6656322
<< end >>
