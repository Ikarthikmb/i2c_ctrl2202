/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pnp_05v5/sky130_fd_pr__pnp_05v5_W3p40L3p40.spice