magic
tech sky130A
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_0
timestamp 1644511149
transform 1 0 120 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_1
timestamp 1644511149
transform 1 0 296 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_2
timestamp 1644511149
transform 1 0 472 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_3
timestamp 1644511149
transform 1 0 648 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_4
timestamp 1644511149
transform 1 0 824 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd2__example_5595914180869  sky130_fd_pr__dfl1sd2__example_5595914180869_5
timestamp 1644511149
transform 1 0 1000 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180868  sky130_fd_pr__dfl1sd__example_5595914180868_1
timestamp 1644511149
transform 1 0 1176 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 1204 29 1204 29 0 FreeSans 300 0 0 0 D
flabel comment s 1028 29 1028 29 0 FreeSans 300 0 0 0 S
flabel comment s 852 29 852 29 0 FreeSans 300 0 0 0 D
flabel comment s 676 29 676 29 0 FreeSans 300 0 0 0 S
flabel comment s 500 29 500 29 0 FreeSans 300 0 0 0 D
flabel comment s 324 29 324 29 0 FreeSans 300 0 0 0 S
flabel comment s 148 29 148 29 0 FreeSans 300 0 0 0 D
flabel comment s -28 29 -28 29 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 8185280
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8181274
<< end >>
