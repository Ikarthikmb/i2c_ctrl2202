magic
tech sky130B
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_0
timestamp 1644511149
transform 1 0 581 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_1
timestamp 1644511149
transform 1 0 1501 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_2
timestamp 1644511149
transform 1 0 2421 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_3
timestamp 1644511149
transform 1 0 3341 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_4
timestamp 1644511149
transform 1 0 4261 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_5
timestamp 1644511149
transform 1 0 5181 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_6
timestamp 1644511149
transform 1 0 6101 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_7
timestamp 1644511149
transform 1 0 7021 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_8
timestamp 1644511149
transform 1 0 7941 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s2__example_55959141808672  sky130_fd_pr__hvdftpl1s2__example_55959141808672_9
timestamp 1644511149
transform 1 0 8861 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s__example_55959141808671  sky130_fd_pr__hvdftpl1s__example_55959141808671_0
timestamp 1644511149
transform -1 0 -79 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdftpl1s__example_55959141808671  sky130_fd_pr__hvdftpl1s__example_55959141808671_1
timestamp 1644511149
transform 1 0 9781 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 9843 1973 9843 1973 0 FreeSans 300 0 0 0 S
flabel comment s 9451 2000 9451 2000 0 FreeSans 300 0 0 0 D
flabel comment s 8991 1967 8991 1967 0 FreeSans 300 0 0 0 S
flabel comment s 8531 2000 8531 2000 0 FreeSans 300 0 0 0 D
flabel comment s 8071 1967 8071 1967 0 FreeSans 300 0 0 0 S
flabel comment s 7611 2000 7611 2000 0 FreeSans 300 0 0 0 D
flabel comment s 7151 1967 7151 1967 0 FreeSans 300 0 0 0 S
flabel comment s 6691 2000 6691 2000 0 FreeSans 300 0 0 0 D
flabel comment s 6231 1967 6231 1967 0 FreeSans 300 0 0 0 S
flabel comment s 5771 2000 5771 2000 0 FreeSans 300 0 0 0 D
flabel comment s 5311 1967 5311 1967 0 FreeSans 300 0 0 0 S
flabel comment s 4851 2000 4851 2000 0 FreeSans 300 0 0 0 D
flabel comment s 4391 1967 4391 1967 0 FreeSans 300 0 0 0 S
flabel comment s 3931 2000 3931 2000 0 FreeSans 300 0 0 0 D
flabel comment s 3471 1967 3471 1967 0 FreeSans 300 0 0 0 S
flabel comment s 3011 2000 3011 2000 0 FreeSans 300 0 0 0 D
flabel comment s 2551 1967 2551 1967 0 FreeSans 300 0 0 0 S
flabel comment s 2091 2000 2091 2000 0 FreeSans 300 0 0 0 D
flabel comment s 1631 1967 1631 1967 0 FreeSans 300 0 0 0 S
flabel comment s 1171 2000 1171 2000 0 FreeSans 300 0 0 0 D
flabel comment s 711 1967 711 1967 0 FreeSans 300 0 0 0 S
flabel comment s 251 2000 251 2000 0 FreeSans 300 0 0 0 D
flabel comment s -141 1973 -141 1973 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 11273402
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 11261682
<< end >>
