/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield/sky130_fd_pr__cap_vpp_11p5x11p7_pol1m1m2m3m4m5_noshield.spice