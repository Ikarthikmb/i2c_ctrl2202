magic
tech sky130B
timestamp 1644511149
<< properties >>
string GDS_END 30691476
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30688144
<< end >>
