magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< locali >>
rect 50 4758 84 4824
<< obsli1 >>
rect 0 2272 2282 2338
rect 0 2166 66 2272
rect 100 2200 2181 2238
rect 0 2132 1080 2166
rect 0 2026 66 2132
rect 1114 2098 1168 2200
rect 2216 2166 2282 2272
rect 1202 2132 2282 2166
rect 100 2060 2181 2098
rect 0 1992 1080 2026
rect 0 1886 66 1992
rect 1114 1958 1168 2060
rect 2216 2026 2282 2132
rect 1202 1992 2282 2026
rect 100 1920 2181 1958
rect 0 1852 1080 1886
rect 0 1746 66 1852
rect 1114 1818 1168 1920
rect 2216 1886 2282 1992
rect 1202 1852 2282 1886
rect 100 1780 2181 1818
rect 0 1712 1080 1746
rect 0 1606 66 1712
rect 1114 1678 1168 1780
rect 2216 1746 2282 1852
rect 1202 1712 2282 1746
rect 100 1640 2181 1678
rect 0 1572 1080 1606
rect 0 1466 66 1572
rect 1114 1538 1168 1640
rect 2216 1606 2282 1712
rect 1202 1572 2282 1606
rect 100 1500 2181 1538
rect 0 1430 1080 1466
rect 0 1326 66 1430
rect 1114 1398 1168 1500
rect 2216 1466 2282 1572
rect 1202 1432 2282 1466
rect 1114 1396 2181 1398
rect 100 1360 2181 1396
rect 0 1292 1080 1326
rect 0 1186 66 1292
rect 1114 1258 1168 1360
rect 2216 1326 2282 1432
rect 1202 1292 2282 1326
rect 100 1220 2181 1258
rect 0 1152 1080 1186
rect 0 1046 66 1152
rect 1114 1118 1168 1220
rect 2216 1186 2282 1292
rect 1202 1152 2282 1186
rect 100 1080 2181 1118
rect 0 1012 1080 1046
rect 0 906 66 1012
rect 1114 978 1168 1080
rect 2216 1046 2282 1152
rect 1202 1012 2282 1046
rect 100 940 2181 978
rect 0 872 1080 906
rect 0 766 66 872
rect 1114 838 1168 940
rect 2216 906 2282 1012
rect 1202 872 2282 906
rect 100 800 2181 838
rect 0 732 1080 766
rect 0 626 66 732
rect 1114 698 1168 800
rect 2216 766 2282 872
rect 1202 732 2282 766
rect 100 660 2181 698
rect 0 592 1080 626
rect 0 486 66 592
rect 1114 558 1168 660
rect 2216 626 2282 732
rect 1202 592 2282 626
rect 100 520 2181 558
rect 0 452 1080 486
rect 0 346 66 452
rect 1114 418 1168 520
rect 2216 486 2282 592
rect 1202 452 2282 486
rect 100 380 2181 418
rect 0 312 1080 346
rect 0 206 66 312
rect 1114 278 1168 380
rect 2216 346 2282 452
rect 1202 312 2282 346
rect 100 240 2181 278
rect 0 172 1080 206
rect 0 66 66 172
rect 1114 138 1168 240
rect 2216 206 2282 312
rect 1202 172 2282 206
rect 100 100 2181 138
rect 2216 66 2282 172
rect 0 0 2282 66
<< obsm1 >>
rect 0 2272 2282 2338
rect 0 66 66 2272
rect 100 1201 128 2244
rect 156 1229 184 2272
rect 212 1201 240 2244
rect 268 1229 296 2272
rect 324 1201 352 2244
rect 380 1229 408 2272
rect 436 1201 464 2244
rect 492 1229 520 2272
rect 548 1201 576 2244
rect 604 1229 632 2272
rect 660 1201 688 2244
rect 716 1229 744 2272
rect 772 1201 800 2244
rect 828 1229 856 2272
rect 884 1201 912 2244
rect 940 1229 968 2272
rect 996 1201 1024 2244
rect 1052 1229 1080 2272
rect 1114 1201 1168 2244
rect 1202 1229 1230 2272
rect 1258 1201 1286 2244
rect 1314 1229 1342 2272
rect 1370 1201 1398 2244
rect 1426 1229 1454 2272
rect 1482 1201 1510 2244
rect 1538 1229 1566 2272
rect 1594 1201 1622 2244
rect 1650 1229 1678 2272
rect 1706 1201 1734 2244
rect 1762 1229 1790 2272
rect 1818 1201 1846 2244
rect 1874 1229 1902 2272
rect 1930 1201 1958 2244
rect 1986 1229 2014 2272
rect 2042 1201 2070 2244
rect 2098 1229 2126 2272
rect 2154 1201 2182 2244
rect 100 1137 2182 1201
rect 100 94 128 1137
rect 156 66 184 1109
rect 212 94 240 1137
rect 268 66 296 1109
rect 324 94 352 1137
rect 380 66 408 1109
rect 436 94 464 1137
rect 492 66 520 1109
rect 548 94 576 1137
rect 604 66 632 1109
rect 660 94 688 1137
rect 716 66 744 1109
rect 772 94 800 1137
rect 828 66 856 1109
rect 884 94 912 1137
rect 940 66 968 1109
rect 996 94 1024 1137
rect 1052 66 1080 1109
rect 1114 94 1168 1137
rect 1202 66 1230 1109
rect 1258 94 1286 1137
rect 1314 66 1342 1109
rect 1370 94 1398 1137
rect 1426 66 1454 1109
rect 1482 94 1510 1137
rect 1538 66 1566 1109
rect 1594 94 1622 1137
rect 1650 66 1678 1109
rect 1706 94 1734 1137
rect 1762 66 1790 1109
rect 1818 94 1846 1137
rect 1874 66 1902 1109
rect 1930 94 1958 1137
rect 1986 66 2014 1109
rect 2042 94 2070 1137
rect 2098 66 2126 1109
rect 2154 94 2182 1137
rect 2216 66 2282 2272
rect 0 0 2282 66
<< obsm2 >>
rect 0 2272 1086 2338
rect 0 2188 66 2272
rect 1114 2244 1168 2338
rect 1196 2272 2282 2338
rect 94 2216 2188 2244
rect 0 2160 1085 2188
rect 0 2076 66 2160
rect 1113 2132 1169 2216
rect 2216 2188 2282 2272
rect 1197 2160 2282 2188
rect 94 2104 2188 2132
rect 0 2048 1085 2076
rect 0 1964 66 2048
rect 1113 2020 1169 2104
rect 2216 2076 2282 2160
rect 1197 2048 2282 2076
rect 94 1992 2188 2020
rect 0 1936 1085 1964
rect 0 1852 66 1936
rect 1113 1908 1169 1992
rect 2216 1964 2282 2048
rect 1197 1936 2282 1964
rect 94 1880 2188 1908
rect 0 1824 1085 1852
rect 0 1740 66 1824
rect 1113 1796 1169 1880
rect 2216 1852 2282 1936
rect 1197 1824 2282 1852
rect 94 1768 2188 1796
rect 0 1712 1085 1740
rect 0 1628 66 1712
rect 1113 1684 1169 1768
rect 2216 1740 2282 1824
rect 1197 1712 2282 1740
rect 94 1656 2188 1684
rect 0 1600 1085 1628
rect 0 1516 66 1600
rect 1113 1572 1169 1656
rect 2216 1628 2282 1712
rect 1197 1600 2282 1628
rect 94 1544 2188 1572
rect 0 1488 1085 1516
rect 0 1404 66 1488
rect 1113 1460 1169 1544
rect 2216 1516 2282 1600
rect 1197 1488 2282 1516
rect 94 1432 2188 1460
rect 0 1376 1085 1404
rect 0 1292 66 1376
rect 1113 1348 1169 1432
rect 2216 1404 2282 1488
rect 1197 1376 2282 1404
rect 94 1320 2188 1348
rect 0 1225 1085 1292
rect 0 1224 66 1225
rect 1113 1197 1169 1320
rect 2216 1292 2282 1376
rect 1197 1225 2282 1292
rect 2216 1224 2282 1225
rect 74 1196 2208 1197
rect 0 1142 2282 1196
rect 74 1141 2208 1142
rect 0 1113 66 1114
rect 0 1046 1085 1113
rect 0 962 66 1046
rect 1113 1018 1169 1141
rect 2216 1113 2282 1114
rect 1197 1046 2282 1113
rect 94 990 2188 1018
rect 0 934 1085 962
rect 0 850 66 934
rect 1113 906 1169 990
rect 2216 962 2282 1046
rect 1197 934 2282 962
rect 94 878 2188 906
rect 0 822 1085 850
rect 0 738 66 822
rect 1113 794 1169 878
rect 2216 850 2282 934
rect 1197 822 2282 850
rect 94 766 2188 794
rect 0 710 1085 738
rect 0 626 66 710
rect 1113 682 1169 766
rect 2216 738 2282 822
rect 1197 710 2282 738
rect 94 654 2188 682
rect 0 598 1085 626
rect 0 514 66 598
rect 1113 570 1169 654
rect 2216 626 2282 710
rect 1197 598 2282 626
rect 94 542 2188 570
rect 0 486 1085 514
rect 0 402 66 486
rect 1113 458 1169 542
rect 2216 514 2282 598
rect 1197 486 2282 514
rect 94 430 2188 458
rect 0 374 1085 402
rect 0 290 66 374
rect 1113 346 1169 430
rect 2216 402 2282 486
rect 1197 374 2282 402
rect 94 318 2188 346
rect 0 262 1085 290
rect 0 178 66 262
rect 1113 234 1169 318
rect 2216 290 2282 374
rect 1197 262 2282 290
rect 94 206 2188 234
rect 0 150 1085 178
rect 0 66 66 150
rect 1113 122 1169 206
rect 2216 178 2282 262
rect 1197 150 2282 178
rect 94 94 2188 122
rect 0 0 1086 66
rect 1114 0 1168 94
rect 2216 66 2282 150
rect 1196 0 2282 66
<< obsm3 >>
rect 0 2272 2282 2338
rect 0 66 66 2272
rect 126 1202 186 2212
rect 246 1262 306 2272
rect 366 1202 426 2212
rect 486 1262 546 2272
rect 606 1202 666 2212
rect 726 1262 786 2272
rect 846 1202 906 2212
rect 966 1262 1048 2272
rect 1108 1202 1174 2212
rect 1234 1262 1316 2272
rect 1376 1202 1436 2212
rect 1496 1262 1556 2272
rect 1616 1202 1676 2212
rect 1736 1262 1796 2272
rect 1856 1202 1916 2212
rect 1976 1262 2036 2272
rect 2096 1202 2156 2212
rect 126 1136 2156 1202
rect 126 126 186 1136
rect 246 66 306 1076
rect 366 126 426 1136
rect 486 66 546 1076
rect 606 126 666 1136
rect 726 66 786 1076
rect 846 126 906 1136
rect 966 66 1048 1076
rect 1108 126 1174 1136
rect 1234 66 1316 1076
rect 1376 126 1436 1136
rect 1496 66 1556 1076
rect 1616 126 1676 1136
rect 1736 66 1796 1076
rect 1856 126 1916 1136
rect 1976 66 2036 1076
rect 2096 126 2156 1136
rect 2216 66 2282 2272
rect 0 0 2282 66
<< metal4 >>
rect -4370 2272 6652 4059
rect -4370 2092 66 2272
rect 126 2152 2156 2212
rect -4370 2032 1048 2092
rect -4370 1852 66 2032
rect 1108 1972 1174 2152
rect 2216 2092 6652 2272
rect 1234 2032 6652 2092
rect 126 1912 2156 1972
rect -4370 1792 1048 1852
rect -4370 1612 66 1792
rect 1108 1732 1174 1912
rect 2216 1852 6652 2032
rect 1234 1792 6652 1852
rect 126 1672 2156 1732
rect -4370 1532 1048 1612
rect -4370 1352 66 1532
rect 1108 1472 1174 1672
rect 2216 1612 6652 1792
rect 1234 1532 6652 1612
rect 126 1412 2156 1472
rect -4370 1262 1048 1352
rect -4370 1076 66 1262
rect 1108 1202 1174 1412
rect 2216 1352 6652 1532
rect 1234 1262 6652 1352
rect 126 1136 2156 1202
rect -4370 986 1048 1076
rect -4370 806 66 986
rect 1108 926 1174 1136
rect 2216 1076 6652 1262
rect 1234 986 6652 1076
rect 126 866 2156 926
rect -4370 726 1048 806
rect -4370 546 66 726
rect 1108 666 1174 866
rect 2216 806 6652 986
rect 1234 726 6652 806
rect 126 606 2156 666
rect -4370 486 1048 546
rect -4370 306 66 486
rect 1108 426 1174 606
rect 2216 546 6652 726
rect 1234 486 6652 546
rect 126 366 2156 426
rect -4370 246 1048 306
rect -4370 66 66 246
rect 1108 186 1174 366
rect 2216 306 6652 486
rect 1234 246 6652 306
rect 126 126 2156 186
rect 2216 66 6652 246
rect -4370 -1721 6652 66
<< metal5 >>
rect 0 0 2282 2338
<< labels >>
rlabel metal4 s 2216 2092 6652 2272 6 C0
port 1 nsew
rlabel metal4 s 2216 1852 6652 2032 6 C0
port 1 nsew
rlabel metal4 s 2216 1612 6652 1792 6 C0
port 1 nsew
rlabel metal4 s 2216 1352 6652 1532 6 C0
port 1 nsew
rlabel metal4 s 2216 1076 6652 1262 6 C0
port 1 nsew
rlabel metal4 s 2216 806 6652 986 6 C0
port 1 nsew
rlabel metal4 s 2216 546 6652 726 6 C0
port 1 nsew
rlabel metal4 s 2216 306 6652 486 6 C0
port 1 nsew
rlabel metal4 s 2216 66 6652 246 6 C0
port 1 nsew
rlabel metal4 s 1234 2032 6652 2092 6 C0
port 1 nsew
rlabel metal4 s 1234 1792 6652 1852 6 C0
port 1 nsew
rlabel metal4 s 1234 1532 6652 1612 6 C0
port 1 nsew
rlabel metal4 s 1234 1262 6652 1352 6 C0
port 1 nsew
rlabel metal4 s 1234 986 6652 1076 6 C0
port 1 nsew
rlabel metal4 s 1234 726 6652 806 6 C0
port 1 nsew
rlabel metal4 s 1234 486 6652 546 6 C0
port 1 nsew
rlabel metal4 s 1234 246 6652 306 6 C0
port 1 nsew
rlabel metal4 s -4370 2272 6652 4059 6 C0
port 1 nsew
rlabel metal4 s -4370 2092 66 2272 4 C0
port 1 nsew
rlabel metal4 s -4370 2032 1048 2092 4 C0
port 1 nsew
rlabel metal4 s -4370 1852 66 2032 4 C0
port 1 nsew
rlabel metal4 s -4370 1792 1048 1852 4 C0
port 1 nsew
rlabel metal4 s -4370 1612 66 1792 4 C0
port 1 nsew
rlabel metal4 s -4370 1532 1048 1612 4 C0
port 1 nsew
rlabel metal4 s -4370 1352 66 1532 4 C0
port 1 nsew
rlabel metal4 s -4370 1262 1048 1352 4 C0
port 1 nsew
rlabel metal4 s -4370 1076 66 1262 4 C0
port 1 nsew
rlabel metal4 s -4370 986 1048 1076 4 C0
port 1 nsew
rlabel metal4 s -4370 806 66 986 4 C0
port 1 nsew
rlabel metal4 s -4370 726 1048 806 4 C0
port 1 nsew
rlabel metal4 s -4370 546 66 726 4 C0
port 1 nsew
rlabel metal4 s -4370 486 1048 546 4 C0
port 1 nsew
rlabel metal4 s -4370 306 66 486 4 C0
port 1 nsew
rlabel metal4 s -4370 246 1048 306 4 C0
port 1 nsew
rlabel metal4 s -4370 66 66 246 4 C0
port 1 nsew
rlabel metal4 s -4370 -1721 6652 66 8 C0
port 1 nsew
rlabel metal4 s 1108 1972 1174 2152 6 C1
port 2 nsew
rlabel metal4 s 1108 1732 1174 1912 6 C1
port 2 nsew
rlabel metal4 s 1108 1472 1174 1672 6 C1
port 2 nsew
rlabel metal4 s 1108 1202 1174 1412 6 C1
port 2 nsew
rlabel metal4 s 1108 926 1174 1136 6 C1
port 2 nsew
rlabel metal4 s 1108 666 1174 866 6 C1
port 2 nsew
rlabel metal4 s 1108 426 1174 606 6 C1
port 2 nsew
rlabel metal4 s 1108 186 1174 366 6 C1
port 2 nsew
rlabel metal4 s 126 2152 2156 2212 6 C1
port 2 nsew
rlabel metal4 s 126 1912 2156 1972 6 C1
port 2 nsew
rlabel metal4 s 126 1672 2156 1732 6 C1
port 2 nsew
rlabel metal4 s 126 1412 2156 1472 6 C1
port 2 nsew
rlabel metal4 s 126 1136 2156 1202 6 C1
port 2 nsew
rlabel metal4 s 126 866 2156 926 6 C1
port 2 nsew
rlabel metal4 s 126 606 2156 666 6 C1
port 2 nsew
rlabel metal4 s 126 366 2156 426 6 C1
port 2 nsew
rlabel metal4 s 126 126 2156 186 6 C1
port 2 nsew
rlabel metal5 s 0 0 2282 2338 6 M5A
port 3 nsew
rlabel locali s 50 4758 84 4824 6 SUB
port 4 nsew
<< properties >>
string FIXED_BBOX -4370 -1721 6652 4832
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1168618
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 1167444
<< end >>
