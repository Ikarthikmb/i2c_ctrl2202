/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/rf_pfet_01v8_mvt/sky130_fd_pr__rf_pfet_01v8_mvt_aF02W0p84L0p15.spice