magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 879 203
rect 30 -17 64 21
<< locali >>
rect 19 331 69 493
rect 187 331 253 425
rect 355 331 432 425
rect 19 297 432 331
rect 30 215 156 255
rect 214 215 340 255
rect 374 169 432 297
rect 489 215 620 255
rect 678 215 900 255
rect 271 135 609 169
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 103 459 525 493
rect 103 365 153 459
rect 287 365 321 459
rect 475 331 525 459
rect 559 365 593 527
rect 627 331 693 493
rect 727 365 761 527
rect 795 331 861 493
rect 475 297 861 331
rect 19 136 237 170
rect 19 51 69 136
rect 103 17 169 102
rect 203 101 237 136
rect 643 136 875 170
rect 643 101 677 136
rect 203 51 421 101
rect 459 51 677 101
rect 711 17 777 102
rect 811 51 875 136
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 489 215 620 255 6 A1
port 1 nsew signal input
rlabel locali s 678 215 900 255 6 A2
port 2 nsew signal input
rlabel locali s 214 215 340 255 6 B1
port 3 nsew signal input
rlabel locali s 30 215 156 255 6 B2
port 4 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 879 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 271 135 609 169 6 Y
port 9 nsew signal output
rlabel locali s 374 169 432 297 6 Y
port 9 nsew signal output
rlabel locali s 19 297 432 331 6 Y
port 9 nsew signal output
rlabel locali s 355 331 432 425 6 Y
port 9 nsew signal output
rlabel locali s 187 331 253 425 6 Y
port 9 nsew signal output
rlabel locali s 19 331 69 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 920 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 4079362
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4070876
<< end >>
