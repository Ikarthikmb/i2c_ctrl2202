magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 98 163 369 203
rect 98 157 634 163
rect 1 27 634 157
rect 1 21 369 27
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 176 47 206 177
rect 260 47 290 177
rect 358 53 388 137
rect 442 53 472 137
rect 526 53 556 137
<< scpmoshvt >>
rect 79 360 109 444
rect 176 297 206 497
rect 260 297 290 497
rect 358 297 388 381
rect 442 297 472 381
rect 526 297 556 381
<< ndiff >>
rect 124 131 176 177
rect 27 108 79 131
rect 27 74 35 108
rect 69 74 79 108
rect 27 47 79 74
rect 109 97 176 131
rect 109 63 119 97
rect 153 63 176 97
rect 109 47 176 63
rect 206 103 260 177
rect 206 69 216 103
rect 250 69 260 103
rect 206 47 260 69
rect 290 137 343 177
rect 290 97 358 137
rect 290 63 304 97
rect 338 63 358 97
rect 290 53 358 63
rect 388 111 442 137
rect 388 77 398 111
rect 432 77 442 111
rect 388 53 442 77
rect 472 97 526 137
rect 472 63 482 97
rect 516 63 526 97
rect 472 53 526 63
rect 556 111 608 137
rect 556 77 566 111
rect 600 77 608 111
rect 556 53 608 77
rect 290 47 343 53
<< pdiff >>
rect 124 476 176 497
rect 124 444 132 476
rect 27 412 79 444
rect 27 378 35 412
rect 69 378 79 412
rect 27 360 79 378
rect 109 442 132 444
rect 166 442 176 476
rect 109 360 176 442
rect 124 297 176 360
rect 206 340 260 497
rect 206 306 216 340
rect 250 306 260 340
rect 206 297 260 306
rect 290 476 343 497
rect 290 442 301 476
rect 335 442 343 476
rect 290 381 343 442
rect 290 297 358 381
rect 388 297 442 381
rect 472 297 526 381
rect 556 354 608 381
rect 556 320 566 354
rect 600 320 608 354
rect 556 297 608 320
<< ndiffc >>
rect 35 74 69 108
rect 119 63 153 97
rect 216 69 250 103
rect 304 63 338 97
rect 398 77 432 111
rect 482 63 516 97
rect 566 77 600 111
<< pdiffc >>
rect 35 378 69 412
rect 132 442 166 476
rect 216 306 250 340
rect 301 442 335 476
rect 566 320 600 354
<< poly >>
rect 176 497 206 523
rect 260 497 290 523
rect 79 444 109 470
rect 79 265 109 360
rect 424 473 490 483
rect 424 439 440 473
rect 474 439 490 473
rect 424 429 490 439
rect 358 381 388 407
rect 442 381 472 429
rect 526 381 556 407
rect 22 249 109 265
rect 22 215 35 249
rect 69 215 109 249
rect 22 199 109 215
rect 79 131 109 199
rect 176 265 206 297
rect 260 265 290 297
rect 358 265 388 297
rect 176 249 299 265
rect 176 215 255 249
rect 289 215 299 249
rect 176 199 299 215
rect 346 249 400 265
rect 346 215 356 249
rect 390 215 400 249
rect 346 199 400 215
rect 176 177 206 199
rect 260 177 290 199
rect 358 137 388 199
rect 442 137 472 297
rect 526 265 556 297
rect 514 249 568 265
rect 514 215 524 249
rect 558 215 568 249
rect 514 199 568 215
rect 526 137 556 199
rect 79 21 109 47
rect 176 21 206 47
rect 260 21 290 47
rect 358 27 388 53
rect 442 27 472 53
rect 526 27 556 53
<< polycont >>
rect 440 439 474 473
rect 35 215 69 249
rect 255 215 289 249
rect 356 215 390 249
rect 524 215 558 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 110 476 182 527
rect 17 412 69 444
rect 110 442 132 476
rect 166 442 182 476
rect 285 476 351 527
rect 285 442 301 476
rect 335 442 351 476
rect 387 439 440 473
rect 474 439 627 473
rect 387 425 627 439
rect 17 378 35 412
rect 69 391 344 408
rect 69 378 532 391
rect 17 374 532 378
rect 17 362 153 374
rect 17 249 85 328
rect 17 215 35 249
rect 69 215 85 249
rect 119 181 153 362
rect 310 357 532 374
rect 17 147 153 181
rect 187 306 216 340
rect 250 306 266 340
rect 187 299 266 306
rect 17 108 69 147
rect 187 119 221 299
rect 255 249 289 265
rect 339 249 446 323
rect 339 215 356 249
rect 390 215 446 249
rect 498 265 532 357
rect 566 354 627 385
rect 600 320 627 354
rect 566 299 627 320
rect 498 249 558 265
rect 498 215 524 249
rect 255 187 289 215
rect 498 199 558 215
rect 255 181 319 187
rect 255 165 432 181
rect 593 165 627 299
rect 255 153 627 165
rect 285 147 627 153
rect 398 131 627 147
rect 17 74 35 108
rect 17 58 69 74
rect 119 97 153 113
rect 119 17 153 63
rect 187 103 257 119
rect 187 69 216 103
rect 250 69 257 103
rect 187 53 257 69
rect 304 97 338 113
rect 304 17 338 63
rect 398 111 432 131
rect 566 121 627 131
rect 566 111 617 121
rect 398 61 432 77
rect 466 63 482 97
rect 516 63 532 97
rect 466 17 532 63
rect 600 77 617 111
rect 566 61 617 77
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 398 221 432 255 0 FreeSans 400 0 0 0 A
port 1 nsew signal input
flabel locali s 490 425 524 459 0 FreeSans 400 180 0 0 B
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 C_N
port 3 nsew signal input
flabel locali s 214 85 248 119 0 FreeSans 200 180 0 0 X
port 8 nsew signal output
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 or3b_2
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 1051096
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1045306
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 2.720 3.220 2.720 
<< end >>
