magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< locali >>
rect 6000 5458 6034 5474
rect 6000 5408 6034 5424
<< viali >>
rect 6000 5424 6034 5458
<< metal1 >>
rect 5985 5415 5991 5467
rect 6043 5415 6049 5467
rect 13141 3609 13147 3661
rect 13199 3609 13205 3661
rect 14389 3609 14395 3661
rect 14447 3609 14453 3661
rect 15637 3609 15643 3661
rect 15695 3609 15701 3661
rect 16885 3609 16891 3661
rect 16943 3609 16949 3661
rect 18133 3609 18139 3661
rect 18191 3609 18197 3661
rect 19381 3609 19387 3661
rect 19439 3609 19445 3661
rect 20629 3609 20635 3661
rect 20687 3609 20693 3661
rect 21877 3609 21883 3661
rect 21935 3609 21941 3661
rect 23125 3609 23131 3661
rect 23183 3609 23189 3661
rect 24373 3609 24379 3661
rect 24431 3609 24437 3661
rect 25621 3609 25627 3661
rect 25679 3609 25685 3661
rect 26869 3609 26875 3661
rect 26927 3609 26933 3661
rect 28117 3609 28123 3661
rect 28175 3609 28181 3661
rect 29365 3609 29371 3661
rect 29423 3609 29429 3661
rect 30613 3609 30619 3661
rect 30671 3609 30677 3661
rect 31861 3609 31867 3661
rect 31919 3609 31925 3661
rect 33109 3609 33115 3661
rect 33167 3609 33173 3661
rect 34357 3609 34363 3661
rect 34415 3609 34421 3661
rect 35605 3609 35611 3661
rect 35663 3609 35669 3661
rect 36853 3609 36859 3661
rect 36911 3609 36917 3661
rect 38101 3609 38107 3661
rect 38159 3609 38165 3661
rect 39349 3609 39355 3661
rect 39407 3609 39413 3661
rect 40597 3609 40603 3661
rect 40655 3609 40661 3661
rect 41845 3609 41851 3661
rect 41903 3609 41909 3661
rect 43093 3609 43099 3661
rect 43151 3609 43157 3661
rect 44341 3609 44347 3661
rect 44399 3609 44405 3661
rect 45589 3609 45595 3661
rect 45647 3609 45653 3661
rect 46837 3609 46843 3661
rect 46895 3609 46901 3661
rect 48085 3609 48091 3661
rect 48143 3609 48149 3661
rect 49333 3609 49339 3661
rect 49391 3609 49397 3661
rect 50581 3609 50587 3661
rect 50639 3609 50645 3661
rect 51829 3609 51835 3661
rect 51887 3609 51893 3661
rect 13299 1350 13305 1402
rect 13357 1350 13363 1402
rect 14547 1350 14553 1402
rect 14605 1350 14611 1402
rect 15795 1350 15801 1402
rect 15853 1350 15859 1402
rect 17043 1350 17049 1402
rect 17101 1350 17107 1402
rect 18291 1350 18297 1402
rect 18349 1350 18355 1402
rect 19539 1350 19545 1402
rect 19597 1350 19603 1402
rect 20787 1350 20793 1402
rect 20845 1350 20851 1402
rect 22035 1350 22041 1402
rect 22093 1350 22099 1402
rect 23283 1350 23289 1402
rect 23341 1350 23347 1402
rect 24531 1350 24537 1402
rect 24589 1350 24595 1402
rect 25779 1350 25785 1402
rect 25837 1350 25843 1402
rect 27027 1350 27033 1402
rect 27085 1350 27091 1402
rect 28275 1350 28281 1402
rect 28333 1350 28339 1402
rect 29523 1350 29529 1402
rect 29581 1350 29587 1402
rect 30771 1350 30777 1402
rect 30829 1350 30835 1402
rect 32019 1350 32025 1402
rect 32077 1350 32083 1402
rect 33267 1350 33273 1402
rect 33325 1350 33331 1402
rect 34515 1350 34521 1402
rect 34573 1350 34579 1402
rect 35763 1350 35769 1402
rect 35821 1350 35827 1402
rect 37011 1350 37017 1402
rect 37069 1350 37075 1402
rect 38259 1350 38265 1402
rect 38317 1350 38323 1402
rect 39507 1350 39513 1402
rect 39565 1350 39571 1402
rect 40755 1350 40761 1402
rect 40813 1350 40819 1402
rect 42003 1350 42009 1402
rect 42061 1350 42067 1402
rect 43251 1350 43257 1402
rect 43309 1350 43315 1402
rect 44499 1350 44505 1402
rect 44557 1350 44563 1402
rect 45747 1350 45753 1402
rect 45805 1350 45811 1402
rect 46995 1350 47001 1402
rect 47053 1350 47059 1402
rect 48243 1350 48249 1402
rect 48301 1350 48307 1402
rect 49491 1350 49497 1402
rect 49549 1350 49555 1402
rect 50739 1350 50745 1402
rect 50797 1350 50803 1402
rect 51987 1350 51993 1402
rect 52045 1350 52051 1402
<< via1 >>
rect 5991 5458 6043 5467
rect 5991 5424 6000 5458
rect 6000 5424 6034 5458
rect 6034 5424 6043 5458
rect 5991 5415 6043 5424
rect 13147 3609 13199 3661
rect 14395 3609 14447 3661
rect 15643 3609 15695 3661
rect 16891 3609 16943 3661
rect 18139 3609 18191 3661
rect 19387 3609 19439 3661
rect 20635 3609 20687 3661
rect 21883 3609 21935 3661
rect 23131 3609 23183 3661
rect 24379 3609 24431 3661
rect 25627 3609 25679 3661
rect 26875 3609 26927 3661
rect 28123 3609 28175 3661
rect 29371 3609 29423 3661
rect 30619 3609 30671 3661
rect 31867 3609 31919 3661
rect 33115 3609 33167 3661
rect 34363 3609 34415 3661
rect 35611 3609 35663 3661
rect 36859 3609 36911 3661
rect 38107 3609 38159 3661
rect 39355 3609 39407 3661
rect 40603 3609 40655 3661
rect 41851 3609 41903 3661
rect 43099 3609 43151 3661
rect 44347 3609 44399 3661
rect 45595 3609 45647 3661
rect 46843 3609 46895 3661
rect 48091 3609 48143 3661
rect 49339 3609 49391 3661
rect 50587 3609 50639 3661
rect 51835 3609 51887 3661
rect 13305 1350 13357 1402
rect 14553 1350 14605 1402
rect 15801 1350 15853 1402
rect 17049 1350 17101 1402
rect 18297 1350 18349 1402
rect 19545 1350 19597 1402
rect 20793 1350 20845 1402
rect 22041 1350 22093 1402
rect 23289 1350 23341 1402
rect 24537 1350 24589 1402
rect 25785 1350 25837 1402
rect 27033 1350 27085 1402
rect 28281 1350 28333 1402
rect 29529 1350 29581 1402
rect 30777 1350 30829 1402
rect 32025 1350 32077 1402
rect 33273 1350 33325 1402
rect 34521 1350 34573 1402
rect 35769 1350 35821 1402
rect 37017 1350 37069 1402
rect 38265 1350 38317 1402
rect 39513 1350 39565 1402
rect 40761 1350 40813 1402
rect 42009 1350 42061 1402
rect 43257 1350 43309 1402
rect 44505 1350 44557 1402
rect 45753 1350 45805 1402
rect 47001 1350 47053 1402
rect 48249 1350 48301 1402
rect 49497 1350 49549 1402
rect 50745 1350 50797 1402
rect 51993 1350 52045 1402
<< metal2 >>
rect 5989 5469 6045 5478
rect 5989 5404 6045 5413
rect 13145 3663 13201 3672
rect 13145 3598 13201 3607
rect 14393 3663 14449 3672
rect 14393 3598 14449 3607
rect 15641 3663 15697 3672
rect 15641 3598 15697 3607
rect 16889 3663 16945 3672
rect 16889 3598 16945 3607
rect 18137 3663 18193 3672
rect 18137 3598 18193 3607
rect 19385 3663 19441 3672
rect 19385 3598 19441 3607
rect 20633 3663 20689 3672
rect 20633 3598 20689 3607
rect 21881 3663 21937 3672
rect 21881 3598 21937 3607
rect 23129 3663 23185 3672
rect 23129 3598 23185 3607
rect 24377 3663 24433 3672
rect 24377 3598 24433 3607
rect 25625 3663 25681 3672
rect 25625 3598 25681 3607
rect 26873 3663 26929 3672
rect 26873 3598 26929 3607
rect 28121 3663 28177 3672
rect 28121 3598 28177 3607
rect 29369 3663 29425 3672
rect 29369 3598 29425 3607
rect 30617 3663 30673 3672
rect 30617 3598 30673 3607
rect 31865 3663 31921 3672
rect 31865 3598 31921 3607
rect 33113 3663 33169 3672
rect 33113 3598 33169 3607
rect 34361 3663 34417 3672
rect 34361 3598 34417 3607
rect 35609 3663 35665 3672
rect 35609 3598 35665 3607
rect 36857 3663 36913 3672
rect 36857 3598 36913 3607
rect 38105 3663 38161 3672
rect 38105 3598 38161 3607
rect 39353 3663 39409 3672
rect 39353 3598 39409 3607
rect 40601 3663 40657 3672
rect 40601 3598 40657 3607
rect 41849 3663 41905 3672
rect 41849 3598 41905 3607
rect 43097 3663 43153 3672
rect 43097 3598 43153 3607
rect 44345 3663 44401 3672
rect 44345 3598 44401 3607
rect 45593 3663 45649 3672
rect 45593 3598 45649 3607
rect 46841 3663 46897 3672
rect 46841 3598 46897 3607
rect 48089 3663 48145 3672
rect 48089 3598 48145 3607
rect 49337 3663 49393 3672
rect 49337 3598 49393 3607
rect 50585 3663 50641 3672
rect 50585 3598 50641 3607
rect 51833 3663 51889 3672
rect 51833 3598 51889 3607
rect 13303 1404 13359 1413
rect 13303 1339 13359 1348
rect 14551 1404 14607 1413
rect 14551 1339 14607 1348
rect 15799 1404 15855 1413
rect 15799 1339 15855 1348
rect 17047 1404 17103 1413
rect 17047 1339 17103 1348
rect 18295 1404 18351 1413
rect 18295 1339 18351 1348
rect 19543 1404 19599 1413
rect 19543 1339 19599 1348
rect 20791 1404 20847 1413
rect 20791 1339 20847 1348
rect 22039 1404 22095 1413
rect 22039 1339 22095 1348
rect 23287 1404 23343 1413
rect 23287 1339 23343 1348
rect 24535 1404 24591 1413
rect 24535 1339 24591 1348
rect 25783 1404 25839 1413
rect 25783 1339 25839 1348
rect 27031 1404 27087 1413
rect 27031 1339 27087 1348
rect 28279 1404 28335 1413
rect 28279 1339 28335 1348
rect 29527 1404 29583 1413
rect 29527 1339 29583 1348
rect 30775 1404 30831 1413
rect 30775 1339 30831 1348
rect 32023 1404 32079 1413
rect 32023 1339 32079 1348
rect 33271 1404 33327 1413
rect 33271 1339 33327 1348
rect 34519 1404 34575 1413
rect 34519 1339 34575 1348
rect 35767 1404 35823 1413
rect 35767 1339 35823 1348
rect 37015 1404 37071 1413
rect 37015 1339 37071 1348
rect 38263 1404 38319 1413
rect 38263 1339 38319 1348
rect 39511 1404 39567 1413
rect 39511 1339 39567 1348
rect 40759 1404 40815 1413
rect 40759 1339 40815 1348
rect 42007 1404 42063 1413
rect 42007 1339 42063 1348
rect 43255 1404 43311 1413
rect 43255 1339 43311 1348
rect 44503 1404 44559 1413
rect 44503 1339 44559 1348
rect 45751 1404 45807 1413
rect 45751 1339 45807 1348
rect 46999 1404 47055 1413
rect 46999 1339 47055 1348
rect 48247 1404 48303 1413
rect 48247 1339 48303 1348
rect 49495 1404 49551 1413
rect 49495 1339 49551 1348
rect 50743 1404 50799 1413
rect 50743 1339 50799 1348
rect 51991 1404 52047 1413
rect 51991 1339 52047 1348
rect 13018 284 13074 293
rect 13018 219 13074 228
rect 23002 284 23058 293
rect 23002 219 23058 228
rect 32986 284 33042 293
rect 32986 219 33042 228
rect 42970 284 43026 293
rect 42970 219 43026 228
rect 2087 -18293 2143 -18284
rect 2087 -18358 2143 -18349
rect 3255 -18293 3311 -18284
rect 3255 -18358 3311 -18349
rect 4423 -18293 4479 -18284
rect 4423 -18358 4479 -18349
rect 5591 -18293 5647 -18284
rect 5591 -18358 5647 -18349
rect 6759 -18293 6815 -18284
rect 6759 -18358 6815 -18349
rect 7927 -18293 7983 -18284
rect 7927 -18358 7983 -18349
rect 9095 -18293 9151 -18284
rect 9095 -18358 9151 -18349
rect 10263 -18293 10319 -18284
rect 10263 -18358 10319 -18349
rect 11431 -18293 11487 -18284
rect 11431 -18358 11487 -18349
rect 12599 -18293 12655 -18284
rect 12599 -18358 12655 -18349
rect 13767 -18293 13823 -18284
rect 13767 -18358 13823 -18349
rect 14935 -18293 14991 -18284
rect 14935 -18358 14991 -18349
rect 16103 -18293 16159 -18284
rect 16103 -18358 16159 -18349
rect 17271 -18293 17327 -18284
rect 17271 -18358 17327 -18349
rect 18439 -18293 18495 -18284
rect 18439 -18358 18495 -18349
rect 19607 -18293 19663 -18284
rect 19607 -18358 19663 -18349
rect 20775 -18293 20831 -18284
rect 20775 -18358 20831 -18349
rect 21943 -18293 21999 -18284
rect 21943 -18358 21999 -18349
rect 23111 -18293 23167 -18284
rect 23111 -18358 23167 -18349
rect 24279 -18293 24335 -18284
rect 24279 -18358 24335 -18349
rect 25447 -18293 25503 -18284
rect 25447 -18358 25503 -18349
rect 26615 -18293 26671 -18284
rect 26615 -18358 26671 -18349
rect 27783 -18293 27839 -18284
rect 27783 -18358 27839 -18349
rect 28951 -18293 29007 -18284
rect 28951 -18358 29007 -18349
rect 30119 -18293 30175 -18284
rect 30119 -18358 30175 -18349
rect 31287 -18293 31343 -18284
rect 31287 -18358 31343 -18349
rect 32455 -18293 32511 -18284
rect 32455 -18358 32511 -18349
rect 33623 -18293 33679 -18284
rect 33623 -18358 33679 -18349
rect 34791 -18293 34847 -18284
rect 34791 -18358 34847 -18349
rect 35959 -18293 36015 -18284
rect 35959 -18358 36015 -18349
rect 37127 -18293 37183 -18284
rect 37127 -18358 37183 -18349
rect 38295 -18293 38351 -18284
rect 38295 -18358 38351 -18349
rect 39463 -18293 39519 -18284
rect 39463 -18358 39519 -18349
rect 40631 -18293 40687 -18284
rect 40631 -18358 40687 -18349
rect 41799 -18293 41855 -18284
rect 41799 -18358 41855 -18349
rect 42967 -18293 43023 -18284
rect 42967 -18358 43023 -18349
rect 44135 -18293 44191 -18284
rect 44135 -18358 44191 -18349
<< via2 >>
rect 5989 5467 6045 5469
rect 5989 5415 5991 5467
rect 5991 5415 6043 5467
rect 6043 5415 6045 5467
rect 5989 5413 6045 5415
rect 13145 3661 13201 3663
rect 13145 3609 13147 3661
rect 13147 3609 13199 3661
rect 13199 3609 13201 3661
rect 13145 3607 13201 3609
rect 14393 3661 14449 3663
rect 14393 3609 14395 3661
rect 14395 3609 14447 3661
rect 14447 3609 14449 3661
rect 14393 3607 14449 3609
rect 15641 3661 15697 3663
rect 15641 3609 15643 3661
rect 15643 3609 15695 3661
rect 15695 3609 15697 3661
rect 15641 3607 15697 3609
rect 16889 3661 16945 3663
rect 16889 3609 16891 3661
rect 16891 3609 16943 3661
rect 16943 3609 16945 3661
rect 16889 3607 16945 3609
rect 18137 3661 18193 3663
rect 18137 3609 18139 3661
rect 18139 3609 18191 3661
rect 18191 3609 18193 3661
rect 18137 3607 18193 3609
rect 19385 3661 19441 3663
rect 19385 3609 19387 3661
rect 19387 3609 19439 3661
rect 19439 3609 19441 3661
rect 19385 3607 19441 3609
rect 20633 3661 20689 3663
rect 20633 3609 20635 3661
rect 20635 3609 20687 3661
rect 20687 3609 20689 3661
rect 20633 3607 20689 3609
rect 21881 3661 21937 3663
rect 21881 3609 21883 3661
rect 21883 3609 21935 3661
rect 21935 3609 21937 3661
rect 21881 3607 21937 3609
rect 23129 3661 23185 3663
rect 23129 3609 23131 3661
rect 23131 3609 23183 3661
rect 23183 3609 23185 3661
rect 23129 3607 23185 3609
rect 24377 3661 24433 3663
rect 24377 3609 24379 3661
rect 24379 3609 24431 3661
rect 24431 3609 24433 3661
rect 24377 3607 24433 3609
rect 25625 3661 25681 3663
rect 25625 3609 25627 3661
rect 25627 3609 25679 3661
rect 25679 3609 25681 3661
rect 25625 3607 25681 3609
rect 26873 3661 26929 3663
rect 26873 3609 26875 3661
rect 26875 3609 26927 3661
rect 26927 3609 26929 3661
rect 26873 3607 26929 3609
rect 28121 3661 28177 3663
rect 28121 3609 28123 3661
rect 28123 3609 28175 3661
rect 28175 3609 28177 3661
rect 28121 3607 28177 3609
rect 29369 3661 29425 3663
rect 29369 3609 29371 3661
rect 29371 3609 29423 3661
rect 29423 3609 29425 3661
rect 29369 3607 29425 3609
rect 30617 3661 30673 3663
rect 30617 3609 30619 3661
rect 30619 3609 30671 3661
rect 30671 3609 30673 3661
rect 30617 3607 30673 3609
rect 31865 3661 31921 3663
rect 31865 3609 31867 3661
rect 31867 3609 31919 3661
rect 31919 3609 31921 3661
rect 31865 3607 31921 3609
rect 33113 3661 33169 3663
rect 33113 3609 33115 3661
rect 33115 3609 33167 3661
rect 33167 3609 33169 3661
rect 33113 3607 33169 3609
rect 34361 3661 34417 3663
rect 34361 3609 34363 3661
rect 34363 3609 34415 3661
rect 34415 3609 34417 3661
rect 34361 3607 34417 3609
rect 35609 3661 35665 3663
rect 35609 3609 35611 3661
rect 35611 3609 35663 3661
rect 35663 3609 35665 3661
rect 35609 3607 35665 3609
rect 36857 3661 36913 3663
rect 36857 3609 36859 3661
rect 36859 3609 36911 3661
rect 36911 3609 36913 3661
rect 36857 3607 36913 3609
rect 38105 3661 38161 3663
rect 38105 3609 38107 3661
rect 38107 3609 38159 3661
rect 38159 3609 38161 3661
rect 38105 3607 38161 3609
rect 39353 3661 39409 3663
rect 39353 3609 39355 3661
rect 39355 3609 39407 3661
rect 39407 3609 39409 3661
rect 39353 3607 39409 3609
rect 40601 3661 40657 3663
rect 40601 3609 40603 3661
rect 40603 3609 40655 3661
rect 40655 3609 40657 3661
rect 40601 3607 40657 3609
rect 41849 3661 41905 3663
rect 41849 3609 41851 3661
rect 41851 3609 41903 3661
rect 41903 3609 41905 3661
rect 41849 3607 41905 3609
rect 43097 3661 43153 3663
rect 43097 3609 43099 3661
rect 43099 3609 43151 3661
rect 43151 3609 43153 3661
rect 43097 3607 43153 3609
rect 44345 3661 44401 3663
rect 44345 3609 44347 3661
rect 44347 3609 44399 3661
rect 44399 3609 44401 3661
rect 44345 3607 44401 3609
rect 45593 3661 45649 3663
rect 45593 3609 45595 3661
rect 45595 3609 45647 3661
rect 45647 3609 45649 3661
rect 45593 3607 45649 3609
rect 46841 3661 46897 3663
rect 46841 3609 46843 3661
rect 46843 3609 46895 3661
rect 46895 3609 46897 3661
rect 46841 3607 46897 3609
rect 48089 3661 48145 3663
rect 48089 3609 48091 3661
rect 48091 3609 48143 3661
rect 48143 3609 48145 3661
rect 48089 3607 48145 3609
rect 49337 3661 49393 3663
rect 49337 3609 49339 3661
rect 49339 3609 49391 3661
rect 49391 3609 49393 3661
rect 49337 3607 49393 3609
rect 50585 3661 50641 3663
rect 50585 3609 50587 3661
rect 50587 3609 50639 3661
rect 50639 3609 50641 3661
rect 50585 3607 50641 3609
rect 51833 3661 51889 3663
rect 51833 3609 51835 3661
rect 51835 3609 51887 3661
rect 51887 3609 51889 3661
rect 51833 3607 51889 3609
rect 13303 1402 13359 1404
rect 13303 1350 13305 1402
rect 13305 1350 13357 1402
rect 13357 1350 13359 1402
rect 13303 1348 13359 1350
rect 14551 1402 14607 1404
rect 14551 1350 14553 1402
rect 14553 1350 14605 1402
rect 14605 1350 14607 1402
rect 14551 1348 14607 1350
rect 15799 1402 15855 1404
rect 15799 1350 15801 1402
rect 15801 1350 15853 1402
rect 15853 1350 15855 1402
rect 15799 1348 15855 1350
rect 17047 1402 17103 1404
rect 17047 1350 17049 1402
rect 17049 1350 17101 1402
rect 17101 1350 17103 1402
rect 17047 1348 17103 1350
rect 18295 1402 18351 1404
rect 18295 1350 18297 1402
rect 18297 1350 18349 1402
rect 18349 1350 18351 1402
rect 18295 1348 18351 1350
rect 19543 1402 19599 1404
rect 19543 1350 19545 1402
rect 19545 1350 19597 1402
rect 19597 1350 19599 1402
rect 19543 1348 19599 1350
rect 20791 1402 20847 1404
rect 20791 1350 20793 1402
rect 20793 1350 20845 1402
rect 20845 1350 20847 1402
rect 20791 1348 20847 1350
rect 22039 1402 22095 1404
rect 22039 1350 22041 1402
rect 22041 1350 22093 1402
rect 22093 1350 22095 1402
rect 22039 1348 22095 1350
rect 23287 1402 23343 1404
rect 23287 1350 23289 1402
rect 23289 1350 23341 1402
rect 23341 1350 23343 1402
rect 23287 1348 23343 1350
rect 24535 1402 24591 1404
rect 24535 1350 24537 1402
rect 24537 1350 24589 1402
rect 24589 1350 24591 1402
rect 24535 1348 24591 1350
rect 25783 1402 25839 1404
rect 25783 1350 25785 1402
rect 25785 1350 25837 1402
rect 25837 1350 25839 1402
rect 25783 1348 25839 1350
rect 27031 1402 27087 1404
rect 27031 1350 27033 1402
rect 27033 1350 27085 1402
rect 27085 1350 27087 1402
rect 27031 1348 27087 1350
rect 28279 1402 28335 1404
rect 28279 1350 28281 1402
rect 28281 1350 28333 1402
rect 28333 1350 28335 1402
rect 28279 1348 28335 1350
rect 29527 1402 29583 1404
rect 29527 1350 29529 1402
rect 29529 1350 29581 1402
rect 29581 1350 29583 1402
rect 29527 1348 29583 1350
rect 30775 1402 30831 1404
rect 30775 1350 30777 1402
rect 30777 1350 30829 1402
rect 30829 1350 30831 1402
rect 30775 1348 30831 1350
rect 32023 1402 32079 1404
rect 32023 1350 32025 1402
rect 32025 1350 32077 1402
rect 32077 1350 32079 1402
rect 32023 1348 32079 1350
rect 33271 1402 33327 1404
rect 33271 1350 33273 1402
rect 33273 1350 33325 1402
rect 33325 1350 33327 1402
rect 33271 1348 33327 1350
rect 34519 1402 34575 1404
rect 34519 1350 34521 1402
rect 34521 1350 34573 1402
rect 34573 1350 34575 1402
rect 34519 1348 34575 1350
rect 35767 1402 35823 1404
rect 35767 1350 35769 1402
rect 35769 1350 35821 1402
rect 35821 1350 35823 1402
rect 35767 1348 35823 1350
rect 37015 1402 37071 1404
rect 37015 1350 37017 1402
rect 37017 1350 37069 1402
rect 37069 1350 37071 1402
rect 37015 1348 37071 1350
rect 38263 1402 38319 1404
rect 38263 1350 38265 1402
rect 38265 1350 38317 1402
rect 38317 1350 38319 1402
rect 38263 1348 38319 1350
rect 39511 1402 39567 1404
rect 39511 1350 39513 1402
rect 39513 1350 39565 1402
rect 39565 1350 39567 1402
rect 39511 1348 39567 1350
rect 40759 1402 40815 1404
rect 40759 1350 40761 1402
rect 40761 1350 40813 1402
rect 40813 1350 40815 1402
rect 40759 1348 40815 1350
rect 42007 1402 42063 1404
rect 42007 1350 42009 1402
rect 42009 1350 42061 1402
rect 42061 1350 42063 1402
rect 42007 1348 42063 1350
rect 43255 1402 43311 1404
rect 43255 1350 43257 1402
rect 43257 1350 43309 1402
rect 43309 1350 43311 1402
rect 43255 1348 43311 1350
rect 44503 1402 44559 1404
rect 44503 1350 44505 1402
rect 44505 1350 44557 1402
rect 44557 1350 44559 1402
rect 44503 1348 44559 1350
rect 45751 1402 45807 1404
rect 45751 1350 45753 1402
rect 45753 1350 45805 1402
rect 45805 1350 45807 1402
rect 45751 1348 45807 1350
rect 46999 1402 47055 1404
rect 46999 1350 47001 1402
rect 47001 1350 47053 1402
rect 47053 1350 47055 1402
rect 46999 1348 47055 1350
rect 48247 1402 48303 1404
rect 48247 1350 48249 1402
rect 48249 1350 48301 1402
rect 48301 1350 48303 1402
rect 48247 1348 48303 1350
rect 49495 1402 49551 1404
rect 49495 1350 49497 1402
rect 49497 1350 49549 1402
rect 49549 1350 49551 1402
rect 49495 1348 49551 1350
rect 50743 1402 50799 1404
rect 50743 1350 50745 1402
rect 50745 1350 50797 1402
rect 50797 1350 50799 1402
rect 50743 1348 50799 1350
rect 51991 1402 52047 1404
rect 51991 1350 51993 1402
rect 51993 1350 52045 1402
rect 52045 1350 52047 1402
rect 51991 1348 52047 1350
rect 13018 228 13074 284
rect 23002 228 23058 284
rect 32986 228 33042 284
rect 42970 228 43026 284
rect 2087 -18349 2143 -18293
rect 3255 -18349 3311 -18293
rect 4423 -18349 4479 -18293
rect 5591 -18349 5647 -18293
rect 6759 -18349 6815 -18293
rect 7927 -18349 7983 -18293
rect 9095 -18349 9151 -18293
rect 10263 -18349 10319 -18293
rect 11431 -18349 11487 -18293
rect 12599 -18349 12655 -18293
rect 13767 -18349 13823 -18293
rect 14935 -18349 14991 -18293
rect 16103 -18349 16159 -18293
rect 17271 -18349 17327 -18293
rect 18439 -18349 18495 -18293
rect 19607 -18349 19663 -18293
rect 20775 -18349 20831 -18293
rect 21943 -18349 21999 -18293
rect 23111 -18349 23167 -18293
rect 24279 -18349 24335 -18293
rect 25447 -18349 25503 -18293
rect 26615 -18349 26671 -18293
rect 27783 -18349 27839 -18293
rect 28951 -18349 29007 -18293
rect 30119 -18349 30175 -18293
rect 31287 -18349 31343 -18293
rect 32455 -18349 32511 -18293
rect 33623 -18349 33679 -18293
rect 34791 -18349 34847 -18293
rect 35959 -18349 36015 -18293
rect 37127 -18349 37183 -18293
rect 38295 -18349 38351 -18293
rect 39463 -18349 39519 -18293
rect 40631 -18349 40687 -18293
rect 41799 -18349 41855 -18293
rect 42967 -18349 43023 -18293
rect 44135 -18349 44191 -18293
<< metal3 >>
rect 5984 5473 6050 5474
rect 5942 5409 5985 5473
rect 6049 5409 6092 5473
rect 5984 5408 6050 5409
rect 13140 3667 13206 3668
rect 14388 3667 14454 3668
rect 15636 3667 15702 3668
rect 16884 3667 16950 3668
rect 18132 3667 18198 3668
rect 19380 3667 19446 3668
rect 20628 3667 20694 3668
rect 21876 3667 21942 3668
rect 23124 3667 23190 3668
rect 24372 3667 24438 3668
rect 25620 3667 25686 3668
rect 26868 3667 26934 3668
rect 28116 3667 28182 3668
rect 29364 3667 29430 3668
rect 30612 3667 30678 3668
rect 31860 3667 31926 3668
rect 33108 3667 33174 3668
rect 34356 3667 34422 3668
rect 35604 3667 35670 3668
rect 36852 3667 36918 3668
rect 38100 3667 38166 3668
rect 39348 3667 39414 3668
rect 40596 3667 40662 3668
rect 41844 3667 41910 3668
rect 43092 3667 43158 3668
rect 44340 3667 44406 3668
rect 45588 3667 45654 3668
rect 46836 3667 46902 3668
rect 48084 3667 48150 3668
rect 49332 3667 49398 3668
rect 50580 3667 50646 3668
rect 51828 3667 51894 3668
rect 13098 3603 13141 3667
rect 13205 3603 13248 3667
rect 14346 3603 14389 3667
rect 14453 3603 14496 3667
rect 15594 3603 15637 3667
rect 15701 3603 15744 3667
rect 16842 3603 16885 3667
rect 16949 3603 16992 3667
rect 18090 3603 18133 3667
rect 18197 3603 18240 3667
rect 19338 3603 19381 3667
rect 19445 3603 19488 3667
rect 20586 3603 20629 3667
rect 20693 3603 20736 3667
rect 21834 3603 21877 3667
rect 21941 3603 21984 3667
rect 23082 3603 23125 3667
rect 23189 3603 23232 3667
rect 24330 3603 24373 3667
rect 24437 3603 24480 3667
rect 25578 3603 25621 3667
rect 25685 3603 25728 3667
rect 26826 3603 26869 3667
rect 26933 3603 26976 3667
rect 28074 3603 28117 3667
rect 28181 3603 28224 3667
rect 29322 3603 29365 3667
rect 29429 3603 29472 3667
rect 30570 3603 30613 3667
rect 30677 3603 30720 3667
rect 31818 3603 31861 3667
rect 31925 3603 31968 3667
rect 33066 3603 33109 3667
rect 33173 3603 33216 3667
rect 34314 3603 34357 3667
rect 34421 3603 34464 3667
rect 35562 3603 35605 3667
rect 35669 3603 35712 3667
rect 36810 3603 36853 3667
rect 36917 3603 36960 3667
rect 38058 3603 38101 3667
rect 38165 3603 38208 3667
rect 39306 3603 39349 3667
rect 39413 3603 39456 3667
rect 40554 3603 40597 3667
rect 40661 3603 40704 3667
rect 41802 3603 41845 3667
rect 41909 3603 41952 3667
rect 43050 3603 43093 3667
rect 43157 3603 43200 3667
rect 44298 3603 44341 3667
rect 44405 3603 44448 3667
rect 45546 3603 45589 3667
rect 45653 3603 45696 3667
rect 46794 3603 46837 3667
rect 46901 3603 46944 3667
rect 48042 3603 48085 3667
rect 48149 3603 48192 3667
rect 49290 3603 49333 3667
rect 49397 3603 49440 3667
rect 50538 3603 50581 3667
rect 50645 3603 50688 3667
rect 51786 3603 51829 3667
rect 51893 3603 51936 3667
rect 13140 3602 13206 3603
rect 14388 3602 14454 3603
rect 15636 3602 15702 3603
rect 16884 3602 16950 3603
rect 18132 3602 18198 3603
rect 19380 3602 19446 3603
rect 20628 3602 20694 3603
rect 21876 3602 21942 3603
rect 23124 3602 23190 3603
rect 24372 3602 24438 3603
rect 25620 3602 25686 3603
rect 26868 3602 26934 3603
rect 28116 3602 28182 3603
rect 29364 3602 29430 3603
rect 30612 3602 30678 3603
rect 31860 3602 31926 3603
rect 33108 3602 33174 3603
rect 34356 3602 34422 3603
rect 35604 3602 35670 3603
rect 36852 3602 36918 3603
rect 38100 3602 38166 3603
rect 39348 3602 39414 3603
rect 40596 3602 40662 3603
rect 41844 3602 41910 3603
rect 43092 3602 43158 3603
rect 44340 3602 44406 3603
rect 45588 3602 45654 3603
rect 46836 3602 46902 3603
rect 48084 3602 48150 3603
rect 49332 3602 49398 3603
rect 50580 3602 50646 3603
rect 51828 3602 51894 3603
rect 13298 1408 13364 1409
rect 14546 1408 14612 1409
rect 15794 1408 15860 1409
rect 17042 1408 17108 1409
rect 18290 1408 18356 1409
rect 19538 1408 19604 1409
rect 20786 1408 20852 1409
rect 22034 1408 22100 1409
rect 23282 1408 23348 1409
rect 24530 1408 24596 1409
rect 25778 1408 25844 1409
rect 27026 1408 27092 1409
rect 28274 1408 28340 1409
rect 29522 1408 29588 1409
rect 30770 1408 30836 1409
rect 32018 1408 32084 1409
rect 33266 1408 33332 1409
rect 34514 1408 34580 1409
rect 35762 1408 35828 1409
rect 37010 1408 37076 1409
rect 38258 1408 38324 1409
rect 39506 1408 39572 1409
rect 40754 1408 40820 1409
rect 42002 1408 42068 1409
rect 43250 1408 43316 1409
rect 44498 1408 44564 1409
rect 45746 1408 45812 1409
rect 46994 1408 47060 1409
rect 48242 1408 48308 1409
rect 49490 1408 49556 1409
rect 50738 1408 50804 1409
rect 51986 1408 52052 1409
rect 13256 1344 13299 1408
rect 13363 1344 13406 1408
rect 14504 1344 14547 1408
rect 14611 1344 14654 1408
rect 15752 1344 15795 1408
rect 15859 1344 15902 1408
rect 17000 1344 17043 1408
rect 17107 1344 17150 1408
rect 18248 1344 18291 1408
rect 18355 1344 18398 1408
rect 19496 1344 19539 1408
rect 19603 1344 19646 1408
rect 20744 1344 20787 1408
rect 20851 1344 20894 1408
rect 21992 1344 22035 1408
rect 22099 1344 22142 1408
rect 23240 1344 23283 1408
rect 23347 1344 23390 1408
rect 24488 1344 24531 1408
rect 24595 1344 24638 1408
rect 25736 1344 25779 1408
rect 25843 1344 25886 1408
rect 26984 1344 27027 1408
rect 27091 1344 27134 1408
rect 28232 1344 28275 1408
rect 28339 1344 28382 1408
rect 29480 1344 29523 1408
rect 29587 1344 29630 1408
rect 30728 1344 30771 1408
rect 30835 1344 30878 1408
rect 31976 1344 32019 1408
rect 32083 1344 32126 1408
rect 33224 1344 33267 1408
rect 33331 1344 33374 1408
rect 34472 1344 34515 1408
rect 34579 1344 34622 1408
rect 35720 1344 35763 1408
rect 35827 1344 35870 1408
rect 36968 1344 37011 1408
rect 37075 1344 37118 1408
rect 38216 1344 38259 1408
rect 38323 1344 38366 1408
rect 39464 1344 39507 1408
rect 39571 1344 39614 1408
rect 40712 1344 40755 1408
rect 40819 1344 40862 1408
rect 41960 1344 42003 1408
rect 42067 1344 42110 1408
rect 43208 1344 43251 1408
rect 43315 1344 43358 1408
rect 44456 1344 44499 1408
rect 44563 1344 44606 1408
rect 45704 1344 45747 1408
rect 45811 1344 45854 1408
rect 46952 1344 46995 1408
rect 47059 1344 47102 1408
rect 48200 1344 48243 1408
rect 48307 1344 48350 1408
rect 49448 1344 49491 1408
rect 49555 1344 49598 1408
rect 50696 1344 50739 1408
rect 50803 1344 50846 1408
rect 51944 1344 51987 1408
rect 52051 1344 52094 1408
rect 13298 1343 13364 1344
rect 14546 1343 14612 1344
rect 15794 1343 15860 1344
rect 17042 1343 17108 1344
rect 18290 1343 18356 1344
rect 19538 1343 19604 1344
rect 20786 1343 20852 1344
rect 22034 1343 22100 1344
rect 23282 1343 23348 1344
rect 24530 1343 24596 1344
rect 25778 1343 25844 1344
rect 27026 1343 27092 1344
rect 28274 1343 28340 1344
rect 29522 1343 29588 1344
rect 30770 1343 30836 1344
rect 32018 1343 32084 1344
rect 33266 1343 33332 1344
rect 34514 1343 34580 1344
rect 35762 1343 35828 1344
rect 37010 1343 37076 1344
rect 38258 1343 38324 1344
rect 39506 1343 39572 1344
rect 40754 1343 40820 1344
rect 42002 1343 42068 1344
rect 43250 1343 43316 1344
rect 44498 1343 44564 1344
rect 45746 1343 45812 1344
rect 46994 1343 47060 1344
rect 48242 1343 48308 1344
rect 49490 1343 49556 1344
rect 50738 1343 50804 1344
rect 51986 1343 52052 1344
rect 13013 288 13079 289
rect 22997 288 23063 289
rect 32981 288 33047 289
rect 42965 288 43031 289
rect 12971 224 13014 288
rect 13078 224 13121 288
rect 22955 224 22998 288
rect 23062 224 23105 288
rect 32939 224 32982 288
rect 33046 224 33089 288
rect 42923 224 42966 288
rect 43030 224 43073 288
rect 13013 223 13079 224
rect 22997 223 23063 224
rect 32981 223 33047 224
rect 42965 223 43031 224
rect 35128 -848 35134 -784
rect 35198 -786 35204 -784
rect 43087 -786 43093 -784
rect 35198 -846 43093 -786
rect 35198 -848 35204 -846
rect 43087 -848 43093 -846
rect 43157 -848 43163 -784
rect 21112 -1092 21118 -1028
rect 21182 -1030 21188 -1028
rect 28111 -1030 28117 -1028
rect 21182 -1090 28117 -1030
rect 21182 -1092 21188 -1090
rect 28111 -1092 28117 -1090
rect 28181 -1092 28187 -1028
rect 15272 -1336 15278 -1272
rect 15342 -1274 15348 -1272
rect 21871 -1274 21877 -1272
rect 15342 -1334 21877 -1274
rect 15342 -1336 15348 -1334
rect 21871 -1336 21877 -1334
rect 21941 -1336 21947 -1272
rect 16093 -1580 16099 -1516
rect 16163 -1518 16169 -1516
rect 22029 -1518 22035 -1516
rect 16163 -1578 22035 -1518
rect 16163 -1580 16169 -1578
rect 22029 -1580 22035 -1578
rect 22099 -1580 22105 -1516
rect 21933 -1824 21939 -1760
rect 22003 -1762 22009 -1760
rect 28269 -1762 28275 -1760
rect 22003 -1822 28275 -1762
rect 22003 -1824 22009 -1822
rect 28269 -1824 28275 -1822
rect 28339 -1824 28345 -1760
rect 28120 -2068 28126 -2004
rect 28190 -2006 28196 -2004
rect 35599 -2006 35605 -2004
rect 28190 -2066 35605 -2006
rect 28190 -2068 28196 -2066
rect 35599 -2068 35605 -2066
rect 35669 -2068 35675 -2004
rect 28941 -2312 28947 -2248
rect 29011 -2250 29017 -2248
rect 35757 -2250 35763 -2248
rect 29011 -2310 35763 -2250
rect 29011 -2312 29017 -2310
rect 35757 -2312 35763 -2310
rect 35827 -2312 35833 -2248
rect 35949 -2556 35955 -2492
rect 36019 -2494 36025 -2492
rect 43245 -2494 43251 -2492
rect 36019 -2554 43251 -2494
rect 36019 -2556 36025 -2554
rect 43245 -2556 43251 -2554
rect 43315 -2556 43321 -2492
rect 43304 -2800 43310 -2736
rect 43374 -2738 43380 -2736
rect 51823 -2738 51829 -2736
rect 43374 -2798 51829 -2738
rect 43374 -2800 43380 -2798
rect 51823 -2800 51829 -2798
rect 51893 -2800 51899 -2736
rect 33960 -3044 33966 -2980
rect 34030 -2982 34036 -2980
rect 41839 -2982 41845 -2980
rect 34030 -3042 41845 -2982
rect 34030 -3044 34036 -3042
rect 41839 -3044 41845 -3042
rect 41909 -3044 41915 -2980
rect 34781 -3288 34787 -3224
rect 34851 -3226 34857 -3224
rect 41997 -3226 42003 -3224
rect 34851 -3286 42003 -3226
rect 34851 -3288 34857 -3286
rect 41997 -3288 42003 -3286
rect 42067 -3288 42073 -3224
rect 42136 -3532 42142 -3468
rect 42206 -3470 42212 -3468
rect 50575 -3470 50581 -3468
rect 42206 -3530 50581 -3470
rect 42206 -3532 42212 -3530
rect 50575 -3532 50581 -3530
rect 50645 -3532 50651 -3468
rect 18776 -3776 18782 -3712
rect 18846 -3714 18852 -3712
rect 25615 -3714 25621 -3712
rect 18846 -3774 25621 -3714
rect 18846 -3776 18852 -3774
rect 25615 -3776 25621 -3774
rect 25685 -3776 25691 -3712
rect 7096 -4020 7102 -3956
rect 7166 -3958 7172 -3956
rect 13135 -3958 13141 -3956
rect 7166 -4018 13141 -3958
rect 7166 -4020 7172 -4018
rect 13135 -4020 13141 -4018
rect 13205 -4020 13211 -3956
rect 3245 -4264 3251 -4200
rect 3315 -4202 3321 -4200
rect 13008 -4202 13014 -4200
rect 3315 -4262 13014 -4202
rect 3315 -4264 3321 -4262
rect 13008 -4264 13014 -4262
rect 13078 -4264 13084 -4200
rect 12936 -4508 12942 -4444
rect 13006 -4446 13012 -4444
rect 19375 -4446 19381 -4444
rect 13006 -4506 19381 -4446
rect 13006 -4508 13012 -4506
rect 19375 -4508 19381 -4506
rect 19445 -4508 19451 -4444
rect 13757 -4752 13763 -4688
rect 13827 -4690 13833 -4688
rect 19533 -4690 19539 -4688
rect 13827 -4750 19539 -4690
rect 13827 -4752 13833 -4750
rect 19533 -4752 19539 -4750
rect 19603 -4752 19609 -4688
rect 19597 -4996 19603 -4932
rect 19667 -4934 19673 -4932
rect 25773 -4934 25779 -4932
rect 19667 -4994 25779 -4934
rect 19667 -4996 19673 -4994
rect 25773 -4996 25779 -4994
rect 25843 -4996 25849 -4932
rect 25784 -5240 25790 -5176
rect 25854 -5178 25860 -5176
rect 33103 -5178 33109 -5176
rect 25854 -5238 33109 -5178
rect 25854 -5240 25860 -5238
rect 33103 -5240 33109 -5238
rect 33173 -5240 33179 -5176
rect 5581 -5484 5587 -5420
rect 5651 -5422 5657 -5420
rect 32976 -5422 32982 -5420
rect 5651 -5482 32982 -5422
rect 5651 -5484 5657 -5482
rect 32976 -5484 32982 -5482
rect 33046 -5484 33052 -5420
rect 32792 -5728 32798 -5664
rect 32862 -5666 32868 -5664
rect 40591 -5666 40597 -5664
rect 32862 -5726 40597 -5666
rect 32862 -5728 32868 -5726
rect 40591 -5728 40597 -5726
rect 40661 -5728 40667 -5664
rect 33613 -5972 33619 -5908
rect 33683 -5910 33689 -5908
rect 40749 -5910 40755 -5908
rect 33683 -5970 40755 -5910
rect 33683 -5972 33689 -5970
rect 40749 -5972 40755 -5970
rect 40819 -5972 40825 -5908
rect 40968 -6216 40974 -6152
rect 41038 -6154 41044 -6152
rect 49327 -6154 49333 -6152
rect 41038 -6214 49333 -6154
rect 41038 -6216 41044 -6214
rect 49327 -6216 49333 -6214
rect 49397 -6216 49403 -6152
rect 39800 -6460 39806 -6396
rect 39870 -6398 39876 -6396
rect 48079 -6398 48085 -6396
rect 39870 -6458 48085 -6398
rect 39870 -6460 39876 -6458
rect 48079 -6460 48085 -6458
rect 48149 -6460 48155 -6396
rect 38632 -6704 38638 -6640
rect 38702 -6642 38708 -6640
rect 46831 -6642 46837 -6640
rect 38702 -6702 46837 -6642
rect 38702 -6704 38708 -6702
rect 46831 -6704 46837 -6702
rect 46901 -6704 46907 -6640
rect 37464 -6948 37470 -6884
rect 37534 -6886 37540 -6884
rect 45583 -6886 45589 -6884
rect 37534 -6946 45589 -6886
rect 37534 -6948 37540 -6946
rect 45583 -6948 45589 -6946
rect 45653 -6948 45659 -6884
rect 36296 -7192 36302 -7128
rect 36366 -7130 36372 -7128
rect 44335 -7130 44341 -7128
rect 36366 -7190 44341 -7130
rect 36366 -7192 36372 -7190
rect 44335 -7192 44341 -7190
rect 44405 -7192 44411 -7128
rect 17608 -7436 17614 -7372
rect 17678 -7374 17684 -7372
rect 24367 -7374 24373 -7372
rect 17678 -7434 24373 -7374
rect 17678 -7436 17684 -7434
rect 24367 -7436 24373 -7434
rect 24437 -7436 24443 -7372
rect 11768 -7680 11774 -7616
rect 11838 -7618 11844 -7616
rect 18127 -7618 18133 -7616
rect 11838 -7678 18133 -7618
rect 11838 -7680 11844 -7678
rect 18127 -7680 18133 -7678
rect 18197 -7680 18203 -7616
rect 12589 -7924 12595 -7860
rect 12659 -7862 12665 -7860
rect 18285 -7862 18291 -7860
rect 12659 -7922 18291 -7862
rect 12659 -7924 12665 -7922
rect 18285 -7924 18291 -7922
rect 18355 -7924 18361 -7860
rect 18429 -8168 18435 -8104
rect 18499 -8106 18505 -8104
rect 24525 -8106 24531 -8104
rect 18499 -8166 24531 -8106
rect 18499 -8168 18505 -8166
rect 24525 -8168 24531 -8166
rect 24595 -8168 24601 -8104
rect 24616 -8412 24622 -8348
rect 24686 -8350 24692 -8348
rect 31855 -8350 31861 -8348
rect 24686 -8410 31861 -8350
rect 24686 -8412 24692 -8410
rect 31855 -8412 31861 -8410
rect 31925 -8412 31931 -8348
rect 31624 -8656 31630 -8592
rect 31694 -8594 31700 -8592
rect 39343 -8594 39349 -8592
rect 31694 -8654 39349 -8594
rect 31694 -8656 31700 -8654
rect 39343 -8656 39349 -8654
rect 39413 -8656 39419 -8592
rect 16440 -8900 16446 -8836
rect 16510 -8838 16516 -8836
rect 23119 -8838 23125 -8836
rect 16510 -8898 23125 -8838
rect 16510 -8900 16516 -8898
rect 23119 -8900 23125 -8898
rect 23189 -8900 23195 -8836
rect 10600 -9144 10606 -9080
rect 10670 -9082 10676 -9080
rect 16879 -9082 16885 -9080
rect 10670 -9142 16885 -9082
rect 10670 -9144 10676 -9142
rect 16879 -9144 16885 -9142
rect 16949 -9144 16955 -9080
rect 11421 -9388 11427 -9324
rect 11491 -9326 11497 -9324
rect 17037 -9326 17043 -9324
rect 11491 -9386 17043 -9326
rect 11491 -9388 11497 -9386
rect 17037 -9388 17043 -9386
rect 17107 -9388 17113 -9324
rect 17261 -9632 17267 -9568
rect 17331 -9570 17337 -9568
rect 23277 -9570 23283 -9568
rect 17331 -9630 23283 -9570
rect 17331 -9632 17337 -9630
rect 23277 -9632 23283 -9630
rect 23347 -9632 23353 -9568
rect 23448 -9876 23454 -9812
rect 23518 -9814 23524 -9812
rect 30607 -9814 30613 -9812
rect 23518 -9874 30613 -9814
rect 23518 -9876 23524 -9874
rect 30607 -9876 30613 -9874
rect 30677 -9876 30683 -9812
rect 30456 -10120 30462 -10056
rect 30526 -10058 30532 -10056
rect 38095 -10058 38101 -10056
rect 30526 -10118 38101 -10058
rect 30526 -10120 30532 -10118
rect 38095 -10120 38101 -10118
rect 38165 -10120 38171 -10056
rect 22280 -10364 22286 -10300
rect 22350 -10302 22356 -10300
rect 29359 -10302 29365 -10300
rect 22350 -10362 29365 -10302
rect 22350 -10364 22356 -10362
rect 29359 -10364 29365 -10362
rect 29429 -10364 29435 -10300
rect 4413 -10608 4419 -10544
rect 4483 -10546 4489 -10544
rect 22992 -10546 22998 -10544
rect 4483 -10606 22998 -10546
rect 4483 -10608 4489 -10606
rect 22992 -10608 22998 -10606
rect 23062 -10608 23068 -10544
rect 23101 -10852 23107 -10788
rect 23171 -10790 23177 -10788
rect 29517 -10790 29523 -10788
rect 23171 -10850 29523 -10790
rect 23171 -10852 23177 -10850
rect 29517 -10852 29523 -10850
rect 29587 -10852 29593 -10788
rect 29288 -11096 29294 -11032
rect 29358 -11034 29364 -11032
rect 36847 -11034 36853 -11032
rect 29358 -11094 36853 -11034
rect 29358 -11096 29364 -11094
rect 36847 -11096 36853 -11094
rect 36917 -11096 36923 -11032
rect 19944 -11340 19950 -11276
rect 20014 -11278 20020 -11276
rect 26863 -11278 26869 -11276
rect 20014 -11338 26869 -11278
rect 20014 -11340 20020 -11338
rect 26863 -11340 26869 -11338
rect 26933 -11340 26939 -11276
rect 14104 -11584 14110 -11520
rect 14174 -11522 14180 -11520
rect 20623 -11522 20629 -11520
rect 14174 -11582 20629 -11522
rect 14174 -11584 14180 -11582
rect 20623 -11584 20629 -11582
rect 20693 -11584 20699 -11520
rect 14925 -11828 14931 -11764
rect 14995 -11766 15001 -11764
rect 20781 -11766 20787 -11764
rect 14995 -11826 20787 -11766
rect 14995 -11828 15001 -11826
rect 20781 -11828 20787 -11826
rect 20851 -11828 20857 -11764
rect 20765 -12072 20771 -12008
rect 20835 -12010 20841 -12008
rect 27021 -12010 27027 -12008
rect 20835 -12070 27027 -12010
rect 20835 -12072 20841 -12070
rect 27021 -12072 27027 -12070
rect 27091 -12072 27097 -12008
rect 26952 -12316 26958 -12252
rect 27022 -12254 27028 -12252
rect 34351 -12254 34357 -12252
rect 27022 -12314 34357 -12254
rect 27022 -12316 27028 -12314
rect 34351 -12316 34357 -12314
rect 34421 -12316 34427 -12252
rect 9432 -12560 9438 -12496
rect 9502 -12498 9508 -12496
rect 15631 -12498 15637 -12496
rect 9502 -12558 15637 -12498
rect 9502 -12560 9508 -12558
rect 15631 -12560 15637 -12558
rect 15701 -12560 15707 -12496
rect 8264 -12804 8270 -12740
rect 8334 -12742 8340 -12740
rect 14383 -12742 14389 -12740
rect 8334 -12802 14389 -12742
rect 8334 -12804 8340 -12802
rect 14383 -12804 14389 -12802
rect 14453 -12804 14459 -12740
rect 44125 -13048 44131 -12984
rect 44195 -12986 44201 -12984
rect 51981 -12986 51987 -12984
rect 44195 -13046 51987 -12986
rect 44195 -13048 44201 -13046
rect 51981 -13048 51987 -13046
rect 52051 -13048 52057 -12984
rect 6749 -13292 6755 -13228
rect 6819 -13230 6825 -13228
rect 42960 -13230 42966 -13228
rect 6819 -13290 42966 -13230
rect 6819 -13292 6825 -13290
rect 42960 -13292 42966 -13290
rect 43030 -13292 43036 -13228
rect 42957 -13536 42963 -13472
rect 43027 -13474 43033 -13472
rect 50733 -13474 50739 -13472
rect 43027 -13534 50739 -13474
rect 43027 -13536 43033 -13534
rect 50733 -13536 50739 -13534
rect 50803 -13536 50809 -13472
rect 41789 -13780 41795 -13716
rect 41859 -13718 41865 -13716
rect 49485 -13718 49491 -13716
rect 41859 -13778 49491 -13718
rect 41859 -13780 41865 -13778
rect 49485 -13780 49491 -13778
rect 49555 -13780 49561 -13716
rect 40621 -14024 40627 -13960
rect 40691 -13962 40697 -13960
rect 48237 -13962 48243 -13960
rect 40691 -14022 48243 -13962
rect 40691 -14024 40697 -14022
rect 48237 -14024 48243 -14022
rect 48307 -14024 48313 -13960
rect 32445 -14268 32451 -14204
rect 32515 -14206 32521 -14204
rect 39501 -14206 39507 -14204
rect 32515 -14266 39507 -14206
rect 32515 -14268 32521 -14266
rect 39501 -14268 39507 -14266
rect 39571 -14268 39577 -14204
rect 39453 -14512 39459 -14448
rect 39523 -14450 39529 -14448
rect 46989 -14450 46995 -14448
rect 39523 -14510 46995 -14450
rect 39523 -14512 39529 -14510
rect 46989 -14512 46995 -14510
rect 47059 -14512 47065 -14448
rect 31277 -14756 31283 -14692
rect 31347 -14694 31353 -14692
rect 38253 -14694 38259 -14692
rect 31347 -14754 38259 -14694
rect 31347 -14756 31353 -14754
rect 38253 -14756 38259 -14754
rect 38323 -14756 38329 -14692
rect 38285 -15000 38291 -14936
rect 38355 -14938 38361 -14936
rect 45741 -14938 45747 -14936
rect 38355 -14998 45747 -14938
rect 38355 -15000 38361 -14998
rect 45741 -15000 45747 -14998
rect 45811 -15000 45817 -14936
rect 30109 -15244 30115 -15180
rect 30179 -15182 30185 -15180
rect 37005 -15182 37011 -15180
rect 30179 -15242 37011 -15182
rect 30179 -15244 30185 -15242
rect 37005 -15244 37011 -15242
rect 37075 -15244 37081 -15180
rect 37117 -15488 37123 -15424
rect 37187 -15426 37193 -15424
rect 44493 -15426 44499 -15424
rect 37187 -15486 44499 -15426
rect 37187 -15488 37193 -15486
rect 44493 -15488 44499 -15486
rect 44563 -15488 44569 -15424
rect 27773 -15732 27779 -15668
rect 27843 -15670 27849 -15668
rect 34509 -15670 34515 -15668
rect 27843 -15730 34515 -15670
rect 27843 -15732 27849 -15730
rect 34509 -15732 34515 -15730
rect 34579 -15732 34585 -15668
rect 26605 -15976 26611 -15912
rect 26675 -15914 26681 -15912
rect 33261 -15914 33267 -15912
rect 26675 -15974 33267 -15914
rect 26675 -15976 26681 -15974
rect 33261 -15976 33267 -15974
rect 33331 -15976 33337 -15912
rect 25437 -16220 25443 -16156
rect 25507 -16158 25513 -16156
rect 32013 -16158 32019 -16156
rect 25507 -16218 32019 -16158
rect 25507 -16220 25513 -16218
rect 32013 -16220 32019 -16218
rect 32083 -16220 32089 -16156
rect 24269 -16464 24275 -16400
rect 24339 -16402 24345 -16400
rect 30765 -16402 30771 -16400
rect 24339 -16462 30771 -16402
rect 24339 -16464 24345 -16462
rect 30765 -16464 30771 -16462
rect 30835 -16464 30841 -16400
rect 10253 -16708 10259 -16644
rect 10323 -16646 10329 -16644
rect 15789 -16646 15795 -16644
rect 10323 -16706 15795 -16646
rect 10323 -16708 10329 -16706
rect 15789 -16708 15795 -16706
rect 15859 -16708 15865 -16644
rect 9085 -16952 9091 -16888
rect 9155 -16890 9161 -16888
rect 14541 -16890 14547 -16888
rect 9155 -16950 14547 -16890
rect 9155 -16952 9161 -16950
rect 14541 -16952 14547 -16950
rect 14611 -16952 14617 -16888
rect 7917 -17196 7923 -17132
rect 7987 -17134 7993 -17132
rect 13293 -17134 13299 -17132
rect 7987 -17194 13299 -17134
rect 7987 -17196 7993 -17194
rect 13293 -17196 13299 -17194
rect 13363 -17196 13369 -17132
rect 2077 -17440 2083 -17376
rect 2147 -17378 2153 -17376
rect 5979 -17378 5985 -17376
rect 2147 -17438 5985 -17378
rect 2147 -17440 2153 -17438
rect 5979 -17440 5985 -17438
rect 6049 -17440 6055 -17376
rect 2082 -18289 2148 -18288
rect 3250 -18289 3316 -18288
rect 4418 -18289 4484 -18288
rect 5586 -18289 5652 -18288
rect 6754 -18289 6820 -18288
rect 7922 -18289 7988 -18288
rect 9090 -18289 9156 -18288
rect 10258 -18289 10324 -18288
rect 11426 -18289 11492 -18288
rect 12594 -18289 12660 -18288
rect 13762 -18289 13828 -18288
rect 14930 -18289 14996 -18288
rect 16098 -18289 16164 -18288
rect 17266 -18289 17332 -18288
rect 18434 -18289 18500 -18288
rect 19602 -18289 19668 -18288
rect 20770 -18289 20836 -18288
rect 21938 -18289 22004 -18288
rect 23106 -18289 23172 -18288
rect 24274 -18289 24340 -18288
rect 25442 -18289 25508 -18288
rect 26610 -18289 26676 -18288
rect 27778 -18289 27844 -18288
rect 28946 -18289 29012 -18288
rect 30114 -18289 30180 -18288
rect 31282 -18289 31348 -18288
rect 32450 -18289 32516 -18288
rect 33618 -18289 33684 -18288
rect 34786 -18289 34852 -18288
rect 35954 -18289 36020 -18288
rect 37122 -18289 37188 -18288
rect 38290 -18289 38356 -18288
rect 39458 -18289 39524 -18288
rect 40626 -18289 40692 -18288
rect 41794 -18289 41860 -18288
rect 42962 -18289 43028 -18288
rect 44130 -18289 44196 -18288
rect 2040 -18353 2083 -18289
rect 2147 -18353 2190 -18289
rect 3208 -18353 3251 -18289
rect 3315 -18353 3358 -18289
rect 4376 -18353 4419 -18289
rect 4483 -18353 4526 -18289
rect 5544 -18353 5587 -18289
rect 5651 -18353 5694 -18289
rect 6712 -18353 6755 -18289
rect 6819 -18353 6862 -18289
rect 7880 -18353 7923 -18289
rect 7987 -18353 8030 -18289
rect 9048 -18353 9091 -18289
rect 9155 -18353 9198 -18289
rect 10216 -18353 10259 -18289
rect 10323 -18353 10366 -18289
rect 11384 -18353 11427 -18289
rect 11491 -18353 11534 -18289
rect 12552 -18353 12595 -18289
rect 12659 -18353 12702 -18289
rect 13720 -18353 13763 -18289
rect 13827 -18353 13870 -18289
rect 14888 -18353 14931 -18289
rect 14995 -18353 15038 -18289
rect 16056 -18353 16099 -18289
rect 16163 -18353 16206 -18289
rect 17224 -18353 17267 -18289
rect 17331 -18353 17374 -18289
rect 18392 -18353 18435 -18289
rect 18499 -18353 18542 -18289
rect 19560 -18353 19603 -18289
rect 19667 -18353 19710 -18289
rect 20728 -18353 20771 -18289
rect 20835 -18353 20878 -18289
rect 21896 -18353 21939 -18289
rect 22003 -18353 22046 -18289
rect 23064 -18353 23107 -18289
rect 23171 -18353 23214 -18289
rect 24232 -18353 24275 -18289
rect 24339 -18353 24382 -18289
rect 25400 -18353 25443 -18289
rect 25507 -18353 25550 -18289
rect 26568 -18353 26611 -18289
rect 26675 -18353 26718 -18289
rect 27736 -18353 27779 -18289
rect 27843 -18353 27886 -18289
rect 28904 -18353 28947 -18289
rect 29011 -18353 29054 -18289
rect 30072 -18353 30115 -18289
rect 30179 -18353 30222 -18289
rect 31240 -18353 31283 -18289
rect 31347 -18353 31390 -18289
rect 32408 -18353 32451 -18289
rect 32515 -18353 32558 -18289
rect 33576 -18353 33619 -18289
rect 33683 -18353 33726 -18289
rect 34744 -18353 34787 -18289
rect 34851 -18353 34894 -18289
rect 35912 -18353 35955 -18289
rect 36019 -18353 36062 -18289
rect 37080 -18353 37123 -18289
rect 37187 -18353 37230 -18289
rect 38248 -18353 38291 -18289
rect 38355 -18353 38398 -18289
rect 39416 -18353 39459 -18289
rect 39523 -18353 39566 -18289
rect 40584 -18353 40627 -18289
rect 40691 -18353 40734 -18289
rect 41752 -18353 41795 -18289
rect 41859 -18353 41902 -18289
rect 42920 -18353 42963 -18289
rect 43027 -18353 43070 -18289
rect 44088 -18353 44131 -18289
rect 44195 -18353 44238 -18289
rect 2082 -18354 2148 -18353
rect 3250 -18354 3316 -18353
rect 4418 -18354 4484 -18353
rect 5586 -18354 5652 -18353
rect 6754 -18354 6820 -18353
rect 7922 -18354 7988 -18353
rect 9090 -18354 9156 -18353
rect 10258 -18354 10324 -18353
rect 11426 -18354 11492 -18353
rect 12594 -18354 12660 -18353
rect 13762 -18354 13828 -18353
rect 14930 -18354 14996 -18353
rect 16098 -18354 16164 -18353
rect 17266 -18354 17332 -18353
rect 18434 -18354 18500 -18353
rect 19602 -18354 19668 -18353
rect 20770 -18354 20836 -18353
rect 21938 -18354 22004 -18353
rect 23106 -18354 23172 -18353
rect 24274 -18354 24340 -18353
rect 25442 -18354 25508 -18353
rect 26610 -18354 26676 -18353
rect 27778 -18354 27844 -18353
rect 28946 -18354 29012 -18353
rect 30114 -18354 30180 -18353
rect 31282 -18354 31348 -18353
rect 32450 -18354 32516 -18353
rect 33618 -18354 33684 -18353
rect 34786 -18354 34852 -18353
rect 35954 -18354 36020 -18353
rect 37122 -18354 37188 -18353
rect 38290 -18354 38356 -18353
rect 39458 -18354 39524 -18353
rect 40626 -18354 40692 -18353
rect 41794 -18354 41860 -18353
rect 42962 -18354 43028 -18353
rect 44130 -18354 44196 -18353
<< via3 >>
rect 5985 5469 6049 5473
rect 5985 5413 5989 5469
rect 5989 5413 6045 5469
rect 6045 5413 6049 5469
rect 5985 5409 6049 5413
rect 13141 3663 13205 3667
rect 13141 3607 13145 3663
rect 13145 3607 13201 3663
rect 13201 3607 13205 3663
rect 13141 3603 13205 3607
rect 14389 3663 14453 3667
rect 14389 3607 14393 3663
rect 14393 3607 14449 3663
rect 14449 3607 14453 3663
rect 14389 3603 14453 3607
rect 15637 3663 15701 3667
rect 15637 3607 15641 3663
rect 15641 3607 15697 3663
rect 15697 3607 15701 3663
rect 15637 3603 15701 3607
rect 16885 3663 16949 3667
rect 16885 3607 16889 3663
rect 16889 3607 16945 3663
rect 16945 3607 16949 3663
rect 16885 3603 16949 3607
rect 18133 3663 18197 3667
rect 18133 3607 18137 3663
rect 18137 3607 18193 3663
rect 18193 3607 18197 3663
rect 18133 3603 18197 3607
rect 19381 3663 19445 3667
rect 19381 3607 19385 3663
rect 19385 3607 19441 3663
rect 19441 3607 19445 3663
rect 19381 3603 19445 3607
rect 20629 3663 20693 3667
rect 20629 3607 20633 3663
rect 20633 3607 20689 3663
rect 20689 3607 20693 3663
rect 20629 3603 20693 3607
rect 21877 3663 21941 3667
rect 21877 3607 21881 3663
rect 21881 3607 21937 3663
rect 21937 3607 21941 3663
rect 21877 3603 21941 3607
rect 23125 3663 23189 3667
rect 23125 3607 23129 3663
rect 23129 3607 23185 3663
rect 23185 3607 23189 3663
rect 23125 3603 23189 3607
rect 24373 3663 24437 3667
rect 24373 3607 24377 3663
rect 24377 3607 24433 3663
rect 24433 3607 24437 3663
rect 24373 3603 24437 3607
rect 25621 3663 25685 3667
rect 25621 3607 25625 3663
rect 25625 3607 25681 3663
rect 25681 3607 25685 3663
rect 25621 3603 25685 3607
rect 26869 3663 26933 3667
rect 26869 3607 26873 3663
rect 26873 3607 26929 3663
rect 26929 3607 26933 3663
rect 26869 3603 26933 3607
rect 28117 3663 28181 3667
rect 28117 3607 28121 3663
rect 28121 3607 28177 3663
rect 28177 3607 28181 3663
rect 28117 3603 28181 3607
rect 29365 3663 29429 3667
rect 29365 3607 29369 3663
rect 29369 3607 29425 3663
rect 29425 3607 29429 3663
rect 29365 3603 29429 3607
rect 30613 3663 30677 3667
rect 30613 3607 30617 3663
rect 30617 3607 30673 3663
rect 30673 3607 30677 3663
rect 30613 3603 30677 3607
rect 31861 3663 31925 3667
rect 31861 3607 31865 3663
rect 31865 3607 31921 3663
rect 31921 3607 31925 3663
rect 31861 3603 31925 3607
rect 33109 3663 33173 3667
rect 33109 3607 33113 3663
rect 33113 3607 33169 3663
rect 33169 3607 33173 3663
rect 33109 3603 33173 3607
rect 34357 3663 34421 3667
rect 34357 3607 34361 3663
rect 34361 3607 34417 3663
rect 34417 3607 34421 3663
rect 34357 3603 34421 3607
rect 35605 3663 35669 3667
rect 35605 3607 35609 3663
rect 35609 3607 35665 3663
rect 35665 3607 35669 3663
rect 35605 3603 35669 3607
rect 36853 3663 36917 3667
rect 36853 3607 36857 3663
rect 36857 3607 36913 3663
rect 36913 3607 36917 3663
rect 36853 3603 36917 3607
rect 38101 3663 38165 3667
rect 38101 3607 38105 3663
rect 38105 3607 38161 3663
rect 38161 3607 38165 3663
rect 38101 3603 38165 3607
rect 39349 3663 39413 3667
rect 39349 3607 39353 3663
rect 39353 3607 39409 3663
rect 39409 3607 39413 3663
rect 39349 3603 39413 3607
rect 40597 3663 40661 3667
rect 40597 3607 40601 3663
rect 40601 3607 40657 3663
rect 40657 3607 40661 3663
rect 40597 3603 40661 3607
rect 41845 3663 41909 3667
rect 41845 3607 41849 3663
rect 41849 3607 41905 3663
rect 41905 3607 41909 3663
rect 41845 3603 41909 3607
rect 43093 3663 43157 3667
rect 43093 3607 43097 3663
rect 43097 3607 43153 3663
rect 43153 3607 43157 3663
rect 43093 3603 43157 3607
rect 44341 3663 44405 3667
rect 44341 3607 44345 3663
rect 44345 3607 44401 3663
rect 44401 3607 44405 3663
rect 44341 3603 44405 3607
rect 45589 3663 45653 3667
rect 45589 3607 45593 3663
rect 45593 3607 45649 3663
rect 45649 3607 45653 3663
rect 45589 3603 45653 3607
rect 46837 3663 46901 3667
rect 46837 3607 46841 3663
rect 46841 3607 46897 3663
rect 46897 3607 46901 3663
rect 46837 3603 46901 3607
rect 48085 3663 48149 3667
rect 48085 3607 48089 3663
rect 48089 3607 48145 3663
rect 48145 3607 48149 3663
rect 48085 3603 48149 3607
rect 49333 3663 49397 3667
rect 49333 3607 49337 3663
rect 49337 3607 49393 3663
rect 49393 3607 49397 3663
rect 49333 3603 49397 3607
rect 50581 3663 50645 3667
rect 50581 3607 50585 3663
rect 50585 3607 50641 3663
rect 50641 3607 50645 3663
rect 50581 3603 50645 3607
rect 51829 3663 51893 3667
rect 51829 3607 51833 3663
rect 51833 3607 51889 3663
rect 51889 3607 51893 3663
rect 51829 3603 51893 3607
rect 13299 1404 13363 1408
rect 13299 1348 13303 1404
rect 13303 1348 13359 1404
rect 13359 1348 13363 1404
rect 13299 1344 13363 1348
rect 14547 1404 14611 1408
rect 14547 1348 14551 1404
rect 14551 1348 14607 1404
rect 14607 1348 14611 1404
rect 14547 1344 14611 1348
rect 15795 1404 15859 1408
rect 15795 1348 15799 1404
rect 15799 1348 15855 1404
rect 15855 1348 15859 1404
rect 15795 1344 15859 1348
rect 17043 1404 17107 1408
rect 17043 1348 17047 1404
rect 17047 1348 17103 1404
rect 17103 1348 17107 1404
rect 17043 1344 17107 1348
rect 18291 1404 18355 1408
rect 18291 1348 18295 1404
rect 18295 1348 18351 1404
rect 18351 1348 18355 1404
rect 18291 1344 18355 1348
rect 19539 1404 19603 1408
rect 19539 1348 19543 1404
rect 19543 1348 19599 1404
rect 19599 1348 19603 1404
rect 19539 1344 19603 1348
rect 20787 1404 20851 1408
rect 20787 1348 20791 1404
rect 20791 1348 20847 1404
rect 20847 1348 20851 1404
rect 20787 1344 20851 1348
rect 22035 1404 22099 1408
rect 22035 1348 22039 1404
rect 22039 1348 22095 1404
rect 22095 1348 22099 1404
rect 22035 1344 22099 1348
rect 23283 1404 23347 1408
rect 23283 1348 23287 1404
rect 23287 1348 23343 1404
rect 23343 1348 23347 1404
rect 23283 1344 23347 1348
rect 24531 1404 24595 1408
rect 24531 1348 24535 1404
rect 24535 1348 24591 1404
rect 24591 1348 24595 1404
rect 24531 1344 24595 1348
rect 25779 1404 25843 1408
rect 25779 1348 25783 1404
rect 25783 1348 25839 1404
rect 25839 1348 25843 1404
rect 25779 1344 25843 1348
rect 27027 1404 27091 1408
rect 27027 1348 27031 1404
rect 27031 1348 27087 1404
rect 27087 1348 27091 1404
rect 27027 1344 27091 1348
rect 28275 1404 28339 1408
rect 28275 1348 28279 1404
rect 28279 1348 28335 1404
rect 28335 1348 28339 1404
rect 28275 1344 28339 1348
rect 29523 1404 29587 1408
rect 29523 1348 29527 1404
rect 29527 1348 29583 1404
rect 29583 1348 29587 1404
rect 29523 1344 29587 1348
rect 30771 1404 30835 1408
rect 30771 1348 30775 1404
rect 30775 1348 30831 1404
rect 30831 1348 30835 1404
rect 30771 1344 30835 1348
rect 32019 1404 32083 1408
rect 32019 1348 32023 1404
rect 32023 1348 32079 1404
rect 32079 1348 32083 1404
rect 32019 1344 32083 1348
rect 33267 1404 33331 1408
rect 33267 1348 33271 1404
rect 33271 1348 33327 1404
rect 33327 1348 33331 1404
rect 33267 1344 33331 1348
rect 34515 1404 34579 1408
rect 34515 1348 34519 1404
rect 34519 1348 34575 1404
rect 34575 1348 34579 1404
rect 34515 1344 34579 1348
rect 35763 1404 35827 1408
rect 35763 1348 35767 1404
rect 35767 1348 35823 1404
rect 35823 1348 35827 1404
rect 35763 1344 35827 1348
rect 37011 1404 37075 1408
rect 37011 1348 37015 1404
rect 37015 1348 37071 1404
rect 37071 1348 37075 1404
rect 37011 1344 37075 1348
rect 38259 1404 38323 1408
rect 38259 1348 38263 1404
rect 38263 1348 38319 1404
rect 38319 1348 38323 1404
rect 38259 1344 38323 1348
rect 39507 1404 39571 1408
rect 39507 1348 39511 1404
rect 39511 1348 39567 1404
rect 39567 1348 39571 1404
rect 39507 1344 39571 1348
rect 40755 1404 40819 1408
rect 40755 1348 40759 1404
rect 40759 1348 40815 1404
rect 40815 1348 40819 1404
rect 40755 1344 40819 1348
rect 42003 1404 42067 1408
rect 42003 1348 42007 1404
rect 42007 1348 42063 1404
rect 42063 1348 42067 1404
rect 42003 1344 42067 1348
rect 43251 1404 43315 1408
rect 43251 1348 43255 1404
rect 43255 1348 43311 1404
rect 43311 1348 43315 1404
rect 43251 1344 43315 1348
rect 44499 1404 44563 1408
rect 44499 1348 44503 1404
rect 44503 1348 44559 1404
rect 44559 1348 44563 1404
rect 44499 1344 44563 1348
rect 45747 1404 45811 1408
rect 45747 1348 45751 1404
rect 45751 1348 45807 1404
rect 45807 1348 45811 1404
rect 45747 1344 45811 1348
rect 46995 1404 47059 1408
rect 46995 1348 46999 1404
rect 46999 1348 47055 1404
rect 47055 1348 47059 1404
rect 46995 1344 47059 1348
rect 48243 1404 48307 1408
rect 48243 1348 48247 1404
rect 48247 1348 48303 1404
rect 48303 1348 48307 1404
rect 48243 1344 48307 1348
rect 49491 1404 49555 1408
rect 49491 1348 49495 1404
rect 49495 1348 49551 1404
rect 49551 1348 49555 1404
rect 49491 1344 49555 1348
rect 50739 1404 50803 1408
rect 50739 1348 50743 1404
rect 50743 1348 50799 1404
rect 50799 1348 50803 1404
rect 50739 1344 50803 1348
rect 51987 1404 52051 1408
rect 51987 1348 51991 1404
rect 51991 1348 52047 1404
rect 52047 1348 52051 1404
rect 51987 1344 52051 1348
rect 13014 284 13078 288
rect 13014 228 13018 284
rect 13018 228 13074 284
rect 13074 228 13078 284
rect 13014 224 13078 228
rect 22998 284 23062 288
rect 22998 228 23002 284
rect 23002 228 23058 284
rect 23058 228 23062 284
rect 22998 224 23062 228
rect 32982 284 33046 288
rect 32982 228 32986 284
rect 32986 228 33042 284
rect 33042 228 33046 284
rect 32982 224 33046 228
rect 42966 284 43030 288
rect 42966 228 42970 284
rect 42970 228 43026 284
rect 43026 228 43030 284
rect 42966 224 43030 228
rect 35134 -848 35198 -784
rect 43093 -848 43157 -784
rect 21118 -1092 21182 -1028
rect 28117 -1092 28181 -1028
rect 15278 -1336 15342 -1272
rect 21877 -1336 21941 -1272
rect 16099 -1580 16163 -1516
rect 22035 -1580 22099 -1516
rect 21939 -1824 22003 -1760
rect 28275 -1824 28339 -1760
rect 28126 -2068 28190 -2004
rect 35605 -2068 35669 -2004
rect 28947 -2312 29011 -2248
rect 35763 -2312 35827 -2248
rect 35955 -2556 36019 -2492
rect 43251 -2556 43315 -2492
rect 43310 -2800 43374 -2736
rect 51829 -2800 51893 -2736
rect 33966 -3044 34030 -2980
rect 41845 -3044 41909 -2980
rect 34787 -3288 34851 -3224
rect 42003 -3288 42067 -3224
rect 42142 -3532 42206 -3468
rect 50581 -3532 50645 -3468
rect 18782 -3776 18846 -3712
rect 25621 -3776 25685 -3712
rect 7102 -4020 7166 -3956
rect 13141 -4020 13205 -3956
rect 3251 -4264 3315 -4200
rect 13014 -4264 13078 -4200
rect 12942 -4508 13006 -4444
rect 19381 -4508 19445 -4444
rect 13763 -4752 13827 -4688
rect 19539 -4752 19603 -4688
rect 19603 -4996 19667 -4932
rect 25779 -4996 25843 -4932
rect 25790 -5240 25854 -5176
rect 33109 -5240 33173 -5176
rect 5587 -5484 5651 -5420
rect 32982 -5484 33046 -5420
rect 32798 -5728 32862 -5664
rect 40597 -5728 40661 -5664
rect 33619 -5972 33683 -5908
rect 40755 -5972 40819 -5908
rect 40974 -6216 41038 -6152
rect 49333 -6216 49397 -6152
rect 39806 -6460 39870 -6396
rect 48085 -6460 48149 -6396
rect 38638 -6704 38702 -6640
rect 46837 -6704 46901 -6640
rect 37470 -6948 37534 -6884
rect 45589 -6948 45653 -6884
rect 36302 -7192 36366 -7128
rect 44341 -7192 44405 -7128
rect 17614 -7436 17678 -7372
rect 24373 -7436 24437 -7372
rect 11774 -7680 11838 -7616
rect 18133 -7680 18197 -7616
rect 12595 -7924 12659 -7860
rect 18291 -7924 18355 -7860
rect 18435 -8168 18499 -8104
rect 24531 -8168 24595 -8104
rect 24622 -8412 24686 -8348
rect 31861 -8412 31925 -8348
rect 31630 -8656 31694 -8592
rect 39349 -8656 39413 -8592
rect 16446 -8900 16510 -8836
rect 23125 -8900 23189 -8836
rect 10606 -9144 10670 -9080
rect 16885 -9144 16949 -9080
rect 11427 -9388 11491 -9324
rect 17043 -9388 17107 -9324
rect 17267 -9632 17331 -9568
rect 23283 -9632 23347 -9568
rect 23454 -9876 23518 -9812
rect 30613 -9876 30677 -9812
rect 30462 -10120 30526 -10056
rect 38101 -10120 38165 -10056
rect 22286 -10364 22350 -10300
rect 29365 -10364 29429 -10300
rect 4419 -10608 4483 -10544
rect 22998 -10608 23062 -10544
rect 23107 -10852 23171 -10788
rect 29523 -10852 29587 -10788
rect 29294 -11096 29358 -11032
rect 36853 -11096 36917 -11032
rect 19950 -11340 20014 -11276
rect 26869 -11340 26933 -11276
rect 14110 -11584 14174 -11520
rect 20629 -11584 20693 -11520
rect 14931 -11828 14995 -11764
rect 20787 -11828 20851 -11764
rect 20771 -12072 20835 -12008
rect 27027 -12072 27091 -12008
rect 26958 -12316 27022 -12252
rect 34357 -12316 34421 -12252
rect 9438 -12560 9502 -12496
rect 15637 -12560 15701 -12496
rect 8270 -12804 8334 -12740
rect 14389 -12804 14453 -12740
rect 44131 -13048 44195 -12984
rect 51987 -13048 52051 -12984
rect 6755 -13292 6819 -13228
rect 42966 -13292 43030 -13228
rect 42963 -13536 43027 -13472
rect 50739 -13536 50803 -13472
rect 41795 -13780 41859 -13716
rect 49491 -13780 49555 -13716
rect 40627 -14024 40691 -13960
rect 48243 -14024 48307 -13960
rect 32451 -14268 32515 -14204
rect 39507 -14268 39571 -14204
rect 39459 -14512 39523 -14448
rect 46995 -14512 47059 -14448
rect 31283 -14756 31347 -14692
rect 38259 -14756 38323 -14692
rect 38291 -15000 38355 -14936
rect 45747 -15000 45811 -14936
rect 30115 -15244 30179 -15180
rect 37011 -15244 37075 -15180
rect 37123 -15488 37187 -15424
rect 44499 -15488 44563 -15424
rect 27779 -15732 27843 -15668
rect 34515 -15732 34579 -15668
rect 26611 -15976 26675 -15912
rect 33267 -15976 33331 -15912
rect 25443 -16220 25507 -16156
rect 32019 -16220 32083 -16156
rect 24275 -16464 24339 -16400
rect 30771 -16464 30835 -16400
rect 10259 -16708 10323 -16644
rect 15795 -16708 15859 -16644
rect 9091 -16952 9155 -16888
rect 14547 -16952 14611 -16888
rect 7923 -17196 7987 -17132
rect 13299 -17196 13363 -17132
rect 2083 -17440 2147 -17376
rect 5985 -17440 6049 -17376
rect 2083 -18293 2147 -18289
rect 2083 -18349 2087 -18293
rect 2087 -18349 2143 -18293
rect 2143 -18349 2147 -18293
rect 2083 -18353 2147 -18349
rect 3251 -18293 3315 -18289
rect 3251 -18349 3255 -18293
rect 3255 -18349 3311 -18293
rect 3311 -18349 3315 -18293
rect 3251 -18353 3315 -18349
rect 4419 -18293 4483 -18289
rect 4419 -18349 4423 -18293
rect 4423 -18349 4479 -18293
rect 4479 -18349 4483 -18293
rect 4419 -18353 4483 -18349
rect 5587 -18293 5651 -18289
rect 5587 -18349 5591 -18293
rect 5591 -18349 5647 -18293
rect 5647 -18349 5651 -18293
rect 5587 -18353 5651 -18349
rect 6755 -18293 6819 -18289
rect 6755 -18349 6759 -18293
rect 6759 -18349 6815 -18293
rect 6815 -18349 6819 -18293
rect 6755 -18353 6819 -18349
rect 7923 -18293 7987 -18289
rect 7923 -18349 7927 -18293
rect 7927 -18349 7983 -18293
rect 7983 -18349 7987 -18293
rect 7923 -18353 7987 -18349
rect 9091 -18293 9155 -18289
rect 9091 -18349 9095 -18293
rect 9095 -18349 9151 -18293
rect 9151 -18349 9155 -18293
rect 9091 -18353 9155 -18349
rect 10259 -18293 10323 -18289
rect 10259 -18349 10263 -18293
rect 10263 -18349 10319 -18293
rect 10319 -18349 10323 -18293
rect 10259 -18353 10323 -18349
rect 11427 -18293 11491 -18289
rect 11427 -18349 11431 -18293
rect 11431 -18349 11487 -18293
rect 11487 -18349 11491 -18293
rect 11427 -18353 11491 -18349
rect 12595 -18293 12659 -18289
rect 12595 -18349 12599 -18293
rect 12599 -18349 12655 -18293
rect 12655 -18349 12659 -18293
rect 12595 -18353 12659 -18349
rect 13763 -18293 13827 -18289
rect 13763 -18349 13767 -18293
rect 13767 -18349 13823 -18293
rect 13823 -18349 13827 -18293
rect 13763 -18353 13827 -18349
rect 14931 -18293 14995 -18289
rect 14931 -18349 14935 -18293
rect 14935 -18349 14991 -18293
rect 14991 -18349 14995 -18293
rect 14931 -18353 14995 -18349
rect 16099 -18293 16163 -18289
rect 16099 -18349 16103 -18293
rect 16103 -18349 16159 -18293
rect 16159 -18349 16163 -18293
rect 16099 -18353 16163 -18349
rect 17267 -18293 17331 -18289
rect 17267 -18349 17271 -18293
rect 17271 -18349 17327 -18293
rect 17327 -18349 17331 -18293
rect 17267 -18353 17331 -18349
rect 18435 -18293 18499 -18289
rect 18435 -18349 18439 -18293
rect 18439 -18349 18495 -18293
rect 18495 -18349 18499 -18293
rect 18435 -18353 18499 -18349
rect 19603 -18293 19667 -18289
rect 19603 -18349 19607 -18293
rect 19607 -18349 19663 -18293
rect 19663 -18349 19667 -18293
rect 19603 -18353 19667 -18349
rect 20771 -18293 20835 -18289
rect 20771 -18349 20775 -18293
rect 20775 -18349 20831 -18293
rect 20831 -18349 20835 -18293
rect 20771 -18353 20835 -18349
rect 21939 -18293 22003 -18289
rect 21939 -18349 21943 -18293
rect 21943 -18349 21999 -18293
rect 21999 -18349 22003 -18293
rect 21939 -18353 22003 -18349
rect 23107 -18293 23171 -18289
rect 23107 -18349 23111 -18293
rect 23111 -18349 23167 -18293
rect 23167 -18349 23171 -18293
rect 23107 -18353 23171 -18349
rect 24275 -18293 24339 -18289
rect 24275 -18349 24279 -18293
rect 24279 -18349 24335 -18293
rect 24335 -18349 24339 -18293
rect 24275 -18353 24339 -18349
rect 25443 -18293 25507 -18289
rect 25443 -18349 25447 -18293
rect 25447 -18349 25503 -18293
rect 25503 -18349 25507 -18293
rect 25443 -18353 25507 -18349
rect 26611 -18293 26675 -18289
rect 26611 -18349 26615 -18293
rect 26615 -18349 26671 -18293
rect 26671 -18349 26675 -18293
rect 26611 -18353 26675 -18349
rect 27779 -18293 27843 -18289
rect 27779 -18349 27783 -18293
rect 27783 -18349 27839 -18293
rect 27839 -18349 27843 -18293
rect 27779 -18353 27843 -18349
rect 28947 -18293 29011 -18289
rect 28947 -18349 28951 -18293
rect 28951 -18349 29007 -18293
rect 29007 -18349 29011 -18293
rect 28947 -18353 29011 -18349
rect 30115 -18293 30179 -18289
rect 30115 -18349 30119 -18293
rect 30119 -18349 30175 -18293
rect 30175 -18349 30179 -18293
rect 30115 -18353 30179 -18349
rect 31283 -18293 31347 -18289
rect 31283 -18349 31287 -18293
rect 31287 -18349 31343 -18293
rect 31343 -18349 31347 -18293
rect 31283 -18353 31347 -18349
rect 32451 -18293 32515 -18289
rect 32451 -18349 32455 -18293
rect 32455 -18349 32511 -18293
rect 32511 -18349 32515 -18293
rect 32451 -18353 32515 -18349
rect 33619 -18293 33683 -18289
rect 33619 -18349 33623 -18293
rect 33623 -18349 33679 -18293
rect 33679 -18349 33683 -18293
rect 33619 -18353 33683 -18349
rect 34787 -18293 34851 -18289
rect 34787 -18349 34791 -18293
rect 34791 -18349 34847 -18293
rect 34847 -18349 34851 -18293
rect 34787 -18353 34851 -18349
rect 35955 -18293 36019 -18289
rect 35955 -18349 35959 -18293
rect 35959 -18349 36015 -18293
rect 36015 -18349 36019 -18293
rect 35955 -18353 36019 -18349
rect 37123 -18293 37187 -18289
rect 37123 -18349 37127 -18293
rect 37127 -18349 37183 -18293
rect 37183 -18349 37187 -18293
rect 37123 -18353 37187 -18349
rect 38291 -18293 38355 -18289
rect 38291 -18349 38295 -18293
rect 38295 -18349 38351 -18293
rect 38351 -18349 38355 -18293
rect 38291 -18353 38355 -18349
rect 39459 -18293 39523 -18289
rect 39459 -18349 39463 -18293
rect 39463 -18349 39519 -18293
rect 39519 -18349 39523 -18293
rect 39459 -18353 39523 -18349
rect 40627 -18293 40691 -18289
rect 40627 -18349 40631 -18293
rect 40631 -18349 40687 -18293
rect 40687 -18349 40691 -18293
rect 40627 -18353 40691 -18349
rect 41795 -18293 41859 -18289
rect 41795 -18349 41799 -18293
rect 41799 -18349 41855 -18293
rect 41855 -18349 41859 -18293
rect 41795 -18353 41859 -18349
rect 42963 -18293 43027 -18289
rect 42963 -18349 42967 -18293
rect 42967 -18349 43023 -18293
rect 43023 -18349 43027 -18293
rect 42963 -18353 43027 -18349
rect 44131 -18293 44195 -18289
rect 44131 -18349 44135 -18293
rect 44135 -18349 44191 -18293
rect 44191 -18349 44195 -18293
rect 44131 -18353 44195 -18349
<< metal4 >>
rect 5984 5473 6050 5474
rect 5984 5409 5985 5473
rect 6049 5409 6050 5473
rect 5984 5408 6050 5409
rect 3250 -4200 3316 -4199
rect 3250 -4264 3251 -4200
rect 3315 -4264 3316 -4200
rect 3250 -4265 3316 -4264
rect 2082 -17376 2148 -17375
rect 2082 -17440 2083 -17376
rect 2147 -17440 2148 -17376
rect 2082 -17441 2148 -17440
rect 2085 -18288 2145 -17441
rect 3253 -18288 3313 -4265
rect 5586 -5420 5652 -5419
rect 5586 -5484 5587 -5420
rect 5651 -5484 5652 -5420
rect 5586 -5485 5652 -5484
rect 4418 -10544 4484 -10543
rect 4418 -10608 4419 -10544
rect 4483 -10608 4484 -10544
rect 4418 -10609 4484 -10608
rect 4421 -18288 4481 -10609
rect 5589 -18288 5649 -5485
rect 5987 -17375 6047 5408
rect 13140 3667 13206 3668
rect 13140 3603 13141 3667
rect 13205 3603 13206 3667
rect 13140 3602 13206 3603
rect 14388 3667 14454 3668
rect 14388 3603 14389 3667
rect 14453 3603 14454 3667
rect 14388 3602 14454 3603
rect 15636 3667 15702 3668
rect 15636 3603 15637 3667
rect 15701 3603 15702 3667
rect 15636 3602 15702 3603
rect 16884 3667 16950 3668
rect 16884 3603 16885 3667
rect 16949 3603 16950 3667
rect 16884 3602 16950 3603
rect 18132 3667 18198 3668
rect 18132 3603 18133 3667
rect 18197 3603 18198 3667
rect 18132 3602 18198 3603
rect 19380 3667 19446 3668
rect 19380 3603 19381 3667
rect 19445 3603 19446 3667
rect 19380 3602 19446 3603
rect 20628 3667 20694 3668
rect 20628 3603 20629 3667
rect 20693 3603 20694 3667
rect 20628 3602 20694 3603
rect 21876 3667 21942 3668
rect 21876 3603 21877 3667
rect 21941 3603 21942 3667
rect 21876 3602 21942 3603
rect 23124 3667 23190 3668
rect 23124 3603 23125 3667
rect 23189 3603 23190 3667
rect 23124 3602 23190 3603
rect 24372 3667 24438 3668
rect 24372 3603 24373 3667
rect 24437 3603 24438 3667
rect 24372 3602 24438 3603
rect 25620 3667 25686 3668
rect 25620 3603 25621 3667
rect 25685 3603 25686 3667
rect 25620 3602 25686 3603
rect 26868 3667 26934 3668
rect 26868 3603 26869 3667
rect 26933 3603 26934 3667
rect 26868 3602 26934 3603
rect 28116 3667 28182 3668
rect 28116 3603 28117 3667
rect 28181 3603 28182 3667
rect 28116 3602 28182 3603
rect 29364 3667 29430 3668
rect 29364 3603 29365 3667
rect 29429 3603 29430 3667
rect 29364 3602 29430 3603
rect 30612 3667 30678 3668
rect 30612 3603 30613 3667
rect 30677 3603 30678 3667
rect 30612 3602 30678 3603
rect 31860 3667 31926 3668
rect 31860 3603 31861 3667
rect 31925 3603 31926 3667
rect 31860 3602 31926 3603
rect 33108 3667 33174 3668
rect 33108 3603 33109 3667
rect 33173 3603 33174 3667
rect 33108 3602 33174 3603
rect 34356 3667 34422 3668
rect 34356 3603 34357 3667
rect 34421 3603 34422 3667
rect 34356 3602 34422 3603
rect 35604 3667 35670 3668
rect 35604 3603 35605 3667
rect 35669 3603 35670 3667
rect 35604 3602 35670 3603
rect 36852 3667 36918 3668
rect 36852 3603 36853 3667
rect 36917 3603 36918 3667
rect 36852 3602 36918 3603
rect 38100 3667 38166 3668
rect 38100 3603 38101 3667
rect 38165 3603 38166 3667
rect 38100 3602 38166 3603
rect 39348 3667 39414 3668
rect 39348 3603 39349 3667
rect 39413 3603 39414 3667
rect 39348 3602 39414 3603
rect 40596 3667 40662 3668
rect 40596 3603 40597 3667
rect 40661 3603 40662 3667
rect 40596 3602 40662 3603
rect 41844 3667 41910 3668
rect 41844 3603 41845 3667
rect 41909 3603 41910 3667
rect 41844 3602 41910 3603
rect 43092 3667 43158 3668
rect 43092 3603 43093 3667
rect 43157 3603 43158 3667
rect 43092 3602 43158 3603
rect 44340 3667 44406 3668
rect 44340 3603 44341 3667
rect 44405 3603 44406 3667
rect 44340 3602 44406 3603
rect 45588 3667 45654 3668
rect 45588 3603 45589 3667
rect 45653 3603 45654 3667
rect 45588 3602 45654 3603
rect 46836 3667 46902 3668
rect 46836 3603 46837 3667
rect 46901 3603 46902 3667
rect 46836 3602 46902 3603
rect 48084 3667 48150 3668
rect 48084 3603 48085 3667
rect 48149 3603 48150 3667
rect 48084 3602 48150 3603
rect 49332 3667 49398 3668
rect 49332 3603 49333 3667
rect 49397 3603 49398 3667
rect 49332 3602 49398 3603
rect 50580 3667 50646 3668
rect 50580 3603 50581 3667
rect 50645 3603 50646 3667
rect 50580 3602 50646 3603
rect 51828 3667 51894 3668
rect 51828 3603 51829 3667
rect 51893 3603 51894 3667
rect 51828 3602 51894 3603
rect 13013 288 13079 289
rect 13013 224 13014 288
rect 13078 224 13079 288
rect 13013 223 13079 224
rect 7101 -3956 7167 -3955
rect 7101 -4020 7102 -3956
rect 7166 -4020 7167 -3956
rect 7101 -4021 7167 -4020
rect 6754 -13228 6820 -13227
rect 6754 -13292 6755 -13228
rect 6819 -13292 6820 -13228
rect 6754 -13293 6820 -13292
rect 5984 -17376 6050 -17375
rect 5984 -17440 5985 -17376
rect 6049 -17440 6050 -17376
rect 5984 -17441 6050 -17440
rect 6757 -18288 6817 -13293
rect 2082 -18289 2148 -18288
rect 2082 -18353 2083 -18289
rect 2147 -18353 2148 -18289
rect 2082 -18354 2148 -18353
rect 3250 -18289 3316 -18288
rect 3250 -18353 3251 -18289
rect 3315 -18353 3316 -18289
rect 3250 -18354 3316 -18353
rect 4418 -18289 4484 -18288
rect 4418 -18353 4419 -18289
rect 4483 -18353 4484 -18289
rect 4418 -18354 4484 -18353
rect 5586 -18289 5652 -18288
rect 5586 -18353 5587 -18289
rect 5651 -18353 5652 -18289
rect 5586 -18354 5652 -18353
rect 6754 -18289 6820 -18288
rect 6754 -18353 6755 -18289
rect 6819 -18353 6820 -18289
rect 6754 -18354 6820 -18353
rect 7104 -18982 7164 -4021
rect 13016 -4199 13076 223
rect 13143 -3955 13203 3602
rect 13298 1408 13364 1409
rect 13298 1344 13299 1408
rect 13363 1344 13364 1408
rect 13298 1343 13364 1344
rect 13140 -3956 13206 -3955
rect 13140 -4020 13141 -3956
rect 13205 -4020 13206 -3956
rect 13140 -4021 13206 -4020
rect 13013 -4200 13079 -4199
rect 13013 -4264 13014 -4200
rect 13078 -4264 13079 -4200
rect 13013 -4265 13079 -4264
rect 12941 -4444 13007 -4443
rect 12941 -4508 12942 -4444
rect 13006 -4508 13007 -4444
rect 12941 -4509 13007 -4508
rect 11773 -7616 11839 -7615
rect 11773 -7680 11774 -7616
rect 11838 -7680 11839 -7616
rect 11773 -7681 11839 -7680
rect 10605 -9080 10671 -9079
rect 10605 -9144 10606 -9080
rect 10670 -9144 10671 -9080
rect 10605 -9145 10671 -9144
rect 9437 -12496 9503 -12495
rect 9437 -12560 9438 -12496
rect 9502 -12560 9503 -12496
rect 9437 -12561 9503 -12560
rect 8269 -12740 8335 -12739
rect 8269 -12804 8270 -12740
rect 8334 -12804 8335 -12740
rect 8269 -12805 8335 -12804
rect 7922 -17132 7988 -17131
rect 7922 -17196 7923 -17132
rect 7987 -17196 7988 -17132
rect 7922 -17197 7988 -17196
rect 7925 -18288 7985 -17197
rect 7922 -18289 7988 -18288
rect 7922 -18353 7923 -18289
rect 7987 -18353 7988 -18289
rect 7922 -18354 7988 -18353
rect 8272 -18982 8332 -12805
rect 9090 -16888 9156 -16887
rect 9090 -16952 9091 -16888
rect 9155 -16952 9156 -16888
rect 9090 -16953 9156 -16952
rect 9093 -18288 9153 -16953
rect 9090 -18289 9156 -18288
rect 9090 -18353 9091 -18289
rect 9155 -18353 9156 -18289
rect 9090 -18354 9156 -18353
rect 9440 -18982 9500 -12561
rect 10258 -16644 10324 -16643
rect 10258 -16708 10259 -16644
rect 10323 -16708 10324 -16644
rect 10258 -16709 10324 -16708
rect 10261 -18288 10321 -16709
rect 10258 -18289 10324 -18288
rect 10258 -18353 10259 -18289
rect 10323 -18353 10324 -18289
rect 10258 -18354 10324 -18353
rect 10608 -18982 10668 -9145
rect 11426 -9324 11492 -9323
rect 11426 -9388 11427 -9324
rect 11491 -9388 11492 -9324
rect 11426 -9389 11492 -9388
rect 11429 -18288 11489 -9389
rect 11426 -18289 11492 -18288
rect 11426 -18353 11427 -18289
rect 11491 -18353 11492 -18289
rect 11426 -18354 11492 -18353
rect 11776 -18982 11836 -7681
rect 12594 -7860 12660 -7859
rect 12594 -7924 12595 -7860
rect 12659 -7924 12660 -7860
rect 12594 -7925 12660 -7924
rect 12597 -18288 12657 -7925
rect 12594 -18289 12660 -18288
rect 12594 -18353 12595 -18289
rect 12659 -18353 12660 -18289
rect 12594 -18354 12660 -18353
rect 12944 -18982 13004 -4509
rect 13301 -17131 13361 1343
rect 13762 -4688 13828 -4687
rect 13762 -4752 13763 -4688
rect 13827 -4752 13828 -4688
rect 13762 -4753 13828 -4752
rect 13298 -17132 13364 -17131
rect 13298 -17196 13299 -17132
rect 13363 -17196 13364 -17132
rect 13298 -17197 13364 -17196
rect 13765 -18288 13825 -4753
rect 14109 -11520 14175 -11519
rect 14109 -11584 14110 -11520
rect 14174 -11584 14175 -11520
rect 14109 -11585 14175 -11584
rect 13762 -18289 13828 -18288
rect 13762 -18353 13763 -18289
rect 13827 -18353 13828 -18289
rect 13762 -18354 13828 -18353
rect 14112 -18982 14172 -11585
rect 14391 -12739 14451 3602
rect 14546 1408 14612 1409
rect 14546 1344 14547 1408
rect 14611 1344 14612 1408
rect 14546 1343 14612 1344
rect 14388 -12740 14454 -12739
rect 14388 -12804 14389 -12740
rect 14453 -12804 14454 -12740
rect 14388 -12805 14454 -12804
rect 14549 -16887 14609 1343
rect 15277 -1272 15343 -1271
rect 15277 -1336 15278 -1272
rect 15342 -1336 15343 -1272
rect 15277 -1337 15343 -1336
rect 14930 -11764 14996 -11763
rect 14930 -11828 14931 -11764
rect 14995 -11828 14996 -11764
rect 14930 -11829 14996 -11828
rect 14546 -16888 14612 -16887
rect 14546 -16952 14547 -16888
rect 14611 -16952 14612 -16888
rect 14546 -16953 14612 -16952
rect 14933 -18288 14993 -11829
rect 14930 -18289 14996 -18288
rect 14930 -18353 14931 -18289
rect 14995 -18353 14996 -18289
rect 14930 -18354 14996 -18353
rect 15280 -18982 15340 -1337
rect 15639 -12495 15699 3602
rect 15794 1408 15860 1409
rect 15794 1344 15795 1408
rect 15859 1344 15860 1408
rect 15794 1343 15860 1344
rect 15636 -12496 15702 -12495
rect 15636 -12560 15637 -12496
rect 15701 -12560 15702 -12496
rect 15636 -12561 15702 -12560
rect 15797 -16643 15857 1343
rect 16098 -1516 16164 -1515
rect 16098 -1580 16099 -1516
rect 16163 -1580 16164 -1516
rect 16098 -1581 16164 -1580
rect 15794 -16644 15860 -16643
rect 15794 -16708 15795 -16644
rect 15859 -16708 15860 -16644
rect 15794 -16709 15860 -16708
rect 16101 -18288 16161 -1581
rect 16445 -8836 16511 -8835
rect 16445 -8900 16446 -8836
rect 16510 -8900 16511 -8836
rect 16445 -8901 16511 -8900
rect 16098 -18289 16164 -18288
rect 16098 -18353 16099 -18289
rect 16163 -18353 16164 -18289
rect 16098 -18354 16164 -18353
rect 16448 -18982 16508 -8901
rect 16887 -9079 16947 3602
rect 17042 1408 17108 1409
rect 17042 1344 17043 1408
rect 17107 1344 17108 1408
rect 17042 1343 17108 1344
rect 16884 -9080 16950 -9079
rect 16884 -9144 16885 -9080
rect 16949 -9144 16950 -9080
rect 16884 -9145 16950 -9144
rect 17045 -9323 17105 1343
rect 17613 -7372 17679 -7371
rect 17613 -7436 17614 -7372
rect 17678 -7436 17679 -7372
rect 17613 -7437 17679 -7436
rect 17042 -9324 17108 -9323
rect 17042 -9388 17043 -9324
rect 17107 -9388 17108 -9324
rect 17042 -9389 17108 -9388
rect 17266 -9568 17332 -9567
rect 17266 -9632 17267 -9568
rect 17331 -9632 17332 -9568
rect 17266 -9633 17332 -9632
rect 17269 -18288 17329 -9633
rect 17266 -18289 17332 -18288
rect 17266 -18353 17267 -18289
rect 17331 -18353 17332 -18289
rect 17266 -18354 17332 -18353
rect 17616 -18982 17676 -7437
rect 18135 -7615 18195 3602
rect 18290 1408 18356 1409
rect 18290 1344 18291 1408
rect 18355 1344 18356 1408
rect 18290 1343 18356 1344
rect 18132 -7616 18198 -7615
rect 18132 -7680 18133 -7616
rect 18197 -7680 18198 -7616
rect 18132 -7681 18198 -7680
rect 18293 -7859 18353 1343
rect 18781 -3712 18847 -3711
rect 18781 -3776 18782 -3712
rect 18846 -3776 18847 -3712
rect 18781 -3777 18847 -3776
rect 18290 -7860 18356 -7859
rect 18290 -7924 18291 -7860
rect 18355 -7924 18356 -7860
rect 18290 -7925 18356 -7924
rect 18434 -8104 18500 -8103
rect 18434 -8168 18435 -8104
rect 18499 -8168 18500 -8104
rect 18434 -8169 18500 -8168
rect 18437 -18288 18497 -8169
rect 18434 -18289 18500 -18288
rect 18434 -18353 18435 -18289
rect 18499 -18353 18500 -18289
rect 18434 -18354 18500 -18353
rect 18784 -18982 18844 -3777
rect 19383 -4443 19443 3602
rect 19538 1408 19604 1409
rect 19538 1344 19539 1408
rect 19603 1344 19604 1408
rect 19538 1343 19604 1344
rect 19380 -4444 19446 -4443
rect 19380 -4508 19381 -4444
rect 19445 -4508 19446 -4444
rect 19380 -4509 19446 -4508
rect 19541 -4687 19601 1343
rect 19538 -4688 19604 -4687
rect 19538 -4752 19539 -4688
rect 19603 -4752 19604 -4688
rect 19538 -4753 19604 -4752
rect 19602 -4932 19668 -4931
rect 19602 -4996 19603 -4932
rect 19667 -4996 19668 -4932
rect 19602 -4997 19668 -4996
rect 19605 -18288 19665 -4997
rect 19949 -11276 20015 -11275
rect 19949 -11340 19950 -11276
rect 20014 -11340 20015 -11276
rect 19949 -11341 20015 -11340
rect 19602 -18289 19668 -18288
rect 19602 -18353 19603 -18289
rect 19667 -18353 19668 -18289
rect 19602 -18354 19668 -18353
rect 19952 -18982 20012 -11341
rect 20631 -11519 20691 3602
rect 20786 1408 20852 1409
rect 20786 1344 20787 1408
rect 20851 1344 20852 1408
rect 20786 1343 20852 1344
rect 20628 -11520 20694 -11519
rect 20628 -11584 20629 -11520
rect 20693 -11584 20694 -11520
rect 20628 -11585 20694 -11584
rect 20789 -11763 20849 1343
rect 21117 -1028 21183 -1027
rect 21117 -1092 21118 -1028
rect 21182 -1092 21183 -1028
rect 21117 -1093 21183 -1092
rect 20786 -11764 20852 -11763
rect 20786 -11828 20787 -11764
rect 20851 -11828 20852 -11764
rect 20786 -11829 20852 -11828
rect 20770 -12008 20836 -12007
rect 20770 -12072 20771 -12008
rect 20835 -12072 20836 -12008
rect 20770 -12073 20836 -12072
rect 20773 -18288 20833 -12073
rect 20770 -18289 20836 -18288
rect 20770 -18353 20771 -18289
rect 20835 -18353 20836 -18289
rect 20770 -18354 20836 -18353
rect 21120 -18982 21180 -1093
rect 21879 -1271 21939 3602
rect 22034 1408 22100 1409
rect 22034 1344 22035 1408
rect 22099 1344 22100 1408
rect 22034 1343 22100 1344
rect 21876 -1272 21942 -1271
rect 21876 -1336 21877 -1272
rect 21941 -1336 21942 -1272
rect 21876 -1337 21942 -1336
rect 22037 -1515 22097 1343
rect 22997 288 23063 289
rect 22997 224 22998 288
rect 23062 224 23063 288
rect 22997 223 23063 224
rect 22034 -1516 22100 -1515
rect 22034 -1580 22035 -1516
rect 22099 -1580 22100 -1516
rect 22034 -1581 22100 -1580
rect 21938 -1760 22004 -1759
rect 21938 -1824 21939 -1760
rect 22003 -1824 22004 -1760
rect 21938 -1825 22004 -1824
rect 21941 -18288 22001 -1825
rect 22285 -10300 22351 -10299
rect 22285 -10364 22286 -10300
rect 22350 -10364 22351 -10300
rect 22285 -10365 22351 -10364
rect 21938 -18289 22004 -18288
rect 21938 -18353 21939 -18289
rect 22003 -18353 22004 -18289
rect 21938 -18354 22004 -18353
rect 22288 -18982 22348 -10365
rect 23000 -10543 23060 223
rect 23127 -8835 23187 3602
rect 23282 1408 23348 1409
rect 23282 1344 23283 1408
rect 23347 1344 23348 1408
rect 23282 1343 23348 1344
rect 23124 -8836 23190 -8835
rect 23124 -8900 23125 -8836
rect 23189 -8900 23190 -8836
rect 23124 -8901 23190 -8900
rect 23285 -9567 23345 1343
rect 24375 -7371 24435 3602
rect 24530 1408 24596 1409
rect 24530 1344 24531 1408
rect 24595 1344 24596 1408
rect 24530 1343 24596 1344
rect 24372 -7372 24438 -7371
rect 24372 -7436 24373 -7372
rect 24437 -7436 24438 -7372
rect 24372 -7437 24438 -7436
rect 24533 -8103 24593 1343
rect 25623 -3711 25683 3602
rect 25778 1408 25844 1409
rect 25778 1344 25779 1408
rect 25843 1344 25844 1408
rect 25778 1343 25844 1344
rect 25620 -3712 25686 -3711
rect 25620 -3776 25621 -3712
rect 25685 -3776 25686 -3712
rect 25620 -3777 25686 -3776
rect 25781 -4931 25841 1343
rect 25778 -4932 25844 -4931
rect 25778 -4996 25779 -4932
rect 25843 -4996 25844 -4932
rect 25778 -4997 25844 -4996
rect 25789 -5176 25855 -5175
rect 25789 -5240 25790 -5176
rect 25854 -5240 25855 -5176
rect 25789 -5241 25855 -5240
rect 24530 -8104 24596 -8103
rect 24530 -8168 24531 -8104
rect 24595 -8168 24596 -8104
rect 24530 -8169 24596 -8168
rect 24621 -8348 24687 -8347
rect 24621 -8412 24622 -8348
rect 24686 -8412 24687 -8348
rect 24621 -8413 24687 -8412
rect 23282 -9568 23348 -9567
rect 23282 -9632 23283 -9568
rect 23347 -9632 23348 -9568
rect 23282 -9633 23348 -9632
rect 23453 -9812 23519 -9811
rect 23453 -9876 23454 -9812
rect 23518 -9876 23519 -9812
rect 23453 -9877 23519 -9876
rect 22997 -10544 23063 -10543
rect 22997 -10608 22998 -10544
rect 23062 -10608 23063 -10544
rect 22997 -10609 23063 -10608
rect 23106 -10788 23172 -10787
rect 23106 -10852 23107 -10788
rect 23171 -10852 23172 -10788
rect 23106 -10853 23172 -10852
rect 23109 -18288 23169 -10853
rect 23106 -18289 23172 -18288
rect 23106 -18353 23107 -18289
rect 23171 -18353 23172 -18289
rect 23106 -18354 23172 -18353
rect 23456 -18982 23516 -9877
rect 24274 -16400 24340 -16399
rect 24274 -16464 24275 -16400
rect 24339 -16464 24340 -16400
rect 24274 -16465 24340 -16464
rect 24277 -18288 24337 -16465
rect 24274 -18289 24340 -18288
rect 24274 -18353 24275 -18289
rect 24339 -18353 24340 -18289
rect 24274 -18354 24340 -18353
rect 24624 -18982 24684 -8413
rect 25442 -16156 25508 -16155
rect 25442 -16220 25443 -16156
rect 25507 -16220 25508 -16156
rect 25442 -16221 25508 -16220
rect 25445 -18288 25505 -16221
rect 25442 -18289 25508 -18288
rect 25442 -18353 25443 -18289
rect 25507 -18353 25508 -18289
rect 25442 -18354 25508 -18353
rect 25792 -18982 25852 -5241
rect 26871 -11275 26931 3602
rect 27026 1408 27092 1409
rect 27026 1344 27027 1408
rect 27091 1344 27092 1408
rect 27026 1343 27092 1344
rect 26868 -11276 26934 -11275
rect 26868 -11340 26869 -11276
rect 26933 -11340 26934 -11276
rect 26868 -11341 26934 -11340
rect 27029 -12007 27089 1343
rect 28119 -1027 28179 3602
rect 28274 1408 28340 1409
rect 28274 1344 28275 1408
rect 28339 1344 28340 1408
rect 28274 1343 28340 1344
rect 28116 -1028 28182 -1027
rect 28116 -1092 28117 -1028
rect 28181 -1092 28182 -1028
rect 28116 -1093 28182 -1092
rect 28277 -1759 28337 1343
rect 28274 -1760 28340 -1759
rect 28274 -1824 28275 -1760
rect 28339 -1824 28340 -1760
rect 28274 -1825 28340 -1824
rect 28125 -2004 28191 -2003
rect 28125 -2068 28126 -2004
rect 28190 -2068 28191 -2004
rect 28125 -2069 28191 -2068
rect 27026 -12008 27092 -12007
rect 27026 -12072 27027 -12008
rect 27091 -12072 27092 -12008
rect 27026 -12073 27092 -12072
rect 26957 -12252 27023 -12251
rect 26957 -12316 26958 -12252
rect 27022 -12316 27023 -12252
rect 26957 -12317 27023 -12316
rect 26610 -15912 26676 -15911
rect 26610 -15976 26611 -15912
rect 26675 -15976 26676 -15912
rect 26610 -15977 26676 -15976
rect 26613 -18288 26673 -15977
rect 26610 -18289 26676 -18288
rect 26610 -18353 26611 -18289
rect 26675 -18353 26676 -18289
rect 26610 -18354 26676 -18353
rect 26960 -18982 27020 -12317
rect 27778 -15668 27844 -15667
rect 27778 -15732 27779 -15668
rect 27843 -15732 27844 -15668
rect 27778 -15733 27844 -15732
rect 27781 -18288 27841 -15733
rect 27778 -18289 27844 -18288
rect 27778 -18353 27779 -18289
rect 27843 -18353 27844 -18289
rect 27778 -18354 27844 -18353
rect 28128 -18982 28188 -2069
rect 28946 -2248 29012 -2247
rect 28946 -2312 28947 -2248
rect 29011 -2312 29012 -2248
rect 28946 -2313 29012 -2312
rect 28949 -18288 29009 -2313
rect 29367 -10299 29427 3602
rect 29522 1408 29588 1409
rect 29522 1344 29523 1408
rect 29587 1344 29588 1408
rect 29522 1343 29588 1344
rect 29364 -10300 29430 -10299
rect 29364 -10364 29365 -10300
rect 29429 -10364 29430 -10300
rect 29364 -10365 29430 -10364
rect 29525 -10787 29585 1343
rect 30615 -9811 30675 3602
rect 30770 1408 30836 1409
rect 30770 1344 30771 1408
rect 30835 1344 30836 1408
rect 30770 1343 30836 1344
rect 30612 -9812 30678 -9811
rect 30612 -9876 30613 -9812
rect 30677 -9876 30678 -9812
rect 30612 -9877 30678 -9876
rect 30461 -10056 30527 -10055
rect 30461 -10120 30462 -10056
rect 30526 -10120 30527 -10056
rect 30461 -10121 30527 -10120
rect 29522 -10788 29588 -10787
rect 29522 -10852 29523 -10788
rect 29587 -10852 29588 -10788
rect 29522 -10853 29588 -10852
rect 29293 -11032 29359 -11031
rect 29293 -11096 29294 -11032
rect 29358 -11096 29359 -11032
rect 29293 -11097 29359 -11096
rect 28946 -18289 29012 -18288
rect 28946 -18353 28947 -18289
rect 29011 -18353 29012 -18289
rect 28946 -18354 29012 -18353
rect 29296 -18982 29356 -11097
rect 30114 -15180 30180 -15179
rect 30114 -15244 30115 -15180
rect 30179 -15244 30180 -15180
rect 30114 -15245 30180 -15244
rect 30117 -18288 30177 -15245
rect 30114 -18289 30180 -18288
rect 30114 -18353 30115 -18289
rect 30179 -18353 30180 -18289
rect 30114 -18354 30180 -18353
rect 30464 -18982 30524 -10121
rect 30773 -16399 30833 1343
rect 31863 -8347 31923 3602
rect 32018 1408 32084 1409
rect 32018 1344 32019 1408
rect 32083 1344 32084 1408
rect 32018 1343 32084 1344
rect 31860 -8348 31926 -8347
rect 31860 -8412 31861 -8348
rect 31925 -8412 31926 -8348
rect 31860 -8413 31926 -8412
rect 31629 -8592 31695 -8591
rect 31629 -8656 31630 -8592
rect 31694 -8656 31695 -8592
rect 31629 -8657 31695 -8656
rect 31282 -14692 31348 -14691
rect 31282 -14756 31283 -14692
rect 31347 -14756 31348 -14692
rect 31282 -14757 31348 -14756
rect 30770 -16400 30836 -16399
rect 30770 -16464 30771 -16400
rect 30835 -16464 30836 -16400
rect 30770 -16465 30836 -16464
rect 31285 -18288 31345 -14757
rect 31282 -18289 31348 -18288
rect 31282 -18353 31283 -18289
rect 31347 -18353 31348 -18289
rect 31282 -18354 31348 -18353
rect 31632 -18982 31692 -8657
rect 32021 -16155 32081 1343
rect 32981 288 33047 289
rect 32981 224 32982 288
rect 33046 224 33047 288
rect 32981 223 33047 224
rect 32984 -5419 33044 223
rect 33111 -5175 33171 3602
rect 33266 1408 33332 1409
rect 33266 1344 33267 1408
rect 33331 1344 33332 1408
rect 33266 1343 33332 1344
rect 33108 -5176 33174 -5175
rect 33108 -5240 33109 -5176
rect 33173 -5240 33174 -5176
rect 33108 -5241 33174 -5240
rect 32981 -5420 33047 -5419
rect 32981 -5484 32982 -5420
rect 33046 -5484 33047 -5420
rect 32981 -5485 33047 -5484
rect 32797 -5664 32863 -5663
rect 32797 -5728 32798 -5664
rect 32862 -5728 32863 -5664
rect 32797 -5729 32863 -5728
rect 32450 -14204 32516 -14203
rect 32450 -14268 32451 -14204
rect 32515 -14268 32516 -14204
rect 32450 -14269 32516 -14268
rect 32018 -16156 32084 -16155
rect 32018 -16220 32019 -16156
rect 32083 -16220 32084 -16156
rect 32018 -16221 32084 -16220
rect 32453 -18288 32513 -14269
rect 32450 -18289 32516 -18288
rect 32450 -18353 32451 -18289
rect 32515 -18353 32516 -18289
rect 32450 -18354 32516 -18353
rect 32800 -18982 32860 -5729
rect 33269 -15911 33329 1343
rect 33965 -2980 34031 -2979
rect 33965 -3044 33966 -2980
rect 34030 -3044 34031 -2980
rect 33965 -3045 34031 -3044
rect 33618 -5908 33684 -5907
rect 33618 -5972 33619 -5908
rect 33683 -5972 33684 -5908
rect 33618 -5973 33684 -5972
rect 33266 -15912 33332 -15911
rect 33266 -15976 33267 -15912
rect 33331 -15976 33332 -15912
rect 33266 -15977 33332 -15976
rect 33621 -18288 33681 -5973
rect 33618 -18289 33684 -18288
rect 33618 -18353 33619 -18289
rect 33683 -18353 33684 -18289
rect 33618 -18354 33684 -18353
rect 33968 -18982 34028 -3045
rect 34359 -12251 34419 3602
rect 34514 1408 34580 1409
rect 34514 1344 34515 1408
rect 34579 1344 34580 1408
rect 34514 1343 34580 1344
rect 34356 -12252 34422 -12251
rect 34356 -12316 34357 -12252
rect 34421 -12316 34422 -12252
rect 34356 -12317 34422 -12316
rect 34517 -15667 34577 1343
rect 35133 -784 35199 -783
rect 35133 -848 35134 -784
rect 35198 -848 35199 -784
rect 35133 -849 35199 -848
rect 34786 -3224 34852 -3223
rect 34786 -3288 34787 -3224
rect 34851 -3288 34852 -3224
rect 34786 -3289 34852 -3288
rect 34514 -15668 34580 -15667
rect 34514 -15732 34515 -15668
rect 34579 -15732 34580 -15668
rect 34514 -15733 34580 -15732
rect 34789 -18288 34849 -3289
rect 34786 -18289 34852 -18288
rect 34786 -18353 34787 -18289
rect 34851 -18353 34852 -18289
rect 34786 -18354 34852 -18353
rect 35136 -18982 35196 -849
rect 35607 -2003 35667 3602
rect 35762 1408 35828 1409
rect 35762 1344 35763 1408
rect 35827 1344 35828 1408
rect 35762 1343 35828 1344
rect 35604 -2004 35670 -2003
rect 35604 -2068 35605 -2004
rect 35669 -2068 35670 -2004
rect 35604 -2069 35670 -2068
rect 35765 -2247 35825 1343
rect 35762 -2248 35828 -2247
rect 35762 -2312 35763 -2248
rect 35827 -2312 35828 -2248
rect 35762 -2313 35828 -2312
rect 35954 -2492 36020 -2491
rect 35954 -2556 35955 -2492
rect 36019 -2556 36020 -2492
rect 35954 -2557 36020 -2556
rect 35957 -18288 36017 -2557
rect 36301 -7128 36367 -7127
rect 36301 -7192 36302 -7128
rect 36366 -7192 36367 -7128
rect 36301 -7193 36367 -7192
rect 35954 -18289 36020 -18288
rect 35954 -18353 35955 -18289
rect 36019 -18353 36020 -18289
rect 35954 -18354 36020 -18353
rect 36304 -18982 36364 -7193
rect 36855 -11031 36915 3602
rect 37010 1408 37076 1409
rect 37010 1344 37011 1408
rect 37075 1344 37076 1408
rect 37010 1343 37076 1344
rect 36852 -11032 36918 -11031
rect 36852 -11096 36853 -11032
rect 36917 -11096 36918 -11032
rect 36852 -11097 36918 -11096
rect 37013 -15179 37073 1343
rect 37469 -6884 37535 -6883
rect 37469 -6948 37470 -6884
rect 37534 -6948 37535 -6884
rect 37469 -6949 37535 -6948
rect 37010 -15180 37076 -15179
rect 37010 -15244 37011 -15180
rect 37075 -15244 37076 -15180
rect 37010 -15245 37076 -15244
rect 37122 -15424 37188 -15423
rect 37122 -15488 37123 -15424
rect 37187 -15488 37188 -15424
rect 37122 -15489 37188 -15488
rect 37125 -18288 37185 -15489
rect 37122 -18289 37188 -18288
rect 37122 -18353 37123 -18289
rect 37187 -18353 37188 -18289
rect 37122 -18354 37188 -18353
rect 37472 -18982 37532 -6949
rect 38103 -10055 38163 3602
rect 38258 1408 38324 1409
rect 38258 1344 38259 1408
rect 38323 1344 38324 1408
rect 38258 1343 38324 1344
rect 38100 -10056 38166 -10055
rect 38100 -10120 38101 -10056
rect 38165 -10120 38166 -10056
rect 38100 -10121 38166 -10120
rect 38261 -14691 38321 1343
rect 38637 -6640 38703 -6639
rect 38637 -6704 38638 -6640
rect 38702 -6704 38703 -6640
rect 38637 -6705 38703 -6704
rect 38258 -14692 38324 -14691
rect 38258 -14756 38259 -14692
rect 38323 -14756 38324 -14692
rect 38258 -14757 38324 -14756
rect 38290 -14936 38356 -14935
rect 38290 -15000 38291 -14936
rect 38355 -15000 38356 -14936
rect 38290 -15001 38356 -15000
rect 38293 -18288 38353 -15001
rect 38290 -18289 38356 -18288
rect 38290 -18353 38291 -18289
rect 38355 -18353 38356 -18289
rect 38290 -18354 38356 -18353
rect 38640 -18982 38700 -6705
rect 39351 -8591 39411 3602
rect 39506 1408 39572 1409
rect 39506 1344 39507 1408
rect 39571 1344 39572 1408
rect 39506 1343 39572 1344
rect 39348 -8592 39414 -8591
rect 39348 -8656 39349 -8592
rect 39413 -8656 39414 -8592
rect 39348 -8657 39414 -8656
rect 39509 -14203 39569 1343
rect 40599 -5663 40659 3602
rect 40754 1408 40820 1409
rect 40754 1344 40755 1408
rect 40819 1344 40820 1408
rect 40754 1343 40820 1344
rect 40596 -5664 40662 -5663
rect 40596 -5728 40597 -5664
rect 40661 -5728 40662 -5664
rect 40596 -5729 40662 -5728
rect 40757 -5907 40817 1343
rect 41847 -2979 41907 3602
rect 42002 1408 42068 1409
rect 42002 1344 42003 1408
rect 42067 1344 42068 1408
rect 42002 1343 42068 1344
rect 41844 -2980 41910 -2979
rect 41844 -3044 41845 -2980
rect 41909 -3044 41910 -2980
rect 41844 -3045 41910 -3044
rect 42005 -3223 42065 1343
rect 42965 288 43031 289
rect 42965 224 42966 288
rect 43030 224 43031 288
rect 42965 223 43031 224
rect 42002 -3224 42068 -3223
rect 42002 -3288 42003 -3224
rect 42067 -3288 42068 -3224
rect 42002 -3289 42068 -3288
rect 42141 -3468 42207 -3467
rect 42141 -3532 42142 -3468
rect 42206 -3532 42207 -3468
rect 42141 -3533 42207 -3532
rect 40754 -5908 40820 -5907
rect 40754 -5972 40755 -5908
rect 40819 -5972 40820 -5908
rect 40754 -5973 40820 -5972
rect 40973 -6152 41039 -6151
rect 40973 -6216 40974 -6152
rect 41038 -6216 41039 -6152
rect 40973 -6217 41039 -6216
rect 39805 -6396 39871 -6395
rect 39805 -6460 39806 -6396
rect 39870 -6460 39871 -6396
rect 39805 -6461 39871 -6460
rect 39506 -14204 39572 -14203
rect 39506 -14268 39507 -14204
rect 39571 -14268 39572 -14204
rect 39506 -14269 39572 -14268
rect 39458 -14448 39524 -14447
rect 39458 -14512 39459 -14448
rect 39523 -14512 39524 -14448
rect 39458 -14513 39524 -14512
rect 39461 -18288 39521 -14513
rect 39458 -18289 39524 -18288
rect 39458 -18353 39459 -18289
rect 39523 -18353 39524 -18289
rect 39458 -18354 39524 -18353
rect 39808 -18982 39868 -6461
rect 40626 -13960 40692 -13959
rect 40626 -14024 40627 -13960
rect 40691 -14024 40692 -13960
rect 40626 -14025 40692 -14024
rect 40629 -18288 40689 -14025
rect 40626 -18289 40692 -18288
rect 40626 -18353 40627 -18289
rect 40691 -18353 40692 -18289
rect 40626 -18354 40692 -18353
rect 40976 -18982 41036 -6217
rect 41794 -13716 41860 -13715
rect 41794 -13780 41795 -13716
rect 41859 -13780 41860 -13716
rect 41794 -13781 41860 -13780
rect 41797 -18288 41857 -13781
rect 41794 -18289 41860 -18288
rect 41794 -18353 41795 -18289
rect 41859 -18353 41860 -18289
rect 41794 -18354 41860 -18353
rect 42144 -18982 42204 -3533
rect 42968 -13227 43028 223
rect 43095 -783 43155 3602
rect 43250 1408 43316 1409
rect 43250 1344 43251 1408
rect 43315 1344 43316 1408
rect 43250 1343 43316 1344
rect 43092 -784 43158 -783
rect 43092 -848 43093 -784
rect 43157 -848 43158 -784
rect 43092 -849 43158 -848
rect 43253 -2491 43313 1343
rect 43250 -2492 43316 -2491
rect 43250 -2556 43251 -2492
rect 43315 -2556 43316 -2492
rect 43250 -2557 43316 -2556
rect 43309 -2736 43375 -2735
rect 43309 -2800 43310 -2736
rect 43374 -2800 43375 -2736
rect 43309 -2801 43375 -2800
rect 42965 -13228 43031 -13227
rect 42965 -13292 42966 -13228
rect 43030 -13292 43031 -13228
rect 42965 -13293 43031 -13292
rect 42962 -13472 43028 -13471
rect 42962 -13536 42963 -13472
rect 43027 -13536 43028 -13472
rect 42962 -13537 43028 -13536
rect 42965 -18288 43025 -13537
rect 42962 -18289 43028 -18288
rect 42962 -18353 42963 -18289
rect 43027 -18353 43028 -18289
rect 42962 -18354 43028 -18353
rect 43312 -18982 43372 -2801
rect 44343 -7127 44403 3602
rect 44498 1408 44564 1409
rect 44498 1344 44499 1408
rect 44563 1344 44564 1408
rect 44498 1343 44564 1344
rect 44340 -7128 44406 -7127
rect 44340 -7192 44341 -7128
rect 44405 -7192 44406 -7128
rect 44340 -7193 44406 -7192
rect 44130 -12984 44196 -12983
rect 44130 -13048 44131 -12984
rect 44195 -13048 44196 -12984
rect 44130 -13049 44196 -13048
rect 44133 -18288 44193 -13049
rect 44501 -15423 44561 1343
rect 45591 -6883 45651 3602
rect 45746 1408 45812 1409
rect 45746 1344 45747 1408
rect 45811 1344 45812 1408
rect 45746 1343 45812 1344
rect 45588 -6884 45654 -6883
rect 45588 -6948 45589 -6884
rect 45653 -6948 45654 -6884
rect 45588 -6949 45654 -6948
rect 45749 -14935 45809 1343
rect 46839 -6639 46899 3602
rect 46994 1408 47060 1409
rect 46994 1344 46995 1408
rect 47059 1344 47060 1408
rect 46994 1343 47060 1344
rect 46836 -6640 46902 -6639
rect 46836 -6704 46837 -6640
rect 46901 -6704 46902 -6640
rect 46836 -6705 46902 -6704
rect 46997 -14447 47057 1343
rect 48087 -6395 48147 3602
rect 48242 1408 48308 1409
rect 48242 1344 48243 1408
rect 48307 1344 48308 1408
rect 48242 1343 48308 1344
rect 48084 -6396 48150 -6395
rect 48084 -6460 48085 -6396
rect 48149 -6460 48150 -6396
rect 48084 -6461 48150 -6460
rect 48245 -13959 48305 1343
rect 49335 -6151 49395 3602
rect 49490 1408 49556 1409
rect 49490 1344 49491 1408
rect 49555 1344 49556 1408
rect 49490 1343 49556 1344
rect 49332 -6152 49398 -6151
rect 49332 -6216 49333 -6152
rect 49397 -6216 49398 -6152
rect 49332 -6217 49398 -6216
rect 49493 -13715 49553 1343
rect 50583 -3467 50643 3602
rect 50738 1408 50804 1409
rect 50738 1344 50739 1408
rect 50803 1344 50804 1408
rect 50738 1343 50804 1344
rect 50580 -3468 50646 -3467
rect 50580 -3532 50581 -3468
rect 50645 -3532 50646 -3468
rect 50580 -3533 50646 -3532
rect 50741 -13471 50801 1343
rect 51831 -2735 51891 3602
rect 51986 1408 52052 1409
rect 51986 1344 51987 1408
rect 52051 1344 52052 1408
rect 51986 1343 52052 1344
rect 51828 -2736 51894 -2735
rect 51828 -2800 51829 -2736
rect 51893 -2800 51894 -2736
rect 51828 -2801 51894 -2800
rect 51989 -12983 52049 1343
rect 51986 -12984 52052 -12983
rect 51986 -13048 51987 -12984
rect 52051 -13048 52052 -12984
rect 51986 -13049 52052 -13048
rect 50738 -13472 50804 -13471
rect 50738 -13536 50739 -13472
rect 50803 -13536 50804 -13472
rect 50738 -13537 50804 -13536
rect 49490 -13716 49556 -13715
rect 49490 -13780 49491 -13716
rect 49555 -13780 49556 -13716
rect 49490 -13781 49556 -13780
rect 48242 -13960 48308 -13959
rect 48242 -14024 48243 -13960
rect 48307 -14024 48308 -13960
rect 48242 -14025 48308 -14024
rect 46994 -14448 47060 -14447
rect 46994 -14512 46995 -14448
rect 47059 -14512 47060 -14448
rect 46994 -14513 47060 -14512
rect 45746 -14936 45812 -14935
rect 45746 -15000 45747 -14936
rect 45811 -15000 45812 -14936
rect 45746 -15001 45812 -15000
rect 44498 -15424 44564 -15423
rect 44498 -15488 44499 -15424
rect 44563 -15488 44564 -15424
rect 44498 -15489 44564 -15488
rect 44130 -18289 44196 -18288
rect 44130 -18353 44131 -18289
rect 44195 -18353 44196 -18289
rect 44130 -18354 44196 -18353
use contact_7  contact_7_0
timestamp 1644511149
transform 1 0 5988 0 1 5408
box 0 0 1 1
use contact_8  contact_8_0
timestamp 1644511149
transform 1 0 17043 0 1 1344
box 0 0 1 1
use contact_8  contact_8_1
timestamp 1644511149
transform 1 0 23283 0 1 1344
box 0 0 1 1
use contact_8  contact_8_2
timestamp 1644511149
transform 1 0 14547 0 1 1344
box 0 0 1 1
use contact_8  contact_8_3
timestamp 1644511149
transform 1 0 21877 0 1 3603
box 0 0 1 1
use contact_8  contact_8_4
timestamp 1644511149
transform 1 0 22035 0 1 1344
box 0 0 1 1
use contact_8  contact_8_5
timestamp 1644511149
transform 1 0 15637 0 1 3603
box 0 0 1 1
use contact_8  contact_8_6
timestamp 1644511149
transform 1 0 14389 0 1 3603
box 0 0 1 1
use contact_8  contact_8_7
timestamp 1644511149
transform 1 0 13299 0 1 1344
box 0 0 1 1
use contact_8  contact_8_8
timestamp 1644511149
transform 1 0 5985 0 1 5409
box 0 0 1 1
use contact_8  contact_8_9
timestamp 1644511149
transform 1 0 26869 0 1 3603
box 0 0 1 1
use contact_8  contact_8_10
timestamp 1644511149
transform 1 0 20629 0 1 3603
box 0 0 1 1
use contact_8  contact_8_11
timestamp 1644511149
transform 1 0 24373 0 1 3603
box 0 0 1 1
use contact_8  contact_8_12
timestamp 1644511149
transform 1 0 18133 0 1 3603
box 0 0 1 1
use contact_8  contact_8_13
timestamp 1644511149
transform 1 0 18291 0 1 1344
box 0 0 1 1
use contact_8  contact_8_14
timestamp 1644511149
transform 1 0 24531 0 1 1344
box 0 0 1 1
use contact_8  contact_8_15
timestamp 1644511149
transform 1 0 20787 0 1 1344
box 0 0 1 1
use contact_8  contact_8_16
timestamp 1644511149
transform 1 0 15795 0 1 1344
box 0 0 1 1
use contact_8  contact_8_17
timestamp 1644511149
transform 1 0 25621 0 1 3603
box 0 0 1 1
use contact_8  contact_8_18
timestamp 1644511149
transform 1 0 13141 0 1 3603
box 0 0 1 1
use contact_8  contact_8_19
timestamp 1644511149
transform 1 0 19381 0 1 3603
box 0 0 1 1
use contact_8  contact_8_20
timestamp 1644511149
transform 1 0 19539 0 1 1344
box 0 0 1 1
use contact_8  contact_8_21
timestamp 1644511149
transform 1 0 25779 0 1 1344
box 0 0 1 1
use contact_8  contact_8_22
timestamp 1644511149
transform 1 0 23125 0 1 3603
box 0 0 1 1
use contact_8  contact_8_23
timestamp 1644511149
transform 1 0 16885 0 1 3603
box 0 0 1 1
use contact_8  contact_8_24
timestamp 1644511149
transform 1 0 31861 0 1 3603
box 0 0 1 1
use contact_8  contact_8_25
timestamp 1644511149
transform 1 0 28117 0 1 3603
box 0 0 1 1
use contact_8  contact_8_26
timestamp 1644511149
transform 1 0 28275 0 1 1344
box 0 0 1 1
use contact_8  contact_8_27
timestamp 1644511149
transform 1 0 35605 0 1 3603
box 0 0 1 1
use contact_8  contact_8_28
timestamp 1644511149
transform 1 0 35763 0 1 1344
box 0 0 1 1
use contact_8  contact_8_29
timestamp 1644511149
transform 1 0 39349 0 1 3603
box 0 0 1 1
use contact_8  contact_8_30
timestamp 1644511149
transform 1 0 30613 0 1 3603
box 0 0 1 1
use contact_8  contact_8_31
timestamp 1644511149
transform 1 0 38101 0 1 3603
box 0 0 1 1
use contact_8  contact_8_32
timestamp 1644511149
transform 1 0 29365 0 1 3603
box 0 0 1 1
use contact_8  contact_8_33
timestamp 1644511149
transform 1 0 29523 0 1 1344
box 0 0 1 1
use contact_8  contact_8_34
timestamp 1644511149
transform 1 0 33109 0 1 3603
box 0 0 1 1
use contact_8  contact_8_35
timestamp 1644511149
transform 1 0 36853 0 1 3603
box 0 0 1 1
use contact_8  contact_8_36
timestamp 1644511149
transform 1 0 32019 0 1 1344
box 0 0 1 1
use contact_8  contact_8_37
timestamp 1644511149
transform 1 0 30771 0 1 1344
box 0 0 1 1
use contact_8  contact_8_38
timestamp 1644511149
transform 1 0 34357 0 1 3603
box 0 0 1 1
use contact_8  contact_8_39
timestamp 1644511149
transform 1 0 34515 0 1 1344
box 0 0 1 1
use contact_8  contact_8_40
timestamp 1644511149
transform 1 0 37011 0 1 1344
box 0 0 1 1
use contact_8  contact_8_41
timestamp 1644511149
transform 1 0 33267 0 1 1344
box 0 0 1 1
use contact_8  contact_8_42
timestamp 1644511149
transform 1 0 38259 0 1 1344
box 0 0 1 1
use contact_8  contact_8_43
timestamp 1644511149
transform 1 0 43093 0 1 3603
box 0 0 1 1
use contact_8  contact_8_44
timestamp 1644511149
transform 1 0 43251 0 1 1344
box 0 0 1 1
use contact_8  contact_8_45
timestamp 1644511149
transform 1 0 51829 0 1 3603
box 0 0 1 1
use contact_8  contact_8_46
timestamp 1644511149
transform 1 0 41845 0 1 3603
box 0 0 1 1
use contact_8  contact_8_47
timestamp 1644511149
transform 1 0 42003 0 1 1344
box 0 0 1 1
use contact_8  contact_8_48
timestamp 1644511149
transform 1 0 50581 0 1 3603
box 0 0 1 1
use contact_8  contact_8_49
timestamp 1644511149
transform 1 0 40597 0 1 3603
box 0 0 1 1
use contact_8  contact_8_50
timestamp 1644511149
transform 1 0 40755 0 1 1344
box 0 0 1 1
use contact_8  contact_8_51
timestamp 1644511149
transform 1 0 49333 0 1 3603
box 0 0 1 1
use contact_8  contact_8_52
timestamp 1644511149
transform 1 0 48085 0 1 3603
box 0 0 1 1
use contact_8  contact_8_53
timestamp 1644511149
transform 1 0 46837 0 1 3603
box 0 0 1 1
use contact_8  contact_8_54
timestamp 1644511149
transform 1 0 45589 0 1 3603
box 0 0 1 1
use contact_8  contact_8_55
timestamp 1644511149
transform 1 0 44341 0 1 3603
box 0 0 1 1
use contact_8  contact_8_56
timestamp 1644511149
transform 1 0 51987 0 1 1344
box 0 0 1 1
use contact_8  contact_8_57
timestamp 1644511149
transform 1 0 50739 0 1 1344
box 0 0 1 1
use contact_8  contact_8_58
timestamp 1644511149
transform 1 0 49491 0 1 1344
box 0 0 1 1
use contact_8  contact_8_59
timestamp 1644511149
transform 1 0 48243 0 1 1344
box 0 0 1 1
use contact_8  contact_8_60
timestamp 1644511149
transform 1 0 44499 0 1 1344
box 0 0 1 1
use contact_8  contact_8_61
timestamp 1644511149
transform 1 0 46995 0 1 1344
box 0 0 1 1
use contact_8  contact_8_62
timestamp 1644511149
transform 1 0 45747 0 1 1344
box 0 0 1 1
use contact_8  contact_8_63
timestamp 1644511149
transform 1 0 39507 0 1 1344
box 0 0 1 1
use contact_8  contact_8_64
timestamp 1644511149
transform 1 0 27027 0 1 1344
box 0 0 1 1
use contact_9  contact_9_0
timestamp 1644511149
transform 1 0 40626 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_1
timestamp 1644511149
transform 1 0 30114 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_2
timestamp 1644511149
transform 1 0 32450 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_3
timestamp 1644511149
transform 1 0 27778 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_4
timestamp 1644511149
transform 1 0 39458 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_5
timestamp 1644511149
transform 1 0 37122 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_6
timestamp 1644511149
transform 1 0 44130 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_7
timestamp 1644511149
transform 1 0 28946 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_8
timestamp 1644511149
transform 1 0 31282 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_9
timestamp 1644511149
transform 1 0 35954 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_10
timestamp 1644511149
transform 1 0 33618 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_11
timestamp 1644511149
transform 1 0 34786 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_12
timestamp 1644511149
transform 1 0 42962 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_13
timestamp 1644511149
transform 1 0 38290 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_14
timestamp 1644511149
transform 1 0 41794 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_15
timestamp 1644511149
transform 1 0 19602 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_16
timestamp 1644511149
transform 1 0 20770 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_17
timestamp 1644511149
transform 1 0 11426 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_18
timestamp 1644511149
transform 1 0 16098 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_19
timestamp 1644511149
transform 1 0 5586 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_20
timestamp 1644511149
transform 1 0 9090 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_21
timestamp 1644511149
transform 1 0 21938 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_22
timestamp 1644511149
transform 1 0 17266 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_23
timestamp 1644511149
transform 1 0 25442 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_24
timestamp 1644511149
transform 1 0 24274 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_25
timestamp 1644511149
transform 1 0 4418 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_26
timestamp 1644511149
transform 1 0 23106 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_27
timestamp 1644511149
transform 1 0 7922 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_28
timestamp 1644511149
transform 1 0 6754 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_29
timestamp 1644511149
transform 1 0 10258 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_30
timestamp 1644511149
transform 1 0 12594 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_31
timestamp 1644511149
transform 1 0 18434 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_32
timestamp 1644511149
transform 1 0 3250 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_33
timestamp 1644511149
transform 1 0 2082 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_34
timestamp 1644511149
transform 1 0 14930 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_35
timestamp 1644511149
transform 1 0 13762 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_36
timestamp 1644511149
transform 1 0 26610 0 1 -18358
box 0 0 1 1
use contact_9  contact_9_37
timestamp 1644511149
transform 1 0 17042 0 1 1339
box 0 0 1 1
use contact_9  contact_9_38
timestamp 1644511149
transform 1 0 23282 0 1 1339
box 0 0 1 1
use contact_9  contact_9_39
timestamp 1644511149
transform 1 0 13298 0 1 1339
box 0 0 1 1
use contact_9  contact_9_40
timestamp 1644511149
transform 1 0 21876 0 1 3598
box 0 0 1 1
use contact_9  contact_9_41
timestamp 1644511149
transform 1 0 22034 0 1 1339
box 0 0 1 1
use contact_9  contact_9_42
timestamp 1644511149
transform 1 0 15636 0 1 3598
box 0 0 1 1
use contact_9  contact_9_43
timestamp 1644511149
transform 1 0 14388 0 1 3598
box 0 0 1 1
use contact_9  contact_9_44
timestamp 1644511149
transform 1 0 22997 0 1 219
box 0 0 1 1
use contact_9  contact_9_45
timestamp 1644511149
transform 1 0 5984 0 1 5404
box 0 0 1 1
use contact_9  contact_9_46
timestamp 1644511149
transform 1 0 26868 0 1 3598
box 0 0 1 1
use contact_9  contact_9_47
timestamp 1644511149
transform 1 0 20628 0 1 3598
box 0 0 1 1
use contact_9  contact_9_48
timestamp 1644511149
transform 1 0 24372 0 1 3598
box 0 0 1 1
use contact_9  contact_9_49
timestamp 1644511149
transform 1 0 18132 0 1 3598
box 0 0 1 1
use contact_9  contact_9_50
timestamp 1644511149
transform 1 0 18290 0 1 1339
box 0 0 1 1
use contact_9  contact_9_51
timestamp 1644511149
transform 1 0 24530 0 1 1339
box 0 0 1 1
use contact_9  contact_9_52
timestamp 1644511149
transform 1 0 20786 0 1 1339
box 0 0 1 1
use contact_9  contact_9_53
timestamp 1644511149
transform 1 0 15794 0 1 1339
box 0 0 1 1
use contact_9  contact_9_54
timestamp 1644511149
transform 1 0 14546 0 1 1339
box 0 0 1 1
use contact_9  contact_9_55
timestamp 1644511149
transform 1 0 25620 0 1 3598
box 0 0 1 1
use contact_9  contact_9_56
timestamp 1644511149
transform 1 0 13140 0 1 3598
box 0 0 1 1
use contact_9  contact_9_57
timestamp 1644511149
transform 1 0 13013 0 1 219
box 0 0 1 1
use contact_9  contact_9_58
timestamp 1644511149
transform 1 0 19380 0 1 3598
box 0 0 1 1
use contact_9  contact_9_59
timestamp 1644511149
transform 1 0 19538 0 1 1339
box 0 0 1 1
use contact_9  contact_9_60
timestamp 1644511149
transform 1 0 25778 0 1 1339
box 0 0 1 1
use contact_9  contact_9_61
timestamp 1644511149
transform 1 0 23124 0 1 3598
box 0 0 1 1
use contact_9  contact_9_62
timestamp 1644511149
transform 1 0 16884 0 1 3598
box 0 0 1 1
use contact_9  contact_9_63
timestamp 1644511149
transform 1 0 31860 0 1 3598
box 0 0 1 1
use contact_9  contact_9_64
timestamp 1644511149
transform 1 0 28116 0 1 3598
box 0 0 1 1
use contact_9  contact_9_65
timestamp 1644511149
transform 1 0 28274 0 1 1339
box 0 0 1 1
use contact_9  contact_9_66
timestamp 1644511149
transform 1 0 35604 0 1 3598
box 0 0 1 1
use contact_9  contact_9_67
timestamp 1644511149
transform 1 0 35762 0 1 1339
box 0 0 1 1
use contact_9  contact_9_68
timestamp 1644511149
transform 1 0 39348 0 1 3598
box 0 0 1 1
use contact_9  contact_9_69
timestamp 1644511149
transform 1 0 30612 0 1 3598
box 0 0 1 1
use contact_9  contact_9_70
timestamp 1644511149
transform 1 0 38100 0 1 3598
box 0 0 1 1
use contact_9  contact_9_71
timestamp 1644511149
transform 1 0 29364 0 1 3598
box 0 0 1 1
use contact_9  contact_9_72
timestamp 1644511149
transform 1 0 29522 0 1 1339
box 0 0 1 1
use contact_9  contact_9_73
timestamp 1644511149
transform 1 0 33108 0 1 3598
box 0 0 1 1
use contact_9  contact_9_74
timestamp 1644511149
transform 1 0 32981 0 1 219
box 0 0 1 1
use contact_9  contact_9_75
timestamp 1644511149
transform 1 0 36852 0 1 3598
box 0 0 1 1
use contact_9  contact_9_76
timestamp 1644511149
transform 1 0 30770 0 1 1339
box 0 0 1 1
use contact_9  contact_9_77
timestamp 1644511149
transform 1 0 34356 0 1 3598
box 0 0 1 1
use contact_9  contact_9_78
timestamp 1644511149
transform 1 0 34514 0 1 1339
box 0 0 1 1
use contact_9  contact_9_79
timestamp 1644511149
transform 1 0 32018 0 1 1339
box 0 0 1 1
use contact_9  contact_9_80
timestamp 1644511149
transform 1 0 37010 0 1 1339
box 0 0 1 1
use contact_9  contact_9_81
timestamp 1644511149
transform 1 0 33266 0 1 1339
box 0 0 1 1
use contact_9  contact_9_82
timestamp 1644511149
transform 1 0 38258 0 1 1339
box 0 0 1 1
use contact_9  contact_9_83
timestamp 1644511149
transform 1 0 43092 0 1 3598
box 0 0 1 1
use contact_9  contact_9_84
timestamp 1644511149
transform 1 0 43250 0 1 1339
box 0 0 1 1
use contact_9  contact_9_85
timestamp 1644511149
transform 1 0 51828 0 1 3598
box 0 0 1 1
use contact_9  contact_9_86
timestamp 1644511149
transform 1 0 41844 0 1 3598
box 0 0 1 1
use contact_9  contact_9_87
timestamp 1644511149
transform 1 0 42002 0 1 1339
box 0 0 1 1
use contact_9  contact_9_88
timestamp 1644511149
transform 1 0 50580 0 1 3598
box 0 0 1 1
use contact_9  contact_9_89
timestamp 1644511149
transform 1 0 40596 0 1 3598
box 0 0 1 1
use contact_9  contact_9_90
timestamp 1644511149
transform 1 0 40754 0 1 1339
box 0 0 1 1
use contact_9  contact_9_91
timestamp 1644511149
transform 1 0 49332 0 1 3598
box 0 0 1 1
use contact_9  contact_9_92
timestamp 1644511149
transform 1 0 48084 0 1 3598
box 0 0 1 1
use contact_9  contact_9_93
timestamp 1644511149
transform 1 0 46836 0 1 3598
box 0 0 1 1
use contact_9  contact_9_94
timestamp 1644511149
transform 1 0 45588 0 1 3598
box 0 0 1 1
use contact_9  contact_9_95
timestamp 1644511149
transform 1 0 44340 0 1 3598
box 0 0 1 1
use contact_9  contact_9_96
timestamp 1644511149
transform 1 0 51986 0 1 1339
box 0 0 1 1
use contact_9  contact_9_97
timestamp 1644511149
transform 1 0 42965 0 1 219
box 0 0 1 1
use contact_9  contact_9_98
timestamp 1644511149
transform 1 0 50738 0 1 1339
box 0 0 1 1
use contact_9  contact_9_99
timestamp 1644511149
transform 1 0 49490 0 1 1339
box 0 0 1 1
use contact_9  contact_9_100
timestamp 1644511149
transform 1 0 48242 0 1 1339
box 0 0 1 1
use contact_9  contact_9_101
timestamp 1644511149
transform 1 0 44498 0 1 1339
box 0 0 1 1
use contact_9  contact_9_102
timestamp 1644511149
transform 1 0 46994 0 1 1339
box 0 0 1 1
use contact_9  contact_9_103
timestamp 1644511149
transform 1 0 45746 0 1 1339
box 0 0 1 1
use contact_9  contact_9_104
timestamp 1644511149
transform 1 0 39506 0 1 1339
box 0 0 1 1
use contact_9  contact_9_105
timestamp 1644511149
transform 1 0 27026 0 1 1339
box 0 0 1 1
use contact_33  contact_33_0
timestamp 1644511149
transform 1 0 49485 0 1 -13781
box 0 0 1 1
use contact_33  contact_33_1
timestamp 1644511149
transform 1 0 40621 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_2
timestamp 1644511149
transform 1 0 46831 0 1 -6705
box 0 0 1 1
use contact_33  contact_33_3
timestamp 1644511149
transform 1 0 37464 0 1 -6949
box 0 0 1 1
use contact_33  contact_33_4
timestamp 1644511149
transform 1 0 40621 0 1 -14025
box 0 0 1 1
use contact_33  contact_33_5
timestamp 1644511149
transform 1 0 30109 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_6
timestamp 1644511149
transform 1 0 45583 0 1 -6949
box 0 0 1 1
use contact_33  contact_33_7
timestamp 1644511149
transform 1 0 36296 0 1 -7193
box 0 0 1 1
use contact_33  contact_33_8
timestamp 1644511149
transform 1 0 30109 0 1 -15245
box 0 0 1 1
use contact_33  contact_33_9
timestamp 1644511149
transform 1 0 48237 0 1 -14025
box 0 0 1 1
use contact_33  contact_33_10
timestamp 1644511149
transform 1 0 44335 0 1 -7193
box 0 0 1 1
use contact_33  contact_33_11
timestamp 1644511149
transform 1 0 32445 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_12
timestamp 1644511149
transform 1 0 32445 0 1 -14269
box 0 0 1 1
use contact_33  contact_33_13
timestamp 1644511149
transform 1 0 30607 0 1 -9877
box 0 0 1 1
use contact_33  contact_33_14
timestamp 1644511149
transform 1 0 30456 0 1 -10121
box 0 0 1 1
use contact_33  contact_33_15
timestamp 1644511149
transform 1 0 34351 0 1 -12317
box 0 0 1 1
use contact_33  contact_33_16
timestamp 1644511149
transform 1 0 27773 0 1 -15733
box 0 0 1 1
use contact_33  contact_33_17
timestamp 1644511149
transform 1 0 38095 0 1 -10121
box 0 0 1 1
use contact_33  contact_33_18
timestamp 1644511149
transform 1 0 33261 0 1 -15977
box 0 0 1 1
use contact_33  contact_33_19
timestamp 1644511149
transform 1 0 39501 0 1 -14269
box 0 0 1 1
use contact_33  contact_33_20
timestamp 1644511149
transform 1 0 39453 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_21
timestamp 1644511149
transform 1 0 29359 0 1 -10365
box 0 0 1 1
use contact_33  contact_33_22
timestamp 1644511149
transform 1 0 39453 0 1 -14513
box 0 0 1 1
use contact_33  contact_33_23
timestamp 1644511149
transform 1 0 37005 0 1 -15245
box 0 0 1 1
use contact_33  contact_33_24
timestamp 1644511149
transform 1 0 37117 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_25
timestamp 1644511149
transform 1 0 46989 0 1 -14513
box 0 0 1 1
use contact_33  contact_33_26
timestamp 1644511149
transform 1 0 44125 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_27
timestamp 1644511149
transform 1 0 28941 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_28
timestamp 1644511149
transform 1 0 44125 0 1 -13049
box 0 0 1 1
use contact_33  contact_33_29
timestamp 1644511149
transform 1 0 31277 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_30
timestamp 1644511149
transform 1 0 31277 0 1 -14757
box 0 0 1 1
use contact_33  contact_33_31
timestamp 1644511149
transform 1 0 51981 0 1 -13049
box 0 0 1 1
use contact_33  contact_33_32
timestamp 1644511149
transform 1 0 35949 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_33
timestamp 1644511149
transform 1 0 29517 0 1 -10853
box 0 0 1 1
use contact_33  contact_33_34
timestamp 1644511149
transform 1 0 29288 0 1 -11097
box 0 0 1 1
use contact_33  contact_33_35
timestamp 1644511149
transform 1 0 31855 0 1 -8413
box 0 0 1 1
use contact_33  contact_33_36
timestamp 1644511149
transform 1 0 31624 0 1 -8657
box 0 0 1 1
use contact_33  contact_33_37
timestamp 1644511149
transform 1 0 37117 0 1 -15489
box 0 0 1 1
use contact_33  contact_33_38
timestamp 1644511149
transform 1 0 32013 0 1 -16221
box 0 0 1 1
use contact_33  contact_33_39
timestamp 1644511149
transform 1 0 30765 0 1 -16465
box 0 0 1 1
use contact_33  contact_33_40
timestamp 1644511149
transform 1 0 39343 0 1 -8657
box 0 0 1 1
use contact_33  contact_33_41
timestamp 1644511149
transform 1 0 36847 0 1 -11097
box 0 0 1 1
use contact_33  contact_33_42
timestamp 1644511149
transform 1 0 33613 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_43
timestamp 1644511149
transform 1 0 38253 0 1 -14757
box 0 0 1 1
use contact_33  contact_33_44
timestamp 1644511149
transform 1 0 38285 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_45
timestamp 1644511149
transform 1 0 42960 0 1 -13293
box 0 0 1 1
use contact_33  contact_33_46
timestamp 1644511149
transform 1 0 42957 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_47
timestamp 1644511149
transform 1 0 34781 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_48
timestamp 1644511149
transform 1 0 42957 0 1 -13537
box 0 0 1 1
use contact_33  contact_33_49
timestamp 1644511149
transform 1 0 38285 0 1 -15001
box 0 0 1 1
use contact_33  contact_33_50
timestamp 1644511149
transform 1 0 34509 0 1 -15733
box 0 0 1 1
use contact_33  contact_33_51
timestamp 1644511149
transform 1 0 50733 0 1 -13537
box 0 0 1 1
use contact_33  contact_33_52
timestamp 1644511149
transform 1 0 41789 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_53
timestamp 1644511149
transform 1 0 41789 0 1 -13781
box 0 0 1 1
use contact_33  contact_33_54
timestamp 1644511149
transform 1 0 44493 0 1 -15489
box 0 0 1 1
use contact_33  contact_33_55
timestamp 1644511149
transform 1 0 27773 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_56
timestamp 1644511149
transform 1 0 38632 0 1 -6705
box 0 0 1 1
use contact_33  contact_33_57
timestamp 1644511149
transform 1 0 45741 0 1 -15001
box 0 0 1 1
use contact_33  contact_33_58
timestamp 1644511149
transform 1 0 20781 0 1 -11829
box 0 0 1 1
use contact_33  contact_33_59
timestamp 1644511149
transform 1 0 20765 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_60
timestamp 1644511149
transform 1 0 19597 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_61
timestamp 1644511149
transform 1 0 23119 0 1 -8901
box 0 0 1 1
use contact_33  contact_33_62
timestamp 1644511149
transform 1 0 10600 0 1 -9145
box 0 0 1 1
use contact_33  contact_33_63
timestamp 1644511149
transform 1 0 20765 0 1 -12073
box 0 0 1 1
use contact_33  contact_33_64
timestamp 1644511149
transform 1 0 26605 0 1 -15977
box 0 0 1 1
use contact_33  contact_33_65
timestamp 1644511149
transform 1 0 16879 0 1 -9145
box 0 0 1 1
use contact_33  contact_33_66
timestamp 1644511149
transform 1 0 11421 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_67
timestamp 1644511149
transform 1 0 11421 0 1 -9389
box 0 0 1 1
use contact_33  contact_33_68
timestamp 1644511149
transform 1 0 9085 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_69
timestamp 1644511149
transform 1 0 5581 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_70
timestamp 1644511149
transform 1 0 16093 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_71
timestamp 1644511149
transform 1 0 9085 0 1 -16953
box 0 0 1 1
use contact_33  contact_33_72
timestamp 1644511149
transform 1 0 17037 0 1 -9389
box 0 0 1 1
use contact_33  contact_33_73
timestamp 1644511149
transform 1 0 17261 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_74
timestamp 1644511149
transform 1 0 21933 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_75
timestamp 1644511149
transform 1 0 17261 0 1 -9633
box 0 0 1 1
use contact_33  contact_33_76
timestamp 1644511149
transform 1 0 26952 0 1 -12317
box 0 0 1 1
use contact_33  contact_33_77
timestamp 1644511149
transform 1 0 25437 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_78
timestamp 1644511149
transform 1 0 23277 0 1 -9633
box 0 0 1 1
use contact_33  contact_33_79
timestamp 1644511149
transform 1 0 23448 0 1 -9877
box 0 0 1 1
use contact_33  contact_33_80
timestamp 1644511149
transform 1 0 25437 0 1 -16221
box 0 0 1 1
use contact_33  contact_33_81
timestamp 1644511149
transform 1 0 9432 0 1 -12561
box 0 0 1 1
use contact_33  contact_33_82
timestamp 1644511149
transform 1 0 5979 0 1 -17441
box 0 0 1 1
use contact_33  contact_33_83
timestamp 1644511149
transform 1 0 13293 0 1 -17197
box 0 0 1 1
use contact_33  contact_33_84
timestamp 1644511149
transform 1 0 2077 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_85
timestamp 1644511149
transform 1 0 15631 0 1 -12561
box 0 0 1 1
use contact_33  contact_33_86
timestamp 1644511149
transform 1 0 22280 0 1 -10365
box 0 0 1 1
use contact_33  contact_33_87
timestamp 1644511149
transform 1 0 8264 0 1 -12805
box 0 0 1 1
use contact_33  contact_33_88
timestamp 1644511149
transform 1 0 24269 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_89
timestamp 1644511149
transform 1 0 4413 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_90
timestamp 1644511149
transform 1 0 4413 0 1 -10609
box 0 0 1 1
use contact_33  contact_33_91
timestamp 1644511149
transform 1 0 24269 0 1 -16465
box 0 0 1 1
use contact_33  contact_33_92
timestamp 1644511149
transform 1 0 14383 0 1 -12805
box 0 0 1 1
use contact_33  contact_33_93
timestamp 1644511149
transform 1 0 22992 0 1 -10609
box 0 0 1 1
use contact_33  contact_33_94
timestamp 1644511149
transform 1 0 23101 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_95
timestamp 1644511149
transform 1 0 23101 0 1 -10853
box 0 0 1 1
use contact_33  contact_33_96
timestamp 1644511149
transform 1 0 14541 0 1 -16953
box 0 0 1 1
use contact_33  contact_33_97
timestamp 1644511149
transform 1 0 7917 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_98
timestamp 1644511149
transform 1 0 17608 0 1 -7437
box 0 0 1 1
use contact_33  contact_33_99
timestamp 1644511149
transform 1 0 6749 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_100
timestamp 1644511149
transform 1 0 6749 0 1 -13293
box 0 0 1 1
use contact_33  contact_33_101
timestamp 1644511149
transform 1 0 24367 0 1 -7437
box 0 0 1 1
use contact_33  contact_33_102
timestamp 1644511149
transform 1 0 11768 0 1 -7681
box 0 0 1 1
use contact_33  contact_33_103
timestamp 1644511149
transform 1 0 19944 0 1 -11341
box 0 0 1 1
use contact_33  contact_33_104
timestamp 1644511149
transform 1 0 10253 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_105
timestamp 1644511149
transform 1 0 18127 0 1 -7681
box 0 0 1 1
use contact_33  contact_33_106
timestamp 1644511149
transform 1 0 12589 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_107
timestamp 1644511149
transform 1 0 12589 0 1 -7925
box 0 0 1 1
use contact_33  contact_33_108
timestamp 1644511149
transform 1 0 10253 0 1 -16709
box 0 0 1 1
use contact_33  contact_33_109
timestamp 1644511149
transform 1 0 26863 0 1 -11341
box 0 0 1 1
use contact_33  contact_33_110
timestamp 1644511149
transform 1 0 14104 0 1 -11585
box 0 0 1 1
use contact_33  contact_33_111
timestamp 1644511149
transform 1 0 18285 0 1 -7925
box 0 0 1 1
use contact_33  contact_33_112
timestamp 1644511149
transform 1 0 18429 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_113
timestamp 1644511149
transform 1 0 18429 0 1 -8169
box 0 0 1 1
use contact_33  contact_33_114
timestamp 1644511149
transform 1 0 7917 0 1 -17197
box 0 0 1 1
use contact_33  contact_33_115
timestamp 1644511149
transform 1 0 3245 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_116
timestamp 1644511149
transform 1 0 2077 0 1 -17441
box 0 0 1 1
use contact_33  contact_33_117
timestamp 1644511149
transform 1 0 24525 0 1 -8169
box 0 0 1 1
use contact_33  contact_33_118
timestamp 1644511149
transform 1 0 24616 0 1 -8413
box 0 0 1 1
use contact_33  contact_33_119
timestamp 1644511149
transform 1 0 20623 0 1 -11585
box 0 0 1 1
use contact_33  contact_33_120
timestamp 1644511149
transform 1 0 14925 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_121
timestamp 1644511149
transform 1 0 14925 0 1 -11829
box 0 0 1 1
use contact_33  contact_33_122
timestamp 1644511149
transform 1 0 15789 0 1 -16709
box 0 0 1 1
use contact_33  contact_33_123
timestamp 1644511149
transform 1 0 13757 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_124
timestamp 1644511149
transform 1 0 26605 0 1 -18354
box 0 0 1 1
use contact_33  contact_33_125
timestamp 1644511149
transform 1 0 16440 0 1 -8901
box 0 0 1 1
use contact_33  contact_33_126
timestamp 1644511149
transform 1 0 17037 0 1 1343
box 0 0 1 1
use contact_33  contact_33_127
timestamp 1644511149
transform 1 0 23277 0 1 1343
box 0 0 1 1
use contact_33  contact_33_128
timestamp 1644511149
transform 1 0 21112 0 1 -1093
box 0 0 1 1
use contact_33  contact_33_129
timestamp 1644511149
transform 1 0 13293 0 1 1343
box 0 0 1 1
use contact_33  contact_33_130
timestamp 1644511149
transform 1 0 15272 0 1 -1337
box 0 0 1 1
use contact_33  contact_33_131
timestamp 1644511149
transform 1 0 21871 0 1 3602
box 0 0 1 1
use contact_33  contact_33_132
timestamp 1644511149
transform 1 0 21871 0 1 -1337
box 0 0 1 1
use contact_33  contact_33_133
timestamp 1644511149
transform 1 0 16093 0 1 -1581
box 0 0 1 1
use contact_33  contact_33_134
timestamp 1644511149
transform 1 0 22029 0 1 1343
box 0 0 1 1
use contact_33  contact_33_135
timestamp 1644511149
transform 1 0 22029 0 1 -1581
box 0 0 1 1
use contact_33  contact_33_136
timestamp 1644511149
transform 1 0 21933 0 1 -1825
box 0 0 1 1
use contact_33  contact_33_137
timestamp 1644511149
transform 1 0 15631 0 1 3602
box 0 0 1 1
use contact_33  contact_33_138
timestamp 1644511149
transform 1 0 14383 0 1 3602
box 0 0 1 1
use contact_33  contact_33_139
timestamp 1644511149
transform 1 0 22992 0 1 223
box 0 0 1 1
use contact_33  contact_33_140
timestamp 1644511149
transform 1 0 5979 0 1 5408
box 0 0 1 1
use contact_33  contact_33_141
timestamp 1644511149
transform 1 0 15789 0 1 1343
box 0 0 1 1
use contact_33  contact_33_142
timestamp 1644511149
transform 1 0 26863 0 1 3602
box 0 0 1 1
use contact_33  contact_33_143
timestamp 1644511149
transform 1 0 20623 0 1 3602
box 0 0 1 1
use contact_33  contact_33_144
timestamp 1644511149
transform 1 0 20781 0 1 1343
box 0 0 1 1
use contact_33  contact_33_145
timestamp 1644511149
transform 1 0 24367 0 1 3602
box 0 0 1 1
use contact_33  contact_33_146
timestamp 1644511149
transform 1 0 18127 0 1 3602
box 0 0 1 1
use contact_33  contact_33_147
timestamp 1644511149
transform 1 0 18285 0 1 1343
box 0 0 1 1
use contact_33  contact_33_148
timestamp 1644511149
transform 1 0 24525 0 1 1343
box 0 0 1 1
use contact_33  contact_33_149
timestamp 1644511149
transform 1 0 14541 0 1 1343
box 0 0 1 1
use contact_33  contact_33_150
timestamp 1644511149
transform 1 0 18776 0 1 -3777
box 0 0 1 1
use contact_33  contact_33_151
timestamp 1644511149
transform 1 0 25615 0 1 3602
box 0 0 1 1
use contact_33  contact_33_152
timestamp 1644511149
transform 1 0 25615 0 1 -3777
box 0 0 1 1
use contact_33  contact_33_153
timestamp 1644511149
transform 1 0 7096 0 1 -4021
box 0 0 1 1
use contact_33  contact_33_154
timestamp 1644511149
transform 1 0 13135 0 1 3602
box 0 0 1 1
use contact_33  contact_33_155
timestamp 1644511149
transform 1 0 13135 0 1 -4021
box 0 0 1 1
use contact_33  contact_33_156
timestamp 1644511149
transform 1 0 3245 0 1 -4265
box 0 0 1 1
use contact_33  contact_33_157
timestamp 1644511149
transform 1 0 13008 0 1 223
box 0 0 1 1
use contact_33  contact_33_158
timestamp 1644511149
transform 1 0 13008 0 1 -4265
box 0 0 1 1
use contact_33  contact_33_159
timestamp 1644511149
transform 1 0 12936 0 1 -4509
box 0 0 1 1
use contact_33  contact_33_160
timestamp 1644511149
transform 1 0 19375 0 1 3602
box 0 0 1 1
use contact_33  contact_33_161
timestamp 1644511149
transform 1 0 19375 0 1 -4509
box 0 0 1 1
use contact_33  contact_33_162
timestamp 1644511149
transform 1 0 13757 0 1 -4753
box 0 0 1 1
use contact_33  contact_33_163
timestamp 1644511149
transform 1 0 19533 0 1 1343
box 0 0 1 1
use contact_33  contact_33_164
timestamp 1644511149
transform 1 0 19533 0 1 -4753
box 0 0 1 1
use contact_33  contact_33_165
timestamp 1644511149
transform 1 0 19597 0 1 -4997
box 0 0 1 1
use contact_33  contact_33_166
timestamp 1644511149
transform 1 0 25773 0 1 1343
box 0 0 1 1
use contact_33  contact_33_167
timestamp 1644511149
transform 1 0 25773 0 1 -4997
box 0 0 1 1
use contact_33  contact_33_168
timestamp 1644511149
transform 1 0 25784 0 1 -5241
box 0 0 1 1
use contact_33  contact_33_169
timestamp 1644511149
transform 1 0 23119 0 1 3602
box 0 0 1 1
use contact_33  contact_33_170
timestamp 1644511149
transform 1 0 16879 0 1 3602
box 0 0 1 1
use contact_33  contact_33_171
timestamp 1644511149
transform 1 0 5581 0 1 -5485
box 0 0 1 1
use contact_33  contact_33_172
timestamp 1644511149
transform 1 0 41997 0 1 -3289
box 0 0 1 1
use contact_33  contact_33_173
timestamp 1644511149
transform 1 0 42136 0 1 -3533
box 0 0 1 1
use contact_33  contact_33_174
timestamp 1644511149
transform 1 0 40749 0 1 -5973
box 0 0 1 1
use contact_33  contact_33_175
timestamp 1644511149
transform 1 0 41839 0 1 -3045
box 0 0 1 1
use contact_33  contact_33_176
timestamp 1644511149
transform 1 0 43087 0 1 -849
box 0 0 1 1
use contact_33  contact_33_177
timestamp 1644511149
transform 1 0 43245 0 1 -2557
box 0 0 1 1
use contact_33  contact_33_178
timestamp 1644511149
transform 1 0 43304 0 1 -2801
box 0 0 1 1
use contact_33  contact_33_179
timestamp 1644511149
transform 1 0 40968 0 1 -6217
box 0 0 1 1
use contact_33  contact_33_180
timestamp 1644511149
transform 1 0 40591 0 1 -5729
box 0 0 1 1
use contact_33  contact_33_181
timestamp 1644511149
transform 1 0 50575 0 1 -3533
box 0 0 1 1
use contact_33  contact_33_182
timestamp 1644511149
transform 1 0 51823 0 1 -2801
box 0 0 1 1
use contact_33  contact_33_183
timestamp 1644511149
transform 1 0 49327 0 1 -6217
box 0 0 1 1
use contact_33  contact_33_184
timestamp 1644511149
transform 1 0 35128 0 1 -849
box 0 0 1 1
use contact_33  contact_33_185
timestamp 1644511149
transform 1 0 33103 0 1 -5241
box 0 0 1 1
use contact_33  contact_33_186
timestamp 1644511149
transform 1 0 32792 0 1 -5729
box 0 0 1 1
use contact_33  contact_33_187
timestamp 1644511149
transform 1 0 35599 0 1 -2069
box 0 0 1 1
use contact_33  contact_33_188
timestamp 1644511149
transform 1 0 28941 0 1 -2313
box 0 0 1 1
use contact_33  contact_33_189
timestamp 1644511149
transform 1 0 33613 0 1 -5973
box 0 0 1 1
use contact_33  contact_33_190
timestamp 1644511149
transform 1 0 34781 0 1 -3289
box 0 0 1 1
use contact_33  contact_33_191
timestamp 1644511149
transform 1 0 28111 0 1 -1093
box 0 0 1 1
use contact_33  contact_33_192
timestamp 1644511149
transform 1 0 32976 0 1 -5485
box 0 0 1 1
use contact_33  contact_33_193
timestamp 1644511149
transform 1 0 35757 0 1 -2313
box 0 0 1 1
use contact_33  contact_33_194
timestamp 1644511149
transform 1 0 35949 0 1 -2557
box 0 0 1 1
use contact_33  contact_33_195
timestamp 1644511149
transform 1 0 28269 0 1 -1825
box 0 0 1 1
use contact_33  contact_33_196
timestamp 1644511149
transform 1 0 28120 0 1 -2069
box 0 0 1 1
use contact_33  contact_33_197
timestamp 1644511149
transform 1 0 33960 0 1 -3045
box 0 0 1 1
use contact_33  contact_33_198
timestamp 1644511149
transform 1 0 39343 0 1 3602
box 0 0 1 1
use contact_33  contact_33_199
timestamp 1644511149
transform 1 0 28111 0 1 3602
box 0 0 1 1
use contact_33  contact_33_200
timestamp 1644511149
transform 1 0 28269 0 1 1343
box 0 0 1 1
use contact_33  contact_33_201
timestamp 1644511149
transform 1 0 35599 0 1 3602
box 0 0 1 1
use contact_33  contact_33_202
timestamp 1644511149
transform 1 0 35757 0 1 1343
box 0 0 1 1
use contact_33  contact_33_203
timestamp 1644511149
transform 1 0 30607 0 1 3602
box 0 0 1 1
use contact_33  contact_33_204
timestamp 1644511149
transform 1 0 38095 0 1 3602
box 0 0 1 1
use contact_33  contact_33_205
timestamp 1644511149
transform 1 0 29359 0 1 3602
box 0 0 1 1
use contact_33  contact_33_206
timestamp 1644511149
transform 1 0 29517 0 1 1343
box 0 0 1 1
use contact_33  contact_33_207
timestamp 1644511149
transform 1 0 36847 0 1 3602
box 0 0 1 1
use contact_33  contact_33_208
timestamp 1644511149
transform 1 0 33103 0 1 3602
box 0 0 1 1
use contact_33  contact_33_209
timestamp 1644511149
transform 1 0 32976 0 1 223
box 0 0 1 1
use contact_33  contact_33_210
timestamp 1644511149
transform 1 0 30765 0 1 1343
box 0 0 1 1
use contact_33  contact_33_211
timestamp 1644511149
transform 1 0 34351 0 1 3602
box 0 0 1 1
use contact_33  contact_33_212
timestamp 1644511149
transform 1 0 32013 0 1 1343
box 0 0 1 1
use contact_33  contact_33_213
timestamp 1644511149
transform 1 0 37005 0 1 1343
box 0 0 1 1
use contact_33  contact_33_214
timestamp 1644511149
transform 1 0 33261 0 1 1343
box 0 0 1 1
use contact_33  contact_33_215
timestamp 1644511149
transform 1 0 38253 0 1 1343
box 0 0 1 1
use contact_33  contact_33_216
timestamp 1644511149
transform 1 0 34509 0 1 1343
box 0 0 1 1
use contact_33  contact_33_217
timestamp 1644511149
transform 1 0 31855 0 1 3602
box 0 0 1 1
use contact_33  contact_33_218
timestamp 1644511149
transform 1 0 43087 0 1 3602
box 0 0 1 1
use contact_33  contact_33_219
timestamp 1644511149
transform 1 0 43245 0 1 1343
box 0 0 1 1
use contact_33  contact_33_220
timestamp 1644511149
transform 1 0 51823 0 1 3602
box 0 0 1 1
use contact_33  contact_33_221
timestamp 1644511149
transform 1 0 41839 0 1 3602
box 0 0 1 1
use contact_33  contact_33_222
timestamp 1644511149
transform 1 0 41997 0 1 1343
box 0 0 1 1
use contact_33  contact_33_223
timestamp 1644511149
transform 1 0 50575 0 1 3602
box 0 0 1 1
use contact_33  contact_33_224
timestamp 1644511149
transform 1 0 40591 0 1 3602
box 0 0 1 1
use contact_33  contact_33_225
timestamp 1644511149
transform 1 0 40749 0 1 1343
box 0 0 1 1
use contact_33  contact_33_226
timestamp 1644511149
transform 1 0 49327 0 1 3602
box 0 0 1 1
use contact_33  contact_33_227
timestamp 1644511149
transform 1 0 48079 0 1 3602
box 0 0 1 1
use contact_33  contact_33_228
timestamp 1644511149
transform 1 0 46831 0 1 3602
box 0 0 1 1
use contact_33  contact_33_229
timestamp 1644511149
transform 1 0 45583 0 1 3602
box 0 0 1 1
use contact_33  contact_33_230
timestamp 1644511149
transform 1 0 44335 0 1 3602
box 0 0 1 1
use contact_33  contact_33_231
timestamp 1644511149
transform 1 0 51981 0 1 1343
box 0 0 1 1
use contact_33  contact_33_232
timestamp 1644511149
transform 1 0 42960 0 1 223
box 0 0 1 1
use contact_33  contact_33_233
timestamp 1644511149
transform 1 0 50733 0 1 1343
box 0 0 1 1
use contact_33  contact_33_234
timestamp 1644511149
transform 1 0 49485 0 1 1343
box 0 0 1 1
use contact_33  contact_33_235
timestamp 1644511149
transform 1 0 48237 0 1 1343
box 0 0 1 1
use contact_33  contact_33_236
timestamp 1644511149
transform 1 0 44493 0 1 1343
box 0 0 1 1
use contact_33  contact_33_237
timestamp 1644511149
transform 1 0 46989 0 1 1343
box 0 0 1 1
use contact_33  contact_33_238
timestamp 1644511149
transform 1 0 45741 0 1 1343
box 0 0 1 1
use contact_33  contact_33_239
timestamp 1644511149
transform 1 0 39501 0 1 1343
box 0 0 1 1
use contact_33  contact_33_240
timestamp 1644511149
transform 1 0 39800 0 1 -6461
box 0 0 1 1
use contact_33  contact_33_241
timestamp 1644511149
transform 1 0 48079 0 1 -6461
box 0 0 1 1
use contact_33  contact_33_242
timestamp 1644511149
transform 1 0 27021 0 1 1343
box 0 0 1 1
use contact_33  contact_33_243
timestamp 1644511149
transform 1 0 27021 0 1 -12073
box 0 0 1 1
<< properties >>
string FIXED_BBOX 2040 -18982 52094 5478
string GDS_END 5301308
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 5260728
<< end >>
