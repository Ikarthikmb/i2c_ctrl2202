magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< dnwell >>
rect 612 9680 14392 36196
<< nwell >>
rect 532 35932 14474 36278
rect 532 9944 818 35932
rect 14128 9944 14474 35932
rect 532 9598 14474 9944
<< nsubdiff >>
rect 569 36191 14437 36241
rect 569 36157 719 36191
rect 753 36157 787 36191
rect 821 36157 855 36191
rect 889 36157 923 36191
rect 957 36157 991 36191
rect 1025 36157 1059 36191
rect 1093 36157 1127 36191
rect 1161 36157 1195 36191
rect 1229 36157 1263 36191
rect 1297 36157 1331 36191
rect 1365 36157 1399 36191
rect 1433 36157 1467 36191
rect 1501 36157 1535 36191
rect 1569 36157 1603 36191
rect 1637 36157 1671 36191
rect 1705 36157 1739 36191
rect 1773 36157 1807 36191
rect 1841 36157 1875 36191
rect 1909 36157 1943 36191
rect 1977 36157 2011 36191
rect 2045 36157 2079 36191
rect 2113 36157 2147 36191
rect 2181 36157 2215 36191
rect 2249 36157 2283 36191
rect 2317 36157 2351 36191
rect 2385 36157 2419 36191
rect 2453 36157 2487 36191
rect 2521 36157 2555 36191
rect 2589 36157 2623 36191
rect 2657 36157 2691 36191
rect 2725 36157 2759 36191
rect 2793 36157 2827 36191
rect 2861 36157 2895 36191
rect 2929 36157 2963 36191
rect 2997 36157 3031 36191
rect 3065 36157 3099 36191
rect 3133 36157 3167 36191
rect 3201 36157 3235 36191
rect 3269 36157 3303 36191
rect 3337 36157 3371 36191
rect 3405 36157 3439 36191
rect 3473 36157 3507 36191
rect 3541 36157 3575 36191
rect 3609 36157 3643 36191
rect 3677 36157 3711 36191
rect 3745 36157 3779 36191
rect 3813 36157 3847 36191
rect 3881 36157 3915 36191
rect 3949 36157 3983 36191
rect 4017 36157 4051 36191
rect 4085 36157 4119 36191
rect 4153 36157 4187 36191
rect 4221 36157 4255 36191
rect 4289 36157 4323 36191
rect 4357 36157 4391 36191
rect 4425 36157 4459 36191
rect 4493 36157 4527 36191
rect 4561 36157 4595 36191
rect 4629 36157 4663 36191
rect 4697 36157 4731 36191
rect 4765 36157 4799 36191
rect 4833 36157 4867 36191
rect 4901 36157 4935 36191
rect 4969 36157 5003 36191
rect 5037 36157 5071 36191
rect 5105 36157 5139 36191
rect 5173 36157 5207 36191
rect 5241 36157 5275 36191
rect 5309 36157 5343 36191
rect 5377 36157 5411 36191
rect 5445 36157 5479 36191
rect 5513 36157 5547 36191
rect 5581 36157 5615 36191
rect 5649 36157 5683 36191
rect 5717 36157 5751 36191
rect 5785 36157 5819 36191
rect 5853 36157 5887 36191
rect 5921 36157 5955 36191
rect 5989 36157 6023 36191
rect 6057 36157 6091 36191
rect 6125 36157 6159 36191
rect 6193 36157 6227 36191
rect 6261 36157 6295 36191
rect 6329 36157 6363 36191
rect 6397 36157 6431 36191
rect 6465 36157 6499 36191
rect 6533 36157 6567 36191
rect 6601 36157 6635 36191
rect 6669 36157 6703 36191
rect 6737 36157 6771 36191
rect 6805 36157 6839 36191
rect 6873 36157 6907 36191
rect 6941 36157 6975 36191
rect 7009 36157 7043 36191
rect 7077 36157 7111 36191
rect 7145 36157 7179 36191
rect 7213 36157 7247 36191
rect 7281 36157 7315 36191
rect 7349 36157 7383 36191
rect 7417 36157 7451 36191
rect 7485 36157 7519 36191
rect 7553 36157 7587 36191
rect 7621 36157 7655 36191
rect 7689 36157 7723 36191
rect 7757 36157 7791 36191
rect 7825 36157 7859 36191
rect 7893 36157 7927 36191
rect 7961 36157 7995 36191
rect 8029 36157 8063 36191
rect 8097 36157 8131 36191
rect 8165 36157 8199 36191
rect 8233 36157 8267 36191
rect 8301 36157 8335 36191
rect 8369 36157 8403 36191
rect 8437 36157 8471 36191
rect 8505 36157 8539 36191
rect 8573 36157 8607 36191
rect 8641 36157 8675 36191
rect 8709 36157 8743 36191
rect 8777 36157 8811 36191
rect 8845 36157 8879 36191
rect 8913 36157 8947 36191
rect 8981 36157 9015 36191
rect 9049 36157 9083 36191
rect 9117 36157 9151 36191
rect 9185 36157 9219 36191
rect 9253 36157 9287 36191
rect 9321 36157 9355 36191
rect 9389 36157 9423 36191
rect 9457 36157 9491 36191
rect 9525 36157 9559 36191
rect 9593 36157 9627 36191
rect 9661 36157 9695 36191
rect 9729 36157 9763 36191
rect 9797 36157 9831 36191
rect 9865 36157 9899 36191
rect 9933 36157 9967 36191
rect 10001 36157 10035 36191
rect 10069 36157 10103 36191
rect 10137 36157 10171 36191
rect 10205 36157 10239 36191
rect 10273 36157 10307 36191
rect 10341 36157 10375 36191
rect 10409 36157 10443 36191
rect 10477 36157 10511 36191
rect 10545 36157 10579 36191
rect 10613 36157 10647 36191
rect 10681 36157 10715 36191
rect 10749 36157 10783 36191
rect 10817 36157 10851 36191
rect 10885 36157 10919 36191
rect 10953 36157 10987 36191
rect 11021 36157 11055 36191
rect 11089 36157 11123 36191
rect 11157 36157 11191 36191
rect 11225 36157 11259 36191
rect 11293 36157 11327 36191
rect 11361 36157 11395 36191
rect 11429 36157 11463 36191
rect 11497 36157 11531 36191
rect 11565 36157 11599 36191
rect 11633 36157 11667 36191
rect 11701 36157 11735 36191
rect 11769 36157 11803 36191
rect 11837 36157 11871 36191
rect 11905 36157 11939 36191
rect 11973 36157 12007 36191
rect 12041 36157 12075 36191
rect 12109 36157 12143 36191
rect 12177 36157 12211 36191
rect 12245 36157 12279 36191
rect 12313 36157 12347 36191
rect 12381 36157 12415 36191
rect 12449 36157 12483 36191
rect 12517 36157 12551 36191
rect 12585 36157 12619 36191
rect 12653 36157 12687 36191
rect 12721 36157 12755 36191
rect 12789 36157 12823 36191
rect 12857 36157 12891 36191
rect 12925 36157 12959 36191
rect 12993 36157 13027 36191
rect 13061 36157 13095 36191
rect 13129 36157 13163 36191
rect 13197 36157 13231 36191
rect 13265 36157 13299 36191
rect 13333 36157 13367 36191
rect 13401 36157 13435 36191
rect 13469 36157 13503 36191
rect 13537 36157 13571 36191
rect 13605 36157 13639 36191
rect 13673 36157 13707 36191
rect 13741 36157 13775 36191
rect 13809 36157 13843 36191
rect 13877 36157 13911 36191
rect 13945 36157 13979 36191
rect 14013 36157 14047 36191
rect 14081 36157 14115 36191
rect 14149 36157 14183 36191
rect 14217 36157 14251 36191
rect 14285 36157 14437 36191
rect 569 36107 14437 36157
rect 569 36079 701 36107
rect 569 36045 618 36079
rect 652 36045 701 36079
rect 569 36011 701 36045
rect 569 35977 618 36011
rect 652 35977 701 36011
rect 569 35943 701 35977
rect 569 35909 618 35943
rect 652 35909 701 35943
rect 569 35875 701 35909
rect 569 35841 618 35875
rect 652 35841 701 35875
rect 569 35807 701 35841
rect 569 35773 618 35807
rect 652 35773 701 35807
rect 569 35739 701 35773
rect 569 35705 618 35739
rect 652 35705 701 35739
rect 569 35671 701 35705
rect 569 35637 618 35671
rect 652 35637 701 35671
rect 569 35603 701 35637
rect 569 35569 618 35603
rect 652 35569 701 35603
rect 569 35535 701 35569
rect 569 35501 618 35535
rect 652 35501 701 35535
rect 569 35467 701 35501
rect 569 35433 618 35467
rect 652 35433 701 35467
rect 569 35399 701 35433
rect 569 35365 618 35399
rect 652 35365 701 35399
rect 569 35331 701 35365
rect 569 35297 618 35331
rect 652 35297 701 35331
rect 569 35263 701 35297
rect 569 35229 618 35263
rect 652 35229 701 35263
rect 569 35195 701 35229
rect 569 35161 618 35195
rect 652 35161 701 35195
rect 569 35127 701 35161
rect 569 35093 618 35127
rect 652 35093 701 35127
rect 569 35059 701 35093
rect 569 35025 618 35059
rect 652 35025 701 35059
rect 569 34991 701 35025
rect 569 34957 618 34991
rect 652 34957 701 34991
rect 569 34923 701 34957
rect 569 34889 618 34923
rect 652 34889 701 34923
rect 569 34855 701 34889
rect 569 34821 618 34855
rect 652 34821 701 34855
rect 569 34787 701 34821
rect 569 34753 618 34787
rect 652 34753 701 34787
rect 569 34719 701 34753
rect 569 34685 618 34719
rect 652 34685 701 34719
rect 569 34651 701 34685
rect 569 34617 618 34651
rect 652 34617 701 34651
rect 569 34583 701 34617
rect 569 34549 618 34583
rect 652 34549 701 34583
rect 569 34515 701 34549
rect 569 34481 618 34515
rect 652 34481 701 34515
rect 569 34447 701 34481
rect 569 34413 618 34447
rect 652 34413 701 34447
rect 569 34379 701 34413
rect 569 34345 618 34379
rect 652 34345 701 34379
rect 569 34311 701 34345
rect 569 34277 618 34311
rect 652 34277 701 34311
rect 569 34243 701 34277
rect 569 34209 618 34243
rect 652 34209 701 34243
rect 569 34175 701 34209
rect 569 34141 618 34175
rect 652 34141 701 34175
rect 569 34107 701 34141
rect 569 34073 618 34107
rect 652 34073 701 34107
rect 569 34039 701 34073
rect 569 34005 618 34039
rect 652 34005 701 34039
rect 569 33971 701 34005
rect 569 33937 618 33971
rect 652 33937 701 33971
rect 569 33903 701 33937
rect 569 33869 618 33903
rect 652 33869 701 33903
rect 569 33835 701 33869
rect 569 33801 618 33835
rect 652 33801 701 33835
rect 569 33767 701 33801
rect 569 33733 618 33767
rect 652 33733 701 33767
rect 569 33699 701 33733
rect 569 33665 618 33699
rect 652 33665 701 33699
rect 569 33631 701 33665
rect 569 33597 618 33631
rect 652 33597 701 33631
rect 569 33563 701 33597
rect 569 33529 618 33563
rect 652 33529 701 33563
rect 569 33495 701 33529
rect 569 33461 618 33495
rect 652 33461 701 33495
rect 569 33427 701 33461
rect 569 33393 618 33427
rect 652 33393 701 33427
rect 569 33359 701 33393
rect 569 33325 618 33359
rect 652 33325 701 33359
rect 569 33291 701 33325
rect 569 33257 618 33291
rect 652 33257 701 33291
rect 569 33223 701 33257
rect 569 33189 618 33223
rect 652 33189 701 33223
rect 569 33155 701 33189
rect 569 33121 618 33155
rect 652 33121 701 33155
rect 569 33087 701 33121
rect 569 33053 618 33087
rect 652 33053 701 33087
rect 569 33019 701 33053
rect 569 32985 618 33019
rect 652 32985 701 33019
rect 569 32951 701 32985
rect 569 32917 618 32951
rect 652 32917 701 32951
rect 569 32883 701 32917
rect 569 32849 618 32883
rect 652 32849 701 32883
rect 569 32815 701 32849
rect 569 32781 618 32815
rect 652 32781 701 32815
rect 569 32747 701 32781
rect 569 32713 618 32747
rect 652 32713 701 32747
rect 569 32679 701 32713
rect 569 32645 618 32679
rect 652 32645 701 32679
rect 569 32611 701 32645
rect 569 32577 618 32611
rect 652 32577 701 32611
rect 569 32543 701 32577
rect 569 32509 618 32543
rect 652 32509 701 32543
rect 569 32475 701 32509
rect 569 32441 618 32475
rect 652 32441 701 32475
rect 569 32407 701 32441
rect 569 32373 618 32407
rect 652 32373 701 32407
rect 569 32339 701 32373
rect 569 32305 618 32339
rect 652 32305 701 32339
rect 569 32271 701 32305
rect 569 32237 618 32271
rect 652 32237 701 32271
rect 569 32203 701 32237
rect 569 32169 618 32203
rect 652 32169 701 32203
rect 569 32135 701 32169
rect 569 32101 618 32135
rect 652 32101 701 32135
rect 569 32067 701 32101
rect 569 32033 618 32067
rect 652 32033 701 32067
rect 569 31999 701 32033
rect 569 31965 618 31999
rect 652 31965 701 31999
rect 569 31931 701 31965
rect 569 31897 618 31931
rect 652 31897 701 31931
rect 569 31863 701 31897
rect 569 31829 618 31863
rect 652 31829 701 31863
rect 569 31795 701 31829
rect 569 31761 618 31795
rect 652 31761 701 31795
rect 569 31727 701 31761
rect 569 31693 618 31727
rect 652 31693 701 31727
rect 569 31659 701 31693
rect 569 31625 618 31659
rect 652 31625 701 31659
rect 569 31591 701 31625
rect 569 31557 618 31591
rect 652 31557 701 31591
rect 569 31523 701 31557
rect 569 31489 618 31523
rect 652 31489 701 31523
rect 569 31455 701 31489
rect 569 31421 618 31455
rect 652 31421 701 31455
rect 569 31387 701 31421
rect 569 31353 618 31387
rect 652 31353 701 31387
rect 569 31319 701 31353
rect 569 31285 618 31319
rect 652 31285 701 31319
rect 569 31251 701 31285
rect 569 31217 618 31251
rect 652 31217 701 31251
rect 569 31183 701 31217
rect 569 31149 618 31183
rect 652 31149 701 31183
rect 569 31115 701 31149
rect 569 31081 618 31115
rect 652 31081 701 31115
rect 569 31047 701 31081
rect 569 31013 618 31047
rect 652 31013 701 31047
rect 569 30979 701 31013
rect 569 30945 618 30979
rect 652 30945 701 30979
rect 569 30911 701 30945
rect 569 30877 618 30911
rect 652 30877 701 30911
rect 569 30843 701 30877
rect 569 30809 618 30843
rect 652 30809 701 30843
rect 569 30775 701 30809
rect 569 30741 618 30775
rect 652 30741 701 30775
rect 569 30707 701 30741
rect 569 30673 618 30707
rect 652 30673 701 30707
rect 569 30639 701 30673
rect 569 30605 618 30639
rect 652 30605 701 30639
rect 569 30571 701 30605
rect 569 30537 618 30571
rect 652 30537 701 30571
rect 569 30503 701 30537
rect 569 30469 618 30503
rect 652 30469 701 30503
rect 569 30435 701 30469
rect 569 30401 618 30435
rect 652 30401 701 30435
rect 569 30367 701 30401
rect 569 30333 618 30367
rect 652 30333 701 30367
rect 569 30299 701 30333
rect 569 30265 618 30299
rect 652 30265 701 30299
rect 569 30231 701 30265
rect 569 30197 618 30231
rect 652 30197 701 30231
rect 569 30163 701 30197
rect 569 30129 618 30163
rect 652 30129 701 30163
rect 569 30095 701 30129
rect 569 30061 618 30095
rect 652 30061 701 30095
rect 569 30027 701 30061
rect 569 29993 618 30027
rect 652 29993 701 30027
rect 569 29959 701 29993
rect 569 29925 618 29959
rect 652 29925 701 29959
rect 569 29891 701 29925
rect 569 29857 618 29891
rect 652 29857 701 29891
rect 569 29823 701 29857
rect 569 29789 618 29823
rect 652 29789 701 29823
rect 569 29755 701 29789
rect 569 29721 618 29755
rect 652 29721 701 29755
rect 569 29687 701 29721
rect 569 29653 618 29687
rect 652 29653 701 29687
rect 569 29619 701 29653
rect 569 29585 618 29619
rect 652 29585 701 29619
rect 569 29551 701 29585
rect 569 29517 618 29551
rect 652 29517 701 29551
rect 569 29483 701 29517
rect 569 29449 618 29483
rect 652 29449 701 29483
rect 569 29415 701 29449
rect 569 29381 618 29415
rect 652 29381 701 29415
rect 569 29347 701 29381
rect 569 29313 618 29347
rect 652 29313 701 29347
rect 569 29279 701 29313
rect 569 29245 618 29279
rect 652 29245 701 29279
rect 569 29211 701 29245
rect 569 29177 618 29211
rect 652 29177 701 29211
rect 569 29143 701 29177
rect 569 29109 618 29143
rect 652 29109 701 29143
rect 569 29075 701 29109
rect 569 29041 618 29075
rect 652 29041 701 29075
rect 569 29007 701 29041
rect 569 28973 618 29007
rect 652 28973 701 29007
rect 569 28939 701 28973
rect 569 28905 618 28939
rect 652 28905 701 28939
rect 569 28871 701 28905
rect 569 28837 618 28871
rect 652 28837 701 28871
rect 569 28803 701 28837
rect 569 28769 618 28803
rect 652 28769 701 28803
rect 569 28735 701 28769
rect 569 28701 618 28735
rect 652 28701 701 28735
rect 569 28667 701 28701
rect 569 28633 618 28667
rect 652 28633 701 28667
rect 569 28599 701 28633
rect 569 28565 618 28599
rect 652 28565 701 28599
rect 569 28531 701 28565
rect 569 28497 618 28531
rect 652 28497 701 28531
rect 569 28463 701 28497
rect 569 28429 618 28463
rect 652 28429 701 28463
rect 569 28395 701 28429
rect 569 28361 618 28395
rect 652 28361 701 28395
rect 569 28327 701 28361
rect 569 28293 618 28327
rect 652 28293 701 28327
rect 569 28259 701 28293
rect 569 28225 618 28259
rect 652 28225 701 28259
rect 569 28191 701 28225
rect 569 28157 618 28191
rect 652 28157 701 28191
rect 569 28123 701 28157
rect 569 28089 618 28123
rect 652 28089 701 28123
rect 569 28055 701 28089
rect 569 28021 618 28055
rect 652 28021 701 28055
rect 569 27987 701 28021
rect 569 27953 618 27987
rect 652 27953 701 27987
rect 569 27919 701 27953
rect 569 27885 618 27919
rect 652 27885 701 27919
rect 569 27851 701 27885
rect 569 27817 618 27851
rect 652 27817 701 27851
rect 569 27783 701 27817
rect 569 27749 618 27783
rect 652 27749 701 27783
rect 569 27715 701 27749
rect 569 27681 618 27715
rect 652 27681 701 27715
rect 569 27647 701 27681
rect 569 27613 618 27647
rect 652 27613 701 27647
rect 569 27579 701 27613
rect 569 27545 618 27579
rect 652 27545 701 27579
rect 569 27511 701 27545
rect 569 27477 618 27511
rect 652 27477 701 27511
rect 569 27443 701 27477
rect 569 27409 618 27443
rect 652 27409 701 27443
rect 569 27375 701 27409
rect 569 27341 618 27375
rect 652 27341 701 27375
rect 569 27307 701 27341
rect 569 27273 618 27307
rect 652 27273 701 27307
rect 569 27239 701 27273
rect 569 27205 618 27239
rect 652 27205 701 27239
rect 569 27171 701 27205
rect 569 27137 618 27171
rect 652 27137 701 27171
rect 569 27103 701 27137
rect 569 27069 618 27103
rect 652 27069 701 27103
rect 569 27035 701 27069
rect 569 27001 618 27035
rect 652 27001 701 27035
rect 569 26967 701 27001
rect 569 26933 618 26967
rect 652 26933 701 26967
rect 569 26899 701 26933
rect 569 26865 618 26899
rect 652 26865 701 26899
rect 569 26831 701 26865
rect 569 26797 618 26831
rect 652 26797 701 26831
rect 569 26763 701 26797
rect 569 26729 618 26763
rect 652 26729 701 26763
rect 569 26695 701 26729
rect 569 26661 618 26695
rect 652 26661 701 26695
rect 569 26627 701 26661
rect 569 26593 618 26627
rect 652 26593 701 26627
rect 569 26559 701 26593
rect 569 26525 618 26559
rect 652 26525 701 26559
rect 569 26491 701 26525
rect 569 26457 618 26491
rect 652 26457 701 26491
rect 569 26423 701 26457
rect 569 26389 618 26423
rect 652 26389 701 26423
rect 569 26355 701 26389
rect 569 26321 618 26355
rect 652 26321 701 26355
rect 569 26287 701 26321
rect 569 26253 618 26287
rect 652 26253 701 26287
rect 569 26219 701 26253
rect 569 26185 618 26219
rect 652 26185 701 26219
rect 569 26151 701 26185
rect 569 26117 618 26151
rect 652 26117 701 26151
rect 569 26083 701 26117
rect 569 26049 618 26083
rect 652 26049 701 26083
rect 569 26015 701 26049
rect 569 25981 618 26015
rect 652 25981 701 26015
rect 569 25947 701 25981
rect 569 25913 618 25947
rect 652 25913 701 25947
rect 569 25879 701 25913
rect 569 25845 618 25879
rect 652 25845 701 25879
rect 569 25811 701 25845
rect 569 25777 618 25811
rect 652 25777 701 25811
rect 569 25743 701 25777
rect 569 25709 618 25743
rect 652 25709 701 25743
rect 569 25675 701 25709
rect 569 25641 618 25675
rect 652 25641 701 25675
rect 569 25607 701 25641
rect 569 25573 618 25607
rect 652 25573 701 25607
rect 569 25539 701 25573
rect 569 25505 618 25539
rect 652 25505 701 25539
rect 569 25471 701 25505
rect 569 25437 618 25471
rect 652 25437 701 25471
rect 569 25403 701 25437
rect 569 25369 618 25403
rect 652 25369 701 25403
rect 569 25335 701 25369
rect 569 25301 618 25335
rect 652 25301 701 25335
rect 569 25267 701 25301
rect 569 25233 618 25267
rect 652 25233 701 25267
rect 569 25199 701 25233
rect 569 25165 618 25199
rect 652 25165 701 25199
rect 569 25131 701 25165
rect 569 25097 618 25131
rect 652 25097 701 25131
rect 569 25063 701 25097
rect 569 25029 618 25063
rect 652 25029 701 25063
rect 569 24995 701 25029
rect 569 24961 618 24995
rect 652 24961 701 24995
rect 569 24927 701 24961
rect 569 24893 618 24927
rect 652 24893 701 24927
rect 569 24859 701 24893
rect 569 24825 618 24859
rect 652 24825 701 24859
rect 569 24791 701 24825
rect 569 24757 618 24791
rect 652 24757 701 24791
rect 569 24723 701 24757
rect 569 24689 618 24723
rect 652 24689 701 24723
rect 569 24655 701 24689
rect 569 24621 618 24655
rect 652 24621 701 24655
rect 569 24587 701 24621
rect 569 24553 618 24587
rect 652 24553 701 24587
rect 569 24519 701 24553
rect 569 24485 618 24519
rect 652 24485 701 24519
rect 569 24451 701 24485
rect 569 24417 618 24451
rect 652 24417 701 24451
rect 569 24383 701 24417
rect 569 24349 618 24383
rect 652 24349 701 24383
rect 569 24315 701 24349
rect 569 24281 618 24315
rect 652 24281 701 24315
rect 569 24247 701 24281
rect 569 24213 618 24247
rect 652 24213 701 24247
rect 569 24179 701 24213
rect 569 24145 618 24179
rect 652 24145 701 24179
rect 569 24111 701 24145
rect 569 24077 618 24111
rect 652 24077 701 24111
rect 569 24043 701 24077
rect 569 24009 618 24043
rect 652 24009 701 24043
rect 569 23975 701 24009
rect 569 23941 618 23975
rect 652 23941 701 23975
rect 569 23907 701 23941
rect 569 23873 618 23907
rect 652 23873 701 23907
rect 569 23839 701 23873
rect 569 23805 618 23839
rect 652 23805 701 23839
rect 569 23771 701 23805
rect 569 23737 618 23771
rect 652 23737 701 23771
rect 569 23703 701 23737
rect 569 23669 618 23703
rect 652 23669 701 23703
rect 569 23635 701 23669
rect 569 23601 618 23635
rect 652 23601 701 23635
rect 569 23567 701 23601
rect 569 23533 618 23567
rect 652 23533 701 23567
rect 569 23499 701 23533
rect 569 23465 618 23499
rect 652 23465 701 23499
rect 569 23431 701 23465
rect 569 23397 618 23431
rect 652 23397 701 23431
rect 569 23363 701 23397
rect 569 23329 618 23363
rect 652 23329 701 23363
rect 569 23295 701 23329
rect 569 23261 618 23295
rect 652 23261 701 23295
rect 569 23227 701 23261
rect 569 23193 618 23227
rect 652 23193 701 23227
rect 569 23159 701 23193
rect 569 23125 618 23159
rect 652 23125 701 23159
rect 569 23091 701 23125
rect 569 23057 618 23091
rect 652 23057 701 23091
rect 569 23023 701 23057
rect 569 22989 618 23023
rect 652 22989 701 23023
rect 569 22955 701 22989
rect 569 22921 618 22955
rect 652 22921 701 22955
rect 569 22887 701 22921
rect 569 22853 618 22887
rect 652 22853 701 22887
rect 569 22819 701 22853
rect 569 22785 618 22819
rect 652 22785 701 22819
rect 569 22751 701 22785
rect 569 22717 618 22751
rect 652 22717 701 22751
rect 569 22683 701 22717
rect 569 22649 618 22683
rect 652 22649 701 22683
rect 569 22615 701 22649
rect 569 22581 618 22615
rect 652 22581 701 22615
rect 569 22547 701 22581
rect 569 22513 618 22547
rect 652 22513 701 22547
rect 569 22479 701 22513
rect 569 22445 618 22479
rect 652 22445 701 22479
rect 569 22411 701 22445
rect 569 22377 618 22411
rect 652 22377 701 22411
rect 569 22343 701 22377
rect 569 22309 618 22343
rect 652 22309 701 22343
rect 569 22275 701 22309
rect 569 22241 618 22275
rect 652 22241 701 22275
rect 569 22207 701 22241
rect 569 22173 618 22207
rect 652 22173 701 22207
rect 569 22139 701 22173
rect 569 22105 618 22139
rect 652 22105 701 22139
rect 569 22071 701 22105
rect 569 22037 618 22071
rect 652 22037 701 22071
rect 569 22003 701 22037
rect 569 21969 618 22003
rect 652 21969 701 22003
rect 569 21935 701 21969
rect 569 21901 618 21935
rect 652 21901 701 21935
rect 569 21867 701 21901
rect 569 21833 618 21867
rect 652 21833 701 21867
rect 569 21799 701 21833
rect 569 21765 618 21799
rect 652 21765 701 21799
rect 569 21731 701 21765
rect 569 21697 618 21731
rect 652 21697 701 21731
rect 569 21663 701 21697
rect 569 21629 618 21663
rect 652 21629 701 21663
rect 569 21595 701 21629
rect 569 21561 618 21595
rect 652 21561 701 21595
rect 569 21527 701 21561
rect 569 21493 618 21527
rect 652 21493 701 21527
rect 569 21459 701 21493
rect 569 21425 618 21459
rect 652 21425 701 21459
rect 569 21391 701 21425
rect 569 21357 618 21391
rect 652 21357 701 21391
rect 569 21323 701 21357
rect 569 21289 618 21323
rect 652 21289 701 21323
rect 569 21255 701 21289
rect 569 21221 618 21255
rect 652 21221 701 21255
rect 569 21187 701 21221
rect 569 21153 618 21187
rect 652 21153 701 21187
rect 569 21119 701 21153
rect 569 21085 618 21119
rect 652 21085 701 21119
rect 569 21051 701 21085
rect 569 21017 618 21051
rect 652 21017 701 21051
rect 569 20983 701 21017
rect 569 20949 618 20983
rect 652 20949 701 20983
rect 569 20915 701 20949
rect 569 20881 618 20915
rect 652 20881 701 20915
rect 569 20847 701 20881
rect 569 20813 618 20847
rect 652 20813 701 20847
rect 569 20779 701 20813
rect 569 20745 618 20779
rect 652 20745 701 20779
rect 569 20711 701 20745
rect 569 20677 618 20711
rect 652 20677 701 20711
rect 569 20643 701 20677
rect 569 20609 618 20643
rect 652 20609 701 20643
rect 569 20575 701 20609
rect 569 20541 618 20575
rect 652 20541 701 20575
rect 569 20507 701 20541
rect 569 20473 618 20507
rect 652 20473 701 20507
rect 569 20439 701 20473
rect 569 20405 618 20439
rect 652 20405 701 20439
rect 569 20371 701 20405
rect 569 20337 618 20371
rect 652 20337 701 20371
rect 569 20303 701 20337
rect 569 20269 618 20303
rect 652 20269 701 20303
rect 569 20235 701 20269
rect 569 20201 618 20235
rect 652 20201 701 20235
rect 569 20167 701 20201
rect 569 20133 618 20167
rect 652 20133 701 20167
rect 569 20099 701 20133
rect 569 20065 618 20099
rect 652 20065 701 20099
rect 569 20031 701 20065
rect 569 19997 618 20031
rect 652 19997 701 20031
rect 569 19963 701 19997
rect 569 19929 618 19963
rect 652 19929 701 19963
rect 569 19895 701 19929
rect 569 19861 618 19895
rect 652 19861 701 19895
rect 569 19827 701 19861
rect 569 19793 618 19827
rect 652 19793 701 19827
rect 569 19759 701 19793
rect 569 19725 618 19759
rect 652 19725 701 19759
rect 569 19691 701 19725
rect 569 19657 618 19691
rect 652 19657 701 19691
rect 569 19623 701 19657
rect 569 19589 618 19623
rect 652 19589 701 19623
rect 569 19555 701 19589
rect 569 19521 618 19555
rect 652 19521 701 19555
rect 569 19487 701 19521
rect 569 19453 618 19487
rect 652 19453 701 19487
rect 569 19419 701 19453
rect 569 19385 618 19419
rect 652 19385 701 19419
rect 569 19351 701 19385
rect 569 19317 618 19351
rect 652 19317 701 19351
rect 569 19283 701 19317
rect 569 19249 618 19283
rect 652 19249 701 19283
rect 569 19215 701 19249
rect 569 19181 618 19215
rect 652 19181 701 19215
rect 569 19147 701 19181
rect 569 19113 618 19147
rect 652 19113 701 19147
rect 569 19079 701 19113
rect 569 19045 618 19079
rect 652 19045 701 19079
rect 569 19011 701 19045
rect 569 18977 618 19011
rect 652 18977 701 19011
rect 569 18943 701 18977
rect 569 18909 618 18943
rect 652 18909 701 18943
rect 569 18875 701 18909
rect 569 18841 618 18875
rect 652 18841 701 18875
rect 569 18807 701 18841
rect 569 18773 618 18807
rect 652 18773 701 18807
rect 569 18739 701 18773
rect 569 18705 618 18739
rect 652 18705 701 18739
rect 569 18671 701 18705
rect 569 18637 618 18671
rect 652 18637 701 18671
rect 569 18603 701 18637
rect 569 18569 618 18603
rect 652 18569 701 18603
rect 569 18535 701 18569
rect 569 18501 618 18535
rect 652 18501 701 18535
rect 569 18467 701 18501
rect 569 18433 618 18467
rect 652 18433 701 18467
rect 569 18399 701 18433
rect 569 18365 618 18399
rect 652 18365 701 18399
rect 569 18331 701 18365
rect 569 18297 618 18331
rect 652 18297 701 18331
rect 569 18263 701 18297
rect 569 18229 618 18263
rect 652 18229 701 18263
rect 569 18195 701 18229
rect 569 18161 618 18195
rect 652 18161 701 18195
rect 569 18127 701 18161
rect 569 18093 618 18127
rect 652 18093 701 18127
rect 569 18059 701 18093
rect 569 18025 618 18059
rect 652 18025 701 18059
rect 569 17991 701 18025
rect 569 17957 618 17991
rect 652 17957 701 17991
rect 569 17923 701 17957
rect 569 17889 618 17923
rect 652 17889 701 17923
rect 569 17855 701 17889
rect 569 17821 618 17855
rect 652 17821 701 17855
rect 569 17787 701 17821
rect 569 17753 618 17787
rect 652 17753 701 17787
rect 569 17719 701 17753
rect 569 17685 618 17719
rect 652 17685 701 17719
rect 569 17651 701 17685
rect 569 17617 618 17651
rect 652 17617 701 17651
rect 569 17583 701 17617
rect 569 17549 618 17583
rect 652 17549 701 17583
rect 569 17515 701 17549
rect 569 17481 618 17515
rect 652 17481 701 17515
rect 569 17447 701 17481
rect 569 17413 618 17447
rect 652 17413 701 17447
rect 569 17379 701 17413
rect 569 17345 618 17379
rect 652 17345 701 17379
rect 569 17311 701 17345
rect 569 17277 618 17311
rect 652 17277 701 17311
rect 569 17243 701 17277
rect 569 17209 618 17243
rect 652 17209 701 17243
rect 569 17175 701 17209
rect 569 17141 618 17175
rect 652 17141 701 17175
rect 569 17107 701 17141
rect 569 17073 618 17107
rect 652 17073 701 17107
rect 569 17039 701 17073
rect 569 17005 618 17039
rect 652 17005 701 17039
rect 569 16971 701 17005
rect 569 16937 618 16971
rect 652 16937 701 16971
rect 569 16903 701 16937
rect 569 16869 618 16903
rect 652 16869 701 16903
rect 569 16835 701 16869
rect 569 16801 618 16835
rect 652 16801 701 16835
rect 569 16767 701 16801
rect 569 16733 618 16767
rect 652 16733 701 16767
rect 569 16699 701 16733
rect 569 16665 618 16699
rect 652 16665 701 16699
rect 569 16631 701 16665
rect 569 16597 618 16631
rect 652 16597 701 16631
rect 569 16563 701 16597
rect 569 16529 618 16563
rect 652 16529 701 16563
rect 569 16495 701 16529
rect 569 16461 618 16495
rect 652 16461 701 16495
rect 569 16427 701 16461
rect 569 16393 618 16427
rect 652 16393 701 16427
rect 569 16359 701 16393
rect 569 16325 618 16359
rect 652 16325 701 16359
rect 569 16291 701 16325
rect 569 16257 618 16291
rect 652 16257 701 16291
rect 569 16223 701 16257
rect 569 16189 618 16223
rect 652 16189 701 16223
rect 569 16155 701 16189
rect 569 16121 618 16155
rect 652 16121 701 16155
rect 569 16087 701 16121
rect 569 16053 618 16087
rect 652 16053 701 16087
rect 569 16019 701 16053
rect 569 15985 618 16019
rect 652 15985 701 16019
rect 569 15951 701 15985
rect 569 15917 618 15951
rect 652 15917 701 15951
rect 569 15883 701 15917
rect 569 15849 618 15883
rect 652 15849 701 15883
rect 569 15815 701 15849
rect 569 15781 618 15815
rect 652 15781 701 15815
rect 569 15747 701 15781
rect 569 15713 618 15747
rect 652 15713 701 15747
rect 569 15679 701 15713
rect 569 15645 618 15679
rect 652 15645 701 15679
rect 569 15611 701 15645
rect 569 15577 618 15611
rect 652 15577 701 15611
rect 569 15543 701 15577
rect 569 15509 618 15543
rect 652 15509 701 15543
rect 569 15475 701 15509
rect 569 15441 618 15475
rect 652 15441 701 15475
rect 569 15407 701 15441
rect 569 15373 618 15407
rect 652 15373 701 15407
rect 569 15339 701 15373
rect 569 15305 618 15339
rect 652 15305 701 15339
rect 569 15271 701 15305
rect 569 15237 618 15271
rect 652 15237 701 15271
rect 569 15203 701 15237
rect 569 15169 618 15203
rect 652 15169 701 15203
rect 569 15135 701 15169
rect 569 15101 618 15135
rect 652 15101 701 15135
rect 569 15067 701 15101
rect 569 15033 618 15067
rect 652 15033 701 15067
rect 569 14999 701 15033
rect 569 14965 618 14999
rect 652 14965 701 14999
rect 569 14931 701 14965
rect 569 14897 618 14931
rect 652 14897 701 14931
rect 569 14863 701 14897
rect 569 14829 618 14863
rect 652 14829 701 14863
rect 569 14795 701 14829
rect 569 14761 618 14795
rect 652 14761 701 14795
rect 569 14727 701 14761
rect 569 14693 618 14727
rect 652 14693 701 14727
rect 569 14659 701 14693
rect 569 14625 618 14659
rect 652 14625 701 14659
rect 569 14591 701 14625
rect 569 14557 618 14591
rect 652 14557 701 14591
rect 569 14523 701 14557
rect 569 14489 618 14523
rect 652 14489 701 14523
rect 569 14455 701 14489
rect 569 14421 618 14455
rect 652 14421 701 14455
rect 569 14387 701 14421
rect 569 14353 618 14387
rect 652 14353 701 14387
rect 569 14319 701 14353
rect 569 14285 618 14319
rect 652 14285 701 14319
rect 569 14251 701 14285
rect 569 14217 618 14251
rect 652 14217 701 14251
rect 569 14183 701 14217
rect 569 14149 618 14183
rect 652 14149 701 14183
rect 569 14115 701 14149
rect 569 14081 618 14115
rect 652 14081 701 14115
rect 569 14047 701 14081
rect 569 14013 618 14047
rect 652 14013 701 14047
rect 569 13979 701 14013
rect 569 13945 618 13979
rect 652 13945 701 13979
rect 569 13911 701 13945
rect 569 13877 618 13911
rect 652 13877 701 13911
rect 569 13843 701 13877
rect 569 13809 618 13843
rect 652 13809 701 13843
rect 569 13775 701 13809
rect 569 13741 618 13775
rect 652 13741 701 13775
rect 569 13707 701 13741
rect 569 13673 618 13707
rect 652 13673 701 13707
rect 569 13639 701 13673
rect 569 13605 618 13639
rect 652 13605 701 13639
rect 569 13571 701 13605
rect 569 13537 618 13571
rect 652 13537 701 13571
rect 569 13503 701 13537
rect 569 13469 618 13503
rect 652 13469 701 13503
rect 569 13435 701 13469
rect 569 13401 618 13435
rect 652 13401 701 13435
rect 569 13367 701 13401
rect 569 13333 618 13367
rect 652 13333 701 13367
rect 569 13299 701 13333
rect 569 13265 618 13299
rect 652 13265 701 13299
rect 569 13231 701 13265
rect 569 13197 618 13231
rect 652 13197 701 13231
rect 569 13163 701 13197
rect 569 13129 618 13163
rect 652 13129 701 13163
rect 569 13095 701 13129
rect 569 13061 618 13095
rect 652 13061 701 13095
rect 569 13027 701 13061
rect 569 12993 618 13027
rect 652 12993 701 13027
rect 569 12959 701 12993
rect 569 12925 618 12959
rect 652 12925 701 12959
rect 569 12891 701 12925
rect 569 12857 618 12891
rect 652 12857 701 12891
rect 569 12823 701 12857
rect 569 12789 618 12823
rect 652 12789 701 12823
rect 569 12755 701 12789
rect 569 12721 618 12755
rect 652 12721 701 12755
rect 569 12687 701 12721
rect 569 12653 618 12687
rect 652 12653 701 12687
rect 569 12619 701 12653
rect 569 12585 618 12619
rect 652 12585 701 12619
rect 569 12551 701 12585
rect 569 12517 618 12551
rect 652 12517 701 12551
rect 569 12483 701 12517
rect 569 12449 618 12483
rect 652 12449 701 12483
rect 569 12415 701 12449
rect 569 12381 618 12415
rect 652 12381 701 12415
rect 569 12347 701 12381
rect 569 12313 618 12347
rect 652 12313 701 12347
rect 569 12279 701 12313
rect 569 12245 618 12279
rect 652 12245 701 12279
rect 569 12211 701 12245
rect 569 12177 618 12211
rect 652 12177 701 12211
rect 569 12143 701 12177
rect 569 12109 618 12143
rect 652 12109 701 12143
rect 569 12075 701 12109
rect 569 12041 618 12075
rect 652 12041 701 12075
rect 569 12007 701 12041
rect 569 11973 618 12007
rect 652 11973 701 12007
rect 569 11939 701 11973
rect 569 11905 618 11939
rect 652 11905 701 11939
rect 569 11871 701 11905
rect 569 11837 618 11871
rect 652 11837 701 11871
rect 569 11803 701 11837
rect 569 11769 618 11803
rect 652 11769 701 11803
rect 569 11735 701 11769
rect 569 11701 618 11735
rect 652 11701 701 11735
rect 569 11667 701 11701
rect 569 11633 618 11667
rect 652 11633 701 11667
rect 569 11599 701 11633
rect 569 11565 618 11599
rect 652 11565 701 11599
rect 569 11531 701 11565
rect 569 11497 618 11531
rect 652 11497 701 11531
rect 569 11463 701 11497
rect 569 11429 618 11463
rect 652 11429 701 11463
rect 569 11395 701 11429
rect 569 11361 618 11395
rect 652 11361 701 11395
rect 569 11327 701 11361
rect 569 11293 618 11327
rect 652 11293 701 11327
rect 569 11259 701 11293
rect 569 11225 618 11259
rect 652 11225 701 11259
rect 569 11191 701 11225
rect 569 11157 618 11191
rect 652 11157 701 11191
rect 569 11123 701 11157
rect 569 11089 618 11123
rect 652 11089 701 11123
rect 569 11055 701 11089
rect 569 11021 618 11055
rect 652 11021 701 11055
rect 569 10987 701 11021
rect 569 10953 618 10987
rect 652 10953 701 10987
rect 569 10919 701 10953
rect 569 10885 618 10919
rect 652 10885 701 10919
rect 569 10851 701 10885
rect 569 10817 618 10851
rect 652 10817 701 10851
rect 569 10783 701 10817
rect 569 10749 618 10783
rect 652 10749 701 10783
rect 569 10715 701 10749
rect 569 10681 618 10715
rect 652 10681 701 10715
rect 569 10647 701 10681
rect 569 10613 618 10647
rect 652 10613 701 10647
rect 569 10579 701 10613
rect 569 10545 618 10579
rect 652 10545 701 10579
rect 569 10511 701 10545
rect 569 10477 618 10511
rect 652 10477 701 10511
rect 569 10443 701 10477
rect 569 10409 618 10443
rect 652 10409 701 10443
rect 569 10375 701 10409
rect 569 10341 618 10375
rect 652 10341 701 10375
rect 569 10307 701 10341
rect 569 10273 618 10307
rect 652 10273 701 10307
rect 569 10239 701 10273
rect 569 10205 618 10239
rect 652 10205 701 10239
rect 569 10171 701 10205
rect 569 10137 618 10171
rect 652 10137 701 10171
rect 569 10103 701 10137
rect 569 10069 618 10103
rect 652 10069 701 10103
rect 569 10035 701 10069
rect 569 10001 618 10035
rect 652 10001 701 10035
rect 569 9967 701 10001
rect 569 9933 618 9967
rect 652 9933 701 9967
rect 569 9899 701 9933
rect 569 9865 618 9899
rect 652 9865 701 9899
rect 569 9831 701 9865
rect 569 9797 618 9831
rect 652 9797 701 9831
rect 569 9769 701 9797
rect 14303 36079 14437 36107
rect 14303 36045 14353 36079
rect 14387 36045 14437 36079
rect 14303 36011 14437 36045
rect 14303 35977 14353 36011
rect 14387 35977 14437 36011
rect 14303 35943 14437 35977
rect 14303 35909 14353 35943
rect 14387 35909 14437 35943
rect 14303 35875 14437 35909
rect 14303 35841 14353 35875
rect 14387 35841 14437 35875
rect 14303 35807 14437 35841
rect 14303 35773 14353 35807
rect 14387 35773 14437 35807
rect 14303 35739 14437 35773
rect 14303 35705 14353 35739
rect 14387 35705 14437 35739
rect 14303 35671 14437 35705
rect 14303 35637 14353 35671
rect 14387 35637 14437 35671
rect 14303 35603 14437 35637
rect 14303 35569 14353 35603
rect 14387 35569 14437 35603
rect 14303 35535 14437 35569
rect 14303 35501 14353 35535
rect 14387 35501 14437 35535
rect 14303 35467 14437 35501
rect 14303 35433 14353 35467
rect 14387 35433 14437 35467
rect 14303 35399 14437 35433
rect 14303 35365 14353 35399
rect 14387 35365 14437 35399
rect 14303 35331 14437 35365
rect 14303 35297 14353 35331
rect 14387 35297 14437 35331
rect 14303 35263 14437 35297
rect 14303 35229 14353 35263
rect 14387 35229 14437 35263
rect 14303 35195 14437 35229
rect 14303 35161 14353 35195
rect 14387 35161 14437 35195
rect 14303 35127 14437 35161
rect 14303 35093 14353 35127
rect 14387 35093 14437 35127
rect 14303 35059 14437 35093
rect 14303 35025 14353 35059
rect 14387 35025 14437 35059
rect 14303 34991 14437 35025
rect 14303 34957 14353 34991
rect 14387 34957 14437 34991
rect 14303 34923 14437 34957
rect 14303 34889 14353 34923
rect 14387 34889 14437 34923
rect 14303 34855 14437 34889
rect 14303 34821 14353 34855
rect 14387 34821 14437 34855
rect 14303 34787 14437 34821
rect 14303 34753 14353 34787
rect 14387 34753 14437 34787
rect 14303 34719 14437 34753
rect 14303 34685 14353 34719
rect 14387 34685 14437 34719
rect 14303 34651 14437 34685
rect 14303 34617 14353 34651
rect 14387 34617 14437 34651
rect 14303 34583 14437 34617
rect 14303 34549 14353 34583
rect 14387 34549 14437 34583
rect 14303 34515 14437 34549
rect 14303 34481 14353 34515
rect 14387 34481 14437 34515
rect 14303 34447 14437 34481
rect 14303 34413 14353 34447
rect 14387 34413 14437 34447
rect 14303 34379 14437 34413
rect 14303 34345 14353 34379
rect 14387 34345 14437 34379
rect 14303 34311 14437 34345
rect 14303 34277 14353 34311
rect 14387 34277 14437 34311
rect 14303 34243 14437 34277
rect 14303 34209 14353 34243
rect 14387 34209 14437 34243
rect 14303 34175 14437 34209
rect 14303 34141 14353 34175
rect 14387 34141 14437 34175
rect 14303 34107 14437 34141
rect 14303 34073 14353 34107
rect 14387 34073 14437 34107
rect 14303 34039 14437 34073
rect 14303 34005 14353 34039
rect 14387 34005 14437 34039
rect 14303 33971 14437 34005
rect 14303 33937 14353 33971
rect 14387 33937 14437 33971
rect 14303 33903 14437 33937
rect 14303 33869 14353 33903
rect 14387 33869 14437 33903
rect 14303 33835 14437 33869
rect 14303 33801 14353 33835
rect 14387 33801 14437 33835
rect 14303 33767 14437 33801
rect 14303 33733 14353 33767
rect 14387 33733 14437 33767
rect 14303 33699 14437 33733
rect 14303 33665 14353 33699
rect 14387 33665 14437 33699
rect 14303 33631 14437 33665
rect 14303 33597 14353 33631
rect 14387 33597 14437 33631
rect 14303 33563 14437 33597
rect 14303 33529 14353 33563
rect 14387 33529 14437 33563
rect 14303 33495 14437 33529
rect 14303 33461 14353 33495
rect 14387 33461 14437 33495
rect 14303 33427 14437 33461
rect 14303 33393 14353 33427
rect 14387 33393 14437 33427
rect 14303 33359 14437 33393
rect 14303 33325 14353 33359
rect 14387 33325 14437 33359
rect 14303 33291 14437 33325
rect 14303 33257 14353 33291
rect 14387 33257 14437 33291
rect 14303 33223 14437 33257
rect 14303 33189 14353 33223
rect 14387 33189 14437 33223
rect 14303 33155 14437 33189
rect 14303 33121 14353 33155
rect 14387 33121 14437 33155
rect 14303 33087 14437 33121
rect 14303 33053 14353 33087
rect 14387 33053 14437 33087
rect 14303 33019 14437 33053
rect 14303 32985 14353 33019
rect 14387 32985 14437 33019
rect 14303 32951 14437 32985
rect 14303 32917 14353 32951
rect 14387 32917 14437 32951
rect 14303 32883 14437 32917
rect 14303 32849 14353 32883
rect 14387 32849 14437 32883
rect 14303 32815 14437 32849
rect 14303 32781 14353 32815
rect 14387 32781 14437 32815
rect 14303 32747 14437 32781
rect 14303 32713 14353 32747
rect 14387 32713 14437 32747
rect 14303 32679 14437 32713
rect 14303 32645 14353 32679
rect 14387 32645 14437 32679
rect 14303 32611 14437 32645
rect 14303 32577 14353 32611
rect 14387 32577 14437 32611
rect 14303 32543 14437 32577
rect 14303 32509 14353 32543
rect 14387 32509 14437 32543
rect 14303 32475 14437 32509
rect 14303 32441 14353 32475
rect 14387 32441 14437 32475
rect 14303 32407 14437 32441
rect 14303 32373 14353 32407
rect 14387 32373 14437 32407
rect 14303 32339 14437 32373
rect 14303 32305 14353 32339
rect 14387 32305 14437 32339
rect 14303 32271 14437 32305
rect 14303 32237 14353 32271
rect 14387 32237 14437 32271
rect 14303 32203 14437 32237
rect 14303 32169 14353 32203
rect 14387 32169 14437 32203
rect 14303 32135 14437 32169
rect 14303 32101 14353 32135
rect 14387 32101 14437 32135
rect 14303 32067 14437 32101
rect 14303 32033 14353 32067
rect 14387 32033 14437 32067
rect 14303 31999 14437 32033
rect 14303 31965 14353 31999
rect 14387 31965 14437 31999
rect 14303 31931 14437 31965
rect 14303 31897 14353 31931
rect 14387 31897 14437 31931
rect 14303 31863 14437 31897
rect 14303 31829 14353 31863
rect 14387 31829 14437 31863
rect 14303 31795 14437 31829
rect 14303 31761 14353 31795
rect 14387 31761 14437 31795
rect 14303 31727 14437 31761
rect 14303 31693 14353 31727
rect 14387 31693 14437 31727
rect 14303 31659 14437 31693
rect 14303 31625 14353 31659
rect 14387 31625 14437 31659
rect 14303 31591 14437 31625
rect 14303 31557 14353 31591
rect 14387 31557 14437 31591
rect 14303 31523 14437 31557
rect 14303 31489 14353 31523
rect 14387 31489 14437 31523
rect 14303 31455 14437 31489
rect 14303 31421 14353 31455
rect 14387 31421 14437 31455
rect 14303 31387 14437 31421
rect 14303 31353 14353 31387
rect 14387 31353 14437 31387
rect 14303 31319 14437 31353
rect 14303 31285 14353 31319
rect 14387 31285 14437 31319
rect 14303 31251 14437 31285
rect 14303 31217 14353 31251
rect 14387 31217 14437 31251
rect 14303 31183 14437 31217
rect 14303 31149 14353 31183
rect 14387 31149 14437 31183
rect 14303 31115 14437 31149
rect 14303 31081 14353 31115
rect 14387 31081 14437 31115
rect 14303 31047 14437 31081
rect 14303 31013 14353 31047
rect 14387 31013 14437 31047
rect 14303 30979 14437 31013
rect 14303 30945 14353 30979
rect 14387 30945 14437 30979
rect 14303 30911 14437 30945
rect 14303 30877 14353 30911
rect 14387 30877 14437 30911
rect 14303 30843 14437 30877
rect 14303 30809 14353 30843
rect 14387 30809 14437 30843
rect 14303 30775 14437 30809
rect 14303 30741 14353 30775
rect 14387 30741 14437 30775
rect 14303 30707 14437 30741
rect 14303 30673 14353 30707
rect 14387 30673 14437 30707
rect 14303 30639 14437 30673
rect 14303 30605 14353 30639
rect 14387 30605 14437 30639
rect 14303 30571 14437 30605
rect 14303 30537 14353 30571
rect 14387 30537 14437 30571
rect 14303 30503 14437 30537
rect 14303 30469 14353 30503
rect 14387 30469 14437 30503
rect 14303 30435 14437 30469
rect 14303 30401 14353 30435
rect 14387 30401 14437 30435
rect 14303 30367 14437 30401
rect 14303 30333 14353 30367
rect 14387 30333 14437 30367
rect 14303 30299 14437 30333
rect 14303 30265 14353 30299
rect 14387 30265 14437 30299
rect 14303 30231 14437 30265
rect 14303 30197 14353 30231
rect 14387 30197 14437 30231
rect 14303 30163 14437 30197
rect 14303 30129 14353 30163
rect 14387 30129 14437 30163
rect 14303 30095 14437 30129
rect 14303 30061 14353 30095
rect 14387 30061 14437 30095
rect 14303 30027 14437 30061
rect 14303 29993 14353 30027
rect 14387 29993 14437 30027
rect 14303 29959 14437 29993
rect 14303 29925 14353 29959
rect 14387 29925 14437 29959
rect 14303 29891 14437 29925
rect 14303 29857 14353 29891
rect 14387 29857 14437 29891
rect 14303 29823 14437 29857
rect 14303 29789 14353 29823
rect 14387 29789 14437 29823
rect 14303 29755 14437 29789
rect 14303 29721 14353 29755
rect 14387 29721 14437 29755
rect 14303 29687 14437 29721
rect 14303 29653 14353 29687
rect 14387 29653 14437 29687
rect 14303 29619 14437 29653
rect 14303 29585 14353 29619
rect 14387 29585 14437 29619
rect 14303 29551 14437 29585
rect 14303 29517 14353 29551
rect 14387 29517 14437 29551
rect 14303 29483 14437 29517
rect 14303 29449 14353 29483
rect 14387 29449 14437 29483
rect 14303 29415 14437 29449
rect 14303 29381 14353 29415
rect 14387 29381 14437 29415
rect 14303 29347 14437 29381
rect 14303 29313 14353 29347
rect 14387 29313 14437 29347
rect 14303 29279 14437 29313
rect 14303 29245 14353 29279
rect 14387 29245 14437 29279
rect 14303 29211 14437 29245
rect 14303 29177 14353 29211
rect 14387 29177 14437 29211
rect 14303 29143 14437 29177
rect 14303 29109 14353 29143
rect 14387 29109 14437 29143
rect 14303 29075 14437 29109
rect 14303 29041 14353 29075
rect 14387 29041 14437 29075
rect 14303 29007 14437 29041
rect 14303 28973 14353 29007
rect 14387 28973 14437 29007
rect 14303 28939 14437 28973
rect 14303 28905 14353 28939
rect 14387 28905 14437 28939
rect 14303 28871 14437 28905
rect 14303 28837 14353 28871
rect 14387 28837 14437 28871
rect 14303 28803 14437 28837
rect 14303 28769 14353 28803
rect 14387 28769 14437 28803
rect 14303 28735 14437 28769
rect 14303 28701 14353 28735
rect 14387 28701 14437 28735
rect 14303 28667 14437 28701
rect 14303 28633 14353 28667
rect 14387 28633 14437 28667
rect 14303 28599 14437 28633
rect 14303 28565 14353 28599
rect 14387 28565 14437 28599
rect 14303 28531 14437 28565
rect 14303 28497 14353 28531
rect 14387 28497 14437 28531
rect 14303 28463 14437 28497
rect 14303 28429 14353 28463
rect 14387 28429 14437 28463
rect 14303 28395 14437 28429
rect 14303 28361 14353 28395
rect 14387 28361 14437 28395
rect 14303 28327 14437 28361
rect 14303 28293 14353 28327
rect 14387 28293 14437 28327
rect 14303 28259 14437 28293
rect 14303 28225 14353 28259
rect 14387 28225 14437 28259
rect 14303 28191 14437 28225
rect 14303 28157 14353 28191
rect 14387 28157 14437 28191
rect 14303 28123 14437 28157
rect 14303 28089 14353 28123
rect 14387 28089 14437 28123
rect 14303 28055 14437 28089
rect 14303 28021 14353 28055
rect 14387 28021 14437 28055
rect 14303 27987 14437 28021
rect 14303 27953 14353 27987
rect 14387 27953 14437 27987
rect 14303 27919 14437 27953
rect 14303 27885 14353 27919
rect 14387 27885 14437 27919
rect 14303 27851 14437 27885
rect 14303 27817 14353 27851
rect 14387 27817 14437 27851
rect 14303 27783 14437 27817
rect 14303 27749 14353 27783
rect 14387 27749 14437 27783
rect 14303 27715 14437 27749
rect 14303 27681 14353 27715
rect 14387 27681 14437 27715
rect 14303 27647 14437 27681
rect 14303 27613 14353 27647
rect 14387 27613 14437 27647
rect 14303 27579 14437 27613
rect 14303 27545 14353 27579
rect 14387 27545 14437 27579
rect 14303 27511 14437 27545
rect 14303 27477 14353 27511
rect 14387 27477 14437 27511
rect 14303 27443 14437 27477
rect 14303 27409 14353 27443
rect 14387 27409 14437 27443
rect 14303 27375 14437 27409
rect 14303 27341 14353 27375
rect 14387 27341 14437 27375
rect 14303 27307 14437 27341
rect 14303 27273 14353 27307
rect 14387 27273 14437 27307
rect 14303 27239 14437 27273
rect 14303 27205 14353 27239
rect 14387 27205 14437 27239
rect 14303 27171 14437 27205
rect 14303 27137 14353 27171
rect 14387 27137 14437 27171
rect 14303 27103 14437 27137
rect 14303 27069 14353 27103
rect 14387 27069 14437 27103
rect 14303 27035 14437 27069
rect 14303 27001 14353 27035
rect 14387 27001 14437 27035
rect 14303 26967 14437 27001
rect 14303 26933 14353 26967
rect 14387 26933 14437 26967
rect 14303 26899 14437 26933
rect 14303 26865 14353 26899
rect 14387 26865 14437 26899
rect 14303 26831 14437 26865
rect 14303 26797 14353 26831
rect 14387 26797 14437 26831
rect 14303 26763 14437 26797
rect 14303 26729 14353 26763
rect 14387 26729 14437 26763
rect 14303 26695 14437 26729
rect 14303 26661 14353 26695
rect 14387 26661 14437 26695
rect 14303 26627 14437 26661
rect 14303 26593 14353 26627
rect 14387 26593 14437 26627
rect 14303 26559 14437 26593
rect 14303 26525 14353 26559
rect 14387 26525 14437 26559
rect 14303 26491 14437 26525
rect 14303 26457 14353 26491
rect 14387 26457 14437 26491
rect 14303 26423 14437 26457
rect 14303 26389 14353 26423
rect 14387 26389 14437 26423
rect 14303 26355 14437 26389
rect 14303 26321 14353 26355
rect 14387 26321 14437 26355
rect 14303 26287 14437 26321
rect 14303 26253 14353 26287
rect 14387 26253 14437 26287
rect 14303 26219 14437 26253
rect 14303 26185 14353 26219
rect 14387 26185 14437 26219
rect 14303 26151 14437 26185
rect 14303 26117 14353 26151
rect 14387 26117 14437 26151
rect 14303 26083 14437 26117
rect 14303 26049 14353 26083
rect 14387 26049 14437 26083
rect 14303 26015 14437 26049
rect 14303 25981 14353 26015
rect 14387 25981 14437 26015
rect 14303 25947 14437 25981
rect 14303 25913 14353 25947
rect 14387 25913 14437 25947
rect 14303 25879 14437 25913
rect 14303 25845 14353 25879
rect 14387 25845 14437 25879
rect 14303 25811 14437 25845
rect 14303 25777 14353 25811
rect 14387 25777 14437 25811
rect 14303 25743 14437 25777
rect 14303 25709 14353 25743
rect 14387 25709 14437 25743
rect 14303 25675 14437 25709
rect 14303 25641 14353 25675
rect 14387 25641 14437 25675
rect 14303 25607 14437 25641
rect 14303 25573 14353 25607
rect 14387 25573 14437 25607
rect 14303 25539 14437 25573
rect 14303 25505 14353 25539
rect 14387 25505 14437 25539
rect 14303 25471 14437 25505
rect 14303 25437 14353 25471
rect 14387 25437 14437 25471
rect 14303 25403 14437 25437
rect 14303 25369 14353 25403
rect 14387 25369 14437 25403
rect 14303 25335 14437 25369
rect 14303 25301 14353 25335
rect 14387 25301 14437 25335
rect 14303 25267 14437 25301
rect 14303 25233 14353 25267
rect 14387 25233 14437 25267
rect 14303 25199 14437 25233
rect 14303 25165 14353 25199
rect 14387 25165 14437 25199
rect 14303 25131 14437 25165
rect 14303 25097 14353 25131
rect 14387 25097 14437 25131
rect 14303 25063 14437 25097
rect 14303 25029 14353 25063
rect 14387 25029 14437 25063
rect 14303 24995 14437 25029
rect 14303 24961 14353 24995
rect 14387 24961 14437 24995
rect 14303 24927 14437 24961
rect 14303 24893 14353 24927
rect 14387 24893 14437 24927
rect 14303 24859 14437 24893
rect 14303 24825 14353 24859
rect 14387 24825 14437 24859
rect 14303 24791 14437 24825
rect 14303 24757 14353 24791
rect 14387 24757 14437 24791
rect 14303 24723 14437 24757
rect 14303 24689 14353 24723
rect 14387 24689 14437 24723
rect 14303 24655 14437 24689
rect 14303 24621 14353 24655
rect 14387 24621 14437 24655
rect 14303 24587 14437 24621
rect 14303 24553 14353 24587
rect 14387 24553 14437 24587
rect 14303 24519 14437 24553
rect 14303 24485 14353 24519
rect 14387 24485 14437 24519
rect 14303 24451 14437 24485
rect 14303 24417 14353 24451
rect 14387 24417 14437 24451
rect 14303 24383 14437 24417
rect 14303 24349 14353 24383
rect 14387 24349 14437 24383
rect 14303 24315 14437 24349
rect 14303 24281 14353 24315
rect 14387 24281 14437 24315
rect 14303 24247 14437 24281
rect 14303 24213 14353 24247
rect 14387 24213 14437 24247
rect 14303 24179 14437 24213
rect 14303 24145 14353 24179
rect 14387 24145 14437 24179
rect 14303 24111 14437 24145
rect 14303 24077 14353 24111
rect 14387 24077 14437 24111
rect 14303 24043 14437 24077
rect 14303 24009 14353 24043
rect 14387 24009 14437 24043
rect 14303 23975 14437 24009
rect 14303 23941 14353 23975
rect 14387 23941 14437 23975
rect 14303 23907 14437 23941
rect 14303 23873 14353 23907
rect 14387 23873 14437 23907
rect 14303 23839 14437 23873
rect 14303 23805 14353 23839
rect 14387 23805 14437 23839
rect 14303 23771 14437 23805
rect 14303 23737 14353 23771
rect 14387 23737 14437 23771
rect 14303 23703 14437 23737
rect 14303 23669 14353 23703
rect 14387 23669 14437 23703
rect 14303 23635 14437 23669
rect 14303 23601 14353 23635
rect 14387 23601 14437 23635
rect 14303 23567 14437 23601
rect 14303 23533 14353 23567
rect 14387 23533 14437 23567
rect 14303 23499 14437 23533
rect 14303 23465 14353 23499
rect 14387 23465 14437 23499
rect 14303 23431 14437 23465
rect 14303 23397 14353 23431
rect 14387 23397 14437 23431
rect 14303 23363 14437 23397
rect 14303 23329 14353 23363
rect 14387 23329 14437 23363
rect 14303 23295 14437 23329
rect 14303 23261 14353 23295
rect 14387 23261 14437 23295
rect 14303 23227 14437 23261
rect 14303 23193 14353 23227
rect 14387 23193 14437 23227
rect 14303 23159 14437 23193
rect 14303 23125 14353 23159
rect 14387 23125 14437 23159
rect 14303 23091 14437 23125
rect 14303 23057 14353 23091
rect 14387 23057 14437 23091
rect 14303 23023 14437 23057
rect 14303 22989 14353 23023
rect 14387 22989 14437 23023
rect 14303 22955 14437 22989
rect 14303 22921 14353 22955
rect 14387 22921 14437 22955
rect 14303 22887 14437 22921
rect 14303 22853 14353 22887
rect 14387 22853 14437 22887
rect 14303 22819 14437 22853
rect 14303 22785 14353 22819
rect 14387 22785 14437 22819
rect 14303 22751 14437 22785
rect 14303 22717 14353 22751
rect 14387 22717 14437 22751
rect 14303 22683 14437 22717
rect 14303 22649 14353 22683
rect 14387 22649 14437 22683
rect 14303 22615 14437 22649
rect 14303 22581 14353 22615
rect 14387 22581 14437 22615
rect 14303 22547 14437 22581
rect 14303 22513 14353 22547
rect 14387 22513 14437 22547
rect 14303 22479 14437 22513
rect 14303 22445 14353 22479
rect 14387 22445 14437 22479
rect 14303 22411 14437 22445
rect 14303 22377 14353 22411
rect 14387 22377 14437 22411
rect 14303 22343 14437 22377
rect 14303 22309 14353 22343
rect 14387 22309 14437 22343
rect 14303 22275 14437 22309
rect 14303 22241 14353 22275
rect 14387 22241 14437 22275
rect 14303 22207 14437 22241
rect 14303 22173 14353 22207
rect 14387 22173 14437 22207
rect 14303 22139 14437 22173
rect 14303 22105 14353 22139
rect 14387 22105 14437 22139
rect 14303 22071 14437 22105
rect 14303 22037 14353 22071
rect 14387 22037 14437 22071
rect 14303 22003 14437 22037
rect 14303 21969 14353 22003
rect 14387 21969 14437 22003
rect 14303 21935 14437 21969
rect 14303 21901 14353 21935
rect 14387 21901 14437 21935
rect 14303 21867 14437 21901
rect 14303 21833 14353 21867
rect 14387 21833 14437 21867
rect 14303 21799 14437 21833
rect 14303 21765 14353 21799
rect 14387 21765 14437 21799
rect 14303 21731 14437 21765
rect 14303 21697 14353 21731
rect 14387 21697 14437 21731
rect 14303 21663 14437 21697
rect 14303 21629 14353 21663
rect 14387 21629 14437 21663
rect 14303 21595 14437 21629
rect 14303 21561 14353 21595
rect 14387 21561 14437 21595
rect 14303 21527 14437 21561
rect 14303 21493 14353 21527
rect 14387 21493 14437 21527
rect 14303 21459 14437 21493
rect 14303 21425 14353 21459
rect 14387 21425 14437 21459
rect 14303 21391 14437 21425
rect 14303 21357 14353 21391
rect 14387 21357 14437 21391
rect 14303 21323 14437 21357
rect 14303 21289 14353 21323
rect 14387 21289 14437 21323
rect 14303 21255 14437 21289
rect 14303 21221 14353 21255
rect 14387 21221 14437 21255
rect 14303 21187 14437 21221
rect 14303 21153 14353 21187
rect 14387 21153 14437 21187
rect 14303 21119 14437 21153
rect 14303 21085 14353 21119
rect 14387 21085 14437 21119
rect 14303 21051 14437 21085
rect 14303 21017 14353 21051
rect 14387 21017 14437 21051
rect 14303 20983 14437 21017
rect 14303 20949 14353 20983
rect 14387 20949 14437 20983
rect 14303 20915 14437 20949
rect 14303 20881 14353 20915
rect 14387 20881 14437 20915
rect 14303 20847 14437 20881
rect 14303 20813 14353 20847
rect 14387 20813 14437 20847
rect 14303 20779 14437 20813
rect 14303 20745 14353 20779
rect 14387 20745 14437 20779
rect 14303 20711 14437 20745
rect 14303 20677 14353 20711
rect 14387 20677 14437 20711
rect 14303 20643 14437 20677
rect 14303 20609 14353 20643
rect 14387 20609 14437 20643
rect 14303 20575 14437 20609
rect 14303 20541 14353 20575
rect 14387 20541 14437 20575
rect 14303 20507 14437 20541
rect 14303 20473 14353 20507
rect 14387 20473 14437 20507
rect 14303 20439 14437 20473
rect 14303 20405 14353 20439
rect 14387 20405 14437 20439
rect 14303 20371 14437 20405
rect 14303 20337 14353 20371
rect 14387 20337 14437 20371
rect 14303 20303 14437 20337
rect 14303 20269 14353 20303
rect 14387 20269 14437 20303
rect 14303 20235 14437 20269
rect 14303 20201 14353 20235
rect 14387 20201 14437 20235
rect 14303 20167 14437 20201
rect 14303 20133 14353 20167
rect 14387 20133 14437 20167
rect 14303 20099 14437 20133
rect 14303 20065 14353 20099
rect 14387 20065 14437 20099
rect 14303 20031 14437 20065
rect 14303 19997 14353 20031
rect 14387 19997 14437 20031
rect 14303 19963 14437 19997
rect 14303 19929 14353 19963
rect 14387 19929 14437 19963
rect 14303 19895 14437 19929
rect 14303 19861 14353 19895
rect 14387 19861 14437 19895
rect 14303 19827 14437 19861
rect 14303 19793 14353 19827
rect 14387 19793 14437 19827
rect 14303 19759 14437 19793
rect 14303 19725 14353 19759
rect 14387 19725 14437 19759
rect 14303 19691 14437 19725
rect 14303 19657 14353 19691
rect 14387 19657 14437 19691
rect 14303 19623 14437 19657
rect 14303 19589 14353 19623
rect 14387 19589 14437 19623
rect 14303 19555 14437 19589
rect 14303 19521 14353 19555
rect 14387 19521 14437 19555
rect 14303 19487 14437 19521
rect 14303 19453 14353 19487
rect 14387 19453 14437 19487
rect 14303 19419 14437 19453
rect 14303 19385 14353 19419
rect 14387 19385 14437 19419
rect 14303 19351 14437 19385
rect 14303 19317 14353 19351
rect 14387 19317 14437 19351
rect 14303 19283 14437 19317
rect 14303 19249 14353 19283
rect 14387 19249 14437 19283
rect 14303 19215 14437 19249
rect 14303 19181 14353 19215
rect 14387 19181 14437 19215
rect 14303 19147 14437 19181
rect 14303 19113 14353 19147
rect 14387 19113 14437 19147
rect 14303 19079 14437 19113
rect 14303 19045 14353 19079
rect 14387 19045 14437 19079
rect 14303 19011 14437 19045
rect 14303 18977 14353 19011
rect 14387 18977 14437 19011
rect 14303 18943 14437 18977
rect 14303 18909 14353 18943
rect 14387 18909 14437 18943
rect 14303 18875 14437 18909
rect 14303 18841 14353 18875
rect 14387 18841 14437 18875
rect 14303 18807 14437 18841
rect 14303 18773 14353 18807
rect 14387 18773 14437 18807
rect 14303 18739 14437 18773
rect 14303 18705 14353 18739
rect 14387 18705 14437 18739
rect 14303 18671 14437 18705
rect 14303 18637 14353 18671
rect 14387 18637 14437 18671
rect 14303 18603 14437 18637
rect 14303 18569 14353 18603
rect 14387 18569 14437 18603
rect 14303 18535 14437 18569
rect 14303 18501 14353 18535
rect 14387 18501 14437 18535
rect 14303 18467 14437 18501
rect 14303 18433 14353 18467
rect 14387 18433 14437 18467
rect 14303 18399 14437 18433
rect 14303 18365 14353 18399
rect 14387 18365 14437 18399
rect 14303 18331 14437 18365
rect 14303 18297 14353 18331
rect 14387 18297 14437 18331
rect 14303 18263 14437 18297
rect 14303 18229 14353 18263
rect 14387 18229 14437 18263
rect 14303 18195 14437 18229
rect 14303 18161 14353 18195
rect 14387 18161 14437 18195
rect 14303 18127 14437 18161
rect 14303 18093 14353 18127
rect 14387 18093 14437 18127
rect 14303 18059 14437 18093
rect 14303 18025 14353 18059
rect 14387 18025 14437 18059
rect 14303 17991 14437 18025
rect 14303 17957 14353 17991
rect 14387 17957 14437 17991
rect 14303 17923 14437 17957
rect 14303 17889 14353 17923
rect 14387 17889 14437 17923
rect 14303 17855 14437 17889
rect 14303 17821 14353 17855
rect 14387 17821 14437 17855
rect 14303 17787 14437 17821
rect 14303 17753 14353 17787
rect 14387 17753 14437 17787
rect 14303 17719 14437 17753
rect 14303 17685 14353 17719
rect 14387 17685 14437 17719
rect 14303 17651 14437 17685
rect 14303 17617 14353 17651
rect 14387 17617 14437 17651
rect 14303 17583 14437 17617
rect 14303 17549 14353 17583
rect 14387 17549 14437 17583
rect 14303 17515 14437 17549
rect 14303 17481 14353 17515
rect 14387 17481 14437 17515
rect 14303 17447 14437 17481
rect 14303 17413 14353 17447
rect 14387 17413 14437 17447
rect 14303 17379 14437 17413
rect 14303 17345 14353 17379
rect 14387 17345 14437 17379
rect 14303 17311 14437 17345
rect 14303 17277 14353 17311
rect 14387 17277 14437 17311
rect 14303 17243 14437 17277
rect 14303 17209 14353 17243
rect 14387 17209 14437 17243
rect 14303 17175 14437 17209
rect 14303 17141 14353 17175
rect 14387 17141 14437 17175
rect 14303 17107 14437 17141
rect 14303 17073 14353 17107
rect 14387 17073 14437 17107
rect 14303 17039 14437 17073
rect 14303 17005 14353 17039
rect 14387 17005 14437 17039
rect 14303 16971 14437 17005
rect 14303 16937 14353 16971
rect 14387 16937 14437 16971
rect 14303 16903 14437 16937
rect 14303 16869 14353 16903
rect 14387 16869 14437 16903
rect 14303 16835 14437 16869
rect 14303 16801 14353 16835
rect 14387 16801 14437 16835
rect 14303 16767 14437 16801
rect 14303 16733 14353 16767
rect 14387 16733 14437 16767
rect 14303 16699 14437 16733
rect 14303 16665 14353 16699
rect 14387 16665 14437 16699
rect 14303 16631 14437 16665
rect 14303 16597 14353 16631
rect 14387 16597 14437 16631
rect 14303 16563 14437 16597
rect 14303 16529 14353 16563
rect 14387 16529 14437 16563
rect 14303 16495 14437 16529
rect 14303 16461 14353 16495
rect 14387 16461 14437 16495
rect 14303 16427 14437 16461
rect 14303 16393 14353 16427
rect 14387 16393 14437 16427
rect 14303 16359 14437 16393
rect 14303 16325 14353 16359
rect 14387 16325 14437 16359
rect 14303 16291 14437 16325
rect 14303 16257 14353 16291
rect 14387 16257 14437 16291
rect 14303 16223 14437 16257
rect 14303 16189 14353 16223
rect 14387 16189 14437 16223
rect 14303 16155 14437 16189
rect 14303 16121 14353 16155
rect 14387 16121 14437 16155
rect 14303 16087 14437 16121
rect 14303 16053 14353 16087
rect 14387 16053 14437 16087
rect 14303 16019 14437 16053
rect 14303 15985 14353 16019
rect 14387 15985 14437 16019
rect 14303 15951 14437 15985
rect 14303 15917 14353 15951
rect 14387 15917 14437 15951
rect 14303 15883 14437 15917
rect 14303 15849 14353 15883
rect 14387 15849 14437 15883
rect 14303 15815 14437 15849
rect 14303 15781 14353 15815
rect 14387 15781 14437 15815
rect 14303 15747 14437 15781
rect 14303 15713 14353 15747
rect 14387 15713 14437 15747
rect 14303 15679 14437 15713
rect 14303 15645 14353 15679
rect 14387 15645 14437 15679
rect 14303 15611 14437 15645
rect 14303 15577 14353 15611
rect 14387 15577 14437 15611
rect 14303 15543 14437 15577
rect 14303 15509 14353 15543
rect 14387 15509 14437 15543
rect 14303 15475 14437 15509
rect 14303 15441 14353 15475
rect 14387 15441 14437 15475
rect 14303 15407 14437 15441
rect 14303 15373 14353 15407
rect 14387 15373 14437 15407
rect 14303 15339 14437 15373
rect 14303 15305 14353 15339
rect 14387 15305 14437 15339
rect 14303 15271 14437 15305
rect 14303 15237 14353 15271
rect 14387 15237 14437 15271
rect 14303 15203 14437 15237
rect 14303 15169 14353 15203
rect 14387 15169 14437 15203
rect 14303 15135 14437 15169
rect 14303 15101 14353 15135
rect 14387 15101 14437 15135
rect 14303 15067 14437 15101
rect 14303 15033 14353 15067
rect 14387 15033 14437 15067
rect 14303 14999 14437 15033
rect 14303 14965 14353 14999
rect 14387 14965 14437 14999
rect 14303 14931 14437 14965
rect 14303 14897 14353 14931
rect 14387 14897 14437 14931
rect 14303 14863 14437 14897
rect 14303 14829 14353 14863
rect 14387 14829 14437 14863
rect 14303 14795 14437 14829
rect 14303 14761 14353 14795
rect 14387 14761 14437 14795
rect 14303 14727 14437 14761
rect 14303 14693 14353 14727
rect 14387 14693 14437 14727
rect 14303 14659 14437 14693
rect 14303 14625 14353 14659
rect 14387 14625 14437 14659
rect 14303 14591 14437 14625
rect 14303 14557 14353 14591
rect 14387 14557 14437 14591
rect 14303 14523 14437 14557
rect 14303 14489 14353 14523
rect 14387 14489 14437 14523
rect 14303 14455 14437 14489
rect 14303 14421 14353 14455
rect 14387 14421 14437 14455
rect 14303 14387 14437 14421
rect 14303 14353 14353 14387
rect 14387 14353 14437 14387
rect 14303 14319 14437 14353
rect 14303 14285 14353 14319
rect 14387 14285 14437 14319
rect 14303 14251 14437 14285
rect 14303 14217 14353 14251
rect 14387 14217 14437 14251
rect 14303 14183 14437 14217
rect 14303 14149 14353 14183
rect 14387 14149 14437 14183
rect 14303 14115 14437 14149
rect 14303 14081 14353 14115
rect 14387 14081 14437 14115
rect 14303 14047 14437 14081
rect 14303 14013 14353 14047
rect 14387 14013 14437 14047
rect 14303 13979 14437 14013
rect 14303 13945 14353 13979
rect 14387 13945 14437 13979
rect 14303 13911 14437 13945
rect 14303 13877 14353 13911
rect 14387 13877 14437 13911
rect 14303 13843 14437 13877
rect 14303 13809 14353 13843
rect 14387 13809 14437 13843
rect 14303 13775 14437 13809
rect 14303 13741 14353 13775
rect 14387 13741 14437 13775
rect 14303 13707 14437 13741
rect 14303 13673 14353 13707
rect 14387 13673 14437 13707
rect 14303 13639 14437 13673
rect 14303 13605 14353 13639
rect 14387 13605 14437 13639
rect 14303 13571 14437 13605
rect 14303 13537 14353 13571
rect 14387 13537 14437 13571
rect 14303 13503 14437 13537
rect 14303 13469 14353 13503
rect 14387 13469 14437 13503
rect 14303 13435 14437 13469
rect 14303 13401 14353 13435
rect 14387 13401 14437 13435
rect 14303 13367 14437 13401
rect 14303 13333 14353 13367
rect 14387 13333 14437 13367
rect 14303 13299 14437 13333
rect 14303 13265 14353 13299
rect 14387 13265 14437 13299
rect 14303 13231 14437 13265
rect 14303 13197 14353 13231
rect 14387 13197 14437 13231
rect 14303 13163 14437 13197
rect 14303 13129 14353 13163
rect 14387 13129 14437 13163
rect 14303 13095 14437 13129
rect 14303 13061 14353 13095
rect 14387 13061 14437 13095
rect 14303 13027 14437 13061
rect 14303 12993 14353 13027
rect 14387 12993 14437 13027
rect 14303 12959 14437 12993
rect 14303 12925 14353 12959
rect 14387 12925 14437 12959
rect 14303 12891 14437 12925
rect 14303 12857 14353 12891
rect 14387 12857 14437 12891
rect 14303 12823 14437 12857
rect 14303 12789 14353 12823
rect 14387 12789 14437 12823
rect 14303 12755 14437 12789
rect 14303 12721 14353 12755
rect 14387 12721 14437 12755
rect 14303 12687 14437 12721
rect 14303 12653 14353 12687
rect 14387 12653 14437 12687
rect 14303 12619 14437 12653
rect 14303 12585 14353 12619
rect 14387 12585 14437 12619
rect 14303 12551 14437 12585
rect 14303 12517 14353 12551
rect 14387 12517 14437 12551
rect 14303 12483 14437 12517
rect 14303 12449 14353 12483
rect 14387 12449 14437 12483
rect 14303 12415 14437 12449
rect 14303 12381 14353 12415
rect 14387 12381 14437 12415
rect 14303 12347 14437 12381
rect 14303 12313 14353 12347
rect 14387 12313 14437 12347
rect 14303 12279 14437 12313
rect 14303 12245 14353 12279
rect 14387 12245 14437 12279
rect 14303 12211 14437 12245
rect 14303 12177 14353 12211
rect 14387 12177 14437 12211
rect 14303 12143 14437 12177
rect 14303 12109 14353 12143
rect 14387 12109 14437 12143
rect 14303 12075 14437 12109
rect 14303 12041 14353 12075
rect 14387 12041 14437 12075
rect 14303 12007 14437 12041
rect 14303 11973 14353 12007
rect 14387 11973 14437 12007
rect 14303 11939 14437 11973
rect 14303 11905 14353 11939
rect 14387 11905 14437 11939
rect 14303 11871 14437 11905
rect 14303 11837 14353 11871
rect 14387 11837 14437 11871
rect 14303 11803 14437 11837
rect 14303 11769 14353 11803
rect 14387 11769 14437 11803
rect 14303 11735 14437 11769
rect 14303 11701 14353 11735
rect 14387 11701 14437 11735
rect 14303 11667 14437 11701
rect 14303 11633 14353 11667
rect 14387 11633 14437 11667
rect 14303 11599 14437 11633
rect 14303 11565 14353 11599
rect 14387 11565 14437 11599
rect 14303 11531 14437 11565
rect 14303 11497 14353 11531
rect 14387 11497 14437 11531
rect 14303 11463 14437 11497
rect 14303 11429 14353 11463
rect 14387 11429 14437 11463
rect 14303 11395 14437 11429
rect 14303 11361 14353 11395
rect 14387 11361 14437 11395
rect 14303 11327 14437 11361
rect 14303 11293 14353 11327
rect 14387 11293 14437 11327
rect 14303 11259 14437 11293
rect 14303 11225 14353 11259
rect 14387 11225 14437 11259
rect 14303 11191 14437 11225
rect 14303 11157 14353 11191
rect 14387 11157 14437 11191
rect 14303 11123 14437 11157
rect 14303 11089 14353 11123
rect 14387 11089 14437 11123
rect 14303 11055 14437 11089
rect 14303 11021 14353 11055
rect 14387 11021 14437 11055
rect 14303 10987 14437 11021
rect 14303 10953 14353 10987
rect 14387 10953 14437 10987
rect 14303 10919 14437 10953
rect 14303 10885 14353 10919
rect 14387 10885 14437 10919
rect 14303 10851 14437 10885
rect 14303 10817 14353 10851
rect 14387 10817 14437 10851
rect 14303 10783 14437 10817
rect 14303 10749 14353 10783
rect 14387 10749 14437 10783
rect 14303 10715 14437 10749
rect 14303 10681 14353 10715
rect 14387 10681 14437 10715
rect 14303 10647 14437 10681
rect 14303 10613 14353 10647
rect 14387 10613 14437 10647
rect 14303 10579 14437 10613
rect 14303 10545 14353 10579
rect 14387 10545 14437 10579
rect 14303 10511 14437 10545
rect 14303 10477 14353 10511
rect 14387 10477 14437 10511
rect 14303 10443 14437 10477
rect 14303 10409 14353 10443
rect 14387 10409 14437 10443
rect 14303 10375 14437 10409
rect 14303 10341 14353 10375
rect 14387 10341 14437 10375
rect 14303 10307 14437 10341
rect 14303 10273 14353 10307
rect 14387 10273 14437 10307
rect 14303 10239 14437 10273
rect 14303 10205 14353 10239
rect 14387 10205 14437 10239
rect 14303 10171 14437 10205
rect 14303 10137 14353 10171
rect 14387 10137 14437 10171
rect 14303 10103 14437 10137
rect 14303 10069 14353 10103
rect 14387 10069 14437 10103
rect 14303 10035 14437 10069
rect 14303 10001 14353 10035
rect 14387 10001 14437 10035
rect 14303 9967 14437 10001
rect 14303 9933 14353 9967
rect 14387 9933 14437 9967
rect 14303 9899 14437 9933
rect 14303 9865 14353 9899
rect 14387 9865 14437 9899
rect 14303 9831 14437 9865
rect 14303 9797 14353 9831
rect 14387 9797 14437 9831
rect 14303 9769 14437 9797
rect 569 9719 14437 9769
rect 569 9685 719 9719
rect 753 9685 787 9719
rect 821 9685 855 9719
rect 889 9685 923 9719
rect 957 9685 991 9719
rect 1025 9685 1059 9719
rect 1093 9685 1127 9719
rect 1161 9685 1195 9719
rect 1229 9685 1263 9719
rect 1297 9685 1331 9719
rect 1365 9685 1399 9719
rect 1433 9685 1467 9719
rect 1501 9685 1535 9719
rect 1569 9685 1603 9719
rect 1637 9685 1671 9719
rect 1705 9685 1739 9719
rect 1773 9685 1807 9719
rect 1841 9685 1875 9719
rect 1909 9685 1943 9719
rect 1977 9685 2011 9719
rect 2045 9685 2079 9719
rect 2113 9685 2147 9719
rect 2181 9685 2215 9719
rect 2249 9685 2283 9719
rect 2317 9685 2351 9719
rect 2385 9685 2419 9719
rect 2453 9685 2487 9719
rect 2521 9685 2555 9719
rect 2589 9685 2623 9719
rect 2657 9685 2691 9719
rect 2725 9685 2759 9719
rect 2793 9685 2827 9719
rect 2861 9685 2895 9719
rect 2929 9685 2963 9719
rect 2997 9685 3031 9719
rect 3065 9685 3099 9719
rect 3133 9685 3167 9719
rect 3201 9685 3235 9719
rect 3269 9685 3303 9719
rect 3337 9685 3371 9719
rect 3405 9685 3439 9719
rect 3473 9685 3507 9719
rect 3541 9685 3575 9719
rect 3609 9685 3643 9719
rect 3677 9685 3711 9719
rect 3745 9685 3779 9719
rect 3813 9685 3847 9719
rect 3881 9685 3915 9719
rect 3949 9685 3983 9719
rect 4017 9685 4051 9719
rect 4085 9685 4119 9719
rect 4153 9685 4187 9719
rect 4221 9685 4255 9719
rect 4289 9685 4323 9719
rect 4357 9685 4391 9719
rect 4425 9685 4459 9719
rect 4493 9685 4527 9719
rect 4561 9685 4595 9719
rect 4629 9685 4663 9719
rect 4697 9685 4731 9719
rect 4765 9685 4799 9719
rect 4833 9685 4867 9719
rect 4901 9685 4935 9719
rect 4969 9685 5003 9719
rect 5037 9685 5071 9719
rect 5105 9685 5139 9719
rect 5173 9685 5207 9719
rect 5241 9685 5275 9719
rect 5309 9685 5343 9719
rect 5377 9685 5411 9719
rect 5445 9685 5479 9719
rect 5513 9685 5547 9719
rect 5581 9685 5615 9719
rect 5649 9685 5683 9719
rect 5717 9685 5751 9719
rect 5785 9685 5819 9719
rect 5853 9685 5887 9719
rect 5921 9685 5955 9719
rect 5989 9685 6023 9719
rect 6057 9685 6091 9719
rect 6125 9685 6159 9719
rect 6193 9685 6227 9719
rect 6261 9685 6295 9719
rect 6329 9685 6363 9719
rect 6397 9685 6431 9719
rect 6465 9685 6499 9719
rect 6533 9685 6567 9719
rect 6601 9685 6635 9719
rect 6669 9685 6703 9719
rect 6737 9685 6771 9719
rect 6805 9685 6839 9719
rect 6873 9685 6907 9719
rect 6941 9685 6975 9719
rect 7009 9685 7043 9719
rect 7077 9685 7111 9719
rect 7145 9685 7179 9719
rect 7213 9685 7247 9719
rect 7281 9685 7315 9719
rect 7349 9685 7383 9719
rect 7417 9685 7451 9719
rect 7485 9685 7519 9719
rect 7553 9685 7587 9719
rect 7621 9685 7655 9719
rect 7689 9685 7723 9719
rect 7757 9685 7791 9719
rect 7825 9685 7859 9719
rect 7893 9685 7927 9719
rect 7961 9685 7995 9719
rect 8029 9685 8063 9719
rect 8097 9685 8131 9719
rect 8165 9685 8199 9719
rect 8233 9685 8267 9719
rect 8301 9685 8335 9719
rect 8369 9685 8403 9719
rect 8437 9685 8471 9719
rect 8505 9685 8539 9719
rect 8573 9685 8607 9719
rect 8641 9685 8675 9719
rect 8709 9685 8743 9719
rect 8777 9685 8811 9719
rect 8845 9685 8879 9719
rect 8913 9685 8947 9719
rect 8981 9685 9015 9719
rect 9049 9685 9083 9719
rect 9117 9685 9151 9719
rect 9185 9685 9219 9719
rect 9253 9685 9287 9719
rect 9321 9685 9355 9719
rect 9389 9685 9423 9719
rect 9457 9685 9491 9719
rect 9525 9685 9559 9719
rect 9593 9685 9627 9719
rect 9661 9685 9695 9719
rect 9729 9685 9763 9719
rect 9797 9685 9831 9719
rect 9865 9685 9899 9719
rect 9933 9685 9967 9719
rect 10001 9685 10035 9719
rect 10069 9685 10103 9719
rect 10137 9685 10171 9719
rect 10205 9685 10239 9719
rect 10273 9685 10307 9719
rect 10341 9685 10375 9719
rect 10409 9685 10443 9719
rect 10477 9685 10511 9719
rect 10545 9685 10579 9719
rect 10613 9685 10647 9719
rect 10681 9685 10715 9719
rect 10749 9685 10783 9719
rect 10817 9685 10851 9719
rect 10885 9685 10919 9719
rect 10953 9685 10987 9719
rect 11021 9685 11055 9719
rect 11089 9685 11123 9719
rect 11157 9685 11191 9719
rect 11225 9685 11259 9719
rect 11293 9685 11327 9719
rect 11361 9685 11395 9719
rect 11429 9685 11463 9719
rect 11497 9685 11531 9719
rect 11565 9685 11599 9719
rect 11633 9685 11667 9719
rect 11701 9685 11735 9719
rect 11769 9685 11803 9719
rect 11837 9685 11871 9719
rect 11905 9685 11939 9719
rect 11973 9685 12007 9719
rect 12041 9685 12075 9719
rect 12109 9685 12143 9719
rect 12177 9685 12211 9719
rect 12245 9685 12279 9719
rect 12313 9685 12347 9719
rect 12381 9685 12415 9719
rect 12449 9685 12483 9719
rect 12517 9685 12551 9719
rect 12585 9685 12619 9719
rect 12653 9685 12687 9719
rect 12721 9685 12755 9719
rect 12789 9685 12823 9719
rect 12857 9685 12891 9719
rect 12925 9685 12959 9719
rect 12993 9685 13027 9719
rect 13061 9685 13095 9719
rect 13129 9685 13163 9719
rect 13197 9685 13231 9719
rect 13265 9685 13299 9719
rect 13333 9685 13367 9719
rect 13401 9685 13435 9719
rect 13469 9685 13503 9719
rect 13537 9685 13571 9719
rect 13605 9685 13639 9719
rect 13673 9685 13707 9719
rect 13741 9685 13775 9719
rect 13809 9685 13843 9719
rect 13877 9685 13911 9719
rect 13945 9685 13979 9719
rect 14013 9685 14047 9719
rect 14081 9685 14115 9719
rect 14149 9685 14183 9719
rect 14217 9685 14251 9719
rect 14285 9685 14437 9719
rect 569 9635 14437 9685
<< nsubdiffcont >>
rect 719 36157 753 36191
rect 787 36157 821 36191
rect 855 36157 889 36191
rect 923 36157 957 36191
rect 991 36157 1025 36191
rect 1059 36157 1093 36191
rect 1127 36157 1161 36191
rect 1195 36157 1229 36191
rect 1263 36157 1297 36191
rect 1331 36157 1365 36191
rect 1399 36157 1433 36191
rect 1467 36157 1501 36191
rect 1535 36157 1569 36191
rect 1603 36157 1637 36191
rect 1671 36157 1705 36191
rect 1739 36157 1773 36191
rect 1807 36157 1841 36191
rect 1875 36157 1909 36191
rect 1943 36157 1977 36191
rect 2011 36157 2045 36191
rect 2079 36157 2113 36191
rect 2147 36157 2181 36191
rect 2215 36157 2249 36191
rect 2283 36157 2317 36191
rect 2351 36157 2385 36191
rect 2419 36157 2453 36191
rect 2487 36157 2521 36191
rect 2555 36157 2589 36191
rect 2623 36157 2657 36191
rect 2691 36157 2725 36191
rect 2759 36157 2793 36191
rect 2827 36157 2861 36191
rect 2895 36157 2929 36191
rect 2963 36157 2997 36191
rect 3031 36157 3065 36191
rect 3099 36157 3133 36191
rect 3167 36157 3201 36191
rect 3235 36157 3269 36191
rect 3303 36157 3337 36191
rect 3371 36157 3405 36191
rect 3439 36157 3473 36191
rect 3507 36157 3541 36191
rect 3575 36157 3609 36191
rect 3643 36157 3677 36191
rect 3711 36157 3745 36191
rect 3779 36157 3813 36191
rect 3847 36157 3881 36191
rect 3915 36157 3949 36191
rect 3983 36157 4017 36191
rect 4051 36157 4085 36191
rect 4119 36157 4153 36191
rect 4187 36157 4221 36191
rect 4255 36157 4289 36191
rect 4323 36157 4357 36191
rect 4391 36157 4425 36191
rect 4459 36157 4493 36191
rect 4527 36157 4561 36191
rect 4595 36157 4629 36191
rect 4663 36157 4697 36191
rect 4731 36157 4765 36191
rect 4799 36157 4833 36191
rect 4867 36157 4901 36191
rect 4935 36157 4969 36191
rect 5003 36157 5037 36191
rect 5071 36157 5105 36191
rect 5139 36157 5173 36191
rect 5207 36157 5241 36191
rect 5275 36157 5309 36191
rect 5343 36157 5377 36191
rect 5411 36157 5445 36191
rect 5479 36157 5513 36191
rect 5547 36157 5581 36191
rect 5615 36157 5649 36191
rect 5683 36157 5717 36191
rect 5751 36157 5785 36191
rect 5819 36157 5853 36191
rect 5887 36157 5921 36191
rect 5955 36157 5989 36191
rect 6023 36157 6057 36191
rect 6091 36157 6125 36191
rect 6159 36157 6193 36191
rect 6227 36157 6261 36191
rect 6295 36157 6329 36191
rect 6363 36157 6397 36191
rect 6431 36157 6465 36191
rect 6499 36157 6533 36191
rect 6567 36157 6601 36191
rect 6635 36157 6669 36191
rect 6703 36157 6737 36191
rect 6771 36157 6805 36191
rect 6839 36157 6873 36191
rect 6907 36157 6941 36191
rect 6975 36157 7009 36191
rect 7043 36157 7077 36191
rect 7111 36157 7145 36191
rect 7179 36157 7213 36191
rect 7247 36157 7281 36191
rect 7315 36157 7349 36191
rect 7383 36157 7417 36191
rect 7451 36157 7485 36191
rect 7519 36157 7553 36191
rect 7587 36157 7621 36191
rect 7655 36157 7689 36191
rect 7723 36157 7757 36191
rect 7791 36157 7825 36191
rect 7859 36157 7893 36191
rect 7927 36157 7961 36191
rect 7995 36157 8029 36191
rect 8063 36157 8097 36191
rect 8131 36157 8165 36191
rect 8199 36157 8233 36191
rect 8267 36157 8301 36191
rect 8335 36157 8369 36191
rect 8403 36157 8437 36191
rect 8471 36157 8505 36191
rect 8539 36157 8573 36191
rect 8607 36157 8641 36191
rect 8675 36157 8709 36191
rect 8743 36157 8777 36191
rect 8811 36157 8845 36191
rect 8879 36157 8913 36191
rect 8947 36157 8981 36191
rect 9015 36157 9049 36191
rect 9083 36157 9117 36191
rect 9151 36157 9185 36191
rect 9219 36157 9253 36191
rect 9287 36157 9321 36191
rect 9355 36157 9389 36191
rect 9423 36157 9457 36191
rect 9491 36157 9525 36191
rect 9559 36157 9593 36191
rect 9627 36157 9661 36191
rect 9695 36157 9729 36191
rect 9763 36157 9797 36191
rect 9831 36157 9865 36191
rect 9899 36157 9933 36191
rect 9967 36157 10001 36191
rect 10035 36157 10069 36191
rect 10103 36157 10137 36191
rect 10171 36157 10205 36191
rect 10239 36157 10273 36191
rect 10307 36157 10341 36191
rect 10375 36157 10409 36191
rect 10443 36157 10477 36191
rect 10511 36157 10545 36191
rect 10579 36157 10613 36191
rect 10647 36157 10681 36191
rect 10715 36157 10749 36191
rect 10783 36157 10817 36191
rect 10851 36157 10885 36191
rect 10919 36157 10953 36191
rect 10987 36157 11021 36191
rect 11055 36157 11089 36191
rect 11123 36157 11157 36191
rect 11191 36157 11225 36191
rect 11259 36157 11293 36191
rect 11327 36157 11361 36191
rect 11395 36157 11429 36191
rect 11463 36157 11497 36191
rect 11531 36157 11565 36191
rect 11599 36157 11633 36191
rect 11667 36157 11701 36191
rect 11735 36157 11769 36191
rect 11803 36157 11837 36191
rect 11871 36157 11905 36191
rect 11939 36157 11973 36191
rect 12007 36157 12041 36191
rect 12075 36157 12109 36191
rect 12143 36157 12177 36191
rect 12211 36157 12245 36191
rect 12279 36157 12313 36191
rect 12347 36157 12381 36191
rect 12415 36157 12449 36191
rect 12483 36157 12517 36191
rect 12551 36157 12585 36191
rect 12619 36157 12653 36191
rect 12687 36157 12721 36191
rect 12755 36157 12789 36191
rect 12823 36157 12857 36191
rect 12891 36157 12925 36191
rect 12959 36157 12993 36191
rect 13027 36157 13061 36191
rect 13095 36157 13129 36191
rect 13163 36157 13197 36191
rect 13231 36157 13265 36191
rect 13299 36157 13333 36191
rect 13367 36157 13401 36191
rect 13435 36157 13469 36191
rect 13503 36157 13537 36191
rect 13571 36157 13605 36191
rect 13639 36157 13673 36191
rect 13707 36157 13741 36191
rect 13775 36157 13809 36191
rect 13843 36157 13877 36191
rect 13911 36157 13945 36191
rect 13979 36157 14013 36191
rect 14047 36157 14081 36191
rect 14115 36157 14149 36191
rect 14183 36157 14217 36191
rect 14251 36157 14285 36191
rect 618 36045 652 36079
rect 618 35977 652 36011
rect 618 35909 652 35943
rect 618 35841 652 35875
rect 618 35773 652 35807
rect 618 35705 652 35739
rect 618 35637 652 35671
rect 618 35569 652 35603
rect 618 35501 652 35535
rect 618 35433 652 35467
rect 618 35365 652 35399
rect 618 35297 652 35331
rect 618 35229 652 35263
rect 618 35161 652 35195
rect 618 35093 652 35127
rect 618 35025 652 35059
rect 618 34957 652 34991
rect 618 34889 652 34923
rect 618 34821 652 34855
rect 618 34753 652 34787
rect 618 34685 652 34719
rect 618 34617 652 34651
rect 618 34549 652 34583
rect 618 34481 652 34515
rect 618 34413 652 34447
rect 618 34345 652 34379
rect 618 34277 652 34311
rect 618 34209 652 34243
rect 618 34141 652 34175
rect 618 34073 652 34107
rect 618 34005 652 34039
rect 618 33937 652 33971
rect 618 33869 652 33903
rect 618 33801 652 33835
rect 618 33733 652 33767
rect 618 33665 652 33699
rect 618 33597 652 33631
rect 618 33529 652 33563
rect 618 33461 652 33495
rect 618 33393 652 33427
rect 618 33325 652 33359
rect 618 33257 652 33291
rect 618 33189 652 33223
rect 618 33121 652 33155
rect 618 33053 652 33087
rect 618 32985 652 33019
rect 618 32917 652 32951
rect 618 32849 652 32883
rect 618 32781 652 32815
rect 618 32713 652 32747
rect 618 32645 652 32679
rect 618 32577 652 32611
rect 618 32509 652 32543
rect 618 32441 652 32475
rect 618 32373 652 32407
rect 618 32305 652 32339
rect 618 32237 652 32271
rect 618 32169 652 32203
rect 618 32101 652 32135
rect 618 32033 652 32067
rect 618 31965 652 31999
rect 618 31897 652 31931
rect 618 31829 652 31863
rect 618 31761 652 31795
rect 618 31693 652 31727
rect 618 31625 652 31659
rect 618 31557 652 31591
rect 618 31489 652 31523
rect 618 31421 652 31455
rect 618 31353 652 31387
rect 618 31285 652 31319
rect 618 31217 652 31251
rect 618 31149 652 31183
rect 618 31081 652 31115
rect 618 31013 652 31047
rect 618 30945 652 30979
rect 618 30877 652 30911
rect 618 30809 652 30843
rect 618 30741 652 30775
rect 618 30673 652 30707
rect 618 30605 652 30639
rect 618 30537 652 30571
rect 618 30469 652 30503
rect 618 30401 652 30435
rect 618 30333 652 30367
rect 618 30265 652 30299
rect 618 30197 652 30231
rect 618 30129 652 30163
rect 618 30061 652 30095
rect 618 29993 652 30027
rect 618 29925 652 29959
rect 618 29857 652 29891
rect 618 29789 652 29823
rect 618 29721 652 29755
rect 618 29653 652 29687
rect 618 29585 652 29619
rect 618 29517 652 29551
rect 618 29449 652 29483
rect 618 29381 652 29415
rect 618 29313 652 29347
rect 618 29245 652 29279
rect 618 29177 652 29211
rect 618 29109 652 29143
rect 618 29041 652 29075
rect 618 28973 652 29007
rect 618 28905 652 28939
rect 618 28837 652 28871
rect 618 28769 652 28803
rect 618 28701 652 28735
rect 618 28633 652 28667
rect 618 28565 652 28599
rect 618 28497 652 28531
rect 618 28429 652 28463
rect 618 28361 652 28395
rect 618 28293 652 28327
rect 618 28225 652 28259
rect 618 28157 652 28191
rect 618 28089 652 28123
rect 618 28021 652 28055
rect 618 27953 652 27987
rect 618 27885 652 27919
rect 618 27817 652 27851
rect 618 27749 652 27783
rect 618 27681 652 27715
rect 618 27613 652 27647
rect 618 27545 652 27579
rect 618 27477 652 27511
rect 618 27409 652 27443
rect 618 27341 652 27375
rect 618 27273 652 27307
rect 618 27205 652 27239
rect 618 27137 652 27171
rect 618 27069 652 27103
rect 618 27001 652 27035
rect 618 26933 652 26967
rect 618 26865 652 26899
rect 618 26797 652 26831
rect 618 26729 652 26763
rect 618 26661 652 26695
rect 618 26593 652 26627
rect 618 26525 652 26559
rect 618 26457 652 26491
rect 618 26389 652 26423
rect 618 26321 652 26355
rect 618 26253 652 26287
rect 618 26185 652 26219
rect 618 26117 652 26151
rect 618 26049 652 26083
rect 618 25981 652 26015
rect 618 25913 652 25947
rect 618 25845 652 25879
rect 618 25777 652 25811
rect 618 25709 652 25743
rect 618 25641 652 25675
rect 618 25573 652 25607
rect 618 25505 652 25539
rect 618 25437 652 25471
rect 618 25369 652 25403
rect 618 25301 652 25335
rect 618 25233 652 25267
rect 618 25165 652 25199
rect 618 25097 652 25131
rect 618 25029 652 25063
rect 618 24961 652 24995
rect 618 24893 652 24927
rect 618 24825 652 24859
rect 618 24757 652 24791
rect 618 24689 652 24723
rect 618 24621 652 24655
rect 618 24553 652 24587
rect 618 24485 652 24519
rect 618 24417 652 24451
rect 618 24349 652 24383
rect 618 24281 652 24315
rect 618 24213 652 24247
rect 618 24145 652 24179
rect 618 24077 652 24111
rect 618 24009 652 24043
rect 618 23941 652 23975
rect 618 23873 652 23907
rect 618 23805 652 23839
rect 618 23737 652 23771
rect 618 23669 652 23703
rect 618 23601 652 23635
rect 618 23533 652 23567
rect 618 23465 652 23499
rect 618 23397 652 23431
rect 618 23329 652 23363
rect 618 23261 652 23295
rect 618 23193 652 23227
rect 618 23125 652 23159
rect 618 23057 652 23091
rect 618 22989 652 23023
rect 618 22921 652 22955
rect 618 22853 652 22887
rect 618 22785 652 22819
rect 618 22717 652 22751
rect 618 22649 652 22683
rect 618 22581 652 22615
rect 618 22513 652 22547
rect 618 22445 652 22479
rect 618 22377 652 22411
rect 618 22309 652 22343
rect 618 22241 652 22275
rect 618 22173 652 22207
rect 618 22105 652 22139
rect 618 22037 652 22071
rect 618 21969 652 22003
rect 618 21901 652 21935
rect 618 21833 652 21867
rect 618 21765 652 21799
rect 618 21697 652 21731
rect 618 21629 652 21663
rect 618 21561 652 21595
rect 618 21493 652 21527
rect 618 21425 652 21459
rect 618 21357 652 21391
rect 618 21289 652 21323
rect 618 21221 652 21255
rect 618 21153 652 21187
rect 618 21085 652 21119
rect 618 21017 652 21051
rect 618 20949 652 20983
rect 618 20881 652 20915
rect 618 20813 652 20847
rect 618 20745 652 20779
rect 618 20677 652 20711
rect 618 20609 652 20643
rect 618 20541 652 20575
rect 618 20473 652 20507
rect 618 20405 652 20439
rect 618 20337 652 20371
rect 618 20269 652 20303
rect 618 20201 652 20235
rect 618 20133 652 20167
rect 618 20065 652 20099
rect 618 19997 652 20031
rect 618 19929 652 19963
rect 618 19861 652 19895
rect 618 19793 652 19827
rect 618 19725 652 19759
rect 618 19657 652 19691
rect 618 19589 652 19623
rect 618 19521 652 19555
rect 618 19453 652 19487
rect 618 19385 652 19419
rect 618 19317 652 19351
rect 618 19249 652 19283
rect 618 19181 652 19215
rect 618 19113 652 19147
rect 618 19045 652 19079
rect 618 18977 652 19011
rect 618 18909 652 18943
rect 618 18841 652 18875
rect 618 18773 652 18807
rect 618 18705 652 18739
rect 618 18637 652 18671
rect 618 18569 652 18603
rect 618 18501 652 18535
rect 618 18433 652 18467
rect 618 18365 652 18399
rect 618 18297 652 18331
rect 618 18229 652 18263
rect 618 18161 652 18195
rect 618 18093 652 18127
rect 618 18025 652 18059
rect 618 17957 652 17991
rect 618 17889 652 17923
rect 618 17821 652 17855
rect 618 17753 652 17787
rect 618 17685 652 17719
rect 618 17617 652 17651
rect 618 17549 652 17583
rect 618 17481 652 17515
rect 618 17413 652 17447
rect 618 17345 652 17379
rect 618 17277 652 17311
rect 618 17209 652 17243
rect 618 17141 652 17175
rect 618 17073 652 17107
rect 618 17005 652 17039
rect 618 16937 652 16971
rect 618 16869 652 16903
rect 618 16801 652 16835
rect 618 16733 652 16767
rect 618 16665 652 16699
rect 618 16597 652 16631
rect 618 16529 652 16563
rect 618 16461 652 16495
rect 618 16393 652 16427
rect 618 16325 652 16359
rect 618 16257 652 16291
rect 618 16189 652 16223
rect 618 16121 652 16155
rect 618 16053 652 16087
rect 618 15985 652 16019
rect 618 15917 652 15951
rect 618 15849 652 15883
rect 618 15781 652 15815
rect 618 15713 652 15747
rect 618 15645 652 15679
rect 618 15577 652 15611
rect 618 15509 652 15543
rect 618 15441 652 15475
rect 618 15373 652 15407
rect 618 15305 652 15339
rect 618 15237 652 15271
rect 618 15169 652 15203
rect 618 15101 652 15135
rect 618 15033 652 15067
rect 618 14965 652 14999
rect 618 14897 652 14931
rect 618 14829 652 14863
rect 618 14761 652 14795
rect 618 14693 652 14727
rect 618 14625 652 14659
rect 618 14557 652 14591
rect 618 14489 652 14523
rect 618 14421 652 14455
rect 618 14353 652 14387
rect 618 14285 652 14319
rect 618 14217 652 14251
rect 618 14149 652 14183
rect 618 14081 652 14115
rect 618 14013 652 14047
rect 618 13945 652 13979
rect 618 13877 652 13911
rect 618 13809 652 13843
rect 618 13741 652 13775
rect 618 13673 652 13707
rect 618 13605 652 13639
rect 618 13537 652 13571
rect 618 13469 652 13503
rect 618 13401 652 13435
rect 618 13333 652 13367
rect 618 13265 652 13299
rect 618 13197 652 13231
rect 618 13129 652 13163
rect 618 13061 652 13095
rect 618 12993 652 13027
rect 618 12925 652 12959
rect 618 12857 652 12891
rect 618 12789 652 12823
rect 618 12721 652 12755
rect 618 12653 652 12687
rect 618 12585 652 12619
rect 618 12517 652 12551
rect 618 12449 652 12483
rect 618 12381 652 12415
rect 618 12313 652 12347
rect 618 12245 652 12279
rect 618 12177 652 12211
rect 618 12109 652 12143
rect 618 12041 652 12075
rect 618 11973 652 12007
rect 618 11905 652 11939
rect 618 11837 652 11871
rect 618 11769 652 11803
rect 618 11701 652 11735
rect 618 11633 652 11667
rect 618 11565 652 11599
rect 618 11497 652 11531
rect 618 11429 652 11463
rect 618 11361 652 11395
rect 618 11293 652 11327
rect 618 11225 652 11259
rect 618 11157 652 11191
rect 618 11089 652 11123
rect 618 11021 652 11055
rect 618 10953 652 10987
rect 618 10885 652 10919
rect 618 10817 652 10851
rect 618 10749 652 10783
rect 618 10681 652 10715
rect 618 10613 652 10647
rect 618 10545 652 10579
rect 618 10477 652 10511
rect 618 10409 652 10443
rect 618 10341 652 10375
rect 618 10273 652 10307
rect 618 10205 652 10239
rect 618 10137 652 10171
rect 618 10069 652 10103
rect 618 10001 652 10035
rect 618 9933 652 9967
rect 618 9865 652 9899
rect 618 9797 652 9831
rect 14353 36045 14387 36079
rect 14353 35977 14387 36011
rect 14353 35909 14387 35943
rect 14353 35841 14387 35875
rect 14353 35773 14387 35807
rect 14353 35705 14387 35739
rect 14353 35637 14387 35671
rect 14353 35569 14387 35603
rect 14353 35501 14387 35535
rect 14353 35433 14387 35467
rect 14353 35365 14387 35399
rect 14353 35297 14387 35331
rect 14353 35229 14387 35263
rect 14353 35161 14387 35195
rect 14353 35093 14387 35127
rect 14353 35025 14387 35059
rect 14353 34957 14387 34991
rect 14353 34889 14387 34923
rect 14353 34821 14387 34855
rect 14353 34753 14387 34787
rect 14353 34685 14387 34719
rect 14353 34617 14387 34651
rect 14353 34549 14387 34583
rect 14353 34481 14387 34515
rect 14353 34413 14387 34447
rect 14353 34345 14387 34379
rect 14353 34277 14387 34311
rect 14353 34209 14387 34243
rect 14353 34141 14387 34175
rect 14353 34073 14387 34107
rect 14353 34005 14387 34039
rect 14353 33937 14387 33971
rect 14353 33869 14387 33903
rect 14353 33801 14387 33835
rect 14353 33733 14387 33767
rect 14353 33665 14387 33699
rect 14353 33597 14387 33631
rect 14353 33529 14387 33563
rect 14353 33461 14387 33495
rect 14353 33393 14387 33427
rect 14353 33325 14387 33359
rect 14353 33257 14387 33291
rect 14353 33189 14387 33223
rect 14353 33121 14387 33155
rect 14353 33053 14387 33087
rect 14353 32985 14387 33019
rect 14353 32917 14387 32951
rect 14353 32849 14387 32883
rect 14353 32781 14387 32815
rect 14353 32713 14387 32747
rect 14353 32645 14387 32679
rect 14353 32577 14387 32611
rect 14353 32509 14387 32543
rect 14353 32441 14387 32475
rect 14353 32373 14387 32407
rect 14353 32305 14387 32339
rect 14353 32237 14387 32271
rect 14353 32169 14387 32203
rect 14353 32101 14387 32135
rect 14353 32033 14387 32067
rect 14353 31965 14387 31999
rect 14353 31897 14387 31931
rect 14353 31829 14387 31863
rect 14353 31761 14387 31795
rect 14353 31693 14387 31727
rect 14353 31625 14387 31659
rect 14353 31557 14387 31591
rect 14353 31489 14387 31523
rect 14353 31421 14387 31455
rect 14353 31353 14387 31387
rect 14353 31285 14387 31319
rect 14353 31217 14387 31251
rect 14353 31149 14387 31183
rect 14353 31081 14387 31115
rect 14353 31013 14387 31047
rect 14353 30945 14387 30979
rect 14353 30877 14387 30911
rect 14353 30809 14387 30843
rect 14353 30741 14387 30775
rect 14353 30673 14387 30707
rect 14353 30605 14387 30639
rect 14353 30537 14387 30571
rect 14353 30469 14387 30503
rect 14353 30401 14387 30435
rect 14353 30333 14387 30367
rect 14353 30265 14387 30299
rect 14353 30197 14387 30231
rect 14353 30129 14387 30163
rect 14353 30061 14387 30095
rect 14353 29993 14387 30027
rect 14353 29925 14387 29959
rect 14353 29857 14387 29891
rect 14353 29789 14387 29823
rect 14353 29721 14387 29755
rect 14353 29653 14387 29687
rect 14353 29585 14387 29619
rect 14353 29517 14387 29551
rect 14353 29449 14387 29483
rect 14353 29381 14387 29415
rect 14353 29313 14387 29347
rect 14353 29245 14387 29279
rect 14353 29177 14387 29211
rect 14353 29109 14387 29143
rect 14353 29041 14387 29075
rect 14353 28973 14387 29007
rect 14353 28905 14387 28939
rect 14353 28837 14387 28871
rect 14353 28769 14387 28803
rect 14353 28701 14387 28735
rect 14353 28633 14387 28667
rect 14353 28565 14387 28599
rect 14353 28497 14387 28531
rect 14353 28429 14387 28463
rect 14353 28361 14387 28395
rect 14353 28293 14387 28327
rect 14353 28225 14387 28259
rect 14353 28157 14387 28191
rect 14353 28089 14387 28123
rect 14353 28021 14387 28055
rect 14353 27953 14387 27987
rect 14353 27885 14387 27919
rect 14353 27817 14387 27851
rect 14353 27749 14387 27783
rect 14353 27681 14387 27715
rect 14353 27613 14387 27647
rect 14353 27545 14387 27579
rect 14353 27477 14387 27511
rect 14353 27409 14387 27443
rect 14353 27341 14387 27375
rect 14353 27273 14387 27307
rect 14353 27205 14387 27239
rect 14353 27137 14387 27171
rect 14353 27069 14387 27103
rect 14353 27001 14387 27035
rect 14353 26933 14387 26967
rect 14353 26865 14387 26899
rect 14353 26797 14387 26831
rect 14353 26729 14387 26763
rect 14353 26661 14387 26695
rect 14353 26593 14387 26627
rect 14353 26525 14387 26559
rect 14353 26457 14387 26491
rect 14353 26389 14387 26423
rect 14353 26321 14387 26355
rect 14353 26253 14387 26287
rect 14353 26185 14387 26219
rect 14353 26117 14387 26151
rect 14353 26049 14387 26083
rect 14353 25981 14387 26015
rect 14353 25913 14387 25947
rect 14353 25845 14387 25879
rect 14353 25777 14387 25811
rect 14353 25709 14387 25743
rect 14353 25641 14387 25675
rect 14353 25573 14387 25607
rect 14353 25505 14387 25539
rect 14353 25437 14387 25471
rect 14353 25369 14387 25403
rect 14353 25301 14387 25335
rect 14353 25233 14387 25267
rect 14353 25165 14387 25199
rect 14353 25097 14387 25131
rect 14353 25029 14387 25063
rect 14353 24961 14387 24995
rect 14353 24893 14387 24927
rect 14353 24825 14387 24859
rect 14353 24757 14387 24791
rect 14353 24689 14387 24723
rect 14353 24621 14387 24655
rect 14353 24553 14387 24587
rect 14353 24485 14387 24519
rect 14353 24417 14387 24451
rect 14353 24349 14387 24383
rect 14353 24281 14387 24315
rect 14353 24213 14387 24247
rect 14353 24145 14387 24179
rect 14353 24077 14387 24111
rect 14353 24009 14387 24043
rect 14353 23941 14387 23975
rect 14353 23873 14387 23907
rect 14353 23805 14387 23839
rect 14353 23737 14387 23771
rect 14353 23669 14387 23703
rect 14353 23601 14387 23635
rect 14353 23533 14387 23567
rect 14353 23465 14387 23499
rect 14353 23397 14387 23431
rect 14353 23329 14387 23363
rect 14353 23261 14387 23295
rect 14353 23193 14387 23227
rect 14353 23125 14387 23159
rect 14353 23057 14387 23091
rect 14353 22989 14387 23023
rect 14353 22921 14387 22955
rect 14353 22853 14387 22887
rect 14353 22785 14387 22819
rect 14353 22717 14387 22751
rect 14353 22649 14387 22683
rect 14353 22581 14387 22615
rect 14353 22513 14387 22547
rect 14353 22445 14387 22479
rect 14353 22377 14387 22411
rect 14353 22309 14387 22343
rect 14353 22241 14387 22275
rect 14353 22173 14387 22207
rect 14353 22105 14387 22139
rect 14353 22037 14387 22071
rect 14353 21969 14387 22003
rect 14353 21901 14387 21935
rect 14353 21833 14387 21867
rect 14353 21765 14387 21799
rect 14353 21697 14387 21731
rect 14353 21629 14387 21663
rect 14353 21561 14387 21595
rect 14353 21493 14387 21527
rect 14353 21425 14387 21459
rect 14353 21357 14387 21391
rect 14353 21289 14387 21323
rect 14353 21221 14387 21255
rect 14353 21153 14387 21187
rect 14353 21085 14387 21119
rect 14353 21017 14387 21051
rect 14353 20949 14387 20983
rect 14353 20881 14387 20915
rect 14353 20813 14387 20847
rect 14353 20745 14387 20779
rect 14353 20677 14387 20711
rect 14353 20609 14387 20643
rect 14353 20541 14387 20575
rect 14353 20473 14387 20507
rect 14353 20405 14387 20439
rect 14353 20337 14387 20371
rect 14353 20269 14387 20303
rect 14353 20201 14387 20235
rect 14353 20133 14387 20167
rect 14353 20065 14387 20099
rect 14353 19997 14387 20031
rect 14353 19929 14387 19963
rect 14353 19861 14387 19895
rect 14353 19793 14387 19827
rect 14353 19725 14387 19759
rect 14353 19657 14387 19691
rect 14353 19589 14387 19623
rect 14353 19521 14387 19555
rect 14353 19453 14387 19487
rect 14353 19385 14387 19419
rect 14353 19317 14387 19351
rect 14353 19249 14387 19283
rect 14353 19181 14387 19215
rect 14353 19113 14387 19147
rect 14353 19045 14387 19079
rect 14353 18977 14387 19011
rect 14353 18909 14387 18943
rect 14353 18841 14387 18875
rect 14353 18773 14387 18807
rect 14353 18705 14387 18739
rect 14353 18637 14387 18671
rect 14353 18569 14387 18603
rect 14353 18501 14387 18535
rect 14353 18433 14387 18467
rect 14353 18365 14387 18399
rect 14353 18297 14387 18331
rect 14353 18229 14387 18263
rect 14353 18161 14387 18195
rect 14353 18093 14387 18127
rect 14353 18025 14387 18059
rect 14353 17957 14387 17991
rect 14353 17889 14387 17923
rect 14353 17821 14387 17855
rect 14353 17753 14387 17787
rect 14353 17685 14387 17719
rect 14353 17617 14387 17651
rect 14353 17549 14387 17583
rect 14353 17481 14387 17515
rect 14353 17413 14387 17447
rect 14353 17345 14387 17379
rect 14353 17277 14387 17311
rect 14353 17209 14387 17243
rect 14353 17141 14387 17175
rect 14353 17073 14387 17107
rect 14353 17005 14387 17039
rect 14353 16937 14387 16971
rect 14353 16869 14387 16903
rect 14353 16801 14387 16835
rect 14353 16733 14387 16767
rect 14353 16665 14387 16699
rect 14353 16597 14387 16631
rect 14353 16529 14387 16563
rect 14353 16461 14387 16495
rect 14353 16393 14387 16427
rect 14353 16325 14387 16359
rect 14353 16257 14387 16291
rect 14353 16189 14387 16223
rect 14353 16121 14387 16155
rect 14353 16053 14387 16087
rect 14353 15985 14387 16019
rect 14353 15917 14387 15951
rect 14353 15849 14387 15883
rect 14353 15781 14387 15815
rect 14353 15713 14387 15747
rect 14353 15645 14387 15679
rect 14353 15577 14387 15611
rect 14353 15509 14387 15543
rect 14353 15441 14387 15475
rect 14353 15373 14387 15407
rect 14353 15305 14387 15339
rect 14353 15237 14387 15271
rect 14353 15169 14387 15203
rect 14353 15101 14387 15135
rect 14353 15033 14387 15067
rect 14353 14965 14387 14999
rect 14353 14897 14387 14931
rect 14353 14829 14387 14863
rect 14353 14761 14387 14795
rect 14353 14693 14387 14727
rect 14353 14625 14387 14659
rect 14353 14557 14387 14591
rect 14353 14489 14387 14523
rect 14353 14421 14387 14455
rect 14353 14353 14387 14387
rect 14353 14285 14387 14319
rect 14353 14217 14387 14251
rect 14353 14149 14387 14183
rect 14353 14081 14387 14115
rect 14353 14013 14387 14047
rect 14353 13945 14387 13979
rect 14353 13877 14387 13911
rect 14353 13809 14387 13843
rect 14353 13741 14387 13775
rect 14353 13673 14387 13707
rect 14353 13605 14387 13639
rect 14353 13537 14387 13571
rect 14353 13469 14387 13503
rect 14353 13401 14387 13435
rect 14353 13333 14387 13367
rect 14353 13265 14387 13299
rect 14353 13197 14387 13231
rect 14353 13129 14387 13163
rect 14353 13061 14387 13095
rect 14353 12993 14387 13027
rect 14353 12925 14387 12959
rect 14353 12857 14387 12891
rect 14353 12789 14387 12823
rect 14353 12721 14387 12755
rect 14353 12653 14387 12687
rect 14353 12585 14387 12619
rect 14353 12517 14387 12551
rect 14353 12449 14387 12483
rect 14353 12381 14387 12415
rect 14353 12313 14387 12347
rect 14353 12245 14387 12279
rect 14353 12177 14387 12211
rect 14353 12109 14387 12143
rect 14353 12041 14387 12075
rect 14353 11973 14387 12007
rect 14353 11905 14387 11939
rect 14353 11837 14387 11871
rect 14353 11769 14387 11803
rect 14353 11701 14387 11735
rect 14353 11633 14387 11667
rect 14353 11565 14387 11599
rect 14353 11497 14387 11531
rect 14353 11429 14387 11463
rect 14353 11361 14387 11395
rect 14353 11293 14387 11327
rect 14353 11225 14387 11259
rect 14353 11157 14387 11191
rect 14353 11089 14387 11123
rect 14353 11021 14387 11055
rect 14353 10953 14387 10987
rect 14353 10885 14387 10919
rect 14353 10817 14387 10851
rect 14353 10749 14387 10783
rect 14353 10681 14387 10715
rect 14353 10613 14387 10647
rect 14353 10545 14387 10579
rect 14353 10477 14387 10511
rect 14353 10409 14387 10443
rect 14353 10341 14387 10375
rect 14353 10273 14387 10307
rect 14353 10205 14387 10239
rect 14353 10137 14387 10171
rect 14353 10069 14387 10103
rect 14353 10001 14387 10035
rect 14353 9933 14387 9967
rect 14353 9865 14387 9899
rect 14353 9797 14387 9831
rect 719 9685 753 9719
rect 787 9685 821 9719
rect 855 9685 889 9719
rect 923 9685 957 9719
rect 991 9685 1025 9719
rect 1059 9685 1093 9719
rect 1127 9685 1161 9719
rect 1195 9685 1229 9719
rect 1263 9685 1297 9719
rect 1331 9685 1365 9719
rect 1399 9685 1433 9719
rect 1467 9685 1501 9719
rect 1535 9685 1569 9719
rect 1603 9685 1637 9719
rect 1671 9685 1705 9719
rect 1739 9685 1773 9719
rect 1807 9685 1841 9719
rect 1875 9685 1909 9719
rect 1943 9685 1977 9719
rect 2011 9685 2045 9719
rect 2079 9685 2113 9719
rect 2147 9685 2181 9719
rect 2215 9685 2249 9719
rect 2283 9685 2317 9719
rect 2351 9685 2385 9719
rect 2419 9685 2453 9719
rect 2487 9685 2521 9719
rect 2555 9685 2589 9719
rect 2623 9685 2657 9719
rect 2691 9685 2725 9719
rect 2759 9685 2793 9719
rect 2827 9685 2861 9719
rect 2895 9685 2929 9719
rect 2963 9685 2997 9719
rect 3031 9685 3065 9719
rect 3099 9685 3133 9719
rect 3167 9685 3201 9719
rect 3235 9685 3269 9719
rect 3303 9685 3337 9719
rect 3371 9685 3405 9719
rect 3439 9685 3473 9719
rect 3507 9685 3541 9719
rect 3575 9685 3609 9719
rect 3643 9685 3677 9719
rect 3711 9685 3745 9719
rect 3779 9685 3813 9719
rect 3847 9685 3881 9719
rect 3915 9685 3949 9719
rect 3983 9685 4017 9719
rect 4051 9685 4085 9719
rect 4119 9685 4153 9719
rect 4187 9685 4221 9719
rect 4255 9685 4289 9719
rect 4323 9685 4357 9719
rect 4391 9685 4425 9719
rect 4459 9685 4493 9719
rect 4527 9685 4561 9719
rect 4595 9685 4629 9719
rect 4663 9685 4697 9719
rect 4731 9685 4765 9719
rect 4799 9685 4833 9719
rect 4867 9685 4901 9719
rect 4935 9685 4969 9719
rect 5003 9685 5037 9719
rect 5071 9685 5105 9719
rect 5139 9685 5173 9719
rect 5207 9685 5241 9719
rect 5275 9685 5309 9719
rect 5343 9685 5377 9719
rect 5411 9685 5445 9719
rect 5479 9685 5513 9719
rect 5547 9685 5581 9719
rect 5615 9685 5649 9719
rect 5683 9685 5717 9719
rect 5751 9685 5785 9719
rect 5819 9685 5853 9719
rect 5887 9685 5921 9719
rect 5955 9685 5989 9719
rect 6023 9685 6057 9719
rect 6091 9685 6125 9719
rect 6159 9685 6193 9719
rect 6227 9685 6261 9719
rect 6295 9685 6329 9719
rect 6363 9685 6397 9719
rect 6431 9685 6465 9719
rect 6499 9685 6533 9719
rect 6567 9685 6601 9719
rect 6635 9685 6669 9719
rect 6703 9685 6737 9719
rect 6771 9685 6805 9719
rect 6839 9685 6873 9719
rect 6907 9685 6941 9719
rect 6975 9685 7009 9719
rect 7043 9685 7077 9719
rect 7111 9685 7145 9719
rect 7179 9685 7213 9719
rect 7247 9685 7281 9719
rect 7315 9685 7349 9719
rect 7383 9685 7417 9719
rect 7451 9685 7485 9719
rect 7519 9685 7553 9719
rect 7587 9685 7621 9719
rect 7655 9685 7689 9719
rect 7723 9685 7757 9719
rect 7791 9685 7825 9719
rect 7859 9685 7893 9719
rect 7927 9685 7961 9719
rect 7995 9685 8029 9719
rect 8063 9685 8097 9719
rect 8131 9685 8165 9719
rect 8199 9685 8233 9719
rect 8267 9685 8301 9719
rect 8335 9685 8369 9719
rect 8403 9685 8437 9719
rect 8471 9685 8505 9719
rect 8539 9685 8573 9719
rect 8607 9685 8641 9719
rect 8675 9685 8709 9719
rect 8743 9685 8777 9719
rect 8811 9685 8845 9719
rect 8879 9685 8913 9719
rect 8947 9685 8981 9719
rect 9015 9685 9049 9719
rect 9083 9685 9117 9719
rect 9151 9685 9185 9719
rect 9219 9685 9253 9719
rect 9287 9685 9321 9719
rect 9355 9685 9389 9719
rect 9423 9685 9457 9719
rect 9491 9685 9525 9719
rect 9559 9685 9593 9719
rect 9627 9685 9661 9719
rect 9695 9685 9729 9719
rect 9763 9685 9797 9719
rect 9831 9685 9865 9719
rect 9899 9685 9933 9719
rect 9967 9685 10001 9719
rect 10035 9685 10069 9719
rect 10103 9685 10137 9719
rect 10171 9685 10205 9719
rect 10239 9685 10273 9719
rect 10307 9685 10341 9719
rect 10375 9685 10409 9719
rect 10443 9685 10477 9719
rect 10511 9685 10545 9719
rect 10579 9685 10613 9719
rect 10647 9685 10681 9719
rect 10715 9685 10749 9719
rect 10783 9685 10817 9719
rect 10851 9685 10885 9719
rect 10919 9685 10953 9719
rect 10987 9685 11021 9719
rect 11055 9685 11089 9719
rect 11123 9685 11157 9719
rect 11191 9685 11225 9719
rect 11259 9685 11293 9719
rect 11327 9685 11361 9719
rect 11395 9685 11429 9719
rect 11463 9685 11497 9719
rect 11531 9685 11565 9719
rect 11599 9685 11633 9719
rect 11667 9685 11701 9719
rect 11735 9685 11769 9719
rect 11803 9685 11837 9719
rect 11871 9685 11905 9719
rect 11939 9685 11973 9719
rect 12007 9685 12041 9719
rect 12075 9685 12109 9719
rect 12143 9685 12177 9719
rect 12211 9685 12245 9719
rect 12279 9685 12313 9719
rect 12347 9685 12381 9719
rect 12415 9685 12449 9719
rect 12483 9685 12517 9719
rect 12551 9685 12585 9719
rect 12619 9685 12653 9719
rect 12687 9685 12721 9719
rect 12755 9685 12789 9719
rect 12823 9685 12857 9719
rect 12891 9685 12925 9719
rect 12959 9685 12993 9719
rect 13027 9685 13061 9719
rect 13095 9685 13129 9719
rect 13163 9685 13197 9719
rect 13231 9685 13265 9719
rect 13299 9685 13333 9719
rect 13367 9685 13401 9719
rect 13435 9685 13469 9719
rect 13503 9685 13537 9719
rect 13571 9685 13605 9719
rect 13639 9685 13673 9719
rect 13707 9685 13741 9719
rect 13775 9685 13809 9719
rect 13843 9685 13877 9719
rect 13911 9685 13945 9719
rect 13979 9685 14013 9719
rect 14047 9685 14081 9719
rect 14115 9685 14149 9719
rect 14183 9685 14217 9719
rect 14251 9685 14285 9719
<< locali >>
rect 589 36191 14417 36221
rect 589 36157 719 36191
rect 753 36157 787 36191
rect 821 36157 855 36191
rect 889 36157 923 36191
rect 957 36157 991 36191
rect 1025 36157 1059 36191
rect 1093 36157 1127 36191
rect 1161 36157 1195 36191
rect 1229 36157 1263 36191
rect 1297 36157 1331 36191
rect 1365 36157 1399 36191
rect 1433 36157 1467 36191
rect 1501 36157 1535 36191
rect 1569 36157 1603 36191
rect 1637 36157 1671 36191
rect 1705 36157 1739 36191
rect 1773 36157 1807 36191
rect 1841 36157 1875 36191
rect 1909 36157 1943 36191
rect 1977 36157 2011 36191
rect 2045 36157 2079 36191
rect 2113 36157 2147 36191
rect 2181 36157 2215 36191
rect 2249 36157 2283 36191
rect 2317 36157 2351 36191
rect 2385 36157 2419 36191
rect 2453 36157 2487 36191
rect 2521 36157 2555 36191
rect 2589 36157 2623 36191
rect 2657 36157 2691 36191
rect 2725 36157 2759 36191
rect 2793 36157 2827 36191
rect 2861 36157 2895 36191
rect 2929 36157 2963 36191
rect 2997 36157 3031 36191
rect 3065 36157 3099 36191
rect 3133 36157 3167 36191
rect 3201 36157 3235 36191
rect 3269 36157 3303 36191
rect 3337 36157 3371 36191
rect 3405 36157 3439 36191
rect 3473 36157 3507 36191
rect 3541 36157 3575 36191
rect 3609 36157 3643 36191
rect 3677 36157 3711 36191
rect 3745 36157 3779 36191
rect 3813 36157 3847 36191
rect 3881 36157 3915 36191
rect 3949 36157 3983 36191
rect 4017 36157 4051 36191
rect 4085 36157 4119 36191
rect 4153 36157 4187 36191
rect 4221 36157 4255 36191
rect 4289 36157 4323 36191
rect 4357 36157 4391 36191
rect 4425 36157 4459 36191
rect 4493 36157 4527 36191
rect 4561 36157 4595 36191
rect 4629 36157 4663 36191
rect 4697 36157 4731 36191
rect 4765 36157 4799 36191
rect 4833 36157 4867 36191
rect 4901 36157 4935 36191
rect 4969 36157 5003 36191
rect 5037 36157 5071 36191
rect 5105 36157 5139 36191
rect 5173 36157 5207 36191
rect 5241 36157 5275 36191
rect 5309 36157 5343 36191
rect 5377 36157 5411 36191
rect 5445 36157 5479 36191
rect 5513 36157 5547 36191
rect 5581 36157 5615 36191
rect 5649 36157 5683 36191
rect 5717 36157 5751 36191
rect 5785 36157 5819 36191
rect 5853 36157 5887 36191
rect 5921 36157 5955 36191
rect 5989 36157 6023 36191
rect 6057 36157 6091 36191
rect 6125 36157 6159 36191
rect 6193 36157 6227 36191
rect 6261 36157 6295 36191
rect 6329 36157 6363 36191
rect 6397 36157 6431 36191
rect 6465 36157 6499 36191
rect 6533 36157 6567 36191
rect 6601 36157 6635 36191
rect 6669 36157 6703 36191
rect 6737 36157 6771 36191
rect 6805 36157 6839 36191
rect 6873 36157 6907 36191
rect 6941 36157 6975 36191
rect 7009 36157 7043 36191
rect 7077 36157 7111 36191
rect 7145 36157 7179 36191
rect 7213 36157 7247 36191
rect 7281 36157 7315 36191
rect 7349 36157 7383 36191
rect 7417 36157 7451 36191
rect 7485 36157 7519 36191
rect 7553 36157 7587 36191
rect 7621 36157 7655 36191
rect 7689 36157 7723 36191
rect 7757 36157 7791 36191
rect 7825 36157 7859 36191
rect 7893 36157 7927 36191
rect 7961 36157 7995 36191
rect 8029 36157 8063 36191
rect 8097 36157 8131 36191
rect 8165 36157 8199 36191
rect 8233 36157 8267 36191
rect 8301 36157 8335 36191
rect 8369 36157 8403 36191
rect 8437 36157 8471 36191
rect 8505 36157 8539 36191
rect 8573 36157 8607 36191
rect 8641 36157 8675 36191
rect 8709 36157 8743 36191
rect 8777 36157 8811 36191
rect 8845 36157 8879 36191
rect 8913 36157 8947 36191
rect 8981 36157 9015 36191
rect 9049 36157 9083 36191
rect 9117 36157 9151 36191
rect 9185 36157 9219 36191
rect 9253 36157 9287 36191
rect 9321 36157 9355 36191
rect 9389 36157 9423 36191
rect 9457 36157 9491 36191
rect 9525 36157 9559 36191
rect 9593 36157 9627 36191
rect 9661 36157 9695 36191
rect 9729 36157 9763 36191
rect 9797 36157 9831 36191
rect 9865 36157 9899 36191
rect 9933 36157 9967 36191
rect 10001 36157 10035 36191
rect 10069 36157 10103 36191
rect 10137 36157 10171 36191
rect 10205 36157 10239 36191
rect 10273 36157 10307 36191
rect 10341 36157 10375 36191
rect 10409 36157 10443 36191
rect 10477 36157 10511 36191
rect 10545 36157 10579 36191
rect 10613 36157 10647 36191
rect 10681 36157 10715 36191
rect 10749 36157 10783 36191
rect 10817 36157 10851 36191
rect 10885 36157 10919 36191
rect 10953 36157 10987 36191
rect 11021 36157 11055 36191
rect 11089 36157 11123 36191
rect 11157 36157 11191 36191
rect 11225 36157 11259 36191
rect 11293 36157 11327 36191
rect 11361 36157 11395 36191
rect 11429 36157 11463 36191
rect 11497 36157 11531 36191
rect 11565 36157 11599 36191
rect 11633 36157 11667 36191
rect 11701 36157 11735 36191
rect 11769 36157 11803 36191
rect 11837 36157 11871 36191
rect 11905 36157 11939 36191
rect 11973 36157 12007 36191
rect 12041 36157 12075 36191
rect 12109 36157 12143 36191
rect 12177 36157 12211 36191
rect 12245 36157 12279 36191
rect 12313 36157 12347 36191
rect 12381 36157 12415 36191
rect 12449 36157 12483 36191
rect 12517 36157 12551 36191
rect 12585 36157 12619 36191
rect 12653 36157 12687 36191
rect 12721 36157 12755 36191
rect 12789 36157 12823 36191
rect 12857 36157 12891 36191
rect 12925 36157 12959 36191
rect 12993 36157 13027 36191
rect 13061 36157 13095 36191
rect 13129 36157 13163 36191
rect 13197 36157 13231 36191
rect 13265 36157 13299 36191
rect 13333 36157 13367 36191
rect 13401 36157 13435 36191
rect 13469 36157 13503 36191
rect 13537 36157 13571 36191
rect 13605 36157 13639 36191
rect 13673 36157 13707 36191
rect 13741 36157 13775 36191
rect 13809 36157 13843 36191
rect 13877 36157 13911 36191
rect 13945 36157 13979 36191
rect 14013 36157 14047 36191
rect 14081 36157 14115 36191
rect 14149 36157 14183 36191
rect 14217 36157 14251 36191
rect 14285 36157 14417 36191
rect 589 36127 14417 36157
rect 589 36079 681 36127
rect 589 36045 618 36079
rect 652 36045 681 36079
rect 589 36011 681 36045
rect 589 35977 618 36011
rect 652 35977 681 36011
rect 589 35943 681 35977
rect 589 35909 618 35943
rect 652 35909 681 35943
rect 589 35875 681 35909
rect 589 35841 618 35875
rect 652 35841 681 35875
rect 589 35807 681 35841
rect 589 35773 618 35807
rect 652 35773 681 35807
rect 589 35739 681 35773
rect 589 35705 618 35739
rect 652 35705 681 35739
rect 589 35671 681 35705
rect 589 35637 618 35671
rect 652 35637 681 35671
rect 589 35603 681 35637
rect 589 35569 618 35603
rect 652 35569 681 35603
rect 589 35535 681 35569
rect 589 35501 618 35535
rect 652 35501 681 35535
rect 589 35467 681 35501
rect 589 35433 618 35467
rect 652 35433 681 35467
rect 589 35399 681 35433
rect 589 35365 618 35399
rect 652 35365 681 35399
rect 589 35331 681 35365
rect 589 35297 618 35331
rect 652 35297 681 35331
rect 589 35263 681 35297
rect 589 35229 618 35263
rect 652 35229 681 35263
rect 589 35195 681 35229
rect 589 35161 618 35195
rect 652 35161 681 35195
rect 589 35127 681 35161
rect 589 35093 618 35127
rect 652 35093 681 35127
rect 589 35059 681 35093
rect 589 35025 618 35059
rect 652 35025 681 35059
rect 589 34991 681 35025
rect 589 34957 618 34991
rect 652 34957 681 34991
rect 589 34923 681 34957
rect 589 34889 618 34923
rect 652 34889 681 34923
rect 589 34855 681 34889
rect 589 34821 618 34855
rect 652 34821 681 34855
rect 589 34787 681 34821
rect 589 34753 618 34787
rect 652 34753 681 34787
rect 589 34719 681 34753
rect 589 34685 618 34719
rect 652 34685 681 34719
rect 589 34651 681 34685
rect 589 34617 618 34651
rect 652 34617 681 34651
rect 589 34583 681 34617
rect 589 34549 618 34583
rect 652 34549 681 34583
rect 589 34515 681 34549
rect 589 34481 618 34515
rect 652 34481 681 34515
rect 589 34447 681 34481
rect 589 34413 618 34447
rect 652 34413 681 34447
rect 589 34379 681 34413
rect 589 34345 618 34379
rect 652 34345 681 34379
rect 589 34311 681 34345
rect 589 34277 618 34311
rect 652 34277 681 34311
rect 589 34243 681 34277
rect 589 34209 618 34243
rect 652 34209 681 34243
rect 589 34175 681 34209
rect 589 34141 618 34175
rect 652 34141 681 34175
rect 589 34107 681 34141
rect 589 34073 618 34107
rect 652 34073 681 34107
rect 589 34039 681 34073
rect 589 34005 618 34039
rect 652 34005 681 34039
rect 589 33971 681 34005
rect 589 33937 618 33971
rect 652 33937 681 33971
rect 589 33903 681 33937
rect 589 33869 618 33903
rect 652 33869 681 33903
rect 589 33835 681 33869
rect 589 33801 618 33835
rect 652 33801 681 33835
rect 589 33767 681 33801
rect 589 33733 618 33767
rect 652 33733 681 33767
rect 589 33699 681 33733
rect 589 33665 618 33699
rect 652 33665 681 33699
rect 589 33631 681 33665
rect 589 33597 618 33631
rect 652 33597 681 33631
rect 589 33563 681 33597
rect 589 33529 618 33563
rect 652 33529 681 33563
rect 589 33495 681 33529
rect 589 33461 618 33495
rect 652 33461 681 33495
rect 589 33427 681 33461
rect 589 33393 618 33427
rect 652 33393 681 33427
rect 589 33359 681 33393
rect 589 33325 618 33359
rect 652 33325 681 33359
rect 589 33291 681 33325
rect 589 33257 618 33291
rect 652 33257 681 33291
rect 589 33223 681 33257
rect 589 33189 618 33223
rect 652 33189 681 33223
rect 589 33155 681 33189
rect 589 33121 618 33155
rect 652 33121 681 33155
rect 589 33087 681 33121
rect 589 33053 618 33087
rect 652 33053 681 33087
rect 589 33019 681 33053
rect 589 32985 618 33019
rect 652 32985 681 33019
rect 589 32951 681 32985
rect 589 32917 618 32951
rect 652 32917 681 32951
rect 589 32883 681 32917
rect 589 32849 618 32883
rect 652 32849 681 32883
rect 589 32815 681 32849
rect 589 32781 618 32815
rect 652 32781 681 32815
rect 589 32747 681 32781
rect 589 32713 618 32747
rect 652 32713 681 32747
rect 589 32679 681 32713
rect 589 32645 618 32679
rect 652 32645 681 32679
rect 589 32611 681 32645
rect 589 32577 618 32611
rect 652 32577 681 32611
rect 589 32543 681 32577
rect 589 32509 618 32543
rect 652 32509 681 32543
rect 589 32475 681 32509
rect 589 32441 618 32475
rect 652 32441 681 32475
rect 589 32407 681 32441
rect 589 32373 618 32407
rect 652 32373 681 32407
rect 589 32339 681 32373
rect 589 32305 618 32339
rect 652 32305 681 32339
rect 589 32271 681 32305
rect 589 32237 618 32271
rect 652 32237 681 32271
rect 589 32203 681 32237
rect 589 32169 618 32203
rect 652 32169 681 32203
rect 589 32135 681 32169
rect 589 32101 618 32135
rect 652 32101 681 32135
rect 589 32067 681 32101
rect 589 32033 618 32067
rect 652 32033 681 32067
rect 589 31999 681 32033
rect 589 31965 618 31999
rect 652 31965 681 31999
rect 589 31931 681 31965
rect 589 31897 618 31931
rect 652 31897 681 31931
rect 589 31863 681 31897
rect 589 31829 618 31863
rect 652 31829 681 31863
rect 589 31795 681 31829
rect 589 31761 618 31795
rect 652 31761 681 31795
rect 589 31727 681 31761
rect 589 31693 618 31727
rect 652 31693 681 31727
rect 589 31659 681 31693
rect 589 31625 618 31659
rect 652 31625 681 31659
rect 589 31591 681 31625
rect 589 31557 618 31591
rect 652 31557 681 31591
rect 589 31523 681 31557
rect 589 31489 618 31523
rect 652 31489 681 31523
rect 589 31455 681 31489
rect 589 31421 618 31455
rect 652 31421 681 31455
rect 589 31387 681 31421
rect 589 31353 618 31387
rect 652 31353 681 31387
rect 589 31319 681 31353
rect 589 31285 618 31319
rect 652 31285 681 31319
rect 589 31251 681 31285
rect 589 31217 618 31251
rect 652 31217 681 31251
rect 589 31183 681 31217
rect 589 31149 618 31183
rect 652 31149 681 31183
rect 589 31115 681 31149
rect 589 31081 618 31115
rect 652 31081 681 31115
rect 589 31047 681 31081
rect 589 31013 618 31047
rect 652 31013 681 31047
rect 589 30979 681 31013
rect 589 30945 618 30979
rect 652 30945 681 30979
rect 589 30911 681 30945
rect 589 30877 618 30911
rect 652 30877 681 30911
rect 589 30843 681 30877
rect 589 30809 618 30843
rect 652 30809 681 30843
rect 589 30775 681 30809
rect 589 30741 618 30775
rect 652 30741 681 30775
rect 589 30707 681 30741
rect 589 30673 618 30707
rect 652 30673 681 30707
rect 589 30639 681 30673
rect 589 30605 618 30639
rect 652 30605 681 30639
rect 589 30571 681 30605
rect 589 30537 618 30571
rect 652 30537 681 30571
rect 589 30503 681 30537
rect 589 30469 618 30503
rect 652 30469 681 30503
rect 589 30435 681 30469
rect 589 30401 618 30435
rect 652 30401 681 30435
rect 589 30367 681 30401
rect 589 30333 618 30367
rect 652 30333 681 30367
rect 589 30299 681 30333
rect 589 30265 618 30299
rect 652 30265 681 30299
rect 589 30231 681 30265
rect 589 30197 618 30231
rect 652 30197 681 30231
rect 589 30163 681 30197
rect 589 30129 618 30163
rect 652 30129 681 30163
rect 589 30095 681 30129
rect 589 30061 618 30095
rect 652 30061 681 30095
rect 589 30027 681 30061
rect 589 29993 618 30027
rect 652 29993 681 30027
rect 589 29959 681 29993
rect 589 29925 618 29959
rect 652 29925 681 29959
rect 589 29891 681 29925
rect 589 29857 618 29891
rect 652 29857 681 29891
rect 589 29823 681 29857
rect 589 29789 618 29823
rect 652 29789 681 29823
rect 589 29755 681 29789
rect 589 29721 618 29755
rect 652 29721 681 29755
rect 589 29687 681 29721
rect 589 29653 618 29687
rect 652 29653 681 29687
rect 589 29619 681 29653
rect 589 29585 618 29619
rect 652 29585 681 29619
rect 589 29551 681 29585
rect 589 29517 618 29551
rect 652 29517 681 29551
rect 589 29483 681 29517
rect 589 29449 618 29483
rect 652 29449 681 29483
rect 589 29415 681 29449
rect 589 29381 618 29415
rect 652 29381 681 29415
rect 589 29347 681 29381
rect 589 29313 618 29347
rect 652 29313 681 29347
rect 589 29279 681 29313
rect 589 29245 618 29279
rect 652 29245 681 29279
rect 589 29211 681 29245
rect 589 29177 618 29211
rect 652 29177 681 29211
rect 589 29143 681 29177
rect 589 29109 618 29143
rect 652 29109 681 29143
rect 589 29075 681 29109
rect 589 29041 618 29075
rect 652 29041 681 29075
rect 589 29007 681 29041
rect 589 28973 618 29007
rect 652 28973 681 29007
rect 589 28939 681 28973
rect 589 28905 618 28939
rect 652 28905 681 28939
rect 589 28871 681 28905
rect 589 28837 618 28871
rect 652 28837 681 28871
rect 589 28803 681 28837
rect 589 28769 618 28803
rect 652 28769 681 28803
rect 589 28735 681 28769
rect 589 28701 618 28735
rect 652 28701 681 28735
rect 589 28667 681 28701
rect 589 28633 618 28667
rect 652 28633 681 28667
rect 589 28599 681 28633
rect 589 28565 618 28599
rect 652 28565 681 28599
rect 589 28531 681 28565
rect 589 28497 618 28531
rect 652 28497 681 28531
rect 589 28463 681 28497
rect 589 28429 618 28463
rect 652 28429 681 28463
rect 589 28395 681 28429
rect 589 28361 618 28395
rect 652 28361 681 28395
rect 589 28327 681 28361
rect 589 28293 618 28327
rect 652 28293 681 28327
rect 589 28259 681 28293
rect 589 28225 618 28259
rect 652 28225 681 28259
rect 589 28191 681 28225
rect 589 28157 618 28191
rect 652 28157 681 28191
rect 589 28123 681 28157
rect 589 28089 618 28123
rect 652 28089 681 28123
rect 589 28055 681 28089
rect 589 28021 618 28055
rect 652 28021 681 28055
rect 589 27987 681 28021
rect 589 27953 618 27987
rect 652 27953 681 27987
rect 589 27919 681 27953
rect 589 27885 618 27919
rect 652 27885 681 27919
rect 589 27851 681 27885
rect 589 27817 618 27851
rect 652 27817 681 27851
rect 589 27783 681 27817
rect 589 27749 618 27783
rect 652 27749 681 27783
rect 589 27715 681 27749
rect 589 27681 618 27715
rect 652 27681 681 27715
rect 589 27647 681 27681
rect 589 27613 618 27647
rect 652 27613 681 27647
rect 589 27579 681 27613
rect 589 27545 618 27579
rect 652 27545 681 27579
rect 589 27511 681 27545
rect 589 27477 618 27511
rect 652 27477 681 27511
rect 589 27443 681 27477
rect 589 27409 618 27443
rect 652 27409 681 27443
rect 589 27375 681 27409
rect 589 27341 618 27375
rect 652 27341 681 27375
rect 589 27307 681 27341
rect 589 27273 618 27307
rect 652 27273 681 27307
rect 589 27239 681 27273
rect 589 27205 618 27239
rect 652 27205 681 27239
rect 589 27171 681 27205
rect 589 27137 618 27171
rect 652 27137 681 27171
rect 589 27103 681 27137
rect 589 27069 618 27103
rect 652 27069 681 27103
rect 589 27035 681 27069
rect 589 27001 618 27035
rect 652 27001 681 27035
rect 589 26967 681 27001
rect 589 26933 618 26967
rect 652 26933 681 26967
rect 589 26899 681 26933
rect 589 26865 618 26899
rect 652 26865 681 26899
rect 589 26831 681 26865
rect 589 26797 618 26831
rect 652 26797 681 26831
rect 589 26763 681 26797
rect 589 26729 618 26763
rect 652 26729 681 26763
rect 589 26695 681 26729
rect 589 26661 618 26695
rect 652 26661 681 26695
rect 589 26627 681 26661
rect 589 26593 618 26627
rect 652 26593 681 26627
rect 589 26559 681 26593
rect 589 26525 618 26559
rect 652 26525 681 26559
rect 589 26491 681 26525
rect 589 26457 618 26491
rect 652 26457 681 26491
rect 589 26423 681 26457
rect 589 26389 618 26423
rect 652 26389 681 26423
rect 589 26355 681 26389
rect 589 26321 618 26355
rect 652 26321 681 26355
rect 589 26287 681 26321
rect 589 26253 618 26287
rect 652 26253 681 26287
rect 589 26219 681 26253
rect 589 26185 618 26219
rect 652 26185 681 26219
rect 589 26151 681 26185
rect 589 26117 618 26151
rect 652 26117 681 26151
rect 589 26083 681 26117
rect 589 26049 618 26083
rect 652 26049 681 26083
rect 589 26015 681 26049
rect 589 25981 618 26015
rect 652 25981 681 26015
rect 589 25947 681 25981
rect 589 25913 618 25947
rect 652 25913 681 25947
rect 589 25879 681 25913
rect 589 25845 618 25879
rect 652 25845 681 25879
rect 589 25811 681 25845
rect 589 25777 618 25811
rect 652 25777 681 25811
rect 589 25743 681 25777
rect 589 25709 618 25743
rect 652 25709 681 25743
rect 589 25675 681 25709
rect 589 25641 618 25675
rect 652 25641 681 25675
rect 589 25607 681 25641
rect 589 25573 618 25607
rect 652 25573 681 25607
rect 589 25539 681 25573
rect 589 25505 618 25539
rect 652 25505 681 25539
rect 589 25471 681 25505
rect 589 25437 618 25471
rect 652 25437 681 25471
rect 589 25403 681 25437
rect 589 25369 618 25403
rect 652 25369 681 25403
rect 589 25335 681 25369
rect 589 25301 618 25335
rect 652 25301 681 25335
rect 589 25267 681 25301
rect 589 25233 618 25267
rect 652 25233 681 25267
rect 589 25199 681 25233
rect 589 25165 618 25199
rect 652 25165 681 25199
rect 589 25131 681 25165
rect 589 25097 618 25131
rect 652 25097 681 25131
rect 589 25063 681 25097
rect 589 25029 618 25063
rect 652 25029 681 25063
rect 589 24995 681 25029
rect 589 24961 618 24995
rect 652 24961 681 24995
rect 589 24927 681 24961
rect 589 24893 618 24927
rect 652 24893 681 24927
rect 589 24859 681 24893
rect 589 24825 618 24859
rect 652 24825 681 24859
rect 589 24791 681 24825
rect 589 24757 618 24791
rect 652 24757 681 24791
rect 589 24723 681 24757
rect 589 24689 618 24723
rect 652 24689 681 24723
rect 589 24655 681 24689
rect 589 24621 618 24655
rect 652 24621 681 24655
rect 589 24587 681 24621
rect 589 24553 618 24587
rect 652 24553 681 24587
rect 589 24519 681 24553
rect 589 24485 618 24519
rect 652 24485 681 24519
rect 589 24451 681 24485
rect 589 24417 618 24451
rect 652 24417 681 24451
rect 589 24383 681 24417
rect 589 24349 618 24383
rect 652 24349 681 24383
rect 589 24315 681 24349
rect 589 24281 618 24315
rect 652 24281 681 24315
rect 589 24247 681 24281
rect 589 24213 618 24247
rect 652 24213 681 24247
rect 589 24179 681 24213
rect 589 24145 618 24179
rect 652 24145 681 24179
rect 589 24111 681 24145
rect 589 24077 618 24111
rect 652 24077 681 24111
rect 589 24043 681 24077
rect 589 24009 618 24043
rect 652 24009 681 24043
rect 589 23975 681 24009
rect 589 23941 618 23975
rect 652 23941 681 23975
rect 589 23907 681 23941
rect 589 23873 618 23907
rect 652 23873 681 23907
rect 589 23839 681 23873
rect 589 23805 618 23839
rect 652 23805 681 23839
rect 589 23771 681 23805
rect 589 23737 618 23771
rect 652 23737 681 23771
rect 589 23703 681 23737
rect 589 23669 618 23703
rect 652 23669 681 23703
rect 589 23635 681 23669
rect 589 23601 618 23635
rect 652 23601 681 23635
rect 589 23567 681 23601
rect 589 23533 618 23567
rect 652 23533 681 23567
rect 589 23499 681 23533
rect 589 23465 618 23499
rect 652 23465 681 23499
rect 589 23431 681 23465
rect 589 23397 618 23431
rect 652 23397 681 23431
rect 589 23363 681 23397
rect 589 23329 618 23363
rect 652 23329 681 23363
rect 589 23295 681 23329
rect 589 23261 618 23295
rect 652 23261 681 23295
rect 589 23227 681 23261
rect 589 23193 618 23227
rect 652 23193 681 23227
rect 589 23159 681 23193
rect 589 23125 618 23159
rect 652 23125 681 23159
rect 589 23091 681 23125
rect 589 23057 618 23091
rect 652 23057 681 23091
rect 589 23023 681 23057
rect 589 22989 618 23023
rect 652 22989 681 23023
rect 589 22955 681 22989
rect 589 22921 618 22955
rect 652 22921 681 22955
rect 589 22887 681 22921
rect 589 22853 618 22887
rect 652 22853 681 22887
rect 589 22819 681 22853
rect 589 22785 618 22819
rect 652 22785 681 22819
rect 589 22751 681 22785
rect 589 22717 618 22751
rect 652 22717 681 22751
rect 589 22683 681 22717
rect 589 22649 618 22683
rect 652 22649 681 22683
rect 589 22615 681 22649
rect 589 22581 618 22615
rect 652 22581 681 22615
rect 589 22547 681 22581
rect 589 22513 618 22547
rect 652 22513 681 22547
rect 589 22479 681 22513
rect 589 22445 618 22479
rect 652 22445 681 22479
rect 589 22411 681 22445
rect 589 22377 618 22411
rect 652 22377 681 22411
rect 589 22343 681 22377
rect 589 22309 618 22343
rect 652 22309 681 22343
rect 589 22275 681 22309
rect 589 22241 618 22275
rect 652 22241 681 22275
rect 589 22207 681 22241
rect 589 22173 618 22207
rect 652 22173 681 22207
rect 589 22139 681 22173
rect 589 22105 618 22139
rect 652 22105 681 22139
rect 589 22071 681 22105
rect 589 22037 618 22071
rect 652 22037 681 22071
rect 589 22003 681 22037
rect 589 21969 618 22003
rect 652 21969 681 22003
rect 589 21935 681 21969
rect 589 21901 618 21935
rect 652 21901 681 21935
rect 589 21867 681 21901
rect 589 21833 618 21867
rect 652 21833 681 21867
rect 589 21799 681 21833
rect 589 21765 618 21799
rect 652 21765 681 21799
rect 589 21731 681 21765
rect 589 21697 618 21731
rect 652 21697 681 21731
rect 589 21663 681 21697
rect 589 21629 618 21663
rect 652 21629 681 21663
rect 589 21595 681 21629
rect 589 21561 618 21595
rect 652 21561 681 21595
rect 589 21527 681 21561
rect 589 21493 618 21527
rect 652 21493 681 21527
rect 589 21459 681 21493
rect 589 21425 618 21459
rect 652 21425 681 21459
rect 589 21391 681 21425
rect 589 21357 618 21391
rect 652 21357 681 21391
rect 589 21323 681 21357
rect 589 21289 618 21323
rect 652 21289 681 21323
rect 589 21255 681 21289
rect 589 21221 618 21255
rect 652 21221 681 21255
rect 589 21187 681 21221
rect 589 21153 618 21187
rect 652 21153 681 21187
rect 589 21119 681 21153
rect 589 21085 618 21119
rect 652 21085 681 21119
rect 589 21051 681 21085
rect 589 21017 618 21051
rect 652 21017 681 21051
rect 589 20983 681 21017
rect 589 20949 618 20983
rect 652 20949 681 20983
rect 589 20915 681 20949
rect 589 20881 618 20915
rect 652 20881 681 20915
rect 589 20847 681 20881
rect 589 20813 618 20847
rect 652 20813 681 20847
rect 589 20779 681 20813
rect 589 20745 618 20779
rect 652 20745 681 20779
rect 589 20711 681 20745
rect 589 20677 618 20711
rect 652 20677 681 20711
rect 589 20643 681 20677
rect 589 20609 618 20643
rect 652 20609 681 20643
rect 589 20575 681 20609
rect 589 20541 618 20575
rect 652 20541 681 20575
rect 589 20507 681 20541
rect 589 20473 618 20507
rect 652 20473 681 20507
rect 589 20439 681 20473
rect 589 20405 618 20439
rect 652 20405 681 20439
rect 589 20371 681 20405
rect 589 20337 618 20371
rect 652 20337 681 20371
rect 589 20303 681 20337
rect 589 20269 618 20303
rect 652 20269 681 20303
rect 589 20235 681 20269
rect 589 20201 618 20235
rect 652 20201 681 20235
rect 589 20167 681 20201
rect 589 20133 618 20167
rect 652 20133 681 20167
rect 589 20099 681 20133
rect 589 20065 618 20099
rect 652 20065 681 20099
rect 589 20031 681 20065
rect 589 19997 618 20031
rect 652 19997 681 20031
rect 589 19963 681 19997
rect 589 19929 618 19963
rect 652 19929 681 19963
rect 589 19895 681 19929
rect 589 19861 618 19895
rect 652 19861 681 19895
rect 589 19827 681 19861
rect 589 19793 618 19827
rect 652 19793 681 19827
rect 589 19759 681 19793
rect 589 19725 618 19759
rect 652 19725 681 19759
rect 589 19691 681 19725
rect 589 19657 618 19691
rect 652 19657 681 19691
rect 589 19623 681 19657
rect 589 19589 618 19623
rect 652 19589 681 19623
rect 589 19555 681 19589
rect 589 19521 618 19555
rect 652 19521 681 19555
rect 589 19487 681 19521
rect 589 19453 618 19487
rect 652 19453 681 19487
rect 589 19419 681 19453
rect 589 19385 618 19419
rect 652 19385 681 19419
rect 589 19351 681 19385
rect 589 19317 618 19351
rect 652 19317 681 19351
rect 589 19283 681 19317
rect 589 19249 618 19283
rect 652 19249 681 19283
rect 589 19215 681 19249
rect 589 19181 618 19215
rect 652 19181 681 19215
rect 589 19147 681 19181
rect 589 19113 618 19147
rect 652 19113 681 19147
rect 589 19079 681 19113
rect 589 19045 618 19079
rect 652 19045 681 19079
rect 589 19011 681 19045
rect 589 18977 618 19011
rect 652 18977 681 19011
rect 589 18943 681 18977
rect 589 18909 618 18943
rect 652 18909 681 18943
rect 589 18875 681 18909
rect 589 18841 618 18875
rect 652 18841 681 18875
rect 589 18807 681 18841
rect 589 18773 618 18807
rect 652 18773 681 18807
rect 589 18739 681 18773
rect 589 18705 618 18739
rect 652 18705 681 18739
rect 589 18671 681 18705
rect 589 18637 618 18671
rect 652 18637 681 18671
rect 589 18603 681 18637
rect 589 18569 618 18603
rect 652 18569 681 18603
rect 589 18535 681 18569
rect 589 18501 618 18535
rect 652 18501 681 18535
rect 589 18467 681 18501
rect 589 18433 618 18467
rect 652 18433 681 18467
rect 589 18399 681 18433
rect 589 18365 618 18399
rect 652 18365 681 18399
rect 589 18331 681 18365
rect 589 18297 618 18331
rect 652 18297 681 18331
rect 589 18263 681 18297
rect 589 18229 618 18263
rect 652 18229 681 18263
rect 589 18195 681 18229
rect 589 18161 618 18195
rect 652 18161 681 18195
rect 589 18127 681 18161
rect 589 18093 618 18127
rect 652 18093 681 18127
rect 589 18059 681 18093
rect 589 18025 618 18059
rect 652 18025 681 18059
rect 589 17991 681 18025
rect 589 17957 618 17991
rect 652 17957 681 17991
rect 589 17923 681 17957
rect 589 17889 618 17923
rect 652 17889 681 17923
rect 589 17855 681 17889
rect 589 17821 618 17855
rect 652 17821 681 17855
rect 589 17787 681 17821
rect 589 17753 618 17787
rect 652 17753 681 17787
rect 589 17719 681 17753
rect 589 17685 618 17719
rect 652 17685 681 17719
rect 589 17651 681 17685
rect 589 17617 618 17651
rect 652 17617 681 17651
rect 589 17583 681 17617
rect 589 17549 618 17583
rect 652 17549 681 17583
rect 589 17515 681 17549
rect 589 17481 618 17515
rect 652 17481 681 17515
rect 589 17447 681 17481
rect 589 17413 618 17447
rect 652 17413 681 17447
rect 589 17379 681 17413
rect 589 17345 618 17379
rect 652 17345 681 17379
rect 589 17311 681 17345
rect 589 17277 618 17311
rect 652 17277 681 17311
rect 589 17243 681 17277
rect 589 17209 618 17243
rect 652 17209 681 17243
rect 589 17175 681 17209
rect 589 17141 618 17175
rect 652 17141 681 17175
rect 589 17107 681 17141
rect 589 17073 618 17107
rect 652 17073 681 17107
rect 589 17039 681 17073
rect 589 17005 618 17039
rect 652 17005 681 17039
rect 589 16971 681 17005
rect 589 16937 618 16971
rect 652 16937 681 16971
rect 589 16903 681 16937
rect 589 16869 618 16903
rect 652 16869 681 16903
rect 589 16835 681 16869
rect 589 16801 618 16835
rect 652 16801 681 16835
rect 589 16767 681 16801
rect 589 16733 618 16767
rect 652 16733 681 16767
rect 589 16699 681 16733
rect 589 16665 618 16699
rect 652 16665 681 16699
rect 589 16631 681 16665
rect 589 16597 618 16631
rect 652 16597 681 16631
rect 589 16563 681 16597
rect 589 16529 618 16563
rect 652 16529 681 16563
rect 589 16495 681 16529
rect 589 16461 618 16495
rect 652 16461 681 16495
rect 589 16427 681 16461
rect 589 16393 618 16427
rect 652 16393 681 16427
rect 589 16359 681 16393
rect 589 16325 618 16359
rect 652 16325 681 16359
rect 589 16291 681 16325
rect 589 16257 618 16291
rect 652 16257 681 16291
rect 589 16223 681 16257
rect 589 16189 618 16223
rect 652 16189 681 16223
rect 589 16155 681 16189
rect 589 16121 618 16155
rect 652 16121 681 16155
rect 589 16087 681 16121
rect 589 16053 618 16087
rect 652 16053 681 16087
rect 589 16019 681 16053
rect 589 15985 618 16019
rect 652 15985 681 16019
rect 589 15951 681 15985
rect 589 15917 618 15951
rect 652 15917 681 15951
rect 589 15883 681 15917
rect 589 15849 618 15883
rect 652 15849 681 15883
rect 589 15815 681 15849
rect 589 15781 618 15815
rect 652 15781 681 15815
rect 589 15747 681 15781
rect 589 15713 618 15747
rect 652 15713 681 15747
rect 589 15679 681 15713
rect 589 15645 618 15679
rect 652 15645 681 15679
rect 589 15611 681 15645
rect 589 15577 618 15611
rect 652 15577 681 15611
rect 589 15543 681 15577
rect 589 15509 618 15543
rect 652 15509 681 15543
rect 589 15475 681 15509
rect 589 15441 618 15475
rect 652 15441 681 15475
rect 589 15407 681 15441
rect 589 15373 618 15407
rect 652 15373 681 15407
rect 589 15339 681 15373
rect 589 15305 618 15339
rect 652 15305 681 15339
rect 589 15271 681 15305
rect 589 15237 618 15271
rect 652 15237 681 15271
rect 589 15203 681 15237
rect 589 15169 618 15203
rect 652 15169 681 15203
rect 589 15135 681 15169
rect 589 15101 618 15135
rect 652 15101 681 15135
rect 589 15067 681 15101
rect 589 15033 618 15067
rect 652 15033 681 15067
rect 589 14999 681 15033
rect 589 14965 618 14999
rect 652 14965 681 14999
rect 589 14931 681 14965
rect 589 14897 618 14931
rect 652 14897 681 14931
rect 589 14863 681 14897
rect 589 14829 618 14863
rect 652 14829 681 14863
rect 589 14795 681 14829
rect 589 14761 618 14795
rect 652 14761 681 14795
rect 589 14727 681 14761
rect 589 14693 618 14727
rect 652 14693 681 14727
rect 589 14659 681 14693
rect 589 14625 618 14659
rect 652 14625 681 14659
rect 589 14591 681 14625
rect 589 14557 618 14591
rect 652 14557 681 14591
rect 589 14523 681 14557
rect 589 14489 618 14523
rect 652 14489 681 14523
rect 589 14455 681 14489
rect 589 14421 618 14455
rect 652 14421 681 14455
rect 589 14387 681 14421
rect 589 14353 618 14387
rect 652 14353 681 14387
rect 589 14319 681 14353
rect 589 14285 618 14319
rect 652 14285 681 14319
rect 589 14251 681 14285
rect 589 14217 618 14251
rect 652 14217 681 14251
rect 589 14183 681 14217
rect 589 14149 618 14183
rect 652 14149 681 14183
rect 589 14115 681 14149
rect 589 14081 618 14115
rect 652 14081 681 14115
rect 589 14047 681 14081
rect 589 14013 618 14047
rect 652 14013 681 14047
rect 589 13979 681 14013
rect 589 13945 618 13979
rect 652 13945 681 13979
rect 589 13911 681 13945
rect 589 13877 618 13911
rect 652 13877 681 13911
rect 589 13843 681 13877
rect 589 13809 618 13843
rect 652 13809 681 13843
rect 589 13775 681 13809
rect 589 13741 618 13775
rect 652 13741 681 13775
rect 589 13707 681 13741
rect 589 13673 618 13707
rect 652 13673 681 13707
rect 589 13639 681 13673
rect 589 13605 618 13639
rect 652 13605 681 13639
rect 589 13571 681 13605
rect 589 13537 618 13571
rect 652 13537 681 13571
rect 589 13503 681 13537
rect 589 13469 618 13503
rect 652 13469 681 13503
rect 589 13435 681 13469
rect 589 13401 618 13435
rect 652 13401 681 13435
rect 589 13367 681 13401
rect 589 13333 618 13367
rect 652 13333 681 13367
rect 589 13299 681 13333
rect 589 13265 618 13299
rect 652 13265 681 13299
rect 589 13231 681 13265
rect 589 13197 618 13231
rect 652 13197 681 13231
rect 589 13163 681 13197
rect 589 13129 618 13163
rect 652 13129 681 13163
rect 589 13095 681 13129
rect 589 13061 618 13095
rect 652 13061 681 13095
rect 589 13027 681 13061
rect 589 12993 618 13027
rect 652 12993 681 13027
rect 589 12959 681 12993
rect 589 12925 618 12959
rect 652 12925 681 12959
rect 589 12891 681 12925
rect 589 12857 618 12891
rect 652 12857 681 12891
rect 589 12823 681 12857
rect 589 12789 618 12823
rect 652 12789 681 12823
rect 589 12755 681 12789
rect 589 12721 618 12755
rect 652 12721 681 12755
rect 589 12687 681 12721
rect 589 12653 618 12687
rect 652 12653 681 12687
rect 589 12619 681 12653
rect 589 12585 618 12619
rect 652 12585 681 12619
rect 589 12551 681 12585
rect 589 12517 618 12551
rect 652 12517 681 12551
rect 589 12483 681 12517
rect 589 12449 618 12483
rect 652 12449 681 12483
rect 589 12415 681 12449
rect 589 12381 618 12415
rect 652 12381 681 12415
rect 589 12347 681 12381
rect 589 12313 618 12347
rect 652 12313 681 12347
rect 589 12279 681 12313
rect 589 12245 618 12279
rect 652 12245 681 12279
rect 589 12211 681 12245
rect 589 12177 618 12211
rect 652 12177 681 12211
rect 589 12143 681 12177
rect 589 12109 618 12143
rect 652 12109 681 12143
rect 589 12075 681 12109
rect 589 12041 618 12075
rect 652 12041 681 12075
rect 589 12007 681 12041
rect 589 11973 618 12007
rect 652 11973 681 12007
rect 589 11939 681 11973
rect 589 11905 618 11939
rect 652 11905 681 11939
rect 589 11871 681 11905
rect 589 11837 618 11871
rect 652 11837 681 11871
rect 589 11803 681 11837
rect 589 11769 618 11803
rect 652 11769 681 11803
rect 589 11735 681 11769
rect 589 11701 618 11735
rect 652 11701 681 11735
rect 589 11667 681 11701
rect 589 11633 618 11667
rect 652 11633 681 11667
rect 589 11599 681 11633
rect 589 11565 618 11599
rect 652 11565 681 11599
rect 589 11531 681 11565
rect 589 11497 618 11531
rect 652 11497 681 11531
rect 589 11463 681 11497
rect 589 11429 618 11463
rect 652 11429 681 11463
rect 589 11395 681 11429
rect 589 11361 618 11395
rect 652 11361 681 11395
rect 589 11327 681 11361
rect 589 11293 618 11327
rect 652 11293 681 11327
rect 589 11259 681 11293
rect 589 11225 618 11259
rect 652 11225 681 11259
rect 589 11191 681 11225
rect 589 11157 618 11191
rect 652 11157 681 11191
rect 589 11123 681 11157
rect 589 11089 618 11123
rect 652 11089 681 11123
rect 589 11055 681 11089
rect 589 11021 618 11055
rect 652 11021 681 11055
rect 589 10987 681 11021
rect 589 10953 618 10987
rect 652 10953 681 10987
rect 589 10919 681 10953
rect 589 10885 618 10919
rect 652 10885 681 10919
rect 589 10851 681 10885
rect 589 10817 618 10851
rect 652 10817 681 10851
rect 589 10783 681 10817
rect 589 10749 618 10783
rect 652 10749 681 10783
rect 589 10715 681 10749
rect 589 10681 618 10715
rect 652 10681 681 10715
rect 589 10647 681 10681
rect 589 10613 618 10647
rect 652 10613 681 10647
rect 589 10579 681 10613
rect 589 10545 618 10579
rect 652 10545 681 10579
rect 589 10511 681 10545
rect 589 10477 618 10511
rect 652 10477 681 10511
rect 589 10443 681 10477
rect 589 10409 618 10443
rect 652 10409 681 10443
rect 589 10375 681 10409
rect 589 10341 618 10375
rect 652 10341 681 10375
rect 589 10307 681 10341
rect 589 10273 618 10307
rect 652 10273 681 10307
rect 589 10239 681 10273
rect 589 10205 618 10239
rect 652 10205 681 10239
rect 589 10171 681 10205
rect 589 10137 618 10171
rect 652 10137 681 10171
rect 589 10103 681 10137
rect 589 10069 618 10103
rect 652 10069 681 10103
rect 589 10035 681 10069
rect 589 10001 618 10035
rect 652 10001 681 10035
rect 589 9967 681 10001
rect 589 9933 618 9967
rect 652 9933 681 9967
rect 589 9899 681 9933
rect 589 9865 618 9899
rect 652 9865 681 9899
rect 589 9831 681 9865
rect 589 9797 618 9831
rect 652 9797 681 9831
rect 589 9749 681 9797
rect 14323 36079 14417 36127
rect 14323 36045 14353 36079
rect 14387 36045 14417 36079
rect 14323 36011 14417 36045
rect 14323 35977 14353 36011
rect 14387 35977 14417 36011
rect 14323 35943 14417 35977
rect 14323 35909 14353 35943
rect 14387 35909 14417 35943
rect 14323 35875 14417 35909
rect 14323 35841 14353 35875
rect 14387 35841 14417 35875
rect 14323 35807 14417 35841
rect 14323 35773 14353 35807
rect 14387 35773 14417 35807
rect 14323 35739 14417 35773
rect 14323 35705 14353 35739
rect 14387 35705 14417 35739
rect 14323 35671 14417 35705
rect 14323 35637 14353 35671
rect 14387 35637 14417 35671
rect 14323 35603 14417 35637
rect 14323 35569 14353 35603
rect 14387 35569 14417 35603
rect 14323 35535 14417 35569
rect 14323 35501 14353 35535
rect 14387 35501 14417 35535
rect 14323 35467 14417 35501
rect 14323 35433 14353 35467
rect 14387 35433 14417 35467
rect 14323 35399 14417 35433
rect 14323 35365 14353 35399
rect 14387 35365 14417 35399
rect 14323 35331 14417 35365
rect 14323 35297 14353 35331
rect 14387 35297 14417 35331
rect 14323 35263 14417 35297
rect 14323 35229 14353 35263
rect 14387 35229 14417 35263
rect 14323 35195 14417 35229
rect 14323 35161 14353 35195
rect 14387 35161 14417 35195
rect 14323 35127 14417 35161
rect 14323 35093 14353 35127
rect 14387 35093 14417 35127
rect 14323 35059 14417 35093
rect 14323 35025 14353 35059
rect 14387 35025 14417 35059
rect 14323 34991 14417 35025
rect 14323 34957 14353 34991
rect 14387 34957 14417 34991
rect 14323 34923 14417 34957
rect 14323 34889 14353 34923
rect 14387 34889 14417 34923
rect 14323 34855 14417 34889
rect 14323 34821 14353 34855
rect 14387 34821 14417 34855
rect 14323 34787 14417 34821
rect 14323 34753 14353 34787
rect 14387 34753 14417 34787
rect 14323 34719 14417 34753
rect 14323 34685 14353 34719
rect 14387 34685 14417 34719
rect 14323 34651 14417 34685
rect 14323 34617 14353 34651
rect 14387 34617 14417 34651
rect 14323 34583 14417 34617
rect 14323 34549 14353 34583
rect 14387 34549 14417 34583
rect 14323 34515 14417 34549
rect 14323 34481 14353 34515
rect 14387 34481 14417 34515
rect 14323 34447 14417 34481
rect 14323 34413 14353 34447
rect 14387 34413 14417 34447
rect 14323 34379 14417 34413
rect 14323 34345 14353 34379
rect 14387 34345 14417 34379
rect 14323 34311 14417 34345
rect 14323 34277 14353 34311
rect 14387 34277 14417 34311
rect 14323 34243 14417 34277
rect 14323 34209 14353 34243
rect 14387 34209 14417 34243
rect 14323 34175 14417 34209
rect 14323 34141 14353 34175
rect 14387 34141 14417 34175
rect 14323 34107 14417 34141
rect 14323 34073 14353 34107
rect 14387 34073 14417 34107
rect 14323 34039 14417 34073
rect 14323 34005 14353 34039
rect 14387 34005 14417 34039
rect 14323 33971 14417 34005
rect 14323 33937 14353 33971
rect 14387 33937 14417 33971
rect 14323 33903 14417 33937
rect 14323 33869 14353 33903
rect 14387 33869 14417 33903
rect 14323 33835 14417 33869
rect 14323 33801 14353 33835
rect 14387 33801 14417 33835
rect 14323 33767 14417 33801
rect 14323 33733 14353 33767
rect 14387 33733 14417 33767
rect 14323 33699 14417 33733
rect 14323 33665 14353 33699
rect 14387 33665 14417 33699
rect 14323 33631 14417 33665
rect 14323 33597 14353 33631
rect 14387 33597 14417 33631
rect 14323 33563 14417 33597
rect 14323 33529 14353 33563
rect 14387 33529 14417 33563
rect 14323 33495 14417 33529
rect 14323 33461 14353 33495
rect 14387 33461 14417 33495
rect 14323 33427 14417 33461
rect 14323 33393 14353 33427
rect 14387 33393 14417 33427
rect 14323 33359 14417 33393
rect 14323 33325 14353 33359
rect 14387 33325 14417 33359
rect 14323 33291 14417 33325
rect 14323 33257 14353 33291
rect 14387 33257 14417 33291
rect 14323 33223 14417 33257
rect 14323 33189 14353 33223
rect 14387 33189 14417 33223
rect 14323 33155 14417 33189
rect 14323 33121 14353 33155
rect 14387 33121 14417 33155
rect 14323 33087 14417 33121
rect 14323 33053 14353 33087
rect 14387 33053 14417 33087
rect 14323 33019 14417 33053
rect 14323 32985 14353 33019
rect 14387 32985 14417 33019
rect 14323 32951 14417 32985
rect 14323 32917 14353 32951
rect 14387 32917 14417 32951
rect 14323 32883 14417 32917
rect 14323 32849 14353 32883
rect 14387 32849 14417 32883
rect 14323 32815 14417 32849
rect 14323 32781 14353 32815
rect 14387 32781 14417 32815
rect 14323 32747 14417 32781
rect 14323 32713 14353 32747
rect 14387 32713 14417 32747
rect 14323 32679 14417 32713
rect 14323 32645 14353 32679
rect 14387 32645 14417 32679
rect 14323 32611 14417 32645
rect 14323 32577 14353 32611
rect 14387 32577 14417 32611
rect 14323 32543 14417 32577
rect 14323 32509 14353 32543
rect 14387 32509 14417 32543
rect 14323 32475 14417 32509
rect 14323 32441 14353 32475
rect 14387 32441 14417 32475
rect 14323 32407 14417 32441
rect 14323 32373 14353 32407
rect 14387 32373 14417 32407
rect 14323 32339 14417 32373
rect 14323 32305 14353 32339
rect 14387 32305 14417 32339
rect 14323 32271 14417 32305
rect 14323 32237 14353 32271
rect 14387 32237 14417 32271
rect 14323 32203 14417 32237
rect 14323 32169 14353 32203
rect 14387 32169 14417 32203
rect 14323 32135 14417 32169
rect 14323 32101 14353 32135
rect 14387 32101 14417 32135
rect 14323 32067 14417 32101
rect 14323 32033 14353 32067
rect 14387 32033 14417 32067
rect 14323 31999 14417 32033
rect 14323 31965 14353 31999
rect 14387 31965 14417 31999
rect 14323 31931 14417 31965
rect 14323 31897 14353 31931
rect 14387 31897 14417 31931
rect 14323 31863 14417 31897
rect 14323 31829 14353 31863
rect 14387 31829 14417 31863
rect 14323 31795 14417 31829
rect 14323 31761 14353 31795
rect 14387 31761 14417 31795
rect 14323 31727 14417 31761
rect 14323 31693 14353 31727
rect 14387 31693 14417 31727
rect 14323 31659 14417 31693
rect 14323 31625 14353 31659
rect 14387 31625 14417 31659
rect 14323 31591 14417 31625
rect 14323 31557 14353 31591
rect 14387 31557 14417 31591
rect 14323 31523 14417 31557
rect 14323 31489 14353 31523
rect 14387 31489 14417 31523
rect 14323 31455 14417 31489
rect 14323 31421 14353 31455
rect 14387 31421 14417 31455
rect 14323 31387 14417 31421
rect 14323 31353 14353 31387
rect 14387 31353 14417 31387
rect 14323 31319 14417 31353
rect 14323 31285 14353 31319
rect 14387 31285 14417 31319
rect 14323 31251 14417 31285
rect 14323 31217 14353 31251
rect 14387 31217 14417 31251
rect 14323 31183 14417 31217
rect 14323 31149 14353 31183
rect 14387 31149 14417 31183
rect 14323 31115 14417 31149
rect 14323 31081 14353 31115
rect 14387 31081 14417 31115
rect 14323 31047 14417 31081
rect 14323 31013 14353 31047
rect 14387 31013 14417 31047
rect 14323 30979 14417 31013
rect 14323 30945 14353 30979
rect 14387 30945 14417 30979
rect 14323 30911 14417 30945
rect 14323 30877 14353 30911
rect 14387 30877 14417 30911
rect 14323 30843 14417 30877
rect 14323 30809 14353 30843
rect 14387 30809 14417 30843
rect 14323 30775 14417 30809
rect 14323 30741 14353 30775
rect 14387 30741 14417 30775
rect 14323 30707 14417 30741
rect 14323 30673 14353 30707
rect 14387 30673 14417 30707
rect 14323 30639 14417 30673
rect 14323 30605 14353 30639
rect 14387 30605 14417 30639
rect 14323 30571 14417 30605
rect 14323 30537 14353 30571
rect 14387 30537 14417 30571
rect 14323 30503 14417 30537
rect 14323 30469 14353 30503
rect 14387 30469 14417 30503
rect 14323 30435 14417 30469
rect 14323 30401 14353 30435
rect 14387 30401 14417 30435
rect 14323 30367 14417 30401
rect 14323 30333 14353 30367
rect 14387 30333 14417 30367
rect 14323 30299 14417 30333
rect 14323 30265 14353 30299
rect 14387 30265 14417 30299
rect 14323 30231 14417 30265
rect 14323 30197 14353 30231
rect 14387 30197 14417 30231
rect 14323 30163 14417 30197
rect 14323 30129 14353 30163
rect 14387 30129 14417 30163
rect 14323 30095 14417 30129
rect 14323 30061 14353 30095
rect 14387 30061 14417 30095
rect 14323 30027 14417 30061
rect 14323 29993 14353 30027
rect 14387 29993 14417 30027
rect 14323 29959 14417 29993
rect 14323 29925 14353 29959
rect 14387 29925 14417 29959
rect 14323 29891 14417 29925
rect 14323 29857 14353 29891
rect 14387 29857 14417 29891
rect 14323 29823 14417 29857
rect 14323 29789 14353 29823
rect 14387 29789 14417 29823
rect 14323 29755 14417 29789
rect 14323 29721 14353 29755
rect 14387 29721 14417 29755
rect 14323 29687 14417 29721
rect 14323 29653 14353 29687
rect 14387 29653 14417 29687
rect 14323 29619 14417 29653
rect 14323 29585 14353 29619
rect 14387 29585 14417 29619
rect 14323 29551 14417 29585
rect 14323 29517 14353 29551
rect 14387 29517 14417 29551
rect 14323 29483 14417 29517
rect 14323 29449 14353 29483
rect 14387 29449 14417 29483
rect 14323 29415 14417 29449
rect 14323 29381 14353 29415
rect 14387 29381 14417 29415
rect 14323 29347 14417 29381
rect 14323 29313 14353 29347
rect 14387 29313 14417 29347
rect 14323 29279 14417 29313
rect 14323 29245 14353 29279
rect 14387 29245 14417 29279
rect 14323 29211 14417 29245
rect 14323 29177 14353 29211
rect 14387 29177 14417 29211
rect 14323 29143 14417 29177
rect 14323 29109 14353 29143
rect 14387 29109 14417 29143
rect 14323 29075 14417 29109
rect 14323 29041 14353 29075
rect 14387 29041 14417 29075
rect 14323 29007 14417 29041
rect 14323 28973 14353 29007
rect 14387 28973 14417 29007
rect 14323 28939 14417 28973
rect 14323 28905 14353 28939
rect 14387 28905 14417 28939
rect 14323 28871 14417 28905
rect 14323 28837 14353 28871
rect 14387 28837 14417 28871
rect 14323 28803 14417 28837
rect 14323 28769 14353 28803
rect 14387 28769 14417 28803
rect 14323 28735 14417 28769
rect 14323 28701 14353 28735
rect 14387 28701 14417 28735
rect 14323 28667 14417 28701
rect 14323 28633 14353 28667
rect 14387 28633 14417 28667
rect 14323 28599 14417 28633
rect 14323 28565 14353 28599
rect 14387 28565 14417 28599
rect 14323 28531 14417 28565
rect 14323 28497 14353 28531
rect 14387 28497 14417 28531
rect 14323 28463 14417 28497
rect 14323 28429 14353 28463
rect 14387 28429 14417 28463
rect 14323 28395 14417 28429
rect 14323 28361 14353 28395
rect 14387 28361 14417 28395
rect 14323 28327 14417 28361
rect 14323 28293 14353 28327
rect 14387 28293 14417 28327
rect 14323 28259 14417 28293
rect 14323 28225 14353 28259
rect 14387 28225 14417 28259
rect 14323 28191 14417 28225
rect 14323 28157 14353 28191
rect 14387 28157 14417 28191
rect 14323 28123 14417 28157
rect 14323 28089 14353 28123
rect 14387 28089 14417 28123
rect 14323 28055 14417 28089
rect 14323 28021 14353 28055
rect 14387 28021 14417 28055
rect 14323 27987 14417 28021
rect 14323 27953 14353 27987
rect 14387 27953 14417 27987
rect 14323 27919 14417 27953
rect 14323 27885 14353 27919
rect 14387 27885 14417 27919
rect 14323 27851 14417 27885
rect 14323 27817 14353 27851
rect 14387 27817 14417 27851
rect 14323 27783 14417 27817
rect 14323 27749 14353 27783
rect 14387 27749 14417 27783
rect 14323 27715 14417 27749
rect 14323 27681 14353 27715
rect 14387 27681 14417 27715
rect 14323 27647 14417 27681
rect 14323 27613 14353 27647
rect 14387 27613 14417 27647
rect 14323 27579 14417 27613
rect 14323 27545 14353 27579
rect 14387 27545 14417 27579
rect 14323 27511 14417 27545
rect 14323 27477 14353 27511
rect 14387 27477 14417 27511
rect 14323 27443 14417 27477
rect 14323 27409 14353 27443
rect 14387 27409 14417 27443
rect 14323 27375 14417 27409
rect 14323 27341 14353 27375
rect 14387 27341 14417 27375
rect 14323 27307 14417 27341
rect 14323 27273 14353 27307
rect 14387 27273 14417 27307
rect 14323 27239 14417 27273
rect 14323 27205 14353 27239
rect 14387 27205 14417 27239
rect 14323 27171 14417 27205
rect 14323 27137 14353 27171
rect 14387 27137 14417 27171
rect 14323 27103 14417 27137
rect 14323 27069 14353 27103
rect 14387 27069 14417 27103
rect 14323 27035 14417 27069
rect 14323 27001 14353 27035
rect 14387 27001 14417 27035
rect 14323 26967 14417 27001
rect 14323 26933 14353 26967
rect 14387 26933 14417 26967
rect 14323 26899 14417 26933
rect 14323 26865 14353 26899
rect 14387 26865 14417 26899
rect 14323 26831 14417 26865
rect 14323 26797 14353 26831
rect 14387 26797 14417 26831
rect 14323 26763 14417 26797
rect 14323 26729 14353 26763
rect 14387 26729 14417 26763
rect 14323 26695 14417 26729
rect 14323 26661 14353 26695
rect 14387 26661 14417 26695
rect 14323 26627 14417 26661
rect 14323 26593 14353 26627
rect 14387 26593 14417 26627
rect 14323 26559 14417 26593
rect 14323 26525 14353 26559
rect 14387 26525 14417 26559
rect 14323 26491 14417 26525
rect 14323 26457 14353 26491
rect 14387 26457 14417 26491
rect 14323 26423 14417 26457
rect 14323 26389 14353 26423
rect 14387 26389 14417 26423
rect 14323 26355 14417 26389
rect 14323 26321 14353 26355
rect 14387 26321 14417 26355
rect 14323 26287 14417 26321
rect 14323 26253 14353 26287
rect 14387 26253 14417 26287
rect 14323 26219 14417 26253
rect 14323 26185 14353 26219
rect 14387 26185 14417 26219
rect 14323 26151 14417 26185
rect 14323 26117 14353 26151
rect 14387 26117 14417 26151
rect 14323 26083 14417 26117
rect 14323 26049 14353 26083
rect 14387 26049 14417 26083
rect 14323 26015 14417 26049
rect 14323 25981 14353 26015
rect 14387 25981 14417 26015
rect 14323 25947 14417 25981
rect 14323 25913 14353 25947
rect 14387 25913 14417 25947
rect 14323 25879 14417 25913
rect 14323 25845 14353 25879
rect 14387 25845 14417 25879
rect 14323 25811 14417 25845
rect 14323 25777 14353 25811
rect 14387 25777 14417 25811
rect 14323 25743 14417 25777
rect 14323 25709 14353 25743
rect 14387 25709 14417 25743
rect 14323 25675 14417 25709
rect 14323 25641 14353 25675
rect 14387 25641 14417 25675
rect 14323 25607 14417 25641
rect 14323 25573 14353 25607
rect 14387 25573 14417 25607
rect 14323 25539 14417 25573
rect 14323 25505 14353 25539
rect 14387 25505 14417 25539
rect 14323 25471 14417 25505
rect 14323 25437 14353 25471
rect 14387 25437 14417 25471
rect 14323 25403 14417 25437
rect 14323 25369 14353 25403
rect 14387 25369 14417 25403
rect 14323 25335 14417 25369
rect 14323 25301 14353 25335
rect 14387 25301 14417 25335
rect 14323 25267 14417 25301
rect 14323 25233 14353 25267
rect 14387 25233 14417 25267
rect 14323 25199 14417 25233
rect 14323 25165 14353 25199
rect 14387 25165 14417 25199
rect 14323 25131 14417 25165
rect 14323 25097 14353 25131
rect 14387 25097 14417 25131
rect 14323 25063 14417 25097
rect 14323 25029 14353 25063
rect 14387 25029 14417 25063
rect 14323 24995 14417 25029
rect 14323 24961 14353 24995
rect 14387 24961 14417 24995
rect 14323 24927 14417 24961
rect 14323 24893 14353 24927
rect 14387 24893 14417 24927
rect 14323 24859 14417 24893
rect 14323 24825 14353 24859
rect 14387 24825 14417 24859
rect 14323 24791 14417 24825
rect 14323 24757 14353 24791
rect 14387 24757 14417 24791
rect 14323 24723 14417 24757
rect 14323 24689 14353 24723
rect 14387 24689 14417 24723
rect 14323 24655 14417 24689
rect 14323 24621 14353 24655
rect 14387 24621 14417 24655
rect 14323 24587 14417 24621
rect 14323 24553 14353 24587
rect 14387 24553 14417 24587
rect 14323 24519 14417 24553
rect 14323 24485 14353 24519
rect 14387 24485 14417 24519
rect 14323 24451 14417 24485
rect 14323 24417 14353 24451
rect 14387 24417 14417 24451
rect 14323 24383 14417 24417
rect 14323 24349 14353 24383
rect 14387 24349 14417 24383
rect 14323 24315 14417 24349
rect 14323 24281 14353 24315
rect 14387 24281 14417 24315
rect 14323 24247 14417 24281
rect 14323 24213 14353 24247
rect 14387 24213 14417 24247
rect 14323 24179 14417 24213
rect 14323 24145 14353 24179
rect 14387 24145 14417 24179
rect 14323 24111 14417 24145
rect 14323 24077 14353 24111
rect 14387 24077 14417 24111
rect 14323 24043 14417 24077
rect 14323 24009 14353 24043
rect 14387 24009 14417 24043
rect 14323 23975 14417 24009
rect 14323 23941 14353 23975
rect 14387 23941 14417 23975
rect 14323 23907 14417 23941
rect 14323 23873 14353 23907
rect 14387 23873 14417 23907
rect 14323 23839 14417 23873
rect 14323 23805 14353 23839
rect 14387 23805 14417 23839
rect 14323 23771 14417 23805
rect 14323 23737 14353 23771
rect 14387 23737 14417 23771
rect 14323 23703 14417 23737
rect 14323 23669 14353 23703
rect 14387 23669 14417 23703
rect 14323 23635 14417 23669
rect 14323 23601 14353 23635
rect 14387 23601 14417 23635
rect 14323 23567 14417 23601
rect 14323 23533 14353 23567
rect 14387 23533 14417 23567
rect 14323 23499 14417 23533
rect 14323 23465 14353 23499
rect 14387 23465 14417 23499
rect 14323 23431 14417 23465
rect 14323 23397 14353 23431
rect 14387 23397 14417 23431
rect 14323 23363 14417 23397
rect 14323 23329 14353 23363
rect 14387 23329 14417 23363
rect 14323 23295 14417 23329
rect 14323 23261 14353 23295
rect 14387 23261 14417 23295
rect 14323 23227 14417 23261
rect 14323 23193 14353 23227
rect 14387 23193 14417 23227
rect 14323 23159 14417 23193
rect 14323 23125 14353 23159
rect 14387 23125 14417 23159
rect 14323 23091 14417 23125
rect 14323 23057 14353 23091
rect 14387 23057 14417 23091
rect 14323 23023 14417 23057
rect 14323 22989 14353 23023
rect 14387 22989 14417 23023
rect 14323 22955 14417 22989
rect 14323 22921 14353 22955
rect 14387 22921 14417 22955
rect 14323 22887 14417 22921
rect 14323 22853 14353 22887
rect 14387 22853 14417 22887
rect 14323 22819 14417 22853
rect 14323 22785 14353 22819
rect 14387 22785 14417 22819
rect 14323 22751 14417 22785
rect 14323 22717 14353 22751
rect 14387 22717 14417 22751
rect 14323 22683 14417 22717
rect 14323 22649 14353 22683
rect 14387 22649 14417 22683
rect 14323 22615 14417 22649
rect 14323 22581 14353 22615
rect 14387 22581 14417 22615
rect 14323 22547 14417 22581
rect 14323 22513 14353 22547
rect 14387 22513 14417 22547
rect 14323 22479 14417 22513
rect 14323 22445 14353 22479
rect 14387 22445 14417 22479
rect 14323 22411 14417 22445
rect 14323 22377 14353 22411
rect 14387 22377 14417 22411
rect 14323 22343 14417 22377
rect 14323 22309 14353 22343
rect 14387 22309 14417 22343
rect 14323 22275 14417 22309
rect 14323 22241 14353 22275
rect 14387 22241 14417 22275
rect 14323 22207 14417 22241
rect 14323 22173 14353 22207
rect 14387 22173 14417 22207
rect 14323 22139 14417 22173
rect 14323 22105 14353 22139
rect 14387 22105 14417 22139
rect 14323 22071 14417 22105
rect 14323 22037 14353 22071
rect 14387 22037 14417 22071
rect 14323 22003 14417 22037
rect 14323 21969 14353 22003
rect 14387 21969 14417 22003
rect 14323 21935 14417 21969
rect 14323 21901 14353 21935
rect 14387 21901 14417 21935
rect 14323 21867 14417 21901
rect 14323 21833 14353 21867
rect 14387 21833 14417 21867
rect 14323 21799 14417 21833
rect 14323 21765 14353 21799
rect 14387 21765 14417 21799
rect 14323 21731 14417 21765
rect 14323 21697 14353 21731
rect 14387 21697 14417 21731
rect 14323 21663 14417 21697
rect 14323 21629 14353 21663
rect 14387 21629 14417 21663
rect 14323 21595 14417 21629
rect 14323 21561 14353 21595
rect 14387 21561 14417 21595
rect 14323 21527 14417 21561
rect 14323 21493 14353 21527
rect 14387 21493 14417 21527
rect 14323 21459 14417 21493
rect 14323 21425 14353 21459
rect 14387 21425 14417 21459
rect 14323 21391 14417 21425
rect 14323 21357 14353 21391
rect 14387 21357 14417 21391
rect 14323 21323 14417 21357
rect 14323 21289 14353 21323
rect 14387 21289 14417 21323
rect 14323 21255 14417 21289
rect 14323 21221 14353 21255
rect 14387 21221 14417 21255
rect 14323 21187 14417 21221
rect 14323 21153 14353 21187
rect 14387 21153 14417 21187
rect 14323 21119 14417 21153
rect 14323 21085 14353 21119
rect 14387 21085 14417 21119
rect 14323 21051 14417 21085
rect 14323 21017 14353 21051
rect 14387 21017 14417 21051
rect 14323 20983 14417 21017
rect 14323 20949 14353 20983
rect 14387 20949 14417 20983
rect 14323 20915 14417 20949
rect 14323 20881 14353 20915
rect 14387 20881 14417 20915
rect 14323 20847 14417 20881
rect 14323 20813 14353 20847
rect 14387 20813 14417 20847
rect 14323 20779 14417 20813
rect 14323 20745 14353 20779
rect 14387 20745 14417 20779
rect 14323 20711 14417 20745
rect 14323 20677 14353 20711
rect 14387 20677 14417 20711
rect 14323 20643 14417 20677
rect 14323 20609 14353 20643
rect 14387 20609 14417 20643
rect 14323 20575 14417 20609
rect 14323 20541 14353 20575
rect 14387 20541 14417 20575
rect 14323 20507 14417 20541
rect 14323 20473 14353 20507
rect 14387 20473 14417 20507
rect 14323 20439 14417 20473
rect 14323 20405 14353 20439
rect 14387 20405 14417 20439
rect 14323 20371 14417 20405
rect 14323 20337 14353 20371
rect 14387 20337 14417 20371
rect 14323 20303 14417 20337
rect 14323 20269 14353 20303
rect 14387 20269 14417 20303
rect 14323 20235 14417 20269
rect 14323 20201 14353 20235
rect 14387 20201 14417 20235
rect 14323 20167 14417 20201
rect 14323 20133 14353 20167
rect 14387 20133 14417 20167
rect 14323 20099 14417 20133
rect 14323 20065 14353 20099
rect 14387 20065 14417 20099
rect 14323 20031 14417 20065
rect 14323 19997 14353 20031
rect 14387 19997 14417 20031
rect 14323 19963 14417 19997
rect 14323 19929 14353 19963
rect 14387 19929 14417 19963
rect 14323 19895 14417 19929
rect 14323 19861 14353 19895
rect 14387 19861 14417 19895
rect 14323 19827 14417 19861
rect 14323 19793 14353 19827
rect 14387 19793 14417 19827
rect 14323 19759 14417 19793
rect 14323 19725 14353 19759
rect 14387 19725 14417 19759
rect 14323 19691 14417 19725
rect 14323 19657 14353 19691
rect 14387 19657 14417 19691
rect 14323 19623 14417 19657
rect 14323 19589 14353 19623
rect 14387 19589 14417 19623
rect 14323 19555 14417 19589
rect 14323 19521 14353 19555
rect 14387 19521 14417 19555
rect 14323 19487 14417 19521
rect 14323 19453 14353 19487
rect 14387 19453 14417 19487
rect 14323 19419 14417 19453
rect 14323 19385 14353 19419
rect 14387 19385 14417 19419
rect 14323 19351 14417 19385
rect 14323 19317 14353 19351
rect 14387 19317 14417 19351
rect 14323 19283 14417 19317
rect 14323 19249 14353 19283
rect 14387 19249 14417 19283
rect 14323 19215 14417 19249
rect 14323 19181 14353 19215
rect 14387 19181 14417 19215
rect 14323 19147 14417 19181
rect 14323 19113 14353 19147
rect 14387 19113 14417 19147
rect 14323 19079 14417 19113
rect 14323 19045 14353 19079
rect 14387 19045 14417 19079
rect 14323 19011 14417 19045
rect 14323 18977 14353 19011
rect 14387 18977 14417 19011
rect 14323 18943 14417 18977
rect 14323 18909 14353 18943
rect 14387 18909 14417 18943
rect 14323 18875 14417 18909
rect 14323 18841 14353 18875
rect 14387 18841 14417 18875
rect 14323 18807 14417 18841
rect 14323 18773 14353 18807
rect 14387 18773 14417 18807
rect 14323 18739 14417 18773
rect 14323 18705 14353 18739
rect 14387 18705 14417 18739
rect 14323 18671 14417 18705
rect 14323 18637 14353 18671
rect 14387 18637 14417 18671
rect 14323 18603 14417 18637
rect 14323 18569 14353 18603
rect 14387 18569 14417 18603
rect 14323 18535 14417 18569
rect 14323 18501 14353 18535
rect 14387 18501 14417 18535
rect 14323 18467 14417 18501
rect 14323 18433 14353 18467
rect 14387 18433 14417 18467
rect 14323 18399 14417 18433
rect 14323 18365 14353 18399
rect 14387 18365 14417 18399
rect 14323 18331 14417 18365
rect 14323 18297 14353 18331
rect 14387 18297 14417 18331
rect 14323 18263 14417 18297
rect 14323 18229 14353 18263
rect 14387 18229 14417 18263
rect 14323 18195 14417 18229
rect 14323 18161 14353 18195
rect 14387 18161 14417 18195
rect 14323 18127 14417 18161
rect 14323 18093 14353 18127
rect 14387 18093 14417 18127
rect 14323 18059 14417 18093
rect 14323 18025 14353 18059
rect 14387 18025 14417 18059
rect 14323 17991 14417 18025
rect 14323 17957 14353 17991
rect 14387 17957 14417 17991
rect 14323 17923 14417 17957
rect 14323 17889 14353 17923
rect 14387 17889 14417 17923
rect 14323 17855 14417 17889
rect 14323 17821 14353 17855
rect 14387 17821 14417 17855
rect 14323 17787 14417 17821
rect 14323 17753 14353 17787
rect 14387 17753 14417 17787
rect 14323 17719 14417 17753
rect 14323 17685 14353 17719
rect 14387 17685 14417 17719
rect 14323 17651 14417 17685
rect 14323 17617 14353 17651
rect 14387 17617 14417 17651
rect 14323 17583 14417 17617
rect 14323 17549 14353 17583
rect 14387 17549 14417 17583
rect 14323 17515 14417 17549
rect 14323 17481 14353 17515
rect 14387 17481 14417 17515
rect 14323 17447 14417 17481
rect 14323 17413 14353 17447
rect 14387 17413 14417 17447
rect 14323 17379 14417 17413
rect 14323 17345 14353 17379
rect 14387 17345 14417 17379
rect 14323 17311 14417 17345
rect 14323 17277 14353 17311
rect 14387 17277 14417 17311
rect 14323 17243 14417 17277
rect 14323 17209 14353 17243
rect 14387 17209 14417 17243
rect 14323 17175 14417 17209
rect 14323 17141 14353 17175
rect 14387 17141 14417 17175
rect 14323 17107 14417 17141
rect 14323 17073 14353 17107
rect 14387 17073 14417 17107
rect 14323 17039 14417 17073
rect 14323 17005 14353 17039
rect 14387 17005 14417 17039
rect 14323 16971 14417 17005
rect 14323 16937 14353 16971
rect 14387 16937 14417 16971
rect 14323 16903 14417 16937
rect 14323 16869 14353 16903
rect 14387 16869 14417 16903
rect 14323 16835 14417 16869
rect 14323 16801 14353 16835
rect 14387 16801 14417 16835
rect 14323 16767 14417 16801
rect 14323 16733 14353 16767
rect 14387 16733 14417 16767
rect 14323 16699 14417 16733
rect 14323 16665 14353 16699
rect 14387 16665 14417 16699
rect 14323 16631 14417 16665
rect 14323 16597 14353 16631
rect 14387 16597 14417 16631
rect 14323 16563 14417 16597
rect 14323 16529 14353 16563
rect 14387 16529 14417 16563
rect 14323 16495 14417 16529
rect 14323 16461 14353 16495
rect 14387 16461 14417 16495
rect 14323 16427 14417 16461
rect 14323 16393 14353 16427
rect 14387 16393 14417 16427
rect 14323 16359 14417 16393
rect 14323 16325 14353 16359
rect 14387 16325 14417 16359
rect 14323 16291 14417 16325
rect 14323 16257 14353 16291
rect 14387 16257 14417 16291
rect 14323 16223 14417 16257
rect 14323 16189 14353 16223
rect 14387 16189 14417 16223
rect 14323 16155 14417 16189
rect 14323 16121 14353 16155
rect 14387 16121 14417 16155
rect 14323 16087 14417 16121
rect 14323 16053 14353 16087
rect 14387 16053 14417 16087
rect 14323 16019 14417 16053
rect 14323 15985 14353 16019
rect 14387 15985 14417 16019
rect 14323 15951 14417 15985
rect 14323 15917 14353 15951
rect 14387 15917 14417 15951
rect 14323 15883 14417 15917
rect 14323 15849 14353 15883
rect 14387 15849 14417 15883
rect 14323 15815 14417 15849
rect 14323 15781 14353 15815
rect 14387 15781 14417 15815
rect 14323 15747 14417 15781
rect 14323 15713 14353 15747
rect 14387 15713 14417 15747
rect 14323 15679 14417 15713
rect 14323 15645 14353 15679
rect 14387 15645 14417 15679
rect 14323 15611 14417 15645
rect 14323 15577 14353 15611
rect 14387 15577 14417 15611
rect 14323 15543 14417 15577
rect 14323 15509 14353 15543
rect 14387 15509 14417 15543
rect 14323 15475 14417 15509
rect 14323 15441 14353 15475
rect 14387 15441 14417 15475
rect 14323 15407 14417 15441
rect 14323 15373 14353 15407
rect 14387 15373 14417 15407
rect 14323 15339 14417 15373
rect 14323 15305 14353 15339
rect 14387 15305 14417 15339
rect 14323 15271 14417 15305
rect 14323 15237 14353 15271
rect 14387 15237 14417 15271
rect 14323 15203 14417 15237
rect 14323 15169 14353 15203
rect 14387 15169 14417 15203
rect 14323 15135 14417 15169
rect 14323 15101 14353 15135
rect 14387 15101 14417 15135
rect 14323 15067 14417 15101
rect 14323 15033 14353 15067
rect 14387 15033 14417 15067
rect 14323 14999 14417 15033
rect 14323 14965 14353 14999
rect 14387 14965 14417 14999
rect 14323 14931 14417 14965
rect 14323 14897 14353 14931
rect 14387 14897 14417 14931
rect 14323 14863 14417 14897
rect 14323 14829 14353 14863
rect 14387 14829 14417 14863
rect 14323 14795 14417 14829
rect 14323 14761 14353 14795
rect 14387 14761 14417 14795
rect 14323 14727 14417 14761
rect 14323 14693 14353 14727
rect 14387 14693 14417 14727
rect 14323 14659 14417 14693
rect 14323 14625 14353 14659
rect 14387 14625 14417 14659
rect 14323 14591 14417 14625
rect 14323 14557 14353 14591
rect 14387 14557 14417 14591
rect 14323 14523 14417 14557
rect 14323 14489 14353 14523
rect 14387 14489 14417 14523
rect 14323 14455 14417 14489
rect 14323 14421 14353 14455
rect 14387 14421 14417 14455
rect 14323 14387 14417 14421
rect 14323 14353 14353 14387
rect 14387 14353 14417 14387
rect 14323 14319 14417 14353
rect 14323 14285 14353 14319
rect 14387 14285 14417 14319
rect 14323 14251 14417 14285
rect 14323 14217 14353 14251
rect 14387 14217 14417 14251
rect 14323 14183 14417 14217
rect 14323 14149 14353 14183
rect 14387 14149 14417 14183
rect 14323 14115 14417 14149
rect 14323 14081 14353 14115
rect 14387 14081 14417 14115
rect 14323 14047 14417 14081
rect 14323 14013 14353 14047
rect 14387 14013 14417 14047
rect 14323 13979 14417 14013
rect 14323 13945 14353 13979
rect 14387 13945 14417 13979
rect 14323 13911 14417 13945
rect 14323 13877 14353 13911
rect 14387 13877 14417 13911
rect 14323 13843 14417 13877
rect 14323 13809 14353 13843
rect 14387 13809 14417 13843
rect 14323 13775 14417 13809
rect 14323 13741 14353 13775
rect 14387 13741 14417 13775
rect 14323 13707 14417 13741
rect 14323 13673 14353 13707
rect 14387 13673 14417 13707
rect 14323 13639 14417 13673
rect 14323 13605 14353 13639
rect 14387 13605 14417 13639
rect 14323 13571 14417 13605
rect 14323 13537 14353 13571
rect 14387 13537 14417 13571
rect 14323 13503 14417 13537
rect 14323 13469 14353 13503
rect 14387 13469 14417 13503
rect 14323 13435 14417 13469
rect 14323 13401 14353 13435
rect 14387 13401 14417 13435
rect 14323 13367 14417 13401
rect 14323 13333 14353 13367
rect 14387 13333 14417 13367
rect 14323 13299 14417 13333
rect 14323 13265 14353 13299
rect 14387 13265 14417 13299
rect 14323 13231 14417 13265
rect 14323 13197 14353 13231
rect 14387 13197 14417 13231
rect 14323 13163 14417 13197
rect 14323 13129 14353 13163
rect 14387 13129 14417 13163
rect 14323 13095 14417 13129
rect 14323 13061 14353 13095
rect 14387 13061 14417 13095
rect 14323 13027 14417 13061
rect 14323 12993 14353 13027
rect 14387 12993 14417 13027
rect 14323 12959 14417 12993
rect 14323 12925 14353 12959
rect 14387 12925 14417 12959
rect 14323 12891 14417 12925
rect 14323 12857 14353 12891
rect 14387 12857 14417 12891
rect 14323 12823 14417 12857
rect 14323 12789 14353 12823
rect 14387 12789 14417 12823
rect 14323 12755 14417 12789
rect 14323 12721 14353 12755
rect 14387 12721 14417 12755
rect 14323 12687 14417 12721
rect 14323 12653 14353 12687
rect 14387 12653 14417 12687
rect 14323 12619 14417 12653
rect 14323 12585 14353 12619
rect 14387 12585 14417 12619
rect 14323 12551 14417 12585
rect 14323 12517 14353 12551
rect 14387 12517 14417 12551
rect 14323 12483 14417 12517
rect 14323 12449 14353 12483
rect 14387 12449 14417 12483
rect 14323 12415 14417 12449
rect 14323 12381 14353 12415
rect 14387 12381 14417 12415
rect 14323 12347 14417 12381
rect 14323 12313 14353 12347
rect 14387 12313 14417 12347
rect 14323 12279 14417 12313
rect 14323 12245 14353 12279
rect 14387 12245 14417 12279
rect 14323 12211 14417 12245
rect 14323 12177 14353 12211
rect 14387 12177 14417 12211
rect 14323 12143 14417 12177
rect 14323 12109 14353 12143
rect 14387 12109 14417 12143
rect 14323 12075 14417 12109
rect 14323 12041 14353 12075
rect 14387 12041 14417 12075
rect 14323 12007 14417 12041
rect 14323 11973 14353 12007
rect 14387 11973 14417 12007
rect 14323 11939 14417 11973
rect 14323 11905 14353 11939
rect 14387 11905 14417 11939
rect 14323 11871 14417 11905
rect 14323 11837 14353 11871
rect 14387 11837 14417 11871
rect 14323 11803 14417 11837
rect 14323 11769 14353 11803
rect 14387 11769 14417 11803
rect 14323 11735 14417 11769
rect 14323 11701 14353 11735
rect 14387 11701 14417 11735
rect 14323 11667 14417 11701
rect 14323 11633 14353 11667
rect 14387 11633 14417 11667
rect 14323 11599 14417 11633
rect 14323 11565 14353 11599
rect 14387 11565 14417 11599
rect 14323 11531 14417 11565
rect 14323 11497 14353 11531
rect 14387 11497 14417 11531
rect 14323 11463 14417 11497
rect 14323 11429 14353 11463
rect 14387 11429 14417 11463
rect 14323 11395 14417 11429
rect 14323 11361 14353 11395
rect 14387 11361 14417 11395
rect 14323 11327 14417 11361
rect 14323 11293 14353 11327
rect 14387 11293 14417 11327
rect 14323 11259 14417 11293
rect 14323 11225 14353 11259
rect 14387 11225 14417 11259
rect 14323 11191 14417 11225
rect 14323 11157 14353 11191
rect 14387 11157 14417 11191
rect 14323 11123 14417 11157
rect 14323 11089 14353 11123
rect 14387 11089 14417 11123
rect 14323 11055 14417 11089
rect 14323 11021 14353 11055
rect 14387 11021 14417 11055
rect 14323 10987 14417 11021
rect 14323 10953 14353 10987
rect 14387 10953 14417 10987
rect 14323 10919 14417 10953
rect 14323 10885 14353 10919
rect 14387 10885 14417 10919
rect 14323 10851 14417 10885
rect 14323 10817 14353 10851
rect 14387 10817 14417 10851
rect 14323 10783 14417 10817
rect 14323 10749 14353 10783
rect 14387 10749 14417 10783
rect 14323 10715 14417 10749
rect 14323 10681 14353 10715
rect 14387 10681 14417 10715
rect 14323 10647 14417 10681
rect 14323 10613 14353 10647
rect 14387 10613 14417 10647
rect 14323 10579 14417 10613
rect 14323 10545 14353 10579
rect 14387 10545 14417 10579
rect 14323 10511 14417 10545
rect 14323 10477 14353 10511
rect 14387 10477 14417 10511
rect 14323 10443 14417 10477
rect 14323 10409 14353 10443
rect 14387 10409 14417 10443
rect 14323 10375 14417 10409
rect 14323 10341 14353 10375
rect 14387 10341 14417 10375
rect 14323 10307 14417 10341
rect 14323 10273 14353 10307
rect 14387 10273 14417 10307
rect 14323 10239 14417 10273
rect 14323 10205 14353 10239
rect 14387 10205 14417 10239
rect 14323 10171 14417 10205
rect 14323 10137 14353 10171
rect 14387 10137 14417 10171
rect 14323 10103 14417 10137
rect 14323 10069 14353 10103
rect 14387 10069 14417 10103
rect 14323 10035 14417 10069
rect 14323 10001 14353 10035
rect 14387 10001 14417 10035
rect 14323 9967 14417 10001
rect 14323 9933 14353 9967
rect 14387 9933 14417 9967
rect 14323 9899 14417 9933
rect 14323 9865 14353 9899
rect 14387 9865 14417 9899
rect 14323 9831 14417 9865
rect 14323 9797 14353 9831
rect 14387 9797 14417 9831
rect 14323 9749 14417 9797
rect 589 9719 14417 9749
rect 589 9685 719 9719
rect 753 9685 787 9719
rect 821 9685 855 9719
rect 889 9718 923 9719
rect 957 9718 991 9719
rect 917 9685 923 9718
rect 989 9685 991 9718
rect 1025 9718 1059 9719
rect 1093 9718 1127 9719
rect 1161 9718 1195 9719
rect 1229 9718 1263 9719
rect 1297 9718 1331 9719
rect 1365 9718 1399 9719
rect 1433 9718 1467 9719
rect 1501 9718 1535 9719
rect 1025 9685 1027 9718
rect 1093 9685 1099 9718
rect 1161 9685 1171 9718
rect 1229 9685 1243 9718
rect 1297 9685 1315 9718
rect 1365 9685 1387 9718
rect 1433 9685 1459 9718
rect 1501 9685 1531 9718
rect 1569 9685 1603 9719
rect 1637 9685 1671 9719
rect 1705 9718 1739 9719
rect 1773 9718 1807 9719
rect 1841 9718 1875 9719
rect 1909 9718 1943 9719
rect 1977 9718 2011 9719
rect 2045 9718 2079 9719
rect 1709 9685 1739 9718
rect 1781 9685 1807 9718
rect 1853 9685 1875 9718
rect 1925 9685 1943 9718
rect 1997 9685 2011 9718
rect 2069 9685 2079 9718
rect 2113 9685 2147 9719
rect 2181 9685 2215 9719
rect 2249 9685 2283 9719
rect 2317 9685 2351 9719
rect 2385 9685 2419 9719
rect 2453 9685 2487 9719
rect 2521 9685 2555 9719
rect 2589 9685 2623 9719
rect 2657 9685 2691 9719
rect 2725 9685 2759 9719
rect 2793 9685 2827 9719
rect 2861 9685 2895 9719
rect 2929 9685 2963 9719
rect 2997 9685 3031 9719
rect 3065 9685 3099 9719
rect 3133 9685 3167 9719
rect 3201 9685 3235 9719
rect 3269 9685 3303 9719
rect 3337 9685 3371 9719
rect 3405 9685 3439 9719
rect 3473 9685 3507 9719
rect 3541 9685 3575 9719
rect 3609 9685 3643 9719
rect 3677 9685 3711 9719
rect 3745 9685 3779 9719
rect 3813 9685 3847 9719
rect 3881 9685 3915 9719
rect 3949 9685 3983 9719
rect 4017 9685 4051 9719
rect 4085 9685 4119 9719
rect 4153 9685 4187 9719
rect 4221 9685 4255 9719
rect 4289 9685 4323 9719
rect 4357 9685 4391 9719
rect 4425 9685 4459 9719
rect 4493 9685 4527 9719
rect 4561 9685 4595 9719
rect 4629 9685 4663 9719
rect 4697 9685 4731 9719
rect 4765 9685 4799 9719
rect 4833 9685 4867 9719
rect 4901 9685 4935 9719
rect 4969 9685 5003 9719
rect 5037 9685 5071 9719
rect 5105 9685 5139 9719
rect 5173 9685 5207 9719
rect 5241 9685 5275 9719
rect 5309 9685 5343 9719
rect 5377 9685 5411 9719
rect 5445 9685 5479 9719
rect 5513 9685 5547 9719
rect 5581 9685 5615 9719
rect 5649 9685 5683 9719
rect 5717 9685 5751 9719
rect 5785 9685 5819 9719
rect 5853 9685 5887 9719
rect 5921 9685 5955 9719
rect 5989 9685 6023 9719
rect 6057 9685 6091 9719
rect 6125 9685 6159 9719
rect 6193 9685 6227 9719
rect 6261 9685 6295 9719
rect 6329 9685 6363 9719
rect 6397 9685 6431 9719
rect 6465 9685 6499 9719
rect 6533 9685 6567 9719
rect 6601 9685 6635 9719
rect 6669 9685 6703 9719
rect 6737 9685 6771 9719
rect 6805 9685 6839 9719
rect 6873 9685 6907 9719
rect 6941 9685 6975 9719
rect 7009 9685 7043 9719
rect 7077 9685 7111 9719
rect 7145 9685 7179 9719
rect 7213 9685 7247 9719
rect 7281 9685 7315 9719
rect 7349 9685 7383 9719
rect 7417 9685 7451 9719
rect 7485 9685 7519 9719
rect 7553 9685 7587 9719
rect 7621 9685 7655 9719
rect 7689 9685 7723 9719
rect 7757 9685 7791 9719
rect 7825 9685 7859 9719
rect 7893 9685 7927 9719
rect 7961 9685 7995 9719
rect 8029 9685 8063 9719
rect 8097 9685 8131 9719
rect 8165 9685 8199 9719
rect 8233 9685 8267 9719
rect 8301 9685 8335 9719
rect 8369 9685 8403 9719
rect 8437 9685 8471 9719
rect 8505 9685 8539 9719
rect 8573 9685 8607 9719
rect 8641 9685 8675 9719
rect 8709 9685 8743 9719
rect 8777 9685 8811 9719
rect 8845 9685 8879 9719
rect 8913 9685 8947 9719
rect 8981 9685 9015 9719
rect 9049 9685 9083 9719
rect 9117 9685 9151 9719
rect 9185 9685 9219 9719
rect 9253 9685 9287 9719
rect 9321 9685 9355 9719
rect 9389 9685 9423 9719
rect 9457 9685 9491 9719
rect 9525 9685 9559 9719
rect 9593 9685 9627 9719
rect 9661 9685 9695 9719
rect 9729 9685 9763 9719
rect 9797 9685 9831 9719
rect 9865 9685 9899 9719
rect 9933 9685 9967 9719
rect 10001 9685 10035 9719
rect 10069 9685 10103 9719
rect 10137 9685 10171 9719
rect 10205 9685 10239 9719
rect 10273 9685 10307 9719
rect 10341 9685 10375 9719
rect 10409 9685 10443 9719
rect 10477 9685 10511 9719
rect 10545 9685 10579 9719
rect 10613 9685 10647 9719
rect 10681 9685 10715 9719
rect 10749 9685 10783 9719
rect 10817 9685 10851 9719
rect 10885 9685 10919 9719
rect 10953 9685 10987 9719
rect 11021 9685 11055 9719
rect 11089 9685 11123 9719
rect 11157 9685 11191 9719
rect 11225 9685 11259 9719
rect 11293 9685 11327 9719
rect 11361 9685 11395 9719
rect 11429 9685 11463 9719
rect 11497 9685 11531 9719
rect 11565 9685 11599 9719
rect 11633 9685 11667 9719
rect 11701 9685 11735 9719
rect 11769 9685 11803 9719
rect 11837 9685 11871 9719
rect 11905 9685 11939 9719
rect 11973 9685 12007 9719
rect 12041 9685 12075 9719
rect 12109 9685 12143 9719
rect 12177 9685 12211 9719
rect 12245 9685 12279 9719
rect 12313 9685 12347 9719
rect 12381 9685 12415 9719
rect 12449 9685 12483 9719
rect 12517 9685 12551 9719
rect 12585 9685 12619 9719
rect 12653 9685 12687 9719
rect 12721 9685 12755 9719
rect 12789 9685 12823 9719
rect 12857 9718 12891 9719
rect 12925 9718 12959 9719
rect 12857 9685 12883 9718
rect 12925 9685 12955 9718
rect 12993 9685 13027 9719
rect 13061 9685 13095 9719
rect 13129 9718 13163 9719
rect 13197 9718 13231 9719
rect 13265 9718 13299 9719
rect 13333 9718 13367 9719
rect 13401 9718 13435 9719
rect 13469 9718 13503 9719
rect 13537 9718 13571 9719
rect 13605 9718 13639 9719
rect 13133 9685 13163 9718
rect 13205 9685 13231 9718
rect 13277 9685 13299 9718
rect 13349 9685 13367 9718
rect 13421 9685 13435 9718
rect 13493 9685 13503 9718
rect 13565 9685 13571 9718
rect 13637 9685 13639 9718
rect 13673 9718 13707 9719
rect 13741 9718 13775 9719
rect 13809 9718 13843 9719
rect 13877 9718 13911 9719
rect 13945 9718 13979 9719
rect 14013 9718 14047 9719
rect 13673 9685 13675 9718
rect 13741 9685 13747 9718
rect 13809 9685 13819 9718
rect 13877 9685 13891 9718
rect 13945 9685 13963 9718
rect 14013 9685 14035 9718
rect 14081 9685 14115 9719
rect 14149 9685 14183 9719
rect 14217 9685 14251 9719
rect 14285 9685 14417 9719
rect 589 9684 883 9685
rect 917 9684 955 9685
rect 989 9684 1027 9685
rect 1061 9684 1099 9685
rect 1133 9684 1171 9685
rect 1205 9684 1243 9685
rect 1277 9684 1315 9685
rect 1349 9684 1387 9685
rect 1421 9684 1459 9685
rect 1493 9684 1531 9685
rect 1565 9684 1603 9685
rect 1637 9684 1675 9685
rect 1709 9684 1747 9685
rect 1781 9684 1819 9685
rect 1853 9684 1891 9685
rect 1925 9684 1963 9685
rect 1997 9684 2035 9685
rect 2069 9684 12883 9685
rect 12917 9684 12955 9685
rect 12989 9684 13027 9685
rect 13061 9684 13099 9685
rect 13133 9684 13171 9685
rect 13205 9684 13243 9685
rect 13277 9684 13315 9685
rect 13349 9684 13387 9685
rect 13421 9684 13459 9685
rect 13493 9684 13531 9685
rect 13565 9684 13603 9685
rect 13637 9684 13675 9685
rect 13709 9684 13747 9685
rect 13781 9684 13819 9685
rect 13853 9684 13891 9685
rect 13925 9684 13963 9685
rect 13997 9684 14035 9685
rect 14069 9684 14417 9685
rect 589 9655 14417 9684
rect 882 9654 2070 9655
rect 12882 9654 14070 9655
<< viali >>
rect 883 9685 889 9718
rect 889 9685 917 9718
rect 955 9685 957 9718
rect 957 9685 989 9718
rect 1027 9685 1059 9718
rect 1059 9685 1061 9718
rect 1099 9685 1127 9718
rect 1127 9685 1133 9718
rect 1171 9685 1195 9718
rect 1195 9685 1205 9718
rect 1243 9685 1263 9718
rect 1263 9685 1277 9718
rect 1315 9685 1331 9718
rect 1331 9685 1349 9718
rect 1387 9685 1399 9718
rect 1399 9685 1421 9718
rect 1459 9685 1467 9718
rect 1467 9685 1493 9718
rect 1531 9685 1535 9718
rect 1535 9685 1565 9718
rect 1603 9685 1637 9718
rect 1675 9685 1705 9718
rect 1705 9685 1709 9718
rect 1747 9685 1773 9718
rect 1773 9685 1781 9718
rect 1819 9685 1841 9718
rect 1841 9685 1853 9718
rect 1891 9685 1909 9718
rect 1909 9685 1925 9718
rect 1963 9685 1977 9718
rect 1977 9685 1997 9718
rect 2035 9685 2045 9718
rect 2045 9685 2069 9718
rect 12883 9685 12891 9718
rect 12891 9685 12917 9718
rect 12955 9685 12959 9718
rect 12959 9685 12989 9718
rect 13027 9685 13061 9718
rect 13099 9685 13129 9718
rect 13129 9685 13133 9718
rect 13171 9685 13197 9718
rect 13197 9685 13205 9718
rect 13243 9685 13265 9718
rect 13265 9685 13277 9718
rect 13315 9685 13333 9718
rect 13333 9685 13349 9718
rect 13387 9685 13401 9718
rect 13401 9685 13421 9718
rect 13459 9685 13469 9718
rect 13469 9685 13493 9718
rect 13531 9685 13537 9718
rect 13537 9685 13565 9718
rect 13603 9685 13605 9718
rect 13605 9685 13637 9718
rect 13675 9685 13707 9718
rect 13707 9685 13709 9718
rect 13747 9685 13775 9718
rect 13775 9685 13781 9718
rect 13819 9685 13843 9718
rect 13843 9685 13853 9718
rect 13891 9685 13911 9718
rect 13911 9685 13925 9718
rect 13963 9685 13979 9718
rect 13979 9685 13997 9718
rect 14035 9685 14047 9718
rect 14047 9685 14069 9718
rect 883 9684 917 9685
rect 955 9684 989 9685
rect 1027 9684 1061 9685
rect 1099 9684 1133 9685
rect 1171 9684 1205 9685
rect 1243 9684 1277 9685
rect 1315 9684 1349 9685
rect 1387 9684 1421 9685
rect 1459 9684 1493 9685
rect 1531 9684 1565 9685
rect 1603 9684 1637 9685
rect 1675 9684 1709 9685
rect 1747 9684 1781 9685
rect 1819 9684 1853 9685
rect 1891 9684 1925 9685
rect 1963 9684 1997 9685
rect 2035 9684 2069 9685
rect 12883 9684 12917 9685
rect 12955 9684 12989 9685
rect 13027 9684 13061 9685
rect 13099 9684 13133 9685
rect 13171 9684 13205 9685
rect 13243 9684 13277 9685
rect 13315 9684 13349 9685
rect 13387 9684 13421 9685
rect 13459 9684 13493 9685
rect 13531 9684 13565 9685
rect 13603 9684 13637 9685
rect 13675 9684 13709 9685
rect 13747 9684 13781 9685
rect 13819 9684 13853 9685
rect 13891 9684 13925 9685
rect 13963 9684 13997 9685
rect 14035 9684 14069 9685
<< metal1 >>
rect 858 9731 2096 9772
rect 858 9718 908 9731
rect 2048 9718 2096 9731
rect 858 9684 883 9718
rect 2069 9684 2096 9718
rect 858 9295 908 9684
rect 2048 9295 2096 9684
rect 858 9252 2096 9295
rect 12858 9731 14096 9772
rect 12858 9718 12908 9731
rect 14048 9718 14096 9731
rect 12858 9684 12883 9718
rect 14069 9684 14096 9718
rect 12858 9295 12908 9684
rect 14048 9295 14096 9684
rect 12858 9252 14096 9295
<< via1 >>
rect 908 9718 2048 9731
rect 908 9684 917 9718
rect 917 9684 955 9718
rect 955 9684 989 9718
rect 989 9684 1027 9718
rect 1027 9684 1061 9718
rect 1061 9684 1099 9718
rect 1099 9684 1133 9718
rect 1133 9684 1171 9718
rect 1171 9684 1205 9718
rect 1205 9684 1243 9718
rect 1243 9684 1277 9718
rect 1277 9684 1315 9718
rect 1315 9684 1349 9718
rect 1349 9684 1387 9718
rect 1387 9684 1421 9718
rect 1421 9684 1459 9718
rect 1459 9684 1493 9718
rect 1493 9684 1531 9718
rect 1531 9684 1565 9718
rect 1565 9684 1603 9718
rect 1603 9684 1637 9718
rect 1637 9684 1675 9718
rect 1675 9684 1709 9718
rect 1709 9684 1747 9718
rect 1747 9684 1781 9718
rect 1781 9684 1819 9718
rect 1819 9684 1853 9718
rect 1853 9684 1891 9718
rect 1891 9684 1925 9718
rect 1925 9684 1963 9718
rect 1963 9684 1997 9718
rect 1997 9684 2035 9718
rect 2035 9684 2048 9718
rect 908 9295 2048 9684
rect 12908 9718 14048 9731
rect 12908 9684 12917 9718
rect 12917 9684 12955 9718
rect 12955 9684 12989 9718
rect 12989 9684 13027 9718
rect 13027 9684 13061 9718
rect 13061 9684 13099 9718
rect 13099 9684 13133 9718
rect 13133 9684 13171 9718
rect 13171 9684 13205 9718
rect 13205 9684 13243 9718
rect 13243 9684 13277 9718
rect 13277 9684 13315 9718
rect 13315 9684 13349 9718
rect 13349 9684 13387 9718
rect 13387 9684 13421 9718
rect 13421 9684 13459 9718
rect 13459 9684 13493 9718
rect 13493 9684 13531 9718
rect 13531 9684 13565 9718
rect 13565 9684 13603 9718
rect 13603 9684 13637 9718
rect 13637 9684 13675 9718
rect 13675 9684 13709 9718
rect 13709 9684 13747 9718
rect 13747 9684 13781 9718
rect 13781 9684 13819 9718
rect 13819 9684 13853 9718
rect 13853 9684 13891 9718
rect 13891 9684 13925 9718
rect 13925 9684 13963 9718
rect 13963 9684 13997 9718
rect 13997 9684 14035 9718
rect 14035 9684 14048 9718
rect 12908 9295 14048 9684
<< metal2 >>
rect 858 9741 2096 9772
rect 858 9285 890 9741
rect 2066 9285 2096 9741
rect 858 9252 2096 9285
rect 12858 9741 14096 9772
rect 12858 9285 12890 9741
rect 14066 9285 14096 9741
rect 12858 9252 14096 9285
<< via2 >>
rect 890 9731 2066 9741
rect 890 9295 908 9731
rect 908 9295 2048 9731
rect 2048 9295 2066 9731
rect 890 9285 2066 9295
rect 12890 9731 14066 9741
rect 12890 9295 12908 9731
rect 12908 9295 14048 9731
rect 14048 9295 14066 9731
rect 12890 9285 14066 9295
<< metal3 >>
rect 2700 34631 13802 34664
tri 99 33575 1155 34631 se
rect 1155 34617 13802 34631
rect 1155 34553 2267 34617
rect 2331 34553 2350 34617
rect 2414 34553 2434 34617
rect 2498 34553 2518 34617
rect 2582 34553 2602 34617
rect 2666 34553 12332 34617
rect 12396 34553 12416 34617
rect 12480 34553 12500 34617
rect 12564 34553 12584 34617
rect 12648 34553 12668 34617
rect 12732 34553 13802 34617
rect 1155 34523 13802 34553
rect 1155 34459 2267 34523
rect 2331 34459 2350 34523
rect 2414 34459 2434 34523
rect 2498 34459 2518 34523
rect 2582 34459 2602 34523
rect 2666 34459 12332 34523
rect 12396 34459 12416 34523
rect 12480 34459 12500 34523
rect 12564 34459 12584 34523
rect 12648 34459 12668 34523
rect 12732 34459 13802 34523
rect 1155 34440 13802 34459
rect 1155 34376 2139 34440
rect 2203 34429 12795 34440
rect 2203 34376 2267 34429
rect 1155 34365 2267 34376
rect 2331 34365 2350 34429
rect 2414 34365 2434 34429
rect 2498 34365 2518 34429
rect 2582 34365 2602 34429
rect 2666 34365 12332 34429
rect 12396 34365 12416 34429
rect 12480 34365 12500 34429
rect 12564 34365 12584 34429
rect 12648 34365 12668 34429
rect 12732 34376 12795 34429
rect 12859 34376 13802 34440
rect 12732 34365 13802 34376
rect 1155 34335 13802 34365
rect 1155 34315 2267 34335
rect 1155 34251 1995 34315
rect 2059 34251 2075 34315
rect 2139 34251 2155 34315
rect 2219 34271 2267 34315
rect 2331 34271 2350 34335
rect 2414 34271 2434 34335
rect 2498 34271 2518 34335
rect 2582 34271 2602 34335
rect 2666 34271 12332 34335
rect 12396 34271 12416 34335
rect 12480 34271 12500 34335
rect 12564 34271 12584 34335
rect 12648 34271 12668 34335
rect 12732 34315 13802 34335
rect 12732 34271 12779 34315
rect 2219 34251 12779 34271
rect 12843 34251 12859 34315
rect 12923 34251 12939 34315
rect 13003 34251 13802 34315
rect 1155 34241 13802 34251
rect 1155 34219 2267 34241
rect 1155 34182 1995 34219
rect 1155 34118 1881 34182
rect 1945 34155 1995 34182
rect 2059 34155 2075 34219
rect 2139 34155 2155 34219
rect 2219 34177 2267 34219
rect 2331 34177 2350 34241
rect 2414 34177 2434 34241
rect 2498 34177 2518 34241
rect 2582 34177 2602 34241
rect 2666 34177 12332 34241
rect 12396 34177 12416 34241
rect 12480 34177 12500 34241
rect 12564 34177 12584 34241
rect 12648 34177 12668 34241
rect 12732 34219 13802 34241
rect 12732 34177 12779 34219
rect 2219 34155 12779 34177
rect 12843 34155 12859 34219
rect 12923 34155 12939 34219
rect 13003 34182 13802 34219
rect 13003 34155 13053 34182
rect 1945 34147 13053 34155
rect 1945 34118 2267 34147
rect 1155 34083 2267 34118
rect 2331 34083 2350 34147
rect 2414 34083 2434 34147
rect 2498 34083 2518 34147
rect 2582 34083 2602 34147
rect 2666 34083 12332 34147
rect 12396 34083 12416 34147
rect 12480 34083 12500 34147
rect 12564 34083 12584 34147
rect 12648 34083 12668 34147
rect 12732 34118 13053 34147
rect 13117 34118 13802 34182
rect 12732 34083 13802 34118
rect 1155 34077 13802 34083
rect 1155 34013 1739 34077
rect 1803 34013 1828 34077
rect 1892 34013 1918 34077
rect 1982 34013 2008 34077
rect 2072 34013 2098 34077
rect 2162 34013 12836 34077
rect 12900 34013 12926 34077
rect 12990 34013 13016 34077
rect 13080 34013 13106 34077
rect 13170 34013 13195 34077
rect 13259 34013 13802 34077
rect 1155 34008 13802 34013
rect 1155 33961 2238 34008
rect 1155 33897 1739 33961
rect 1803 33897 1828 33961
rect 1892 33897 1918 33961
rect 1982 33897 2008 33961
rect 2072 33897 2098 33961
rect 2162 33944 2238 33961
rect 2302 33944 12696 34008
rect 12760 33961 13802 34008
rect 12760 33944 12836 33961
rect 2162 33897 12836 33944
rect 12900 33897 12926 33961
rect 12990 33897 13016 33961
rect 13080 33897 13106 33961
rect 13170 33897 13195 33961
rect 13259 33897 13802 33961
rect 1155 33885 13802 33897
rect 1155 33821 1635 33885
rect 1699 33848 13299 33885
rect 1699 33845 2700 33848
rect 1699 33821 1739 33845
rect 1155 33781 1739 33821
rect 1803 33781 1828 33845
rect 1892 33781 1918 33845
rect 1982 33781 2008 33845
rect 2072 33781 2098 33845
rect 2162 33781 2700 33845
rect 1155 33753 2700 33781
rect 1155 33689 1415 33753
rect 1479 33689 1504 33753
rect 1568 33689 1594 33753
rect 1658 33689 1684 33753
rect 1748 33689 1774 33753
rect 1838 33720 2700 33753
rect 1838 33689 1920 33720
rect 1155 33656 1920 33689
rect 1984 33656 2700 33720
rect 1155 33637 2700 33656
rect 1155 33575 1415 33637
rect 99 33573 1415 33575
rect 1479 33573 1504 33637
rect 1568 33573 1594 33637
rect 1658 33573 1684 33637
rect 1748 33573 1774 33637
rect 1838 33573 2700 33637
rect 99 33557 2700 33573
rect 99 33493 1307 33557
rect 1371 33521 2700 33557
rect 1371 33493 1415 33521
rect 99 33457 1415 33493
rect 1479 33457 1504 33521
rect 1568 33457 1594 33521
rect 1658 33457 1684 33521
rect 1748 33457 1774 33521
rect 1838 33457 2700 33521
rect 99 33433 2700 33457
tri 2700 33448 3100 33848 nw
tri 11900 33448 12300 33848 ne
rect 12300 33845 13299 33848
rect 12300 33781 12836 33845
rect 12900 33781 12926 33845
rect 12990 33781 13016 33845
rect 13080 33781 13106 33845
rect 13170 33781 13195 33845
rect 13259 33821 13299 33845
rect 13363 33821 13802 33885
rect 13259 33781 13802 33821
rect 12300 33753 13802 33781
rect 12300 33720 13160 33753
rect 12300 33656 13014 33720
rect 13078 33689 13160 33720
rect 13224 33689 13250 33753
rect 13314 33689 13340 33753
rect 13404 33689 13430 33753
rect 13494 33689 13519 33753
rect 13583 33689 13802 33753
rect 13078 33656 13802 33689
rect 12300 33637 13802 33656
rect 12300 33573 13160 33637
rect 13224 33573 13250 33637
rect 13314 33573 13340 33637
rect 13404 33573 13430 33637
rect 13494 33573 13519 33637
rect 13583 33608 13802 33637
tri 13802 33608 14858 34664 sw
rect 13583 33573 14858 33608
rect 12300 33557 14858 33573
rect 12300 33521 13627 33557
rect 12300 33457 13160 33521
rect 13224 33457 13250 33521
rect 13314 33457 13340 33521
rect 13404 33457 13430 33521
rect 13494 33457 13519 33521
rect 13583 33493 13627 33521
rect 13691 33493 14858 33557
rect 13583 33457 14858 33493
rect 99 33369 1095 33433
rect 1159 33369 1184 33433
rect 1248 33369 1274 33433
rect 1338 33369 1364 33433
rect 1428 33369 1454 33433
rect 1518 33395 2700 33433
rect 1518 33369 1595 33395
rect 99 33331 1595 33369
rect 1659 33331 2700 33395
rect 99 33317 2700 33331
rect 99 33253 1095 33317
rect 1159 33253 1184 33317
rect 1248 33253 1274 33317
rect 1338 33253 1364 33317
rect 1428 33253 1454 33317
rect 1518 33253 2700 33317
rect 99 33201 2700 33253
rect 99 33137 1095 33201
rect 1159 33137 1184 33201
rect 1248 33137 1274 33201
rect 1338 33137 1364 33201
rect 1428 33137 1454 33201
rect 1518 33137 2700 33201
rect 99 33108 2700 33137
rect 99 33044 973 33108
rect 1037 33044 1063 33108
rect 1127 33044 1153 33108
rect 1217 33044 1243 33108
rect 1307 33044 1333 33108
rect 1397 33044 1423 33108
rect 1487 33044 2700 33108
rect 99 33028 2700 33044
rect 99 32964 973 33028
rect 1037 32964 1063 33028
rect 1127 32964 1153 33028
rect 1217 32964 1243 33028
rect 1307 32964 1333 33028
rect 1397 32964 1423 33028
rect 1487 32964 2700 33028
rect 99 32948 2700 32964
rect 99 32884 973 32948
rect 1037 32884 1063 32948
rect 1127 32884 1153 32948
rect 1217 32884 1243 32948
rect 1307 32884 1333 32948
rect 1397 32884 1423 32948
rect 1487 32884 2700 32948
rect 99 32868 2700 32884
rect 99 32804 973 32868
rect 1037 32804 1063 32868
rect 1127 32804 1153 32868
rect 1217 32804 1243 32868
rect 1307 32804 1333 32868
rect 1397 32804 1423 32868
rect 1487 32804 2700 32868
rect 99 32788 2700 32804
rect 99 32724 973 32788
rect 1037 32724 1063 32788
rect 1127 32724 1153 32788
rect 1217 32724 1243 32788
rect 1307 32724 1333 32788
rect 1397 32724 1423 32788
rect 1487 32724 2700 32788
rect 99 32708 2700 32724
rect 99 32644 973 32708
rect 1037 32644 1063 32708
rect 1127 32644 1153 32708
rect 1217 32644 1243 32708
rect 1307 32644 1333 32708
rect 1397 32644 1423 32708
rect 1487 32644 2700 32708
rect 99 32628 2700 32644
rect 99 32564 973 32628
rect 1037 32564 1063 32628
rect 1127 32564 1153 32628
rect 1217 32564 1243 32628
rect 1307 32564 1333 32628
rect 1397 32564 1423 32628
rect 1487 32564 2700 32628
rect 99 32548 2700 32564
rect 99 32484 973 32548
rect 1037 32484 1063 32548
rect 1127 32484 1153 32548
rect 1217 32484 1243 32548
rect 1307 32484 1333 32548
rect 1397 32484 1423 32548
rect 1487 32484 2700 32548
rect 99 32468 2700 32484
rect 99 32404 973 32468
rect 1037 32404 1063 32468
rect 1127 32404 1153 32468
rect 1217 32404 1243 32468
rect 1307 32404 1333 32468
rect 1397 32404 1423 32468
rect 1487 32404 2700 32468
rect 99 32388 2700 32404
rect 99 32324 973 32388
rect 1037 32324 1063 32388
rect 1127 32324 1153 32388
rect 1217 32324 1243 32388
rect 1307 32324 1333 32388
rect 1397 32324 1423 32388
rect 1487 32324 2700 32388
rect 99 32308 2700 32324
rect 99 32244 973 32308
rect 1037 32244 1063 32308
rect 1127 32244 1153 32308
rect 1217 32244 1243 32308
rect 1307 32244 1333 32308
rect 1397 32244 1423 32308
rect 1487 32244 2700 32308
rect 99 32228 2700 32244
rect 99 32164 973 32228
rect 1037 32164 1063 32228
rect 1127 32164 1153 32228
rect 1217 32164 1243 32228
rect 1307 32164 1333 32228
rect 1397 32164 1423 32228
rect 1487 32164 2700 32228
rect 99 32148 2700 32164
rect 99 32084 973 32148
rect 1037 32084 1063 32148
rect 1127 32084 1153 32148
rect 1217 32084 1243 32148
rect 1307 32084 1333 32148
rect 1397 32084 1423 32148
rect 1487 32084 2700 32148
rect 99 32068 2700 32084
rect 99 32004 973 32068
rect 1037 32004 1063 32068
rect 1127 32004 1153 32068
rect 1217 32004 1243 32068
rect 1307 32004 1333 32068
rect 1397 32004 1423 32068
rect 1487 32004 2700 32068
rect 99 31988 2700 32004
rect 99 31924 973 31988
rect 1037 31924 1063 31988
rect 1127 31924 1153 31988
rect 1217 31924 1243 31988
rect 1307 31924 1333 31988
rect 1397 31924 1423 31988
rect 1487 31924 2700 31988
rect 99 31908 2700 31924
rect 99 31844 973 31908
rect 1037 31844 1063 31908
rect 1127 31844 1153 31908
rect 1217 31844 1243 31908
rect 1307 31844 1333 31908
rect 1397 31844 1423 31908
rect 1487 31844 2700 31908
rect 99 31828 2700 31844
rect 99 31764 973 31828
rect 1037 31764 1063 31828
rect 1127 31764 1153 31828
rect 1217 31764 1243 31828
rect 1307 31764 1333 31828
rect 1397 31764 1423 31828
rect 1487 31764 2700 31828
rect 99 31748 2700 31764
rect 99 31684 973 31748
rect 1037 31684 1063 31748
rect 1127 31684 1153 31748
rect 1217 31684 1243 31748
rect 1307 31684 1333 31748
rect 1397 31684 1423 31748
rect 1487 31684 2700 31748
rect 99 31668 2700 31684
rect 99 31604 973 31668
rect 1037 31604 1063 31668
rect 1127 31604 1153 31668
rect 1217 31604 1243 31668
rect 1307 31604 1333 31668
rect 1397 31604 1423 31668
rect 1487 31604 2700 31668
rect 99 31588 2700 31604
rect 99 31524 973 31588
rect 1037 31524 1063 31588
rect 1127 31524 1153 31588
rect 1217 31524 1243 31588
rect 1307 31524 1333 31588
rect 1397 31524 1423 31588
rect 1487 31524 2700 31588
rect 99 31508 2700 31524
rect 99 31444 973 31508
rect 1037 31444 1063 31508
rect 1127 31444 1153 31508
rect 1217 31444 1243 31508
rect 1307 31444 1333 31508
rect 1397 31444 1423 31508
rect 1487 31444 2700 31508
rect 99 31428 2700 31444
rect 99 31364 973 31428
rect 1037 31364 1063 31428
rect 1127 31364 1153 31428
rect 1217 31364 1243 31428
rect 1307 31364 1333 31428
rect 1397 31364 1423 31428
rect 1487 31364 2700 31428
rect 99 31348 2700 31364
rect 99 31284 973 31348
rect 1037 31284 1063 31348
rect 1127 31284 1153 31348
rect 1217 31284 1243 31348
rect 1307 31284 1333 31348
rect 1397 31284 1423 31348
rect 1487 31284 2700 31348
rect 99 31268 2700 31284
rect 99 31204 973 31268
rect 1037 31204 1063 31268
rect 1127 31204 1153 31268
rect 1217 31204 1243 31268
rect 1307 31204 1333 31268
rect 1397 31204 1423 31268
rect 1487 31204 2700 31268
rect 99 31188 2700 31204
rect 99 31124 973 31188
rect 1037 31124 1063 31188
rect 1127 31124 1153 31188
rect 1217 31124 1243 31188
rect 1307 31124 1333 31188
rect 1397 31124 1423 31188
rect 1487 31124 2700 31188
rect 99 31108 2700 31124
rect 99 31044 973 31108
rect 1037 31044 1063 31108
rect 1127 31044 1153 31108
rect 1217 31044 1243 31108
rect 1307 31044 1333 31108
rect 1397 31044 1423 31108
rect 1487 31044 2700 31108
rect 99 31028 2700 31044
rect 99 30964 973 31028
rect 1037 30964 1063 31028
rect 1127 30964 1153 31028
rect 1217 30964 1243 31028
rect 1307 30964 1333 31028
rect 1397 30964 1423 31028
rect 1487 30964 2700 31028
rect 99 30948 2700 30964
rect 99 30884 973 30948
rect 1037 30884 1063 30948
rect 1127 30884 1153 30948
rect 1217 30884 1243 30948
rect 1307 30884 1333 30948
rect 1397 30884 1423 30948
rect 1487 30884 2700 30948
rect 99 30868 2700 30884
rect 99 30804 973 30868
rect 1037 30804 1063 30868
rect 1127 30804 1153 30868
rect 1217 30804 1243 30868
rect 1307 30804 1333 30868
rect 1397 30804 1423 30868
rect 1487 30804 2700 30868
rect 99 30788 2700 30804
rect 99 30724 973 30788
rect 1037 30724 1063 30788
rect 1127 30724 1153 30788
rect 1217 30724 1243 30788
rect 1307 30724 1333 30788
rect 1397 30724 1423 30788
rect 1487 30724 2700 30788
rect 99 30708 2700 30724
rect 99 30644 973 30708
rect 1037 30644 1063 30708
rect 1127 30644 1153 30708
rect 1217 30644 1243 30708
rect 1307 30644 1333 30708
rect 1397 30644 1423 30708
rect 1487 30644 2700 30708
rect 99 30628 2700 30644
rect 99 30564 973 30628
rect 1037 30564 1063 30628
rect 1127 30564 1153 30628
rect 1217 30564 1243 30628
rect 1307 30564 1333 30628
rect 1397 30564 1423 30628
rect 1487 30564 2700 30628
rect 99 30548 2700 30564
rect 99 30484 973 30548
rect 1037 30484 1063 30548
rect 1127 30484 1153 30548
rect 1217 30484 1243 30548
rect 1307 30484 1333 30548
rect 1397 30484 1423 30548
rect 1487 30484 2700 30548
rect 99 30468 2700 30484
rect 99 30404 973 30468
rect 1037 30404 1063 30468
rect 1127 30404 1153 30468
rect 1217 30404 1243 30468
rect 1307 30404 1333 30468
rect 1397 30404 1423 30468
rect 1487 30404 2700 30468
rect 99 30388 2700 30404
rect 99 30324 973 30388
rect 1037 30324 1063 30388
rect 1127 30324 1153 30388
rect 1217 30324 1243 30388
rect 1307 30324 1333 30388
rect 1397 30324 1423 30388
rect 1487 30324 2700 30388
rect 99 30308 2700 30324
rect 99 30244 973 30308
rect 1037 30244 1063 30308
rect 1127 30244 1153 30308
rect 1217 30244 1243 30308
rect 1307 30244 1333 30308
rect 1397 30244 1423 30308
rect 1487 30244 2700 30308
rect 99 30228 2700 30244
rect 99 30164 973 30228
rect 1037 30164 1063 30228
rect 1127 30164 1153 30228
rect 1217 30164 1243 30228
rect 1307 30164 1333 30228
rect 1397 30164 1423 30228
rect 1487 30164 2700 30228
rect 99 30148 2700 30164
rect 99 30084 973 30148
rect 1037 30084 1063 30148
rect 1127 30084 1153 30148
rect 1217 30084 1243 30148
rect 1307 30084 1333 30148
rect 1397 30084 1423 30148
rect 1487 30084 2700 30148
rect 99 30068 2700 30084
rect 99 30004 973 30068
rect 1037 30004 1063 30068
rect 1127 30004 1153 30068
rect 1217 30004 1243 30068
rect 1307 30004 1333 30068
rect 1397 30004 1423 30068
rect 1487 30004 2700 30068
rect 99 29988 2700 30004
rect 99 29924 973 29988
rect 1037 29924 1063 29988
rect 1127 29924 1153 29988
rect 1217 29924 1243 29988
rect 1307 29924 1333 29988
rect 1397 29924 1423 29988
rect 1487 29924 2700 29988
rect 99 29908 2700 29924
rect 99 29844 973 29908
rect 1037 29844 1063 29908
rect 1127 29844 1153 29908
rect 1217 29844 1243 29908
rect 1307 29844 1333 29908
rect 1397 29844 1423 29908
rect 1487 29844 2700 29908
rect 99 29828 2700 29844
rect 99 29764 973 29828
rect 1037 29764 1063 29828
rect 1127 29764 1153 29828
rect 1217 29764 1243 29828
rect 1307 29764 1333 29828
rect 1397 29764 1423 29828
rect 1487 29764 2700 29828
rect 99 29748 2700 29764
rect 99 29684 973 29748
rect 1037 29684 1063 29748
rect 1127 29684 1153 29748
rect 1217 29684 1243 29748
rect 1307 29684 1333 29748
rect 1397 29684 1423 29748
rect 1487 29684 2700 29748
rect 99 29668 2700 29684
rect 99 29604 973 29668
rect 1037 29604 1063 29668
rect 1127 29604 1153 29668
rect 1217 29604 1243 29668
rect 1307 29604 1333 29668
rect 1397 29604 1423 29668
rect 1487 29604 2700 29668
rect 99 29588 2700 29604
rect 99 29524 973 29588
rect 1037 29524 1063 29588
rect 1127 29524 1153 29588
rect 1217 29524 1243 29588
rect 1307 29524 1333 29588
rect 1397 29524 1423 29588
rect 1487 29524 2700 29588
rect 99 29508 2700 29524
rect 99 29444 973 29508
rect 1037 29444 1063 29508
rect 1127 29444 1153 29508
rect 1217 29444 1243 29508
rect 1307 29444 1333 29508
rect 1397 29444 1423 29508
rect 1487 29444 2700 29508
rect 99 29428 2700 29444
rect 99 29364 973 29428
rect 1037 29364 1063 29428
rect 1127 29364 1153 29428
rect 1217 29364 1243 29428
rect 1307 29364 1333 29428
rect 1397 29364 1423 29428
rect 1487 29364 2700 29428
rect 99 29348 2700 29364
rect 99 29284 973 29348
rect 1037 29284 1063 29348
rect 1127 29284 1153 29348
rect 1217 29284 1243 29348
rect 1307 29284 1333 29348
rect 1397 29284 1423 29348
rect 1487 29284 2700 29348
rect 99 29268 2700 29284
rect 99 29204 973 29268
rect 1037 29204 1063 29268
rect 1127 29204 1153 29268
rect 1217 29204 1243 29268
rect 1307 29204 1333 29268
rect 1397 29204 1423 29268
rect 1487 29204 2700 29268
rect 99 29188 2700 29204
rect 99 29124 973 29188
rect 1037 29124 1063 29188
rect 1127 29124 1153 29188
rect 1217 29124 1243 29188
rect 1307 29124 1333 29188
rect 1397 29124 1423 29188
rect 1487 29124 2700 29188
rect 99 29108 2700 29124
rect 99 29044 973 29108
rect 1037 29044 1063 29108
rect 1127 29044 1153 29108
rect 1217 29044 1243 29108
rect 1307 29044 1333 29108
rect 1397 29044 1423 29108
rect 1487 29044 2700 29108
rect 99 29028 2700 29044
rect 99 28964 973 29028
rect 1037 28964 1063 29028
rect 1127 28964 1153 29028
rect 1217 28964 1243 29028
rect 1307 28964 1333 29028
rect 1397 28964 1423 29028
rect 1487 28964 2700 29028
rect 99 28948 2700 28964
rect 99 28884 973 28948
rect 1037 28884 1063 28948
rect 1127 28884 1153 28948
rect 1217 28884 1243 28948
rect 1307 28884 1333 28948
rect 1397 28884 1423 28948
rect 1487 28884 2700 28948
rect 99 28868 2700 28884
rect 99 28804 973 28868
rect 1037 28804 1063 28868
rect 1127 28804 1153 28868
rect 1217 28804 1243 28868
rect 1307 28804 1333 28868
rect 1397 28804 1423 28868
rect 1487 28804 2700 28868
rect 99 28788 2700 28804
rect 99 28724 973 28788
rect 1037 28724 1063 28788
rect 1127 28724 1153 28788
rect 1217 28724 1243 28788
rect 1307 28724 1333 28788
rect 1397 28724 1423 28788
rect 1487 28724 2700 28788
rect 99 28708 2700 28724
rect 99 28644 973 28708
rect 1037 28644 1063 28708
rect 1127 28644 1153 28708
rect 1217 28644 1243 28708
rect 1307 28644 1333 28708
rect 1397 28644 1423 28708
rect 1487 28644 2700 28708
rect 99 28628 2700 28644
rect 99 28564 973 28628
rect 1037 28564 1063 28628
rect 1127 28564 1153 28628
rect 1217 28564 1243 28628
rect 1307 28564 1333 28628
rect 1397 28564 1423 28628
rect 1487 28564 2700 28628
rect 99 28548 2700 28564
rect 99 28484 973 28548
rect 1037 28484 1063 28548
rect 1127 28484 1153 28548
rect 1217 28484 1243 28548
rect 1307 28484 1333 28548
rect 1397 28484 1423 28548
rect 1487 28484 2700 28548
rect 99 28468 2700 28484
rect 99 28404 973 28468
rect 1037 28404 1063 28468
rect 1127 28404 1153 28468
rect 1217 28404 1243 28468
rect 1307 28404 1333 28468
rect 1397 28404 1423 28468
rect 1487 28404 2700 28468
rect 99 28388 2700 28404
rect 99 28324 973 28388
rect 1037 28324 1063 28388
rect 1127 28324 1153 28388
rect 1217 28324 1243 28388
rect 1307 28324 1333 28388
rect 1397 28324 1423 28388
rect 1487 28324 2700 28388
rect 99 28308 2700 28324
rect 99 28244 973 28308
rect 1037 28244 1063 28308
rect 1127 28244 1153 28308
rect 1217 28244 1243 28308
rect 1307 28244 1333 28308
rect 1397 28244 1423 28308
rect 1487 28244 2700 28308
rect 99 28228 2700 28244
rect 99 28164 973 28228
rect 1037 28164 1063 28228
rect 1127 28164 1153 28228
rect 1217 28164 1243 28228
rect 1307 28164 1333 28228
rect 1397 28164 1423 28228
rect 1487 28164 2700 28228
rect 99 28148 2700 28164
rect 99 28084 973 28148
rect 1037 28084 1063 28148
rect 1127 28084 1153 28148
rect 1217 28084 1243 28148
rect 1307 28084 1333 28148
rect 1397 28084 1423 28148
rect 1487 28084 2700 28148
rect 99 28068 2700 28084
rect 99 28004 973 28068
rect 1037 28004 1063 28068
rect 1127 28004 1153 28068
rect 1217 28004 1243 28068
rect 1307 28004 1333 28068
rect 1397 28004 1423 28068
rect 1487 28004 2700 28068
rect 99 27988 2700 28004
rect 99 27924 973 27988
rect 1037 27924 1063 27988
rect 1127 27924 1153 27988
rect 1217 27924 1243 27988
rect 1307 27924 1333 27988
rect 1397 27924 1423 27988
rect 1487 27924 2700 27988
rect 99 27908 2700 27924
rect 99 27844 973 27908
rect 1037 27844 1063 27908
rect 1127 27844 1153 27908
rect 1217 27844 1243 27908
rect 1307 27844 1333 27908
rect 1397 27844 1423 27908
rect 1487 27844 2700 27908
rect 99 27828 2700 27844
rect 99 27764 973 27828
rect 1037 27764 1063 27828
rect 1127 27764 1153 27828
rect 1217 27764 1243 27828
rect 1307 27764 1333 27828
rect 1397 27764 1423 27828
rect 1487 27764 2700 27828
rect 99 27748 2700 27764
rect 99 27684 973 27748
rect 1037 27684 1063 27748
rect 1127 27684 1153 27748
rect 1217 27684 1243 27748
rect 1307 27684 1333 27748
rect 1397 27684 1423 27748
rect 1487 27684 2700 27748
rect 99 27668 2700 27684
rect 99 27604 973 27668
rect 1037 27604 1063 27668
rect 1127 27604 1153 27668
rect 1217 27604 1243 27668
rect 1307 27604 1333 27668
rect 1397 27604 1423 27668
rect 1487 27604 2700 27668
rect 99 27588 2700 27604
rect 99 27524 973 27588
rect 1037 27524 1063 27588
rect 1127 27524 1153 27588
rect 1217 27524 1243 27588
rect 1307 27524 1333 27588
rect 1397 27524 1423 27588
rect 1487 27524 2700 27588
rect 99 27508 2700 27524
rect 99 27444 973 27508
rect 1037 27444 1063 27508
rect 1127 27444 1153 27508
rect 1217 27444 1243 27508
rect 1307 27444 1333 27508
rect 1397 27444 1423 27508
rect 1487 27444 2700 27508
rect 99 27428 2700 27444
rect 99 27364 973 27428
rect 1037 27364 1063 27428
rect 1127 27364 1153 27428
rect 1217 27364 1243 27428
rect 1307 27364 1333 27428
rect 1397 27364 1423 27428
rect 1487 27364 2700 27428
rect 99 27348 2700 27364
rect 99 27284 973 27348
rect 1037 27284 1063 27348
rect 1127 27284 1153 27348
rect 1217 27284 1243 27348
rect 1307 27284 1333 27348
rect 1397 27284 1423 27348
rect 1487 27284 2700 27348
rect 99 27268 2700 27284
rect 99 27204 973 27268
rect 1037 27204 1063 27268
rect 1127 27204 1153 27268
rect 1217 27204 1243 27268
rect 1307 27204 1333 27268
rect 1397 27204 1423 27268
rect 1487 27204 2700 27268
rect 99 27188 2700 27204
rect 99 27124 973 27188
rect 1037 27124 1063 27188
rect 1127 27124 1153 27188
rect 1217 27124 1243 27188
rect 1307 27124 1333 27188
rect 1397 27124 1423 27188
rect 1487 27124 2700 27188
rect 99 27108 2700 27124
rect 99 27044 973 27108
rect 1037 27044 1063 27108
rect 1127 27044 1153 27108
rect 1217 27044 1243 27108
rect 1307 27044 1333 27108
rect 1397 27044 1423 27108
rect 1487 27044 2700 27108
rect 99 27028 2700 27044
rect 99 26964 973 27028
rect 1037 26964 1063 27028
rect 1127 26964 1153 27028
rect 1217 26964 1243 27028
rect 1307 26964 1333 27028
rect 1397 26964 1423 27028
rect 1487 26964 2700 27028
rect 99 26948 2700 26964
rect 99 26884 973 26948
rect 1037 26884 1063 26948
rect 1127 26884 1153 26948
rect 1217 26884 1243 26948
rect 1307 26884 1333 26948
rect 1397 26884 1423 26948
rect 1487 26884 2700 26948
rect 99 26868 2700 26884
rect 99 26804 973 26868
rect 1037 26804 1063 26868
rect 1127 26804 1153 26868
rect 1217 26804 1243 26868
rect 1307 26804 1333 26868
rect 1397 26804 1423 26868
rect 1487 26804 2700 26868
rect 99 26788 2700 26804
rect 99 26724 973 26788
rect 1037 26724 1063 26788
rect 1127 26724 1153 26788
rect 1217 26724 1243 26788
rect 1307 26724 1333 26788
rect 1397 26724 1423 26788
rect 1487 26724 2700 26788
rect 99 26708 2700 26724
rect 99 26644 973 26708
rect 1037 26644 1063 26708
rect 1127 26644 1153 26708
rect 1217 26644 1243 26708
rect 1307 26644 1333 26708
rect 1397 26644 1423 26708
rect 1487 26644 2700 26708
rect 99 26628 2700 26644
rect 99 26564 973 26628
rect 1037 26564 1063 26628
rect 1127 26564 1153 26628
rect 1217 26564 1243 26628
rect 1307 26564 1333 26628
rect 1397 26564 1423 26628
rect 1487 26564 2700 26628
rect 99 26548 2700 26564
rect 99 26484 973 26548
rect 1037 26484 1063 26548
rect 1127 26484 1153 26548
rect 1217 26484 1243 26548
rect 1307 26484 1333 26548
rect 1397 26484 1423 26548
rect 1487 26484 2700 26548
rect 99 26468 2700 26484
rect 99 26404 973 26468
rect 1037 26404 1063 26468
rect 1127 26404 1153 26468
rect 1217 26404 1243 26468
rect 1307 26404 1333 26468
rect 1397 26404 1423 26468
rect 1487 26404 2700 26468
rect 99 26388 2700 26404
rect 99 26324 973 26388
rect 1037 26324 1063 26388
rect 1127 26324 1153 26388
rect 1217 26324 1243 26388
rect 1307 26324 1333 26388
rect 1397 26324 1423 26388
rect 1487 26324 2700 26388
rect 99 26308 2700 26324
rect 99 26244 973 26308
rect 1037 26244 1063 26308
rect 1127 26244 1153 26308
rect 1217 26244 1243 26308
rect 1307 26244 1333 26308
rect 1397 26244 1423 26308
rect 1487 26244 2700 26308
rect 99 26228 2700 26244
rect 99 26164 973 26228
rect 1037 26164 1063 26228
rect 1127 26164 1153 26228
rect 1217 26164 1243 26228
rect 1307 26164 1333 26228
rect 1397 26164 1423 26228
rect 1487 26164 2700 26228
rect 99 26148 2700 26164
rect 99 26084 973 26148
rect 1037 26084 1063 26148
rect 1127 26084 1153 26148
rect 1217 26084 1243 26148
rect 1307 26084 1333 26148
rect 1397 26084 1423 26148
rect 1487 26084 2700 26148
rect 99 26068 2700 26084
rect 99 26004 973 26068
rect 1037 26004 1063 26068
rect 1127 26004 1153 26068
rect 1217 26004 1243 26068
rect 1307 26004 1333 26068
rect 1397 26004 1423 26068
rect 1487 26004 2700 26068
rect 99 25988 2700 26004
rect 99 25924 973 25988
rect 1037 25924 1063 25988
rect 1127 25924 1153 25988
rect 1217 25924 1243 25988
rect 1307 25924 1333 25988
rect 1397 25924 1423 25988
rect 1487 25924 2700 25988
rect 99 25908 2700 25924
rect 99 25844 973 25908
rect 1037 25844 1063 25908
rect 1127 25844 1153 25908
rect 1217 25844 1243 25908
rect 1307 25844 1333 25908
rect 1397 25844 1423 25908
rect 1487 25844 2700 25908
rect 99 25828 2700 25844
rect 99 25764 973 25828
rect 1037 25764 1063 25828
rect 1127 25764 1153 25828
rect 1217 25764 1243 25828
rect 1307 25764 1333 25828
rect 1397 25764 1423 25828
rect 1487 25764 2700 25828
rect 99 25748 2700 25764
rect 99 25684 973 25748
rect 1037 25684 1063 25748
rect 1127 25684 1153 25748
rect 1217 25684 1243 25748
rect 1307 25684 1333 25748
rect 1397 25684 1423 25748
rect 1487 25684 2700 25748
rect 99 25668 2700 25684
rect 99 25604 973 25668
rect 1037 25604 1063 25668
rect 1127 25604 1153 25668
rect 1217 25604 1243 25668
rect 1307 25604 1333 25668
rect 1397 25604 1423 25668
rect 1487 25604 2700 25668
rect 99 25588 2700 25604
rect 99 25524 973 25588
rect 1037 25524 1063 25588
rect 1127 25524 1153 25588
rect 1217 25524 1243 25588
rect 1307 25524 1333 25588
rect 1397 25524 1423 25588
rect 1487 25524 2700 25588
rect 99 25508 2700 25524
rect 99 25444 973 25508
rect 1037 25444 1063 25508
rect 1127 25444 1153 25508
rect 1217 25444 1243 25508
rect 1307 25444 1333 25508
rect 1397 25444 1423 25508
rect 1487 25444 2700 25508
rect 99 25428 2700 25444
rect 99 25364 973 25428
rect 1037 25364 1063 25428
rect 1127 25364 1153 25428
rect 1217 25364 1243 25428
rect 1307 25364 1333 25428
rect 1397 25364 1423 25428
rect 1487 25364 2700 25428
rect 99 25348 2700 25364
rect 99 25284 973 25348
rect 1037 25284 1063 25348
rect 1127 25284 1153 25348
rect 1217 25284 1243 25348
rect 1307 25284 1333 25348
rect 1397 25284 1423 25348
rect 1487 25284 2700 25348
rect 99 25268 2700 25284
rect 99 25204 973 25268
rect 1037 25204 1063 25268
rect 1127 25204 1153 25268
rect 1217 25204 1243 25268
rect 1307 25204 1333 25268
rect 1397 25204 1423 25268
rect 1487 25204 2700 25268
rect 99 25188 2700 25204
rect 99 25124 973 25188
rect 1037 25124 1063 25188
rect 1127 25124 1153 25188
rect 1217 25124 1243 25188
rect 1307 25124 1333 25188
rect 1397 25124 1423 25188
rect 1487 25124 2700 25188
rect 99 25108 2700 25124
rect 99 25044 973 25108
rect 1037 25044 1063 25108
rect 1127 25044 1153 25108
rect 1217 25044 1243 25108
rect 1307 25044 1333 25108
rect 1397 25044 1423 25108
rect 1487 25044 2700 25108
rect 99 25028 2700 25044
rect 99 24964 973 25028
rect 1037 24964 1063 25028
rect 1127 24964 1153 25028
rect 1217 24964 1243 25028
rect 1307 24964 1333 25028
rect 1397 24964 1423 25028
rect 1487 24964 2700 25028
rect 99 24948 2700 24964
rect 99 24884 973 24948
rect 1037 24884 1063 24948
rect 1127 24884 1153 24948
rect 1217 24884 1243 24948
rect 1307 24884 1333 24948
rect 1397 24884 1423 24948
rect 1487 24884 2700 24948
rect 99 24868 2700 24884
rect 99 24804 973 24868
rect 1037 24804 1063 24868
rect 1127 24804 1153 24868
rect 1217 24804 1243 24868
rect 1307 24804 1333 24868
rect 1397 24804 1423 24868
rect 1487 24804 2700 24868
rect 99 24788 2700 24804
rect 99 24724 973 24788
rect 1037 24724 1063 24788
rect 1127 24724 1153 24788
rect 1217 24724 1243 24788
rect 1307 24724 1333 24788
rect 1397 24724 1423 24788
rect 1487 24724 2700 24788
rect 99 24708 2700 24724
rect 99 24644 973 24708
rect 1037 24644 1063 24708
rect 1127 24644 1153 24708
rect 1217 24644 1243 24708
rect 1307 24644 1333 24708
rect 1397 24644 1423 24708
rect 1487 24644 2700 24708
rect 99 24628 2700 24644
rect 99 24564 973 24628
rect 1037 24564 1063 24628
rect 1127 24564 1153 24628
rect 1217 24564 1243 24628
rect 1307 24564 1333 24628
rect 1397 24564 1423 24628
rect 1487 24564 2700 24628
rect 99 24548 2700 24564
rect 99 24484 973 24548
rect 1037 24484 1063 24548
rect 1127 24484 1153 24548
rect 1217 24484 1243 24548
rect 1307 24484 1333 24548
rect 1397 24484 1423 24548
rect 1487 24484 2700 24548
rect 99 24468 2700 24484
rect 99 24404 973 24468
rect 1037 24404 1063 24468
rect 1127 24404 1153 24468
rect 1217 24404 1243 24468
rect 1307 24404 1333 24468
rect 1397 24404 1423 24468
rect 1487 24404 2700 24468
rect 99 24388 2700 24404
rect 99 24324 973 24388
rect 1037 24324 1063 24388
rect 1127 24324 1153 24388
rect 1217 24324 1243 24388
rect 1307 24324 1333 24388
rect 1397 24324 1423 24388
rect 1487 24324 2700 24388
rect 99 24308 2700 24324
rect 99 24244 973 24308
rect 1037 24244 1063 24308
rect 1127 24244 1153 24308
rect 1217 24244 1243 24308
rect 1307 24244 1333 24308
rect 1397 24244 1423 24308
rect 1487 24244 2700 24308
rect 99 24228 2700 24244
rect 99 24164 973 24228
rect 1037 24164 1063 24228
rect 1127 24164 1153 24228
rect 1217 24164 1243 24228
rect 1307 24164 1333 24228
rect 1397 24164 1423 24228
rect 1487 24164 2700 24228
rect 99 24148 2700 24164
rect 99 24084 973 24148
rect 1037 24084 1063 24148
rect 1127 24084 1153 24148
rect 1217 24084 1243 24148
rect 1307 24084 1333 24148
rect 1397 24084 1423 24148
rect 1487 24084 2700 24148
rect 99 24068 2700 24084
rect 99 24004 973 24068
rect 1037 24004 1063 24068
rect 1127 24004 1153 24068
rect 1217 24004 1243 24068
rect 1307 24004 1333 24068
rect 1397 24004 1423 24068
rect 1487 24004 2700 24068
rect 99 23988 2700 24004
rect 99 23924 973 23988
rect 1037 23924 1063 23988
rect 1127 23924 1153 23988
rect 1217 23924 1243 23988
rect 1307 23924 1333 23988
rect 1397 23924 1423 23988
rect 1487 23924 2700 23988
rect 99 23908 2700 23924
rect 99 23844 973 23908
rect 1037 23844 1063 23908
rect 1127 23844 1153 23908
rect 1217 23844 1243 23908
rect 1307 23844 1333 23908
rect 1397 23844 1423 23908
rect 1487 23844 2700 23908
rect 99 23828 2700 23844
rect 99 23764 973 23828
rect 1037 23764 1063 23828
rect 1127 23764 1153 23828
rect 1217 23764 1243 23828
rect 1307 23764 1333 23828
rect 1397 23764 1423 23828
rect 1487 23764 2700 23828
rect 99 23748 2700 23764
rect 99 23684 973 23748
rect 1037 23684 1063 23748
rect 1127 23684 1153 23748
rect 1217 23684 1243 23748
rect 1307 23684 1333 23748
rect 1397 23684 1423 23748
rect 1487 23684 2700 23748
rect 99 23668 2700 23684
rect 99 23604 973 23668
rect 1037 23604 1063 23668
rect 1127 23604 1153 23668
rect 1217 23604 1243 23668
rect 1307 23604 1333 23668
rect 1397 23604 1423 23668
rect 1487 23604 2700 23668
rect 99 23588 2700 23604
rect 99 23524 973 23588
rect 1037 23524 1063 23588
rect 1127 23524 1153 23588
rect 1217 23524 1243 23588
rect 1307 23524 1333 23588
rect 1397 23524 1423 23588
rect 1487 23524 2700 23588
rect 99 23508 2700 23524
rect 99 23444 973 23508
rect 1037 23444 1063 23508
rect 1127 23444 1153 23508
rect 1217 23444 1243 23508
rect 1307 23444 1333 23508
rect 1397 23444 1423 23508
rect 1487 23444 2700 23508
rect 99 23428 2700 23444
rect 99 23364 973 23428
rect 1037 23364 1063 23428
rect 1127 23364 1153 23428
rect 1217 23364 1243 23428
rect 1307 23364 1333 23428
rect 1397 23364 1423 23428
rect 1487 23364 2700 23428
rect 99 23348 2700 23364
rect 99 23284 973 23348
rect 1037 23284 1063 23348
rect 1127 23284 1153 23348
rect 1217 23284 1243 23348
rect 1307 23284 1333 23348
rect 1397 23284 1423 23348
rect 1487 23284 2700 23348
rect 99 23267 2700 23284
rect 99 23203 973 23267
rect 1037 23203 1063 23267
rect 1127 23203 1153 23267
rect 1217 23203 1243 23267
rect 1307 23203 1333 23267
rect 1397 23203 1423 23267
rect 1487 23203 2700 23267
rect 99 23186 2700 23203
rect 99 23122 973 23186
rect 1037 23122 1063 23186
rect 1127 23122 1153 23186
rect 1217 23122 1243 23186
rect 1307 23122 1333 23186
rect 1397 23122 1423 23186
rect 1487 23122 2700 23186
rect 99 23105 2700 23122
rect 99 23041 973 23105
rect 1037 23041 1063 23105
rect 1127 23041 1153 23105
rect 1217 23041 1243 23105
rect 1307 23041 1333 23105
rect 1397 23041 1423 23105
rect 1487 23041 2700 23105
rect 99 23024 2700 23041
rect 99 22960 973 23024
rect 1037 22960 1063 23024
rect 1127 22960 1153 23024
rect 1217 22960 1243 23024
rect 1307 22960 1333 23024
rect 1397 22960 1423 23024
rect 1487 22960 2700 23024
rect 99 22943 2700 22960
rect 99 22879 973 22943
rect 1037 22879 1063 22943
rect 1127 22879 1153 22943
rect 1217 22879 1243 22943
rect 1307 22879 1333 22943
rect 1397 22879 1423 22943
rect 1487 22879 2700 22943
rect 99 22862 2700 22879
rect 99 22798 973 22862
rect 1037 22798 1063 22862
rect 1127 22798 1153 22862
rect 1217 22798 1243 22862
rect 1307 22798 1333 22862
rect 1397 22798 1423 22862
rect 1487 22798 2700 22862
rect 99 22781 2700 22798
rect 99 22717 973 22781
rect 1037 22717 1063 22781
rect 1127 22717 1153 22781
rect 1217 22717 1243 22781
rect 1307 22717 1333 22781
rect 1397 22717 1423 22781
rect 1487 22717 2700 22781
rect 99 22700 2700 22717
rect 99 22636 973 22700
rect 1037 22636 1063 22700
rect 1127 22636 1153 22700
rect 1217 22636 1243 22700
rect 1307 22636 1333 22700
rect 1397 22636 1423 22700
rect 1487 22636 2700 22700
rect 99 22619 2700 22636
rect 99 22555 973 22619
rect 1037 22555 1063 22619
rect 1127 22555 1153 22619
rect 1217 22555 1243 22619
rect 1307 22555 1333 22619
rect 1397 22555 1423 22619
rect 1487 22555 2700 22619
rect 99 22538 2700 22555
rect 99 22474 973 22538
rect 1037 22474 1063 22538
rect 1127 22474 1153 22538
rect 1217 22474 1243 22538
rect 1307 22474 1333 22538
rect 1397 22474 1423 22538
rect 1487 22474 2700 22538
rect 99 22457 2700 22474
rect 99 22393 973 22457
rect 1037 22393 1063 22457
rect 1127 22393 1153 22457
rect 1217 22393 1243 22457
rect 1307 22393 1333 22457
rect 1397 22393 1423 22457
rect 1487 22393 2700 22457
rect 99 22376 2700 22393
rect 99 22312 973 22376
rect 1037 22312 1063 22376
rect 1127 22312 1153 22376
rect 1217 22312 1243 22376
rect 1307 22312 1333 22376
rect 1397 22312 1423 22376
rect 1487 22312 2700 22376
rect 99 22295 2700 22312
rect 99 22231 973 22295
rect 1037 22231 1063 22295
rect 1127 22231 1153 22295
rect 1217 22231 1243 22295
rect 1307 22231 1333 22295
rect 1397 22231 1423 22295
rect 1487 22231 2700 22295
rect 99 22214 2700 22231
rect 99 22150 973 22214
rect 1037 22150 1063 22214
rect 1127 22150 1153 22214
rect 1217 22150 1243 22214
rect 1307 22150 1333 22214
rect 1397 22150 1423 22214
rect 1487 22150 2700 22214
rect 99 22133 2700 22150
rect 99 22069 973 22133
rect 1037 22069 1063 22133
rect 1127 22069 1153 22133
rect 1217 22069 1243 22133
rect 1307 22069 1333 22133
rect 1397 22069 1423 22133
rect 1487 22069 2700 22133
rect 99 22052 2700 22069
rect 99 21988 973 22052
rect 1037 21988 1063 22052
rect 1127 21988 1153 22052
rect 1217 21988 1243 22052
rect 1307 21988 1333 22052
rect 1397 21988 1423 22052
rect 1487 21988 2700 22052
rect 99 21971 2700 21988
rect 99 21907 973 21971
rect 1037 21907 1063 21971
rect 1127 21907 1153 21971
rect 1217 21907 1243 21971
rect 1307 21907 1333 21971
rect 1397 21907 1423 21971
rect 1487 21907 2700 21971
rect 99 21890 2700 21907
rect 99 21826 973 21890
rect 1037 21826 1063 21890
rect 1127 21826 1153 21890
rect 1217 21826 1243 21890
rect 1307 21826 1333 21890
rect 1397 21826 1423 21890
rect 1487 21826 2700 21890
rect 99 21809 2700 21826
rect 99 21745 973 21809
rect 1037 21745 1063 21809
rect 1127 21745 1153 21809
rect 1217 21745 1243 21809
rect 1307 21745 1333 21809
rect 1397 21745 1423 21809
rect 1487 21745 2700 21809
rect 99 21728 2700 21745
rect 99 21664 973 21728
rect 1037 21664 1063 21728
rect 1127 21664 1153 21728
rect 1217 21664 1243 21728
rect 1307 21664 1333 21728
rect 1397 21664 1423 21728
rect 1487 21664 2700 21728
rect 99 21647 2700 21664
rect 99 21583 973 21647
rect 1037 21583 1063 21647
rect 1127 21583 1153 21647
rect 1217 21583 1243 21647
rect 1307 21583 1333 21647
rect 1397 21583 1423 21647
rect 1487 21583 2700 21647
rect 99 21566 2700 21583
rect 99 21502 973 21566
rect 1037 21502 1063 21566
rect 1127 21502 1153 21566
rect 1217 21502 1243 21566
rect 1307 21502 1333 21566
rect 1397 21502 1423 21566
rect 1487 21502 2700 21566
rect 99 21485 2700 21502
rect 99 21421 973 21485
rect 1037 21421 1063 21485
rect 1127 21421 1153 21485
rect 1217 21421 1243 21485
rect 1307 21421 1333 21485
rect 1397 21421 1423 21485
rect 1487 21421 2700 21485
rect 99 21404 2700 21421
rect 99 21340 973 21404
rect 1037 21340 1063 21404
rect 1127 21340 1153 21404
rect 1217 21340 1243 21404
rect 1307 21340 1333 21404
rect 1397 21340 1423 21404
rect 1487 21340 2700 21404
rect 99 21323 2700 21340
rect 99 21259 973 21323
rect 1037 21259 1063 21323
rect 1127 21259 1153 21323
rect 1217 21259 1243 21323
rect 1307 21259 1333 21323
rect 1397 21259 1423 21323
rect 1487 21259 2700 21323
rect 99 21242 2700 21259
rect 99 21178 973 21242
rect 1037 21178 1063 21242
rect 1127 21178 1153 21242
rect 1217 21178 1243 21242
rect 1307 21178 1333 21242
rect 1397 21178 1423 21242
rect 1487 21178 2700 21242
rect 99 21161 2700 21178
rect 99 21097 973 21161
rect 1037 21097 1063 21161
rect 1127 21097 1153 21161
rect 1217 21097 1243 21161
rect 1307 21097 1333 21161
rect 1397 21097 1423 21161
rect 1487 21097 2700 21161
rect 99 21080 2700 21097
rect 99 21016 973 21080
rect 1037 21016 1063 21080
rect 1127 21016 1153 21080
rect 1217 21016 1243 21080
rect 1307 21016 1333 21080
rect 1397 21016 1423 21080
rect 1487 21016 2700 21080
rect 99 20999 2700 21016
rect 99 20935 973 20999
rect 1037 20935 1063 20999
rect 1127 20935 1153 20999
rect 1217 20935 1243 20999
rect 1307 20935 1333 20999
rect 1397 20935 1423 20999
rect 1487 20938 2700 20999
rect 1487 20935 1522 20938
rect 99 20918 1522 20935
rect 99 20854 973 20918
rect 1037 20854 1063 20918
rect 1127 20854 1153 20918
rect 1217 20854 1243 20918
rect 1307 20854 1333 20918
rect 1397 20854 1423 20918
rect 1487 20874 1522 20918
rect 1586 20874 2700 20938
rect 1487 20854 2700 20874
rect 99 20824 2700 20854
rect 99 20782 1303 20824
rect 99 20718 1132 20782
rect 1196 20760 1303 20782
rect 1367 20760 1392 20824
rect 1456 20760 1482 20824
rect 1546 20760 1572 20824
rect 1636 20760 1662 20824
rect 1726 20760 2700 20824
rect 1196 20718 2700 20760
rect 99 20708 2700 20718
rect 99 20644 1303 20708
rect 1367 20644 1392 20708
rect 1456 20644 1482 20708
rect 1546 20644 1572 20708
rect 1636 20644 1662 20708
rect 1726 20644 2700 20708
rect 99 20630 2700 20644
rect 99 20592 1803 20630
rect 99 20528 1303 20592
rect 1367 20528 1392 20592
rect 1456 20528 1482 20592
rect 1546 20528 1572 20592
rect 1636 20528 1662 20592
rect 1726 20566 1803 20592
rect 1867 20566 2700 20630
rect 1726 20528 2700 20566
rect 99 20504 2700 20528
rect 99 20468 1623 20504
rect 99 20404 1515 20468
rect 1579 20440 1623 20468
rect 1687 20440 1712 20504
rect 1776 20440 1802 20504
rect 1866 20440 1892 20504
rect 1956 20440 1982 20504
rect 2046 20440 2700 20504
rect 1579 20404 2700 20440
rect 99 20388 2700 20404
rect 99 20324 1623 20388
rect 1687 20324 1712 20388
rect 1776 20324 1802 20388
rect 1866 20324 1892 20388
rect 1956 20324 1982 20388
rect 2046 20324 2700 20388
rect 99 20305 2700 20324
rect 99 20272 2128 20305
rect 99 20208 1623 20272
rect 1687 20208 1712 20272
rect 1776 20208 1802 20272
rect 1866 20208 1892 20272
rect 1956 20208 1982 20272
rect 2046 20241 2128 20272
rect 2192 20241 2700 20305
rect 12300 33433 14858 33457
rect 12300 33395 13480 33433
rect 12300 33331 13339 33395
rect 13403 33369 13480 33395
rect 13544 33369 13570 33433
rect 13634 33369 13660 33433
rect 13724 33369 13750 33433
rect 13814 33369 13839 33433
rect 13903 33369 14858 33433
rect 13403 33331 14858 33369
rect 12300 33317 14858 33331
rect 12300 33253 13480 33317
rect 13544 33253 13570 33317
rect 13634 33253 13660 33317
rect 13724 33253 13750 33317
rect 13814 33253 13839 33317
rect 13903 33253 14858 33317
rect 12300 33201 14858 33253
rect 12300 33137 13480 33201
rect 13544 33137 13570 33201
rect 13634 33137 13660 33201
rect 13724 33137 13750 33201
rect 13814 33137 13839 33201
rect 13903 33137 14858 33201
rect 12300 33108 14858 33137
rect 12300 33044 13511 33108
rect 13575 33044 13601 33108
rect 13665 33044 13691 33108
rect 13755 33044 13781 33108
rect 13845 33044 13871 33108
rect 13935 33044 13961 33108
rect 14025 33044 14858 33108
rect 12300 33028 14858 33044
rect 12300 32964 13511 33028
rect 13575 32964 13601 33028
rect 13665 32964 13691 33028
rect 13755 32964 13781 33028
rect 13845 32964 13871 33028
rect 13935 32964 13961 33028
rect 14025 32964 14858 33028
rect 12300 32948 14858 32964
rect 12300 32884 13511 32948
rect 13575 32884 13601 32948
rect 13665 32884 13691 32948
rect 13755 32884 13781 32948
rect 13845 32884 13871 32948
rect 13935 32884 13961 32948
rect 14025 32884 14858 32948
rect 12300 32868 14858 32884
rect 12300 32804 13511 32868
rect 13575 32804 13601 32868
rect 13665 32804 13691 32868
rect 13755 32804 13781 32868
rect 13845 32804 13871 32868
rect 13935 32804 13961 32868
rect 14025 32804 14858 32868
rect 12300 32788 14858 32804
rect 12300 32724 13511 32788
rect 13575 32724 13601 32788
rect 13665 32724 13691 32788
rect 13755 32724 13781 32788
rect 13845 32724 13871 32788
rect 13935 32724 13961 32788
rect 14025 32724 14858 32788
rect 12300 32708 14858 32724
rect 12300 32644 13511 32708
rect 13575 32644 13601 32708
rect 13665 32644 13691 32708
rect 13755 32644 13781 32708
rect 13845 32644 13871 32708
rect 13935 32644 13961 32708
rect 14025 32644 14858 32708
rect 12300 32628 14858 32644
rect 12300 32564 13511 32628
rect 13575 32564 13601 32628
rect 13665 32564 13691 32628
rect 13755 32564 13781 32628
rect 13845 32564 13871 32628
rect 13935 32564 13961 32628
rect 14025 32564 14858 32628
rect 12300 32548 14858 32564
rect 12300 32484 13511 32548
rect 13575 32484 13601 32548
rect 13665 32484 13691 32548
rect 13755 32484 13781 32548
rect 13845 32484 13871 32548
rect 13935 32484 13961 32548
rect 14025 32484 14858 32548
rect 12300 32468 14858 32484
rect 12300 32404 13511 32468
rect 13575 32404 13601 32468
rect 13665 32404 13691 32468
rect 13755 32404 13781 32468
rect 13845 32404 13871 32468
rect 13935 32404 13961 32468
rect 14025 32404 14858 32468
rect 12300 32388 14858 32404
rect 12300 32324 13511 32388
rect 13575 32324 13601 32388
rect 13665 32324 13691 32388
rect 13755 32324 13781 32388
rect 13845 32324 13871 32388
rect 13935 32324 13961 32388
rect 14025 32324 14858 32388
rect 12300 32308 14858 32324
rect 12300 32244 13511 32308
rect 13575 32244 13601 32308
rect 13665 32244 13691 32308
rect 13755 32244 13781 32308
rect 13845 32244 13871 32308
rect 13935 32244 13961 32308
rect 14025 32244 14858 32308
rect 12300 32228 14858 32244
rect 12300 32164 13511 32228
rect 13575 32164 13601 32228
rect 13665 32164 13691 32228
rect 13755 32164 13781 32228
rect 13845 32164 13871 32228
rect 13935 32164 13961 32228
rect 14025 32164 14858 32228
rect 12300 32148 14858 32164
rect 12300 32084 13511 32148
rect 13575 32084 13601 32148
rect 13665 32084 13691 32148
rect 13755 32084 13781 32148
rect 13845 32084 13871 32148
rect 13935 32084 13961 32148
rect 14025 32084 14858 32148
rect 12300 32068 14858 32084
rect 12300 32004 13511 32068
rect 13575 32004 13601 32068
rect 13665 32004 13691 32068
rect 13755 32004 13781 32068
rect 13845 32004 13871 32068
rect 13935 32004 13961 32068
rect 14025 32004 14858 32068
rect 12300 31988 14858 32004
rect 12300 31924 13511 31988
rect 13575 31924 13601 31988
rect 13665 31924 13691 31988
rect 13755 31924 13781 31988
rect 13845 31924 13871 31988
rect 13935 31924 13961 31988
rect 14025 31924 14858 31988
rect 12300 31908 14858 31924
rect 12300 31844 13511 31908
rect 13575 31844 13601 31908
rect 13665 31844 13691 31908
rect 13755 31844 13781 31908
rect 13845 31844 13871 31908
rect 13935 31844 13961 31908
rect 14025 31844 14858 31908
rect 12300 31828 14858 31844
rect 12300 31764 13511 31828
rect 13575 31764 13601 31828
rect 13665 31764 13691 31828
rect 13755 31764 13781 31828
rect 13845 31764 13871 31828
rect 13935 31764 13961 31828
rect 14025 31764 14858 31828
rect 12300 31748 14858 31764
rect 12300 31684 13511 31748
rect 13575 31684 13601 31748
rect 13665 31684 13691 31748
rect 13755 31684 13781 31748
rect 13845 31684 13871 31748
rect 13935 31684 13961 31748
rect 14025 31684 14858 31748
rect 12300 31668 14858 31684
rect 12300 31604 13511 31668
rect 13575 31604 13601 31668
rect 13665 31604 13691 31668
rect 13755 31604 13781 31668
rect 13845 31604 13871 31668
rect 13935 31604 13961 31668
rect 14025 31604 14858 31668
rect 12300 31588 14858 31604
rect 12300 31524 13511 31588
rect 13575 31524 13601 31588
rect 13665 31524 13691 31588
rect 13755 31524 13781 31588
rect 13845 31524 13871 31588
rect 13935 31524 13961 31588
rect 14025 31524 14858 31588
rect 12300 31508 14858 31524
rect 12300 31444 13511 31508
rect 13575 31444 13601 31508
rect 13665 31444 13691 31508
rect 13755 31444 13781 31508
rect 13845 31444 13871 31508
rect 13935 31444 13961 31508
rect 14025 31444 14858 31508
rect 12300 31428 14858 31444
rect 12300 31364 13511 31428
rect 13575 31364 13601 31428
rect 13665 31364 13691 31428
rect 13755 31364 13781 31428
rect 13845 31364 13871 31428
rect 13935 31364 13961 31428
rect 14025 31364 14858 31428
rect 12300 31348 14858 31364
rect 12300 31284 13511 31348
rect 13575 31284 13601 31348
rect 13665 31284 13691 31348
rect 13755 31284 13781 31348
rect 13845 31284 13871 31348
rect 13935 31284 13961 31348
rect 14025 31284 14858 31348
rect 12300 31268 14858 31284
rect 12300 31204 13511 31268
rect 13575 31204 13601 31268
rect 13665 31204 13691 31268
rect 13755 31204 13781 31268
rect 13845 31204 13871 31268
rect 13935 31204 13961 31268
rect 14025 31204 14858 31268
rect 12300 31188 14858 31204
rect 12300 31124 13511 31188
rect 13575 31124 13601 31188
rect 13665 31124 13691 31188
rect 13755 31124 13781 31188
rect 13845 31124 13871 31188
rect 13935 31124 13961 31188
rect 14025 31124 14858 31188
rect 12300 31108 14858 31124
rect 12300 31044 13511 31108
rect 13575 31044 13601 31108
rect 13665 31044 13691 31108
rect 13755 31044 13781 31108
rect 13845 31044 13871 31108
rect 13935 31044 13961 31108
rect 14025 31044 14858 31108
rect 12300 31028 14858 31044
rect 12300 30964 13511 31028
rect 13575 30964 13601 31028
rect 13665 30964 13691 31028
rect 13755 30964 13781 31028
rect 13845 30964 13871 31028
rect 13935 30964 13961 31028
rect 14025 30964 14858 31028
rect 12300 30948 14858 30964
rect 12300 30884 13511 30948
rect 13575 30884 13601 30948
rect 13665 30884 13691 30948
rect 13755 30884 13781 30948
rect 13845 30884 13871 30948
rect 13935 30884 13961 30948
rect 14025 30884 14858 30948
rect 12300 30868 14858 30884
rect 12300 30804 13511 30868
rect 13575 30804 13601 30868
rect 13665 30804 13691 30868
rect 13755 30804 13781 30868
rect 13845 30804 13871 30868
rect 13935 30804 13961 30868
rect 14025 30804 14858 30868
rect 12300 30788 14858 30804
rect 12300 30724 13511 30788
rect 13575 30724 13601 30788
rect 13665 30724 13691 30788
rect 13755 30724 13781 30788
rect 13845 30724 13871 30788
rect 13935 30724 13961 30788
rect 14025 30724 14858 30788
rect 12300 30708 14858 30724
rect 12300 30644 13511 30708
rect 13575 30644 13601 30708
rect 13665 30644 13691 30708
rect 13755 30644 13781 30708
rect 13845 30644 13871 30708
rect 13935 30644 13961 30708
rect 14025 30644 14858 30708
rect 12300 30628 14858 30644
rect 12300 30564 13511 30628
rect 13575 30564 13601 30628
rect 13665 30564 13691 30628
rect 13755 30564 13781 30628
rect 13845 30564 13871 30628
rect 13935 30564 13961 30628
rect 14025 30564 14858 30628
rect 12300 30548 14858 30564
rect 12300 30484 13511 30548
rect 13575 30484 13601 30548
rect 13665 30484 13691 30548
rect 13755 30484 13781 30548
rect 13845 30484 13871 30548
rect 13935 30484 13961 30548
rect 14025 30484 14858 30548
rect 12300 30468 14858 30484
rect 12300 30404 13511 30468
rect 13575 30404 13601 30468
rect 13665 30404 13691 30468
rect 13755 30404 13781 30468
rect 13845 30404 13871 30468
rect 13935 30404 13961 30468
rect 14025 30404 14858 30468
rect 12300 30388 14858 30404
rect 12300 30324 13511 30388
rect 13575 30324 13601 30388
rect 13665 30324 13691 30388
rect 13755 30324 13781 30388
rect 13845 30324 13871 30388
rect 13935 30324 13961 30388
rect 14025 30324 14858 30388
rect 12300 30308 14858 30324
rect 12300 30244 13511 30308
rect 13575 30244 13601 30308
rect 13665 30244 13691 30308
rect 13755 30244 13781 30308
rect 13845 30244 13871 30308
rect 13935 30244 13961 30308
rect 14025 30244 14858 30308
rect 12300 30228 14858 30244
rect 12300 30164 13511 30228
rect 13575 30164 13601 30228
rect 13665 30164 13691 30228
rect 13755 30164 13781 30228
rect 13845 30164 13871 30228
rect 13935 30164 13961 30228
rect 14025 30164 14858 30228
rect 12300 30148 14858 30164
rect 12300 30084 13511 30148
rect 13575 30084 13601 30148
rect 13665 30084 13691 30148
rect 13755 30084 13781 30148
rect 13845 30084 13871 30148
rect 13935 30084 13961 30148
rect 14025 30084 14858 30148
rect 12300 30068 14858 30084
rect 12300 30004 13511 30068
rect 13575 30004 13601 30068
rect 13665 30004 13691 30068
rect 13755 30004 13781 30068
rect 13845 30004 13871 30068
rect 13935 30004 13961 30068
rect 14025 30004 14858 30068
rect 12300 29988 14858 30004
rect 12300 29924 13511 29988
rect 13575 29924 13601 29988
rect 13665 29924 13691 29988
rect 13755 29924 13781 29988
rect 13845 29924 13871 29988
rect 13935 29924 13961 29988
rect 14025 29924 14858 29988
rect 12300 29908 14858 29924
rect 12300 29844 13511 29908
rect 13575 29844 13601 29908
rect 13665 29844 13691 29908
rect 13755 29844 13781 29908
rect 13845 29844 13871 29908
rect 13935 29844 13961 29908
rect 14025 29844 14858 29908
rect 12300 29828 14858 29844
rect 12300 29764 13511 29828
rect 13575 29764 13601 29828
rect 13665 29764 13691 29828
rect 13755 29764 13781 29828
rect 13845 29764 13871 29828
rect 13935 29764 13961 29828
rect 14025 29764 14858 29828
rect 12300 29748 14858 29764
rect 12300 29684 13511 29748
rect 13575 29684 13601 29748
rect 13665 29684 13691 29748
rect 13755 29684 13781 29748
rect 13845 29684 13871 29748
rect 13935 29684 13961 29748
rect 14025 29684 14858 29748
rect 12300 29668 14858 29684
rect 12300 29604 13511 29668
rect 13575 29604 13601 29668
rect 13665 29604 13691 29668
rect 13755 29604 13781 29668
rect 13845 29604 13871 29668
rect 13935 29604 13961 29668
rect 14025 29604 14858 29668
rect 12300 29588 14858 29604
rect 12300 29524 13511 29588
rect 13575 29524 13601 29588
rect 13665 29524 13691 29588
rect 13755 29524 13781 29588
rect 13845 29524 13871 29588
rect 13935 29524 13961 29588
rect 14025 29524 14858 29588
rect 12300 29508 14858 29524
rect 12300 29444 13511 29508
rect 13575 29444 13601 29508
rect 13665 29444 13691 29508
rect 13755 29444 13781 29508
rect 13845 29444 13871 29508
rect 13935 29444 13961 29508
rect 14025 29444 14858 29508
rect 12300 29428 14858 29444
rect 12300 29364 13511 29428
rect 13575 29364 13601 29428
rect 13665 29364 13691 29428
rect 13755 29364 13781 29428
rect 13845 29364 13871 29428
rect 13935 29364 13961 29428
rect 14025 29364 14858 29428
rect 12300 29348 14858 29364
rect 12300 29284 13511 29348
rect 13575 29284 13601 29348
rect 13665 29284 13691 29348
rect 13755 29284 13781 29348
rect 13845 29284 13871 29348
rect 13935 29284 13961 29348
rect 14025 29284 14858 29348
rect 12300 29268 14858 29284
rect 12300 29204 13511 29268
rect 13575 29204 13601 29268
rect 13665 29204 13691 29268
rect 13755 29204 13781 29268
rect 13845 29204 13871 29268
rect 13935 29204 13961 29268
rect 14025 29204 14858 29268
rect 12300 29188 14858 29204
rect 12300 29124 13511 29188
rect 13575 29124 13601 29188
rect 13665 29124 13691 29188
rect 13755 29124 13781 29188
rect 13845 29124 13871 29188
rect 13935 29124 13961 29188
rect 14025 29124 14858 29188
rect 12300 29108 14858 29124
rect 12300 29044 13511 29108
rect 13575 29044 13601 29108
rect 13665 29044 13691 29108
rect 13755 29044 13781 29108
rect 13845 29044 13871 29108
rect 13935 29044 13961 29108
rect 14025 29044 14858 29108
rect 12300 29028 14858 29044
rect 12300 28964 13511 29028
rect 13575 28964 13601 29028
rect 13665 28964 13691 29028
rect 13755 28964 13781 29028
rect 13845 28964 13871 29028
rect 13935 28964 13961 29028
rect 14025 28964 14858 29028
rect 12300 28948 14858 28964
rect 12300 28884 13511 28948
rect 13575 28884 13601 28948
rect 13665 28884 13691 28948
rect 13755 28884 13781 28948
rect 13845 28884 13871 28948
rect 13935 28884 13961 28948
rect 14025 28884 14858 28948
rect 12300 28868 14858 28884
rect 12300 28804 13511 28868
rect 13575 28804 13601 28868
rect 13665 28804 13691 28868
rect 13755 28804 13781 28868
rect 13845 28804 13871 28868
rect 13935 28804 13961 28868
rect 14025 28804 14858 28868
rect 12300 28788 14858 28804
rect 12300 28724 13511 28788
rect 13575 28724 13601 28788
rect 13665 28724 13691 28788
rect 13755 28724 13781 28788
rect 13845 28724 13871 28788
rect 13935 28724 13961 28788
rect 14025 28724 14858 28788
rect 12300 28708 14858 28724
rect 12300 28644 13511 28708
rect 13575 28644 13601 28708
rect 13665 28644 13691 28708
rect 13755 28644 13781 28708
rect 13845 28644 13871 28708
rect 13935 28644 13961 28708
rect 14025 28644 14858 28708
rect 12300 28628 14858 28644
rect 12300 28564 13511 28628
rect 13575 28564 13601 28628
rect 13665 28564 13691 28628
rect 13755 28564 13781 28628
rect 13845 28564 13871 28628
rect 13935 28564 13961 28628
rect 14025 28564 14858 28628
rect 12300 28548 14858 28564
rect 12300 28484 13511 28548
rect 13575 28484 13601 28548
rect 13665 28484 13691 28548
rect 13755 28484 13781 28548
rect 13845 28484 13871 28548
rect 13935 28484 13961 28548
rect 14025 28484 14858 28548
rect 12300 28468 14858 28484
rect 12300 28404 13511 28468
rect 13575 28404 13601 28468
rect 13665 28404 13691 28468
rect 13755 28404 13781 28468
rect 13845 28404 13871 28468
rect 13935 28404 13961 28468
rect 14025 28404 14858 28468
rect 12300 28388 14858 28404
rect 12300 28324 13511 28388
rect 13575 28324 13601 28388
rect 13665 28324 13691 28388
rect 13755 28324 13781 28388
rect 13845 28324 13871 28388
rect 13935 28324 13961 28388
rect 14025 28324 14858 28388
rect 12300 28308 14858 28324
rect 12300 28244 13511 28308
rect 13575 28244 13601 28308
rect 13665 28244 13691 28308
rect 13755 28244 13781 28308
rect 13845 28244 13871 28308
rect 13935 28244 13961 28308
rect 14025 28244 14858 28308
rect 12300 28228 14858 28244
rect 12300 28164 13511 28228
rect 13575 28164 13601 28228
rect 13665 28164 13691 28228
rect 13755 28164 13781 28228
rect 13845 28164 13871 28228
rect 13935 28164 13961 28228
rect 14025 28164 14858 28228
rect 12300 28148 14858 28164
rect 12300 28084 13511 28148
rect 13575 28084 13601 28148
rect 13665 28084 13691 28148
rect 13755 28084 13781 28148
rect 13845 28084 13871 28148
rect 13935 28084 13961 28148
rect 14025 28084 14858 28148
rect 12300 28068 14858 28084
rect 12300 28004 13511 28068
rect 13575 28004 13601 28068
rect 13665 28004 13691 28068
rect 13755 28004 13781 28068
rect 13845 28004 13871 28068
rect 13935 28004 13961 28068
rect 14025 28004 14858 28068
rect 12300 27988 14858 28004
rect 12300 27924 13511 27988
rect 13575 27924 13601 27988
rect 13665 27924 13691 27988
rect 13755 27924 13781 27988
rect 13845 27924 13871 27988
rect 13935 27924 13961 27988
rect 14025 27924 14858 27988
rect 12300 27908 14858 27924
rect 12300 27844 13511 27908
rect 13575 27844 13601 27908
rect 13665 27844 13691 27908
rect 13755 27844 13781 27908
rect 13845 27844 13871 27908
rect 13935 27844 13961 27908
rect 14025 27844 14858 27908
rect 12300 27828 14858 27844
rect 12300 27764 13511 27828
rect 13575 27764 13601 27828
rect 13665 27764 13691 27828
rect 13755 27764 13781 27828
rect 13845 27764 13871 27828
rect 13935 27764 13961 27828
rect 14025 27764 14858 27828
rect 12300 27748 14858 27764
rect 12300 27684 13511 27748
rect 13575 27684 13601 27748
rect 13665 27684 13691 27748
rect 13755 27684 13781 27748
rect 13845 27684 13871 27748
rect 13935 27684 13961 27748
rect 14025 27684 14858 27748
rect 12300 27668 14858 27684
rect 12300 27604 13511 27668
rect 13575 27604 13601 27668
rect 13665 27604 13691 27668
rect 13755 27604 13781 27668
rect 13845 27604 13871 27668
rect 13935 27604 13961 27668
rect 14025 27604 14858 27668
rect 12300 27588 14858 27604
rect 12300 27524 13511 27588
rect 13575 27524 13601 27588
rect 13665 27524 13691 27588
rect 13755 27524 13781 27588
rect 13845 27524 13871 27588
rect 13935 27524 13961 27588
rect 14025 27524 14858 27588
rect 12300 27508 14858 27524
rect 12300 27444 13511 27508
rect 13575 27444 13601 27508
rect 13665 27444 13691 27508
rect 13755 27444 13781 27508
rect 13845 27444 13871 27508
rect 13935 27444 13961 27508
rect 14025 27444 14858 27508
rect 12300 27428 14858 27444
rect 12300 27364 13511 27428
rect 13575 27364 13601 27428
rect 13665 27364 13691 27428
rect 13755 27364 13781 27428
rect 13845 27364 13871 27428
rect 13935 27364 13961 27428
rect 14025 27364 14858 27428
rect 12300 27348 14858 27364
rect 12300 27284 13511 27348
rect 13575 27284 13601 27348
rect 13665 27284 13691 27348
rect 13755 27284 13781 27348
rect 13845 27284 13871 27348
rect 13935 27284 13961 27348
rect 14025 27284 14858 27348
rect 12300 27268 14858 27284
rect 12300 27204 13511 27268
rect 13575 27204 13601 27268
rect 13665 27204 13691 27268
rect 13755 27204 13781 27268
rect 13845 27204 13871 27268
rect 13935 27204 13961 27268
rect 14025 27204 14858 27268
rect 12300 27188 14858 27204
rect 12300 27124 13511 27188
rect 13575 27124 13601 27188
rect 13665 27124 13691 27188
rect 13755 27124 13781 27188
rect 13845 27124 13871 27188
rect 13935 27124 13961 27188
rect 14025 27124 14858 27188
rect 12300 27108 14858 27124
rect 12300 27044 13511 27108
rect 13575 27044 13601 27108
rect 13665 27044 13691 27108
rect 13755 27044 13781 27108
rect 13845 27044 13871 27108
rect 13935 27044 13961 27108
rect 14025 27044 14858 27108
rect 12300 27028 14858 27044
rect 12300 26964 13511 27028
rect 13575 26964 13601 27028
rect 13665 26964 13691 27028
rect 13755 26964 13781 27028
rect 13845 26964 13871 27028
rect 13935 26964 13961 27028
rect 14025 26964 14858 27028
rect 12300 26948 14858 26964
rect 12300 26884 13511 26948
rect 13575 26884 13601 26948
rect 13665 26884 13691 26948
rect 13755 26884 13781 26948
rect 13845 26884 13871 26948
rect 13935 26884 13961 26948
rect 14025 26884 14858 26948
rect 12300 26868 14858 26884
rect 12300 26804 13511 26868
rect 13575 26804 13601 26868
rect 13665 26804 13691 26868
rect 13755 26804 13781 26868
rect 13845 26804 13871 26868
rect 13935 26804 13961 26868
rect 14025 26804 14858 26868
rect 12300 26788 14858 26804
rect 12300 26724 13511 26788
rect 13575 26724 13601 26788
rect 13665 26724 13691 26788
rect 13755 26724 13781 26788
rect 13845 26724 13871 26788
rect 13935 26724 13961 26788
rect 14025 26724 14858 26788
rect 12300 26708 14858 26724
rect 12300 26644 13511 26708
rect 13575 26644 13601 26708
rect 13665 26644 13691 26708
rect 13755 26644 13781 26708
rect 13845 26644 13871 26708
rect 13935 26644 13961 26708
rect 14025 26644 14858 26708
rect 12300 26628 14858 26644
rect 12300 26564 13511 26628
rect 13575 26564 13601 26628
rect 13665 26564 13691 26628
rect 13755 26564 13781 26628
rect 13845 26564 13871 26628
rect 13935 26564 13961 26628
rect 14025 26564 14858 26628
rect 12300 26548 14858 26564
rect 12300 26484 13511 26548
rect 13575 26484 13601 26548
rect 13665 26484 13691 26548
rect 13755 26484 13781 26548
rect 13845 26484 13871 26548
rect 13935 26484 13961 26548
rect 14025 26484 14858 26548
rect 12300 26468 14858 26484
rect 12300 26404 13511 26468
rect 13575 26404 13601 26468
rect 13665 26404 13691 26468
rect 13755 26404 13781 26468
rect 13845 26404 13871 26468
rect 13935 26404 13961 26468
rect 14025 26404 14858 26468
rect 12300 26388 14858 26404
rect 12300 26324 13511 26388
rect 13575 26324 13601 26388
rect 13665 26324 13691 26388
rect 13755 26324 13781 26388
rect 13845 26324 13871 26388
rect 13935 26324 13961 26388
rect 14025 26324 14858 26388
rect 12300 26308 14858 26324
rect 12300 26244 13511 26308
rect 13575 26244 13601 26308
rect 13665 26244 13691 26308
rect 13755 26244 13781 26308
rect 13845 26244 13871 26308
rect 13935 26244 13961 26308
rect 14025 26244 14858 26308
rect 12300 26228 14858 26244
rect 12300 26164 13511 26228
rect 13575 26164 13601 26228
rect 13665 26164 13691 26228
rect 13755 26164 13781 26228
rect 13845 26164 13871 26228
rect 13935 26164 13961 26228
rect 14025 26164 14858 26228
rect 12300 26148 14858 26164
rect 12300 26084 13511 26148
rect 13575 26084 13601 26148
rect 13665 26084 13691 26148
rect 13755 26084 13781 26148
rect 13845 26084 13871 26148
rect 13935 26084 13961 26148
rect 14025 26084 14858 26148
rect 12300 26068 14858 26084
rect 12300 26004 13511 26068
rect 13575 26004 13601 26068
rect 13665 26004 13691 26068
rect 13755 26004 13781 26068
rect 13845 26004 13871 26068
rect 13935 26004 13961 26068
rect 14025 26004 14858 26068
rect 12300 25988 14858 26004
rect 12300 25924 13511 25988
rect 13575 25924 13601 25988
rect 13665 25924 13691 25988
rect 13755 25924 13781 25988
rect 13845 25924 13871 25988
rect 13935 25924 13961 25988
rect 14025 25924 14858 25988
rect 12300 25908 14858 25924
rect 12300 25844 13511 25908
rect 13575 25844 13601 25908
rect 13665 25844 13691 25908
rect 13755 25844 13781 25908
rect 13845 25844 13871 25908
rect 13935 25844 13961 25908
rect 14025 25844 14858 25908
rect 12300 25828 14858 25844
rect 12300 25764 13511 25828
rect 13575 25764 13601 25828
rect 13665 25764 13691 25828
rect 13755 25764 13781 25828
rect 13845 25764 13871 25828
rect 13935 25764 13961 25828
rect 14025 25764 14858 25828
rect 12300 25748 14858 25764
rect 12300 25684 13511 25748
rect 13575 25684 13601 25748
rect 13665 25684 13691 25748
rect 13755 25684 13781 25748
rect 13845 25684 13871 25748
rect 13935 25684 13961 25748
rect 14025 25684 14858 25748
rect 12300 25668 14858 25684
rect 12300 25604 13511 25668
rect 13575 25604 13601 25668
rect 13665 25604 13691 25668
rect 13755 25604 13781 25668
rect 13845 25604 13871 25668
rect 13935 25604 13961 25668
rect 14025 25604 14858 25668
rect 12300 25588 14858 25604
rect 12300 25524 13511 25588
rect 13575 25524 13601 25588
rect 13665 25524 13691 25588
rect 13755 25524 13781 25588
rect 13845 25524 13871 25588
rect 13935 25524 13961 25588
rect 14025 25524 14858 25588
rect 12300 25508 14858 25524
rect 12300 25444 13511 25508
rect 13575 25444 13601 25508
rect 13665 25444 13691 25508
rect 13755 25444 13781 25508
rect 13845 25444 13871 25508
rect 13935 25444 13961 25508
rect 14025 25444 14858 25508
rect 12300 25428 14858 25444
rect 12300 25364 13511 25428
rect 13575 25364 13601 25428
rect 13665 25364 13691 25428
rect 13755 25364 13781 25428
rect 13845 25364 13871 25428
rect 13935 25364 13961 25428
rect 14025 25364 14858 25428
rect 12300 25348 14858 25364
rect 12300 25284 13511 25348
rect 13575 25284 13601 25348
rect 13665 25284 13691 25348
rect 13755 25284 13781 25348
rect 13845 25284 13871 25348
rect 13935 25284 13961 25348
rect 14025 25284 14858 25348
rect 12300 25268 14858 25284
rect 12300 25204 13511 25268
rect 13575 25204 13601 25268
rect 13665 25204 13691 25268
rect 13755 25204 13781 25268
rect 13845 25204 13871 25268
rect 13935 25204 13961 25268
rect 14025 25204 14858 25268
rect 12300 25188 14858 25204
rect 12300 25124 13511 25188
rect 13575 25124 13601 25188
rect 13665 25124 13691 25188
rect 13755 25124 13781 25188
rect 13845 25124 13871 25188
rect 13935 25124 13961 25188
rect 14025 25124 14858 25188
rect 12300 25108 14858 25124
rect 12300 25044 13511 25108
rect 13575 25044 13601 25108
rect 13665 25044 13691 25108
rect 13755 25044 13781 25108
rect 13845 25044 13871 25108
rect 13935 25044 13961 25108
rect 14025 25044 14858 25108
rect 12300 25028 14858 25044
rect 12300 24964 13511 25028
rect 13575 24964 13601 25028
rect 13665 24964 13691 25028
rect 13755 24964 13781 25028
rect 13845 24964 13871 25028
rect 13935 24964 13961 25028
rect 14025 24964 14858 25028
rect 12300 24948 14858 24964
rect 12300 24884 13511 24948
rect 13575 24884 13601 24948
rect 13665 24884 13691 24948
rect 13755 24884 13781 24948
rect 13845 24884 13871 24948
rect 13935 24884 13961 24948
rect 14025 24884 14858 24948
rect 12300 24868 14858 24884
rect 12300 24804 13511 24868
rect 13575 24804 13601 24868
rect 13665 24804 13691 24868
rect 13755 24804 13781 24868
rect 13845 24804 13871 24868
rect 13935 24804 13961 24868
rect 14025 24804 14858 24868
rect 12300 24788 14858 24804
rect 12300 24724 13511 24788
rect 13575 24724 13601 24788
rect 13665 24724 13691 24788
rect 13755 24724 13781 24788
rect 13845 24724 13871 24788
rect 13935 24724 13961 24788
rect 14025 24724 14858 24788
rect 12300 24708 14858 24724
rect 12300 24644 13511 24708
rect 13575 24644 13601 24708
rect 13665 24644 13691 24708
rect 13755 24644 13781 24708
rect 13845 24644 13871 24708
rect 13935 24644 13961 24708
rect 14025 24644 14858 24708
rect 12300 24628 14858 24644
rect 12300 24564 13511 24628
rect 13575 24564 13601 24628
rect 13665 24564 13691 24628
rect 13755 24564 13781 24628
rect 13845 24564 13871 24628
rect 13935 24564 13961 24628
rect 14025 24564 14858 24628
rect 12300 24548 14858 24564
rect 12300 24484 13511 24548
rect 13575 24484 13601 24548
rect 13665 24484 13691 24548
rect 13755 24484 13781 24548
rect 13845 24484 13871 24548
rect 13935 24484 13961 24548
rect 14025 24484 14858 24548
rect 12300 24468 14858 24484
rect 12300 24404 13511 24468
rect 13575 24404 13601 24468
rect 13665 24404 13691 24468
rect 13755 24404 13781 24468
rect 13845 24404 13871 24468
rect 13935 24404 13961 24468
rect 14025 24404 14858 24468
rect 12300 24388 14858 24404
rect 12300 24324 13511 24388
rect 13575 24324 13601 24388
rect 13665 24324 13691 24388
rect 13755 24324 13781 24388
rect 13845 24324 13871 24388
rect 13935 24324 13961 24388
rect 14025 24324 14858 24388
rect 12300 24308 14858 24324
rect 12300 24244 13511 24308
rect 13575 24244 13601 24308
rect 13665 24244 13691 24308
rect 13755 24244 13781 24308
rect 13845 24244 13871 24308
rect 13935 24244 13961 24308
rect 14025 24244 14858 24308
rect 12300 24228 14858 24244
rect 12300 24164 13511 24228
rect 13575 24164 13601 24228
rect 13665 24164 13691 24228
rect 13755 24164 13781 24228
rect 13845 24164 13871 24228
rect 13935 24164 13961 24228
rect 14025 24164 14858 24228
rect 12300 24148 14858 24164
rect 12300 24084 13511 24148
rect 13575 24084 13601 24148
rect 13665 24084 13691 24148
rect 13755 24084 13781 24148
rect 13845 24084 13871 24148
rect 13935 24084 13961 24148
rect 14025 24084 14858 24148
rect 12300 24068 14858 24084
rect 12300 24004 13511 24068
rect 13575 24004 13601 24068
rect 13665 24004 13691 24068
rect 13755 24004 13781 24068
rect 13845 24004 13871 24068
rect 13935 24004 13961 24068
rect 14025 24004 14858 24068
rect 12300 23988 14858 24004
rect 12300 23924 13511 23988
rect 13575 23924 13601 23988
rect 13665 23924 13691 23988
rect 13755 23924 13781 23988
rect 13845 23924 13871 23988
rect 13935 23924 13961 23988
rect 14025 23924 14858 23988
rect 12300 23908 14858 23924
rect 12300 23844 13511 23908
rect 13575 23844 13601 23908
rect 13665 23844 13691 23908
rect 13755 23844 13781 23908
rect 13845 23844 13871 23908
rect 13935 23844 13961 23908
rect 14025 23844 14858 23908
rect 12300 23828 14858 23844
rect 12300 23764 13511 23828
rect 13575 23764 13601 23828
rect 13665 23764 13691 23828
rect 13755 23764 13781 23828
rect 13845 23764 13871 23828
rect 13935 23764 13961 23828
rect 14025 23764 14858 23828
rect 12300 23748 14858 23764
rect 12300 23684 13511 23748
rect 13575 23684 13601 23748
rect 13665 23684 13691 23748
rect 13755 23684 13781 23748
rect 13845 23684 13871 23748
rect 13935 23684 13961 23748
rect 14025 23684 14858 23748
rect 12300 23668 14858 23684
rect 12300 23604 13511 23668
rect 13575 23604 13601 23668
rect 13665 23604 13691 23668
rect 13755 23604 13781 23668
rect 13845 23604 13871 23668
rect 13935 23604 13961 23668
rect 14025 23604 14858 23668
rect 12300 23588 14858 23604
rect 12300 23524 13511 23588
rect 13575 23524 13601 23588
rect 13665 23524 13691 23588
rect 13755 23524 13781 23588
rect 13845 23524 13871 23588
rect 13935 23524 13961 23588
rect 14025 23524 14858 23588
rect 12300 23508 14858 23524
rect 12300 23444 13511 23508
rect 13575 23444 13601 23508
rect 13665 23444 13691 23508
rect 13755 23444 13781 23508
rect 13845 23444 13871 23508
rect 13935 23444 13961 23508
rect 14025 23444 14858 23508
rect 12300 23428 14858 23444
rect 12300 23364 13511 23428
rect 13575 23364 13601 23428
rect 13665 23364 13691 23428
rect 13755 23364 13781 23428
rect 13845 23364 13871 23428
rect 13935 23364 13961 23428
rect 14025 23364 14858 23428
rect 12300 23348 14858 23364
rect 12300 23284 13511 23348
rect 13575 23284 13601 23348
rect 13665 23284 13691 23348
rect 13755 23284 13781 23348
rect 13845 23284 13871 23348
rect 13935 23284 13961 23348
rect 14025 23284 14858 23348
rect 12300 23267 14858 23284
rect 12300 23203 13511 23267
rect 13575 23203 13601 23267
rect 13665 23203 13691 23267
rect 13755 23203 13781 23267
rect 13845 23203 13871 23267
rect 13935 23203 13961 23267
rect 14025 23203 14858 23267
rect 12300 23186 14858 23203
rect 12300 23122 13511 23186
rect 13575 23122 13601 23186
rect 13665 23122 13691 23186
rect 13755 23122 13781 23186
rect 13845 23122 13871 23186
rect 13935 23122 13961 23186
rect 14025 23122 14858 23186
rect 12300 23105 14858 23122
rect 12300 23041 13511 23105
rect 13575 23041 13601 23105
rect 13665 23041 13691 23105
rect 13755 23041 13781 23105
rect 13845 23041 13871 23105
rect 13935 23041 13961 23105
rect 14025 23041 14858 23105
rect 12300 23024 14858 23041
rect 12300 22960 13511 23024
rect 13575 22960 13601 23024
rect 13665 22960 13691 23024
rect 13755 22960 13781 23024
rect 13845 22960 13871 23024
rect 13935 22960 13961 23024
rect 14025 22960 14858 23024
rect 12300 22943 14858 22960
rect 12300 22879 13511 22943
rect 13575 22879 13601 22943
rect 13665 22879 13691 22943
rect 13755 22879 13781 22943
rect 13845 22879 13871 22943
rect 13935 22879 13961 22943
rect 14025 22879 14858 22943
rect 12300 22862 14858 22879
rect 12300 22798 13511 22862
rect 13575 22798 13601 22862
rect 13665 22798 13691 22862
rect 13755 22798 13781 22862
rect 13845 22798 13871 22862
rect 13935 22798 13961 22862
rect 14025 22798 14858 22862
rect 12300 22781 14858 22798
rect 12300 22717 13511 22781
rect 13575 22717 13601 22781
rect 13665 22717 13691 22781
rect 13755 22717 13781 22781
rect 13845 22717 13871 22781
rect 13935 22717 13961 22781
rect 14025 22717 14858 22781
rect 12300 22700 14858 22717
rect 12300 22636 13511 22700
rect 13575 22636 13601 22700
rect 13665 22636 13691 22700
rect 13755 22636 13781 22700
rect 13845 22636 13871 22700
rect 13935 22636 13961 22700
rect 14025 22636 14858 22700
rect 12300 22619 14858 22636
rect 12300 22555 13511 22619
rect 13575 22555 13601 22619
rect 13665 22555 13691 22619
rect 13755 22555 13781 22619
rect 13845 22555 13871 22619
rect 13935 22555 13961 22619
rect 14025 22555 14858 22619
rect 12300 22538 14858 22555
rect 12300 22474 13511 22538
rect 13575 22474 13601 22538
rect 13665 22474 13691 22538
rect 13755 22474 13781 22538
rect 13845 22474 13871 22538
rect 13935 22474 13961 22538
rect 14025 22474 14858 22538
rect 12300 22457 14858 22474
rect 12300 22393 13511 22457
rect 13575 22393 13601 22457
rect 13665 22393 13691 22457
rect 13755 22393 13781 22457
rect 13845 22393 13871 22457
rect 13935 22393 13961 22457
rect 14025 22393 14858 22457
rect 12300 22376 14858 22393
rect 12300 22312 13511 22376
rect 13575 22312 13601 22376
rect 13665 22312 13691 22376
rect 13755 22312 13781 22376
rect 13845 22312 13871 22376
rect 13935 22312 13961 22376
rect 14025 22312 14858 22376
rect 12300 22295 14858 22312
rect 12300 22231 13511 22295
rect 13575 22231 13601 22295
rect 13665 22231 13691 22295
rect 13755 22231 13781 22295
rect 13845 22231 13871 22295
rect 13935 22231 13961 22295
rect 14025 22231 14858 22295
rect 12300 22214 14858 22231
rect 12300 22150 13511 22214
rect 13575 22150 13601 22214
rect 13665 22150 13691 22214
rect 13755 22150 13781 22214
rect 13845 22150 13871 22214
rect 13935 22150 13961 22214
rect 14025 22150 14858 22214
rect 12300 22133 14858 22150
rect 12300 22069 13511 22133
rect 13575 22069 13601 22133
rect 13665 22069 13691 22133
rect 13755 22069 13781 22133
rect 13845 22069 13871 22133
rect 13935 22069 13961 22133
rect 14025 22069 14858 22133
rect 12300 22052 14858 22069
rect 12300 21988 13511 22052
rect 13575 21988 13601 22052
rect 13665 21988 13691 22052
rect 13755 21988 13781 22052
rect 13845 21988 13871 22052
rect 13935 21988 13961 22052
rect 14025 21988 14858 22052
rect 12300 21971 14858 21988
rect 12300 21907 13511 21971
rect 13575 21907 13601 21971
rect 13665 21907 13691 21971
rect 13755 21907 13781 21971
rect 13845 21907 13871 21971
rect 13935 21907 13961 21971
rect 14025 21907 14858 21971
rect 12300 21890 14858 21907
rect 12300 21826 13511 21890
rect 13575 21826 13601 21890
rect 13665 21826 13691 21890
rect 13755 21826 13781 21890
rect 13845 21826 13871 21890
rect 13935 21826 13961 21890
rect 14025 21826 14858 21890
rect 12300 21809 14858 21826
rect 12300 21745 13511 21809
rect 13575 21745 13601 21809
rect 13665 21745 13691 21809
rect 13755 21745 13781 21809
rect 13845 21745 13871 21809
rect 13935 21745 13961 21809
rect 14025 21745 14858 21809
rect 12300 21728 14858 21745
rect 12300 21664 13511 21728
rect 13575 21664 13601 21728
rect 13665 21664 13691 21728
rect 13755 21664 13781 21728
rect 13845 21664 13871 21728
rect 13935 21664 13961 21728
rect 14025 21664 14858 21728
rect 12300 21647 14858 21664
rect 12300 21583 13511 21647
rect 13575 21583 13601 21647
rect 13665 21583 13691 21647
rect 13755 21583 13781 21647
rect 13845 21583 13871 21647
rect 13935 21583 13961 21647
rect 14025 21583 14858 21647
rect 12300 21566 14858 21583
rect 12300 21502 13511 21566
rect 13575 21502 13601 21566
rect 13665 21502 13691 21566
rect 13755 21502 13781 21566
rect 13845 21502 13871 21566
rect 13935 21502 13961 21566
rect 14025 21502 14858 21566
rect 12300 21485 14858 21502
rect 12300 21421 13511 21485
rect 13575 21421 13601 21485
rect 13665 21421 13691 21485
rect 13755 21421 13781 21485
rect 13845 21421 13871 21485
rect 13935 21421 13961 21485
rect 14025 21421 14858 21485
rect 12300 21404 14858 21421
rect 12300 21340 13511 21404
rect 13575 21340 13601 21404
rect 13665 21340 13691 21404
rect 13755 21340 13781 21404
rect 13845 21340 13871 21404
rect 13935 21340 13961 21404
rect 14025 21340 14858 21404
rect 12300 21323 14858 21340
rect 12300 21259 13511 21323
rect 13575 21259 13601 21323
rect 13665 21259 13691 21323
rect 13755 21259 13781 21323
rect 13845 21259 13871 21323
rect 13935 21259 13961 21323
rect 14025 21259 14858 21323
rect 12300 21242 14858 21259
rect 12300 21178 13511 21242
rect 13575 21178 13601 21242
rect 13665 21178 13691 21242
rect 13755 21178 13781 21242
rect 13845 21178 13871 21242
rect 13935 21178 13961 21242
rect 14025 21178 14858 21242
rect 12300 21161 14858 21178
rect 12300 21097 13511 21161
rect 13575 21097 13601 21161
rect 13665 21097 13691 21161
rect 13755 21097 13781 21161
rect 13845 21097 13871 21161
rect 13935 21097 13961 21161
rect 14025 21097 14858 21161
rect 12300 21080 14858 21097
rect 12300 21016 13511 21080
rect 13575 21016 13601 21080
rect 13665 21016 13691 21080
rect 13755 21016 13781 21080
rect 13845 21016 13871 21080
rect 13935 21016 13961 21080
rect 14025 21016 14858 21080
rect 12300 20999 14858 21016
rect 12300 20938 13511 20999
rect 12300 20874 13412 20938
rect 13476 20935 13511 20938
rect 13575 20935 13601 20999
rect 13665 20935 13691 20999
rect 13755 20935 13781 20999
rect 13845 20935 13871 20999
rect 13935 20935 13961 20999
rect 14025 20935 14858 20999
rect 13476 20918 14858 20935
rect 13476 20874 13511 20918
rect 12300 20854 13511 20874
rect 13575 20854 13601 20918
rect 13665 20854 13691 20918
rect 13755 20854 13781 20918
rect 13845 20854 13871 20918
rect 13935 20854 13961 20918
rect 14025 20854 14858 20918
rect 12300 20824 14858 20854
rect 12300 20760 13272 20824
rect 13336 20760 13362 20824
rect 13426 20760 13452 20824
rect 13516 20760 13542 20824
rect 13606 20760 13631 20824
rect 13695 20822 14858 20824
rect 13695 20760 13740 20822
rect 12300 20758 13740 20760
rect 13804 20815 14858 20822
rect 13804 20758 13842 20815
rect 12300 20751 13842 20758
rect 13906 20751 14858 20815
rect 12300 20711 14858 20751
rect 12300 20708 13740 20711
rect 12300 20644 13272 20708
rect 13336 20644 13362 20708
rect 13426 20644 13452 20708
rect 13516 20644 13542 20708
rect 13606 20644 13631 20708
rect 13695 20647 13740 20708
rect 13804 20647 14858 20711
rect 13695 20644 14858 20647
rect 12300 20630 14858 20644
rect 12300 20566 13131 20630
rect 13195 20592 14858 20630
rect 13195 20566 13272 20592
rect 12300 20528 13272 20566
rect 13336 20528 13362 20592
rect 13426 20528 13452 20592
rect 13516 20528 13542 20592
rect 13606 20528 13631 20592
rect 13695 20528 14858 20592
rect 12300 20504 14858 20528
rect 12300 20440 12952 20504
rect 13016 20440 13042 20504
rect 13106 20440 13132 20504
rect 13196 20440 13222 20504
rect 13286 20440 13311 20504
rect 13375 20468 14858 20504
rect 13375 20440 13419 20468
rect 12300 20404 13419 20440
rect 13483 20404 14858 20468
rect 12300 20388 14858 20404
rect 12300 20324 12952 20388
rect 13016 20324 13042 20388
rect 13106 20324 13132 20388
rect 13196 20324 13222 20388
rect 13286 20324 13311 20388
rect 13375 20324 14858 20388
rect 12300 20305 14858 20324
rect 2046 20208 2700 20241
rect 99 20180 2700 20208
rect 99 20140 1947 20180
rect 99 20076 1843 20140
rect 1907 20116 1947 20140
rect 2011 20116 2036 20180
rect 2100 20116 2126 20180
rect 2190 20116 2216 20180
rect 2280 20116 2306 20180
rect 2370 20116 2700 20180
rect 1907 20076 2700 20116
rect 99 20064 2700 20076
rect 99 20000 1947 20064
rect 2011 20000 2036 20064
rect 2100 20000 2126 20064
rect 2190 20000 2216 20064
rect 2280 20000 2306 20064
rect 2370 20000 2700 20064
rect 99 19948 2700 20000
rect 99 19884 1947 19948
rect 2011 19884 2036 19948
rect 2100 19884 2126 19948
rect 2190 19884 2216 19948
rect 2280 19884 2306 19948
rect 2370 19884 2700 19948
rect 99 19799 2700 19884
rect 99 19735 2184 19799
rect 2248 19735 2700 19799
rect 99 16575 2700 19735
tri 99 14722 1952 16575 ne
rect 1952 16471 2700 16575
tri 2700 16471 6508 20279 sw
tri 12110 20069 12300 20259 se
rect 12300 20241 12806 20305
rect 12870 20272 14858 20305
rect 12870 20241 12952 20272
rect 12300 20208 12952 20241
rect 13016 20208 13042 20272
rect 13106 20208 13132 20272
rect 13196 20208 13222 20272
rect 13286 20208 13311 20272
rect 13375 20208 14858 20272
rect 12300 20180 14858 20208
rect 12300 20116 12628 20180
rect 12692 20116 12718 20180
rect 12782 20116 12808 20180
rect 12872 20116 12898 20180
rect 12962 20116 12987 20180
rect 13051 20140 14858 20180
rect 13051 20116 13091 20140
rect 12300 20076 13091 20116
rect 13155 20076 14858 20140
rect 12300 20069 14858 20076
tri 12027 19986 12110 20069 se
rect 12110 20005 12141 20069
rect 12205 20005 12257 20069
rect 12321 20005 12372 20069
rect 12436 20005 12487 20069
rect 12551 20064 14858 20069
rect 12551 20005 12628 20064
rect 12110 20000 12628 20005
rect 12692 20000 12718 20064
rect 12782 20000 12808 20064
rect 12872 20000 12898 20064
rect 12962 20000 12987 20064
rect 13051 20000 14858 20064
rect 12110 19986 14858 20000
tri 11885 19844 12027 19986 se
rect 12027 19954 14858 19986
rect 12027 19890 12037 19954
rect 12101 19949 14858 19954
rect 12101 19890 12141 19949
rect 12027 19885 12141 19890
rect 12205 19885 12257 19949
rect 12321 19885 12372 19949
rect 12436 19885 12487 19949
rect 12551 19948 14858 19949
rect 12551 19885 12628 19948
rect 12027 19884 12628 19885
rect 12692 19884 12718 19948
rect 12782 19884 12808 19948
rect 12872 19884 12898 19948
rect 12962 19884 12987 19948
rect 13051 19884 14858 19948
rect 12027 19844 14858 19884
tri 11753 19712 11885 19844 se
rect 11885 19843 14858 19844
rect 11885 19779 11894 19843
rect 11958 19779 11978 19843
rect 12042 19779 12062 19843
rect 12126 19779 12146 19843
rect 12210 19779 12230 19843
rect 12294 19779 12314 19843
rect 12378 19779 12398 19843
rect 12462 19779 12482 19843
rect 12546 19779 12566 19843
rect 12630 19779 12650 19843
rect 12714 19799 14858 19843
rect 12714 19779 12750 19799
rect 11885 19735 12750 19779
rect 12814 19735 14858 19799
rect 11885 19727 14858 19735
rect 11885 19712 11894 19727
tri 11271 19230 11753 19712 se
rect 11753 19706 11894 19712
rect 11753 19642 11790 19706
rect 11854 19663 11894 19706
rect 11958 19663 11978 19727
rect 12042 19663 12062 19727
rect 12126 19663 12146 19727
rect 12210 19663 12230 19727
rect 12294 19663 12314 19727
rect 12378 19663 12398 19727
rect 12462 19663 12482 19727
rect 12546 19663 12566 19727
rect 12630 19663 12650 19727
rect 12714 19663 14858 19727
rect 11854 19642 14858 19663
rect 11753 19613 14858 19642
rect 11753 19549 11790 19613
rect 11854 19611 14858 19613
rect 11854 19549 11894 19611
rect 11753 19547 11894 19549
rect 11958 19547 11978 19611
rect 12042 19547 12062 19611
rect 12126 19547 12146 19611
rect 12210 19547 12230 19611
rect 12294 19547 12314 19611
rect 12378 19547 12398 19611
rect 12462 19547 12482 19611
rect 12546 19547 12566 19611
rect 12630 19547 12650 19611
rect 12714 19547 14858 19611
rect 11753 19230 14858 19547
tri 8512 16471 11271 19230 se
rect 11271 16628 14858 19230
rect 11271 16471 12952 16628
rect 1952 14722 12952 16471
tri 12952 14722 14858 16628 nw
tri 1952 11722 4952 14722 ne
rect 858 9741 2098 9774
rect 858 9285 890 9741
rect 2066 9285 2098 9741
rect 858 3646 2098 9285
rect 858 3022 887 3646
rect 2071 3022 2098 3646
rect 858 2982 2098 3022
rect 4952 1 9952 14722
tri 9952 11722 12952 14722 nw
rect 12858 9741 14098 9774
rect 12858 9285 12890 9741
rect 14066 9285 14098 9741
rect 12858 3646 14098 9285
rect 12858 3022 12887 3646
rect 14071 3022 14098 3646
rect 12858 2982 14098 3022
<< via3 >>
rect 2267 34553 2331 34617
rect 2350 34553 2414 34617
rect 2434 34553 2498 34617
rect 2518 34553 2582 34617
rect 2602 34553 2666 34617
rect 12332 34553 12396 34617
rect 12416 34553 12480 34617
rect 12500 34553 12564 34617
rect 12584 34553 12648 34617
rect 12668 34553 12732 34617
rect 2267 34459 2331 34523
rect 2350 34459 2414 34523
rect 2434 34459 2498 34523
rect 2518 34459 2582 34523
rect 2602 34459 2666 34523
rect 12332 34459 12396 34523
rect 12416 34459 12480 34523
rect 12500 34459 12564 34523
rect 12584 34459 12648 34523
rect 12668 34459 12732 34523
rect 2139 34376 2203 34440
rect 2267 34365 2331 34429
rect 2350 34365 2414 34429
rect 2434 34365 2498 34429
rect 2518 34365 2582 34429
rect 2602 34365 2666 34429
rect 12332 34365 12396 34429
rect 12416 34365 12480 34429
rect 12500 34365 12564 34429
rect 12584 34365 12648 34429
rect 12668 34365 12732 34429
rect 12795 34376 12859 34440
rect 1995 34251 2059 34315
rect 2075 34251 2139 34315
rect 2155 34251 2219 34315
rect 2267 34271 2331 34335
rect 2350 34271 2414 34335
rect 2434 34271 2498 34335
rect 2518 34271 2582 34335
rect 2602 34271 2666 34335
rect 12332 34271 12396 34335
rect 12416 34271 12480 34335
rect 12500 34271 12564 34335
rect 12584 34271 12648 34335
rect 12668 34271 12732 34335
rect 12779 34251 12843 34315
rect 12859 34251 12923 34315
rect 12939 34251 13003 34315
rect 1881 34118 1945 34182
rect 1995 34155 2059 34219
rect 2075 34155 2139 34219
rect 2155 34155 2219 34219
rect 2267 34177 2331 34241
rect 2350 34177 2414 34241
rect 2434 34177 2498 34241
rect 2518 34177 2582 34241
rect 2602 34177 2666 34241
rect 12332 34177 12396 34241
rect 12416 34177 12480 34241
rect 12500 34177 12564 34241
rect 12584 34177 12648 34241
rect 12668 34177 12732 34241
rect 12779 34155 12843 34219
rect 12859 34155 12923 34219
rect 12939 34155 13003 34219
rect 2267 34083 2331 34147
rect 2350 34083 2414 34147
rect 2434 34083 2498 34147
rect 2518 34083 2582 34147
rect 2602 34083 2666 34147
rect 12332 34083 12396 34147
rect 12416 34083 12480 34147
rect 12500 34083 12564 34147
rect 12584 34083 12648 34147
rect 12668 34083 12732 34147
rect 13053 34118 13117 34182
rect 1739 34013 1803 34077
rect 1828 34013 1892 34077
rect 1918 34013 1982 34077
rect 2008 34013 2072 34077
rect 2098 34013 2162 34077
rect 12836 34013 12900 34077
rect 12926 34013 12990 34077
rect 13016 34013 13080 34077
rect 13106 34013 13170 34077
rect 13195 34013 13259 34077
rect 1739 33897 1803 33961
rect 1828 33897 1892 33961
rect 1918 33897 1982 33961
rect 2008 33897 2072 33961
rect 2098 33897 2162 33961
rect 2238 33944 2302 34008
rect 12696 33944 12760 34008
rect 12836 33897 12900 33961
rect 12926 33897 12990 33961
rect 13016 33897 13080 33961
rect 13106 33897 13170 33961
rect 13195 33897 13259 33961
rect 1635 33821 1699 33885
rect 1739 33781 1803 33845
rect 1828 33781 1892 33845
rect 1918 33781 1982 33845
rect 2008 33781 2072 33845
rect 2098 33781 2162 33845
rect 1415 33689 1479 33753
rect 1504 33689 1568 33753
rect 1594 33689 1658 33753
rect 1684 33689 1748 33753
rect 1774 33689 1838 33753
rect 1920 33656 1984 33720
rect 1415 33573 1479 33637
rect 1504 33573 1568 33637
rect 1594 33573 1658 33637
rect 1684 33573 1748 33637
rect 1774 33573 1838 33637
rect 1307 33493 1371 33557
rect 1415 33457 1479 33521
rect 1504 33457 1568 33521
rect 1594 33457 1658 33521
rect 1684 33457 1748 33521
rect 1774 33457 1838 33521
rect 12836 33781 12900 33845
rect 12926 33781 12990 33845
rect 13016 33781 13080 33845
rect 13106 33781 13170 33845
rect 13195 33781 13259 33845
rect 13299 33821 13363 33885
rect 13014 33656 13078 33720
rect 13160 33689 13224 33753
rect 13250 33689 13314 33753
rect 13340 33689 13404 33753
rect 13430 33689 13494 33753
rect 13519 33689 13583 33753
rect 13160 33573 13224 33637
rect 13250 33573 13314 33637
rect 13340 33573 13404 33637
rect 13430 33573 13494 33637
rect 13519 33573 13583 33637
rect 13160 33457 13224 33521
rect 13250 33457 13314 33521
rect 13340 33457 13404 33521
rect 13430 33457 13494 33521
rect 13519 33457 13583 33521
rect 13627 33493 13691 33557
rect 1095 33369 1159 33433
rect 1184 33369 1248 33433
rect 1274 33369 1338 33433
rect 1364 33369 1428 33433
rect 1454 33369 1518 33433
rect 1595 33331 1659 33395
rect 1095 33253 1159 33317
rect 1184 33253 1248 33317
rect 1274 33253 1338 33317
rect 1364 33253 1428 33317
rect 1454 33253 1518 33317
rect 1095 33137 1159 33201
rect 1184 33137 1248 33201
rect 1274 33137 1338 33201
rect 1364 33137 1428 33201
rect 1454 33137 1518 33201
rect 973 33044 1037 33108
rect 1063 33044 1127 33108
rect 1153 33044 1217 33108
rect 1243 33044 1307 33108
rect 1333 33044 1397 33108
rect 1423 33044 1487 33108
rect 973 32964 1037 33028
rect 1063 32964 1127 33028
rect 1153 32964 1217 33028
rect 1243 32964 1307 33028
rect 1333 32964 1397 33028
rect 1423 32964 1487 33028
rect 973 32884 1037 32948
rect 1063 32884 1127 32948
rect 1153 32884 1217 32948
rect 1243 32884 1307 32948
rect 1333 32884 1397 32948
rect 1423 32884 1487 32948
rect 973 32804 1037 32868
rect 1063 32804 1127 32868
rect 1153 32804 1217 32868
rect 1243 32804 1307 32868
rect 1333 32804 1397 32868
rect 1423 32804 1487 32868
rect 973 32724 1037 32788
rect 1063 32724 1127 32788
rect 1153 32724 1217 32788
rect 1243 32724 1307 32788
rect 1333 32724 1397 32788
rect 1423 32724 1487 32788
rect 973 32644 1037 32708
rect 1063 32644 1127 32708
rect 1153 32644 1217 32708
rect 1243 32644 1307 32708
rect 1333 32644 1397 32708
rect 1423 32644 1487 32708
rect 973 32564 1037 32628
rect 1063 32564 1127 32628
rect 1153 32564 1217 32628
rect 1243 32564 1307 32628
rect 1333 32564 1397 32628
rect 1423 32564 1487 32628
rect 973 32484 1037 32548
rect 1063 32484 1127 32548
rect 1153 32484 1217 32548
rect 1243 32484 1307 32548
rect 1333 32484 1397 32548
rect 1423 32484 1487 32548
rect 973 32404 1037 32468
rect 1063 32404 1127 32468
rect 1153 32404 1217 32468
rect 1243 32404 1307 32468
rect 1333 32404 1397 32468
rect 1423 32404 1487 32468
rect 973 32324 1037 32388
rect 1063 32324 1127 32388
rect 1153 32324 1217 32388
rect 1243 32324 1307 32388
rect 1333 32324 1397 32388
rect 1423 32324 1487 32388
rect 973 32244 1037 32308
rect 1063 32244 1127 32308
rect 1153 32244 1217 32308
rect 1243 32244 1307 32308
rect 1333 32244 1397 32308
rect 1423 32244 1487 32308
rect 973 32164 1037 32228
rect 1063 32164 1127 32228
rect 1153 32164 1217 32228
rect 1243 32164 1307 32228
rect 1333 32164 1397 32228
rect 1423 32164 1487 32228
rect 973 32084 1037 32148
rect 1063 32084 1127 32148
rect 1153 32084 1217 32148
rect 1243 32084 1307 32148
rect 1333 32084 1397 32148
rect 1423 32084 1487 32148
rect 973 32004 1037 32068
rect 1063 32004 1127 32068
rect 1153 32004 1217 32068
rect 1243 32004 1307 32068
rect 1333 32004 1397 32068
rect 1423 32004 1487 32068
rect 973 31924 1037 31988
rect 1063 31924 1127 31988
rect 1153 31924 1217 31988
rect 1243 31924 1307 31988
rect 1333 31924 1397 31988
rect 1423 31924 1487 31988
rect 973 31844 1037 31908
rect 1063 31844 1127 31908
rect 1153 31844 1217 31908
rect 1243 31844 1307 31908
rect 1333 31844 1397 31908
rect 1423 31844 1487 31908
rect 973 31764 1037 31828
rect 1063 31764 1127 31828
rect 1153 31764 1217 31828
rect 1243 31764 1307 31828
rect 1333 31764 1397 31828
rect 1423 31764 1487 31828
rect 973 31684 1037 31748
rect 1063 31684 1127 31748
rect 1153 31684 1217 31748
rect 1243 31684 1307 31748
rect 1333 31684 1397 31748
rect 1423 31684 1487 31748
rect 973 31604 1037 31668
rect 1063 31604 1127 31668
rect 1153 31604 1217 31668
rect 1243 31604 1307 31668
rect 1333 31604 1397 31668
rect 1423 31604 1487 31668
rect 973 31524 1037 31588
rect 1063 31524 1127 31588
rect 1153 31524 1217 31588
rect 1243 31524 1307 31588
rect 1333 31524 1397 31588
rect 1423 31524 1487 31588
rect 973 31444 1037 31508
rect 1063 31444 1127 31508
rect 1153 31444 1217 31508
rect 1243 31444 1307 31508
rect 1333 31444 1397 31508
rect 1423 31444 1487 31508
rect 973 31364 1037 31428
rect 1063 31364 1127 31428
rect 1153 31364 1217 31428
rect 1243 31364 1307 31428
rect 1333 31364 1397 31428
rect 1423 31364 1487 31428
rect 973 31284 1037 31348
rect 1063 31284 1127 31348
rect 1153 31284 1217 31348
rect 1243 31284 1307 31348
rect 1333 31284 1397 31348
rect 1423 31284 1487 31348
rect 973 31204 1037 31268
rect 1063 31204 1127 31268
rect 1153 31204 1217 31268
rect 1243 31204 1307 31268
rect 1333 31204 1397 31268
rect 1423 31204 1487 31268
rect 973 31124 1037 31188
rect 1063 31124 1127 31188
rect 1153 31124 1217 31188
rect 1243 31124 1307 31188
rect 1333 31124 1397 31188
rect 1423 31124 1487 31188
rect 973 31044 1037 31108
rect 1063 31044 1127 31108
rect 1153 31044 1217 31108
rect 1243 31044 1307 31108
rect 1333 31044 1397 31108
rect 1423 31044 1487 31108
rect 973 30964 1037 31028
rect 1063 30964 1127 31028
rect 1153 30964 1217 31028
rect 1243 30964 1307 31028
rect 1333 30964 1397 31028
rect 1423 30964 1487 31028
rect 973 30884 1037 30948
rect 1063 30884 1127 30948
rect 1153 30884 1217 30948
rect 1243 30884 1307 30948
rect 1333 30884 1397 30948
rect 1423 30884 1487 30948
rect 973 30804 1037 30868
rect 1063 30804 1127 30868
rect 1153 30804 1217 30868
rect 1243 30804 1307 30868
rect 1333 30804 1397 30868
rect 1423 30804 1487 30868
rect 973 30724 1037 30788
rect 1063 30724 1127 30788
rect 1153 30724 1217 30788
rect 1243 30724 1307 30788
rect 1333 30724 1397 30788
rect 1423 30724 1487 30788
rect 973 30644 1037 30708
rect 1063 30644 1127 30708
rect 1153 30644 1217 30708
rect 1243 30644 1307 30708
rect 1333 30644 1397 30708
rect 1423 30644 1487 30708
rect 973 30564 1037 30628
rect 1063 30564 1127 30628
rect 1153 30564 1217 30628
rect 1243 30564 1307 30628
rect 1333 30564 1397 30628
rect 1423 30564 1487 30628
rect 973 30484 1037 30548
rect 1063 30484 1127 30548
rect 1153 30484 1217 30548
rect 1243 30484 1307 30548
rect 1333 30484 1397 30548
rect 1423 30484 1487 30548
rect 973 30404 1037 30468
rect 1063 30404 1127 30468
rect 1153 30404 1217 30468
rect 1243 30404 1307 30468
rect 1333 30404 1397 30468
rect 1423 30404 1487 30468
rect 973 30324 1037 30388
rect 1063 30324 1127 30388
rect 1153 30324 1217 30388
rect 1243 30324 1307 30388
rect 1333 30324 1397 30388
rect 1423 30324 1487 30388
rect 973 30244 1037 30308
rect 1063 30244 1127 30308
rect 1153 30244 1217 30308
rect 1243 30244 1307 30308
rect 1333 30244 1397 30308
rect 1423 30244 1487 30308
rect 973 30164 1037 30228
rect 1063 30164 1127 30228
rect 1153 30164 1217 30228
rect 1243 30164 1307 30228
rect 1333 30164 1397 30228
rect 1423 30164 1487 30228
rect 973 30084 1037 30148
rect 1063 30084 1127 30148
rect 1153 30084 1217 30148
rect 1243 30084 1307 30148
rect 1333 30084 1397 30148
rect 1423 30084 1487 30148
rect 973 30004 1037 30068
rect 1063 30004 1127 30068
rect 1153 30004 1217 30068
rect 1243 30004 1307 30068
rect 1333 30004 1397 30068
rect 1423 30004 1487 30068
rect 973 29924 1037 29988
rect 1063 29924 1127 29988
rect 1153 29924 1217 29988
rect 1243 29924 1307 29988
rect 1333 29924 1397 29988
rect 1423 29924 1487 29988
rect 973 29844 1037 29908
rect 1063 29844 1127 29908
rect 1153 29844 1217 29908
rect 1243 29844 1307 29908
rect 1333 29844 1397 29908
rect 1423 29844 1487 29908
rect 973 29764 1037 29828
rect 1063 29764 1127 29828
rect 1153 29764 1217 29828
rect 1243 29764 1307 29828
rect 1333 29764 1397 29828
rect 1423 29764 1487 29828
rect 973 29684 1037 29748
rect 1063 29684 1127 29748
rect 1153 29684 1217 29748
rect 1243 29684 1307 29748
rect 1333 29684 1397 29748
rect 1423 29684 1487 29748
rect 973 29604 1037 29668
rect 1063 29604 1127 29668
rect 1153 29604 1217 29668
rect 1243 29604 1307 29668
rect 1333 29604 1397 29668
rect 1423 29604 1487 29668
rect 973 29524 1037 29588
rect 1063 29524 1127 29588
rect 1153 29524 1217 29588
rect 1243 29524 1307 29588
rect 1333 29524 1397 29588
rect 1423 29524 1487 29588
rect 973 29444 1037 29508
rect 1063 29444 1127 29508
rect 1153 29444 1217 29508
rect 1243 29444 1307 29508
rect 1333 29444 1397 29508
rect 1423 29444 1487 29508
rect 973 29364 1037 29428
rect 1063 29364 1127 29428
rect 1153 29364 1217 29428
rect 1243 29364 1307 29428
rect 1333 29364 1397 29428
rect 1423 29364 1487 29428
rect 973 29284 1037 29348
rect 1063 29284 1127 29348
rect 1153 29284 1217 29348
rect 1243 29284 1307 29348
rect 1333 29284 1397 29348
rect 1423 29284 1487 29348
rect 973 29204 1037 29268
rect 1063 29204 1127 29268
rect 1153 29204 1217 29268
rect 1243 29204 1307 29268
rect 1333 29204 1397 29268
rect 1423 29204 1487 29268
rect 973 29124 1037 29188
rect 1063 29124 1127 29188
rect 1153 29124 1217 29188
rect 1243 29124 1307 29188
rect 1333 29124 1397 29188
rect 1423 29124 1487 29188
rect 973 29044 1037 29108
rect 1063 29044 1127 29108
rect 1153 29044 1217 29108
rect 1243 29044 1307 29108
rect 1333 29044 1397 29108
rect 1423 29044 1487 29108
rect 973 28964 1037 29028
rect 1063 28964 1127 29028
rect 1153 28964 1217 29028
rect 1243 28964 1307 29028
rect 1333 28964 1397 29028
rect 1423 28964 1487 29028
rect 973 28884 1037 28948
rect 1063 28884 1127 28948
rect 1153 28884 1217 28948
rect 1243 28884 1307 28948
rect 1333 28884 1397 28948
rect 1423 28884 1487 28948
rect 973 28804 1037 28868
rect 1063 28804 1127 28868
rect 1153 28804 1217 28868
rect 1243 28804 1307 28868
rect 1333 28804 1397 28868
rect 1423 28804 1487 28868
rect 973 28724 1037 28788
rect 1063 28724 1127 28788
rect 1153 28724 1217 28788
rect 1243 28724 1307 28788
rect 1333 28724 1397 28788
rect 1423 28724 1487 28788
rect 973 28644 1037 28708
rect 1063 28644 1127 28708
rect 1153 28644 1217 28708
rect 1243 28644 1307 28708
rect 1333 28644 1397 28708
rect 1423 28644 1487 28708
rect 973 28564 1037 28628
rect 1063 28564 1127 28628
rect 1153 28564 1217 28628
rect 1243 28564 1307 28628
rect 1333 28564 1397 28628
rect 1423 28564 1487 28628
rect 973 28484 1037 28548
rect 1063 28484 1127 28548
rect 1153 28484 1217 28548
rect 1243 28484 1307 28548
rect 1333 28484 1397 28548
rect 1423 28484 1487 28548
rect 973 28404 1037 28468
rect 1063 28404 1127 28468
rect 1153 28404 1217 28468
rect 1243 28404 1307 28468
rect 1333 28404 1397 28468
rect 1423 28404 1487 28468
rect 973 28324 1037 28388
rect 1063 28324 1127 28388
rect 1153 28324 1217 28388
rect 1243 28324 1307 28388
rect 1333 28324 1397 28388
rect 1423 28324 1487 28388
rect 973 28244 1037 28308
rect 1063 28244 1127 28308
rect 1153 28244 1217 28308
rect 1243 28244 1307 28308
rect 1333 28244 1397 28308
rect 1423 28244 1487 28308
rect 973 28164 1037 28228
rect 1063 28164 1127 28228
rect 1153 28164 1217 28228
rect 1243 28164 1307 28228
rect 1333 28164 1397 28228
rect 1423 28164 1487 28228
rect 973 28084 1037 28148
rect 1063 28084 1127 28148
rect 1153 28084 1217 28148
rect 1243 28084 1307 28148
rect 1333 28084 1397 28148
rect 1423 28084 1487 28148
rect 973 28004 1037 28068
rect 1063 28004 1127 28068
rect 1153 28004 1217 28068
rect 1243 28004 1307 28068
rect 1333 28004 1397 28068
rect 1423 28004 1487 28068
rect 973 27924 1037 27988
rect 1063 27924 1127 27988
rect 1153 27924 1217 27988
rect 1243 27924 1307 27988
rect 1333 27924 1397 27988
rect 1423 27924 1487 27988
rect 973 27844 1037 27908
rect 1063 27844 1127 27908
rect 1153 27844 1217 27908
rect 1243 27844 1307 27908
rect 1333 27844 1397 27908
rect 1423 27844 1487 27908
rect 973 27764 1037 27828
rect 1063 27764 1127 27828
rect 1153 27764 1217 27828
rect 1243 27764 1307 27828
rect 1333 27764 1397 27828
rect 1423 27764 1487 27828
rect 973 27684 1037 27748
rect 1063 27684 1127 27748
rect 1153 27684 1217 27748
rect 1243 27684 1307 27748
rect 1333 27684 1397 27748
rect 1423 27684 1487 27748
rect 973 27604 1037 27668
rect 1063 27604 1127 27668
rect 1153 27604 1217 27668
rect 1243 27604 1307 27668
rect 1333 27604 1397 27668
rect 1423 27604 1487 27668
rect 973 27524 1037 27588
rect 1063 27524 1127 27588
rect 1153 27524 1217 27588
rect 1243 27524 1307 27588
rect 1333 27524 1397 27588
rect 1423 27524 1487 27588
rect 973 27444 1037 27508
rect 1063 27444 1127 27508
rect 1153 27444 1217 27508
rect 1243 27444 1307 27508
rect 1333 27444 1397 27508
rect 1423 27444 1487 27508
rect 973 27364 1037 27428
rect 1063 27364 1127 27428
rect 1153 27364 1217 27428
rect 1243 27364 1307 27428
rect 1333 27364 1397 27428
rect 1423 27364 1487 27428
rect 973 27284 1037 27348
rect 1063 27284 1127 27348
rect 1153 27284 1217 27348
rect 1243 27284 1307 27348
rect 1333 27284 1397 27348
rect 1423 27284 1487 27348
rect 973 27204 1037 27268
rect 1063 27204 1127 27268
rect 1153 27204 1217 27268
rect 1243 27204 1307 27268
rect 1333 27204 1397 27268
rect 1423 27204 1487 27268
rect 973 27124 1037 27188
rect 1063 27124 1127 27188
rect 1153 27124 1217 27188
rect 1243 27124 1307 27188
rect 1333 27124 1397 27188
rect 1423 27124 1487 27188
rect 973 27044 1037 27108
rect 1063 27044 1127 27108
rect 1153 27044 1217 27108
rect 1243 27044 1307 27108
rect 1333 27044 1397 27108
rect 1423 27044 1487 27108
rect 973 26964 1037 27028
rect 1063 26964 1127 27028
rect 1153 26964 1217 27028
rect 1243 26964 1307 27028
rect 1333 26964 1397 27028
rect 1423 26964 1487 27028
rect 973 26884 1037 26948
rect 1063 26884 1127 26948
rect 1153 26884 1217 26948
rect 1243 26884 1307 26948
rect 1333 26884 1397 26948
rect 1423 26884 1487 26948
rect 973 26804 1037 26868
rect 1063 26804 1127 26868
rect 1153 26804 1217 26868
rect 1243 26804 1307 26868
rect 1333 26804 1397 26868
rect 1423 26804 1487 26868
rect 973 26724 1037 26788
rect 1063 26724 1127 26788
rect 1153 26724 1217 26788
rect 1243 26724 1307 26788
rect 1333 26724 1397 26788
rect 1423 26724 1487 26788
rect 973 26644 1037 26708
rect 1063 26644 1127 26708
rect 1153 26644 1217 26708
rect 1243 26644 1307 26708
rect 1333 26644 1397 26708
rect 1423 26644 1487 26708
rect 973 26564 1037 26628
rect 1063 26564 1127 26628
rect 1153 26564 1217 26628
rect 1243 26564 1307 26628
rect 1333 26564 1397 26628
rect 1423 26564 1487 26628
rect 973 26484 1037 26548
rect 1063 26484 1127 26548
rect 1153 26484 1217 26548
rect 1243 26484 1307 26548
rect 1333 26484 1397 26548
rect 1423 26484 1487 26548
rect 973 26404 1037 26468
rect 1063 26404 1127 26468
rect 1153 26404 1217 26468
rect 1243 26404 1307 26468
rect 1333 26404 1397 26468
rect 1423 26404 1487 26468
rect 973 26324 1037 26388
rect 1063 26324 1127 26388
rect 1153 26324 1217 26388
rect 1243 26324 1307 26388
rect 1333 26324 1397 26388
rect 1423 26324 1487 26388
rect 973 26244 1037 26308
rect 1063 26244 1127 26308
rect 1153 26244 1217 26308
rect 1243 26244 1307 26308
rect 1333 26244 1397 26308
rect 1423 26244 1487 26308
rect 973 26164 1037 26228
rect 1063 26164 1127 26228
rect 1153 26164 1217 26228
rect 1243 26164 1307 26228
rect 1333 26164 1397 26228
rect 1423 26164 1487 26228
rect 973 26084 1037 26148
rect 1063 26084 1127 26148
rect 1153 26084 1217 26148
rect 1243 26084 1307 26148
rect 1333 26084 1397 26148
rect 1423 26084 1487 26148
rect 973 26004 1037 26068
rect 1063 26004 1127 26068
rect 1153 26004 1217 26068
rect 1243 26004 1307 26068
rect 1333 26004 1397 26068
rect 1423 26004 1487 26068
rect 973 25924 1037 25988
rect 1063 25924 1127 25988
rect 1153 25924 1217 25988
rect 1243 25924 1307 25988
rect 1333 25924 1397 25988
rect 1423 25924 1487 25988
rect 973 25844 1037 25908
rect 1063 25844 1127 25908
rect 1153 25844 1217 25908
rect 1243 25844 1307 25908
rect 1333 25844 1397 25908
rect 1423 25844 1487 25908
rect 973 25764 1037 25828
rect 1063 25764 1127 25828
rect 1153 25764 1217 25828
rect 1243 25764 1307 25828
rect 1333 25764 1397 25828
rect 1423 25764 1487 25828
rect 973 25684 1037 25748
rect 1063 25684 1127 25748
rect 1153 25684 1217 25748
rect 1243 25684 1307 25748
rect 1333 25684 1397 25748
rect 1423 25684 1487 25748
rect 973 25604 1037 25668
rect 1063 25604 1127 25668
rect 1153 25604 1217 25668
rect 1243 25604 1307 25668
rect 1333 25604 1397 25668
rect 1423 25604 1487 25668
rect 973 25524 1037 25588
rect 1063 25524 1127 25588
rect 1153 25524 1217 25588
rect 1243 25524 1307 25588
rect 1333 25524 1397 25588
rect 1423 25524 1487 25588
rect 973 25444 1037 25508
rect 1063 25444 1127 25508
rect 1153 25444 1217 25508
rect 1243 25444 1307 25508
rect 1333 25444 1397 25508
rect 1423 25444 1487 25508
rect 973 25364 1037 25428
rect 1063 25364 1127 25428
rect 1153 25364 1217 25428
rect 1243 25364 1307 25428
rect 1333 25364 1397 25428
rect 1423 25364 1487 25428
rect 973 25284 1037 25348
rect 1063 25284 1127 25348
rect 1153 25284 1217 25348
rect 1243 25284 1307 25348
rect 1333 25284 1397 25348
rect 1423 25284 1487 25348
rect 973 25204 1037 25268
rect 1063 25204 1127 25268
rect 1153 25204 1217 25268
rect 1243 25204 1307 25268
rect 1333 25204 1397 25268
rect 1423 25204 1487 25268
rect 973 25124 1037 25188
rect 1063 25124 1127 25188
rect 1153 25124 1217 25188
rect 1243 25124 1307 25188
rect 1333 25124 1397 25188
rect 1423 25124 1487 25188
rect 973 25044 1037 25108
rect 1063 25044 1127 25108
rect 1153 25044 1217 25108
rect 1243 25044 1307 25108
rect 1333 25044 1397 25108
rect 1423 25044 1487 25108
rect 973 24964 1037 25028
rect 1063 24964 1127 25028
rect 1153 24964 1217 25028
rect 1243 24964 1307 25028
rect 1333 24964 1397 25028
rect 1423 24964 1487 25028
rect 973 24884 1037 24948
rect 1063 24884 1127 24948
rect 1153 24884 1217 24948
rect 1243 24884 1307 24948
rect 1333 24884 1397 24948
rect 1423 24884 1487 24948
rect 973 24804 1037 24868
rect 1063 24804 1127 24868
rect 1153 24804 1217 24868
rect 1243 24804 1307 24868
rect 1333 24804 1397 24868
rect 1423 24804 1487 24868
rect 973 24724 1037 24788
rect 1063 24724 1127 24788
rect 1153 24724 1217 24788
rect 1243 24724 1307 24788
rect 1333 24724 1397 24788
rect 1423 24724 1487 24788
rect 973 24644 1037 24708
rect 1063 24644 1127 24708
rect 1153 24644 1217 24708
rect 1243 24644 1307 24708
rect 1333 24644 1397 24708
rect 1423 24644 1487 24708
rect 973 24564 1037 24628
rect 1063 24564 1127 24628
rect 1153 24564 1217 24628
rect 1243 24564 1307 24628
rect 1333 24564 1397 24628
rect 1423 24564 1487 24628
rect 973 24484 1037 24548
rect 1063 24484 1127 24548
rect 1153 24484 1217 24548
rect 1243 24484 1307 24548
rect 1333 24484 1397 24548
rect 1423 24484 1487 24548
rect 973 24404 1037 24468
rect 1063 24404 1127 24468
rect 1153 24404 1217 24468
rect 1243 24404 1307 24468
rect 1333 24404 1397 24468
rect 1423 24404 1487 24468
rect 973 24324 1037 24388
rect 1063 24324 1127 24388
rect 1153 24324 1217 24388
rect 1243 24324 1307 24388
rect 1333 24324 1397 24388
rect 1423 24324 1487 24388
rect 973 24244 1037 24308
rect 1063 24244 1127 24308
rect 1153 24244 1217 24308
rect 1243 24244 1307 24308
rect 1333 24244 1397 24308
rect 1423 24244 1487 24308
rect 973 24164 1037 24228
rect 1063 24164 1127 24228
rect 1153 24164 1217 24228
rect 1243 24164 1307 24228
rect 1333 24164 1397 24228
rect 1423 24164 1487 24228
rect 973 24084 1037 24148
rect 1063 24084 1127 24148
rect 1153 24084 1217 24148
rect 1243 24084 1307 24148
rect 1333 24084 1397 24148
rect 1423 24084 1487 24148
rect 973 24004 1037 24068
rect 1063 24004 1127 24068
rect 1153 24004 1217 24068
rect 1243 24004 1307 24068
rect 1333 24004 1397 24068
rect 1423 24004 1487 24068
rect 973 23924 1037 23988
rect 1063 23924 1127 23988
rect 1153 23924 1217 23988
rect 1243 23924 1307 23988
rect 1333 23924 1397 23988
rect 1423 23924 1487 23988
rect 973 23844 1037 23908
rect 1063 23844 1127 23908
rect 1153 23844 1217 23908
rect 1243 23844 1307 23908
rect 1333 23844 1397 23908
rect 1423 23844 1487 23908
rect 973 23764 1037 23828
rect 1063 23764 1127 23828
rect 1153 23764 1217 23828
rect 1243 23764 1307 23828
rect 1333 23764 1397 23828
rect 1423 23764 1487 23828
rect 973 23684 1037 23748
rect 1063 23684 1127 23748
rect 1153 23684 1217 23748
rect 1243 23684 1307 23748
rect 1333 23684 1397 23748
rect 1423 23684 1487 23748
rect 973 23604 1037 23668
rect 1063 23604 1127 23668
rect 1153 23604 1217 23668
rect 1243 23604 1307 23668
rect 1333 23604 1397 23668
rect 1423 23604 1487 23668
rect 973 23524 1037 23588
rect 1063 23524 1127 23588
rect 1153 23524 1217 23588
rect 1243 23524 1307 23588
rect 1333 23524 1397 23588
rect 1423 23524 1487 23588
rect 973 23444 1037 23508
rect 1063 23444 1127 23508
rect 1153 23444 1217 23508
rect 1243 23444 1307 23508
rect 1333 23444 1397 23508
rect 1423 23444 1487 23508
rect 973 23364 1037 23428
rect 1063 23364 1127 23428
rect 1153 23364 1217 23428
rect 1243 23364 1307 23428
rect 1333 23364 1397 23428
rect 1423 23364 1487 23428
rect 973 23284 1037 23348
rect 1063 23284 1127 23348
rect 1153 23284 1217 23348
rect 1243 23284 1307 23348
rect 1333 23284 1397 23348
rect 1423 23284 1487 23348
rect 973 23203 1037 23267
rect 1063 23203 1127 23267
rect 1153 23203 1217 23267
rect 1243 23203 1307 23267
rect 1333 23203 1397 23267
rect 1423 23203 1487 23267
rect 973 23122 1037 23186
rect 1063 23122 1127 23186
rect 1153 23122 1217 23186
rect 1243 23122 1307 23186
rect 1333 23122 1397 23186
rect 1423 23122 1487 23186
rect 973 23041 1037 23105
rect 1063 23041 1127 23105
rect 1153 23041 1217 23105
rect 1243 23041 1307 23105
rect 1333 23041 1397 23105
rect 1423 23041 1487 23105
rect 973 22960 1037 23024
rect 1063 22960 1127 23024
rect 1153 22960 1217 23024
rect 1243 22960 1307 23024
rect 1333 22960 1397 23024
rect 1423 22960 1487 23024
rect 973 22879 1037 22943
rect 1063 22879 1127 22943
rect 1153 22879 1217 22943
rect 1243 22879 1307 22943
rect 1333 22879 1397 22943
rect 1423 22879 1487 22943
rect 973 22798 1037 22862
rect 1063 22798 1127 22862
rect 1153 22798 1217 22862
rect 1243 22798 1307 22862
rect 1333 22798 1397 22862
rect 1423 22798 1487 22862
rect 973 22717 1037 22781
rect 1063 22717 1127 22781
rect 1153 22717 1217 22781
rect 1243 22717 1307 22781
rect 1333 22717 1397 22781
rect 1423 22717 1487 22781
rect 973 22636 1037 22700
rect 1063 22636 1127 22700
rect 1153 22636 1217 22700
rect 1243 22636 1307 22700
rect 1333 22636 1397 22700
rect 1423 22636 1487 22700
rect 973 22555 1037 22619
rect 1063 22555 1127 22619
rect 1153 22555 1217 22619
rect 1243 22555 1307 22619
rect 1333 22555 1397 22619
rect 1423 22555 1487 22619
rect 973 22474 1037 22538
rect 1063 22474 1127 22538
rect 1153 22474 1217 22538
rect 1243 22474 1307 22538
rect 1333 22474 1397 22538
rect 1423 22474 1487 22538
rect 973 22393 1037 22457
rect 1063 22393 1127 22457
rect 1153 22393 1217 22457
rect 1243 22393 1307 22457
rect 1333 22393 1397 22457
rect 1423 22393 1487 22457
rect 973 22312 1037 22376
rect 1063 22312 1127 22376
rect 1153 22312 1217 22376
rect 1243 22312 1307 22376
rect 1333 22312 1397 22376
rect 1423 22312 1487 22376
rect 973 22231 1037 22295
rect 1063 22231 1127 22295
rect 1153 22231 1217 22295
rect 1243 22231 1307 22295
rect 1333 22231 1397 22295
rect 1423 22231 1487 22295
rect 973 22150 1037 22214
rect 1063 22150 1127 22214
rect 1153 22150 1217 22214
rect 1243 22150 1307 22214
rect 1333 22150 1397 22214
rect 1423 22150 1487 22214
rect 973 22069 1037 22133
rect 1063 22069 1127 22133
rect 1153 22069 1217 22133
rect 1243 22069 1307 22133
rect 1333 22069 1397 22133
rect 1423 22069 1487 22133
rect 973 21988 1037 22052
rect 1063 21988 1127 22052
rect 1153 21988 1217 22052
rect 1243 21988 1307 22052
rect 1333 21988 1397 22052
rect 1423 21988 1487 22052
rect 973 21907 1037 21971
rect 1063 21907 1127 21971
rect 1153 21907 1217 21971
rect 1243 21907 1307 21971
rect 1333 21907 1397 21971
rect 1423 21907 1487 21971
rect 973 21826 1037 21890
rect 1063 21826 1127 21890
rect 1153 21826 1217 21890
rect 1243 21826 1307 21890
rect 1333 21826 1397 21890
rect 1423 21826 1487 21890
rect 973 21745 1037 21809
rect 1063 21745 1127 21809
rect 1153 21745 1217 21809
rect 1243 21745 1307 21809
rect 1333 21745 1397 21809
rect 1423 21745 1487 21809
rect 973 21664 1037 21728
rect 1063 21664 1127 21728
rect 1153 21664 1217 21728
rect 1243 21664 1307 21728
rect 1333 21664 1397 21728
rect 1423 21664 1487 21728
rect 973 21583 1037 21647
rect 1063 21583 1127 21647
rect 1153 21583 1217 21647
rect 1243 21583 1307 21647
rect 1333 21583 1397 21647
rect 1423 21583 1487 21647
rect 973 21502 1037 21566
rect 1063 21502 1127 21566
rect 1153 21502 1217 21566
rect 1243 21502 1307 21566
rect 1333 21502 1397 21566
rect 1423 21502 1487 21566
rect 973 21421 1037 21485
rect 1063 21421 1127 21485
rect 1153 21421 1217 21485
rect 1243 21421 1307 21485
rect 1333 21421 1397 21485
rect 1423 21421 1487 21485
rect 973 21340 1037 21404
rect 1063 21340 1127 21404
rect 1153 21340 1217 21404
rect 1243 21340 1307 21404
rect 1333 21340 1397 21404
rect 1423 21340 1487 21404
rect 973 21259 1037 21323
rect 1063 21259 1127 21323
rect 1153 21259 1217 21323
rect 1243 21259 1307 21323
rect 1333 21259 1397 21323
rect 1423 21259 1487 21323
rect 973 21178 1037 21242
rect 1063 21178 1127 21242
rect 1153 21178 1217 21242
rect 1243 21178 1307 21242
rect 1333 21178 1397 21242
rect 1423 21178 1487 21242
rect 973 21097 1037 21161
rect 1063 21097 1127 21161
rect 1153 21097 1217 21161
rect 1243 21097 1307 21161
rect 1333 21097 1397 21161
rect 1423 21097 1487 21161
rect 973 21016 1037 21080
rect 1063 21016 1127 21080
rect 1153 21016 1217 21080
rect 1243 21016 1307 21080
rect 1333 21016 1397 21080
rect 1423 21016 1487 21080
rect 973 20935 1037 20999
rect 1063 20935 1127 20999
rect 1153 20935 1217 20999
rect 1243 20935 1307 20999
rect 1333 20935 1397 20999
rect 1423 20935 1487 20999
rect 973 20854 1037 20918
rect 1063 20854 1127 20918
rect 1153 20854 1217 20918
rect 1243 20854 1307 20918
rect 1333 20854 1397 20918
rect 1423 20854 1487 20918
rect 1522 20874 1586 20938
rect 1132 20718 1196 20782
rect 1303 20760 1367 20824
rect 1392 20760 1456 20824
rect 1482 20760 1546 20824
rect 1572 20760 1636 20824
rect 1662 20760 1726 20824
rect 1303 20644 1367 20708
rect 1392 20644 1456 20708
rect 1482 20644 1546 20708
rect 1572 20644 1636 20708
rect 1662 20644 1726 20708
rect 1303 20528 1367 20592
rect 1392 20528 1456 20592
rect 1482 20528 1546 20592
rect 1572 20528 1636 20592
rect 1662 20528 1726 20592
rect 1803 20566 1867 20630
rect 1515 20404 1579 20468
rect 1623 20440 1687 20504
rect 1712 20440 1776 20504
rect 1802 20440 1866 20504
rect 1892 20440 1956 20504
rect 1982 20440 2046 20504
rect 1623 20324 1687 20388
rect 1712 20324 1776 20388
rect 1802 20324 1866 20388
rect 1892 20324 1956 20388
rect 1982 20324 2046 20388
rect 1623 20208 1687 20272
rect 1712 20208 1776 20272
rect 1802 20208 1866 20272
rect 1892 20208 1956 20272
rect 1982 20208 2046 20272
rect 2128 20241 2192 20305
rect 13339 33331 13403 33395
rect 13480 33369 13544 33433
rect 13570 33369 13634 33433
rect 13660 33369 13724 33433
rect 13750 33369 13814 33433
rect 13839 33369 13903 33433
rect 13480 33253 13544 33317
rect 13570 33253 13634 33317
rect 13660 33253 13724 33317
rect 13750 33253 13814 33317
rect 13839 33253 13903 33317
rect 13480 33137 13544 33201
rect 13570 33137 13634 33201
rect 13660 33137 13724 33201
rect 13750 33137 13814 33201
rect 13839 33137 13903 33201
rect 13511 33044 13575 33108
rect 13601 33044 13665 33108
rect 13691 33044 13755 33108
rect 13781 33044 13845 33108
rect 13871 33044 13935 33108
rect 13961 33044 14025 33108
rect 13511 32964 13575 33028
rect 13601 32964 13665 33028
rect 13691 32964 13755 33028
rect 13781 32964 13845 33028
rect 13871 32964 13935 33028
rect 13961 32964 14025 33028
rect 13511 32884 13575 32948
rect 13601 32884 13665 32948
rect 13691 32884 13755 32948
rect 13781 32884 13845 32948
rect 13871 32884 13935 32948
rect 13961 32884 14025 32948
rect 13511 32804 13575 32868
rect 13601 32804 13665 32868
rect 13691 32804 13755 32868
rect 13781 32804 13845 32868
rect 13871 32804 13935 32868
rect 13961 32804 14025 32868
rect 13511 32724 13575 32788
rect 13601 32724 13665 32788
rect 13691 32724 13755 32788
rect 13781 32724 13845 32788
rect 13871 32724 13935 32788
rect 13961 32724 14025 32788
rect 13511 32644 13575 32708
rect 13601 32644 13665 32708
rect 13691 32644 13755 32708
rect 13781 32644 13845 32708
rect 13871 32644 13935 32708
rect 13961 32644 14025 32708
rect 13511 32564 13575 32628
rect 13601 32564 13665 32628
rect 13691 32564 13755 32628
rect 13781 32564 13845 32628
rect 13871 32564 13935 32628
rect 13961 32564 14025 32628
rect 13511 32484 13575 32548
rect 13601 32484 13665 32548
rect 13691 32484 13755 32548
rect 13781 32484 13845 32548
rect 13871 32484 13935 32548
rect 13961 32484 14025 32548
rect 13511 32404 13575 32468
rect 13601 32404 13665 32468
rect 13691 32404 13755 32468
rect 13781 32404 13845 32468
rect 13871 32404 13935 32468
rect 13961 32404 14025 32468
rect 13511 32324 13575 32388
rect 13601 32324 13665 32388
rect 13691 32324 13755 32388
rect 13781 32324 13845 32388
rect 13871 32324 13935 32388
rect 13961 32324 14025 32388
rect 13511 32244 13575 32308
rect 13601 32244 13665 32308
rect 13691 32244 13755 32308
rect 13781 32244 13845 32308
rect 13871 32244 13935 32308
rect 13961 32244 14025 32308
rect 13511 32164 13575 32228
rect 13601 32164 13665 32228
rect 13691 32164 13755 32228
rect 13781 32164 13845 32228
rect 13871 32164 13935 32228
rect 13961 32164 14025 32228
rect 13511 32084 13575 32148
rect 13601 32084 13665 32148
rect 13691 32084 13755 32148
rect 13781 32084 13845 32148
rect 13871 32084 13935 32148
rect 13961 32084 14025 32148
rect 13511 32004 13575 32068
rect 13601 32004 13665 32068
rect 13691 32004 13755 32068
rect 13781 32004 13845 32068
rect 13871 32004 13935 32068
rect 13961 32004 14025 32068
rect 13511 31924 13575 31988
rect 13601 31924 13665 31988
rect 13691 31924 13755 31988
rect 13781 31924 13845 31988
rect 13871 31924 13935 31988
rect 13961 31924 14025 31988
rect 13511 31844 13575 31908
rect 13601 31844 13665 31908
rect 13691 31844 13755 31908
rect 13781 31844 13845 31908
rect 13871 31844 13935 31908
rect 13961 31844 14025 31908
rect 13511 31764 13575 31828
rect 13601 31764 13665 31828
rect 13691 31764 13755 31828
rect 13781 31764 13845 31828
rect 13871 31764 13935 31828
rect 13961 31764 14025 31828
rect 13511 31684 13575 31748
rect 13601 31684 13665 31748
rect 13691 31684 13755 31748
rect 13781 31684 13845 31748
rect 13871 31684 13935 31748
rect 13961 31684 14025 31748
rect 13511 31604 13575 31668
rect 13601 31604 13665 31668
rect 13691 31604 13755 31668
rect 13781 31604 13845 31668
rect 13871 31604 13935 31668
rect 13961 31604 14025 31668
rect 13511 31524 13575 31588
rect 13601 31524 13665 31588
rect 13691 31524 13755 31588
rect 13781 31524 13845 31588
rect 13871 31524 13935 31588
rect 13961 31524 14025 31588
rect 13511 31444 13575 31508
rect 13601 31444 13665 31508
rect 13691 31444 13755 31508
rect 13781 31444 13845 31508
rect 13871 31444 13935 31508
rect 13961 31444 14025 31508
rect 13511 31364 13575 31428
rect 13601 31364 13665 31428
rect 13691 31364 13755 31428
rect 13781 31364 13845 31428
rect 13871 31364 13935 31428
rect 13961 31364 14025 31428
rect 13511 31284 13575 31348
rect 13601 31284 13665 31348
rect 13691 31284 13755 31348
rect 13781 31284 13845 31348
rect 13871 31284 13935 31348
rect 13961 31284 14025 31348
rect 13511 31204 13575 31268
rect 13601 31204 13665 31268
rect 13691 31204 13755 31268
rect 13781 31204 13845 31268
rect 13871 31204 13935 31268
rect 13961 31204 14025 31268
rect 13511 31124 13575 31188
rect 13601 31124 13665 31188
rect 13691 31124 13755 31188
rect 13781 31124 13845 31188
rect 13871 31124 13935 31188
rect 13961 31124 14025 31188
rect 13511 31044 13575 31108
rect 13601 31044 13665 31108
rect 13691 31044 13755 31108
rect 13781 31044 13845 31108
rect 13871 31044 13935 31108
rect 13961 31044 14025 31108
rect 13511 30964 13575 31028
rect 13601 30964 13665 31028
rect 13691 30964 13755 31028
rect 13781 30964 13845 31028
rect 13871 30964 13935 31028
rect 13961 30964 14025 31028
rect 13511 30884 13575 30948
rect 13601 30884 13665 30948
rect 13691 30884 13755 30948
rect 13781 30884 13845 30948
rect 13871 30884 13935 30948
rect 13961 30884 14025 30948
rect 13511 30804 13575 30868
rect 13601 30804 13665 30868
rect 13691 30804 13755 30868
rect 13781 30804 13845 30868
rect 13871 30804 13935 30868
rect 13961 30804 14025 30868
rect 13511 30724 13575 30788
rect 13601 30724 13665 30788
rect 13691 30724 13755 30788
rect 13781 30724 13845 30788
rect 13871 30724 13935 30788
rect 13961 30724 14025 30788
rect 13511 30644 13575 30708
rect 13601 30644 13665 30708
rect 13691 30644 13755 30708
rect 13781 30644 13845 30708
rect 13871 30644 13935 30708
rect 13961 30644 14025 30708
rect 13511 30564 13575 30628
rect 13601 30564 13665 30628
rect 13691 30564 13755 30628
rect 13781 30564 13845 30628
rect 13871 30564 13935 30628
rect 13961 30564 14025 30628
rect 13511 30484 13575 30548
rect 13601 30484 13665 30548
rect 13691 30484 13755 30548
rect 13781 30484 13845 30548
rect 13871 30484 13935 30548
rect 13961 30484 14025 30548
rect 13511 30404 13575 30468
rect 13601 30404 13665 30468
rect 13691 30404 13755 30468
rect 13781 30404 13845 30468
rect 13871 30404 13935 30468
rect 13961 30404 14025 30468
rect 13511 30324 13575 30388
rect 13601 30324 13665 30388
rect 13691 30324 13755 30388
rect 13781 30324 13845 30388
rect 13871 30324 13935 30388
rect 13961 30324 14025 30388
rect 13511 30244 13575 30308
rect 13601 30244 13665 30308
rect 13691 30244 13755 30308
rect 13781 30244 13845 30308
rect 13871 30244 13935 30308
rect 13961 30244 14025 30308
rect 13511 30164 13575 30228
rect 13601 30164 13665 30228
rect 13691 30164 13755 30228
rect 13781 30164 13845 30228
rect 13871 30164 13935 30228
rect 13961 30164 14025 30228
rect 13511 30084 13575 30148
rect 13601 30084 13665 30148
rect 13691 30084 13755 30148
rect 13781 30084 13845 30148
rect 13871 30084 13935 30148
rect 13961 30084 14025 30148
rect 13511 30004 13575 30068
rect 13601 30004 13665 30068
rect 13691 30004 13755 30068
rect 13781 30004 13845 30068
rect 13871 30004 13935 30068
rect 13961 30004 14025 30068
rect 13511 29924 13575 29988
rect 13601 29924 13665 29988
rect 13691 29924 13755 29988
rect 13781 29924 13845 29988
rect 13871 29924 13935 29988
rect 13961 29924 14025 29988
rect 13511 29844 13575 29908
rect 13601 29844 13665 29908
rect 13691 29844 13755 29908
rect 13781 29844 13845 29908
rect 13871 29844 13935 29908
rect 13961 29844 14025 29908
rect 13511 29764 13575 29828
rect 13601 29764 13665 29828
rect 13691 29764 13755 29828
rect 13781 29764 13845 29828
rect 13871 29764 13935 29828
rect 13961 29764 14025 29828
rect 13511 29684 13575 29748
rect 13601 29684 13665 29748
rect 13691 29684 13755 29748
rect 13781 29684 13845 29748
rect 13871 29684 13935 29748
rect 13961 29684 14025 29748
rect 13511 29604 13575 29668
rect 13601 29604 13665 29668
rect 13691 29604 13755 29668
rect 13781 29604 13845 29668
rect 13871 29604 13935 29668
rect 13961 29604 14025 29668
rect 13511 29524 13575 29588
rect 13601 29524 13665 29588
rect 13691 29524 13755 29588
rect 13781 29524 13845 29588
rect 13871 29524 13935 29588
rect 13961 29524 14025 29588
rect 13511 29444 13575 29508
rect 13601 29444 13665 29508
rect 13691 29444 13755 29508
rect 13781 29444 13845 29508
rect 13871 29444 13935 29508
rect 13961 29444 14025 29508
rect 13511 29364 13575 29428
rect 13601 29364 13665 29428
rect 13691 29364 13755 29428
rect 13781 29364 13845 29428
rect 13871 29364 13935 29428
rect 13961 29364 14025 29428
rect 13511 29284 13575 29348
rect 13601 29284 13665 29348
rect 13691 29284 13755 29348
rect 13781 29284 13845 29348
rect 13871 29284 13935 29348
rect 13961 29284 14025 29348
rect 13511 29204 13575 29268
rect 13601 29204 13665 29268
rect 13691 29204 13755 29268
rect 13781 29204 13845 29268
rect 13871 29204 13935 29268
rect 13961 29204 14025 29268
rect 13511 29124 13575 29188
rect 13601 29124 13665 29188
rect 13691 29124 13755 29188
rect 13781 29124 13845 29188
rect 13871 29124 13935 29188
rect 13961 29124 14025 29188
rect 13511 29044 13575 29108
rect 13601 29044 13665 29108
rect 13691 29044 13755 29108
rect 13781 29044 13845 29108
rect 13871 29044 13935 29108
rect 13961 29044 14025 29108
rect 13511 28964 13575 29028
rect 13601 28964 13665 29028
rect 13691 28964 13755 29028
rect 13781 28964 13845 29028
rect 13871 28964 13935 29028
rect 13961 28964 14025 29028
rect 13511 28884 13575 28948
rect 13601 28884 13665 28948
rect 13691 28884 13755 28948
rect 13781 28884 13845 28948
rect 13871 28884 13935 28948
rect 13961 28884 14025 28948
rect 13511 28804 13575 28868
rect 13601 28804 13665 28868
rect 13691 28804 13755 28868
rect 13781 28804 13845 28868
rect 13871 28804 13935 28868
rect 13961 28804 14025 28868
rect 13511 28724 13575 28788
rect 13601 28724 13665 28788
rect 13691 28724 13755 28788
rect 13781 28724 13845 28788
rect 13871 28724 13935 28788
rect 13961 28724 14025 28788
rect 13511 28644 13575 28708
rect 13601 28644 13665 28708
rect 13691 28644 13755 28708
rect 13781 28644 13845 28708
rect 13871 28644 13935 28708
rect 13961 28644 14025 28708
rect 13511 28564 13575 28628
rect 13601 28564 13665 28628
rect 13691 28564 13755 28628
rect 13781 28564 13845 28628
rect 13871 28564 13935 28628
rect 13961 28564 14025 28628
rect 13511 28484 13575 28548
rect 13601 28484 13665 28548
rect 13691 28484 13755 28548
rect 13781 28484 13845 28548
rect 13871 28484 13935 28548
rect 13961 28484 14025 28548
rect 13511 28404 13575 28468
rect 13601 28404 13665 28468
rect 13691 28404 13755 28468
rect 13781 28404 13845 28468
rect 13871 28404 13935 28468
rect 13961 28404 14025 28468
rect 13511 28324 13575 28388
rect 13601 28324 13665 28388
rect 13691 28324 13755 28388
rect 13781 28324 13845 28388
rect 13871 28324 13935 28388
rect 13961 28324 14025 28388
rect 13511 28244 13575 28308
rect 13601 28244 13665 28308
rect 13691 28244 13755 28308
rect 13781 28244 13845 28308
rect 13871 28244 13935 28308
rect 13961 28244 14025 28308
rect 13511 28164 13575 28228
rect 13601 28164 13665 28228
rect 13691 28164 13755 28228
rect 13781 28164 13845 28228
rect 13871 28164 13935 28228
rect 13961 28164 14025 28228
rect 13511 28084 13575 28148
rect 13601 28084 13665 28148
rect 13691 28084 13755 28148
rect 13781 28084 13845 28148
rect 13871 28084 13935 28148
rect 13961 28084 14025 28148
rect 13511 28004 13575 28068
rect 13601 28004 13665 28068
rect 13691 28004 13755 28068
rect 13781 28004 13845 28068
rect 13871 28004 13935 28068
rect 13961 28004 14025 28068
rect 13511 27924 13575 27988
rect 13601 27924 13665 27988
rect 13691 27924 13755 27988
rect 13781 27924 13845 27988
rect 13871 27924 13935 27988
rect 13961 27924 14025 27988
rect 13511 27844 13575 27908
rect 13601 27844 13665 27908
rect 13691 27844 13755 27908
rect 13781 27844 13845 27908
rect 13871 27844 13935 27908
rect 13961 27844 14025 27908
rect 13511 27764 13575 27828
rect 13601 27764 13665 27828
rect 13691 27764 13755 27828
rect 13781 27764 13845 27828
rect 13871 27764 13935 27828
rect 13961 27764 14025 27828
rect 13511 27684 13575 27748
rect 13601 27684 13665 27748
rect 13691 27684 13755 27748
rect 13781 27684 13845 27748
rect 13871 27684 13935 27748
rect 13961 27684 14025 27748
rect 13511 27604 13575 27668
rect 13601 27604 13665 27668
rect 13691 27604 13755 27668
rect 13781 27604 13845 27668
rect 13871 27604 13935 27668
rect 13961 27604 14025 27668
rect 13511 27524 13575 27588
rect 13601 27524 13665 27588
rect 13691 27524 13755 27588
rect 13781 27524 13845 27588
rect 13871 27524 13935 27588
rect 13961 27524 14025 27588
rect 13511 27444 13575 27508
rect 13601 27444 13665 27508
rect 13691 27444 13755 27508
rect 13781 27444 13845 27508
rect 13871 27444 13935 27508
rect 13961 27444 14025 27508
rect 13511 27364 13575 27428
rect 13601 27364 13665 27428
rect 13691 27364 13755 27428
rect 13781 27364 13845 27428
rect 13871 27364 13935 27428
rect 13961 27364 14025 27428
rect 13511 27284 13575 27348
rect 13601 27284 13665 27348
rect 13691 27284 13755 27348
rect 13781 27284 13845 27348
rect 13871 27284 13935 27348
rect 13961 27284 14025 27348
rect 13511 27204 13575 27268
rect 13601 27204 13665 27268
rect 13691 27204 13755 27268
rect 13781 27204 13845 27268
rect 13871 27204 13935 27268
rect 13961 27204 14025 27268
rect 13511 27124 13575 27188
rect 13601 27124 13665 27188
rect 13691 27124 13755 27188
rect 13781 27124 13845 27188
rect 13871 27124 13935 27188
rect 13961 27124 14025 27188
rect 13511 27044 13575 27108
rect 13601 27044 13665 27108
rect 13691 27044 13755 27108
rect 13781 27044 13845 27108
rect 13871 27044 13935 27108
rect 13961 27044 14025 27108
rect 13511 26964 13575 27028
rect 13601 26964 13665 27028
rect 13691 26964 13755 27028
rect 13781 26964 13845 27028
rect 13871 26964 13935 27028
rect 13961 26964 14025 27028
rect 13511 26884 13575 26948
rect 13601 26884 13665 26948
rect 13691 26884 13755 26948
rect 13781 26884 13845 26948
rect 13871 26884 13935 26948
rect 13961 26884 14025 26948
rect 13511 26804 13575 26868
rect 13601 26804 13665 26868
rect 13691 26804 13755 26868
rect 13781 26804 13845 26868
rect 13871 26804 13935 26868
rect 13961 26804 14025 26868
rect 13511 26724 13575 26788
rect 13601 26724 13665 26788
rect 13691 26724 13755 26788
rect 13781 26724 13845 26788
rect 13871 26724 13935 26788
rect 13961 26724 14025 26788
rect 13511 26644 13575 26708
rect 13601 26644 13665 26708
rect 13691 26644 13755 26708
rect 13781 26644 13845 26708
rect 13871 26644 13935 26708
rect 13961 26644 14025 26708
rect 13511 26564 13575 26628
rect 13601 26564 13665 26628
rect 13691 26564 13755 26628
rect 13781 26564 13845 26628
rect 13871 26564 13935 26628
rect 13961 26564 14025 26628
rect 13511 26484 13575 26548
rect 13601 26484 13665 26548
rect 13691 26484 13755 26548
rect 13781 26484 13845 26548
rect 13871 26484 13935 26548
rect 13961 26484 14025 26548
rect 13511 26404 13575 26468
rect 13601 26404 13665 26468
rect 13691 26404 13755 26468
rect 13781 26404 13845 26468
rect 13871 26404 13935 26468
rect 13961 26404 14025 26468
rect 13511 26324 13575 26388
rect 13601 26324 13665 26388
rect 13691 26324 13755 26388
rect 13781 26324 13845 26388
rect 13871 26324 13935 26388
rect 13961 26324 14025 26388
rect 13511 26244 13575 26308
rect 13601 26244 13665 26308
rect 13691 26244 13755 26308
rect 13781 26244 13845 26308
rect 13871 26244 13935 26308
rect 13961 26244 14025 26308
rect 13511 26164 13575 26228
rect 13601 26164 13665 26228
rect 13691 26164 13755 26228
rect 13781 26164 13845 26228
rect 13871 26164 13935 26228
rect 13961 26164 14025 26228
rect 13511 26084 13575 26148
rect 13601 26084 13665 26148
rect 13691 26084 13755 26148
rect 13781 26084 13845 26148
rect 13871 26084 13935 26148
rect 13961 26084 14025 26148
rect 13511 26004 13575 26068
rect 13601 26004 13665 26068
rect 13691 26004 13755 26068
rect 13781 26004 13845 26068
rect 13871 26004 13935 26068
rect 13961 26004 14025 26068
rect 13511 25924 13575 25988
rect 13601 25924 13665 25988
rect 13691 25924 13755 25988
rect 13781 25924 13845 25988
rect 13871 25924 13935 25988
rect 13961 25924 14025 25988
rect 13511 25844 13575 25908
rect 13601 25844 13665 25908
rect 13691 25844 13755 25908
rect 13781 25844 13845 25908
rect 13871 25844 13935 25908
rect 13961 25844 14025 25908
rect 13511 25764 13575 25828
rect 13601 25764 13665 25828
rect 13691 25764 13755 25828
rect 13781 25764 13845 25828
rect 13871 25764 13935 25828
rect 13961 25764 14025 25828
rect 13511 25684 13575 25748
rect 13601 25684 13665 25748
rect 13691 25684 13755 25748
rect 13781 25684 13845 25748
rect 13871 25684 13935 25748
rect 13961 25684 14025 25748
rect 13511 25604 13575 25668
rect 13601 25604 13665 25668
rect 13691 25604 13755 25668
rect 13781 25604 13845 25668
rect 13871 25604 13935 25668
rect 13961 25604 14025 25668
rect 13511 25524 13575 25588
rect 13601 25524 13665 25588
rect 13691 25524 13755 25588
rect 13781 25524 13845 25588
rect 13871 25524 13935 25588
rect 13961 25524 14025 25588
rect 13511 25444 13575 25508
rect 13601 25444 13665 25508
rect 13691 25444 13755 25508
rect 13781 25444 13845 25508
rect 13871 25444 13935 25508
rect 13961 25444 14025 25508
rect 13511 25364 13575 25428
rect 13601 25364 13665 25428
rect 13691 25364 13755 25428
rect 13781 25364 13845 25428
rect 13871 25364 13935 25428
rect 13961 25364 14025 25428
rect 13511 25284 13575 25348
rect 13601 25284 13665 25348
rect 13691 25284 13755 25348
rect 13781 25284 13845 25348
rect 13871 25284 13935 25348
rect 13961 25284 14025 25348
rect 13511 25204 13575 25268
rect 13601 25204 13665 25268
rect 13691 25204 13755 25268
rect 13781 25204 13845 25268
rect 13871 25204 13935 25268
rect 13961 25204 14025 25268
rect 13511 25124 13575 25188
rect 13601 25124 13665 25188
rect 13691 25124 13755 25188
rect 13781 25124 13845 25188
rect 13871 25124 13935 25188
rect 13961 25124 14025 25188
rect 13511 25044 13575 25108
rect 13601 25044 13665 25108
rect 13691 25044 13755 25108
rect 13781 25044 13845 25108
rect 13871 25044 13935 25108
rect 13961 25044 14025 25108
rect 13511 24964 13575 25028
rect 13601 24964 13665 25028
rect 13691 24964 13755 25028
rect 13781 24964 13845 25028
rect 13871 24964 13935 25028
rect 13961 24964 14025 25028
rect 13511 24884 13575 24948
rect 13601 24884 13665 24948
rect 13691 24884 13755 24948
rect 13781 24884 13845 24948
rect 13871 24884 13935 24948
rect 13961 24884 14025 24948
rect 13511 24804 13575 24868
rect 13601 24804 13665 24868
rect 13691 24804 13755 24868
rect 13781 24804 13845 24868
rect 13871 24804 13935 24868
rect 13961 24804 14025 24868
rect 13511 24724 13575 24788
rect 13601 24724 13665 24788
rect 13691 24724 13755 24788
rect 13781 24724 13845 24788
rect 13871 24724 13935 24788
rect 13961 24724 14025 24788
rect 13511 24644 13575 24708
rect 13601 24644 13665 24708
rect 13691 24644 13755 24708
rect 13781 24644 13845 24708
rect 13871 24644 13935 24708
rect 13961 24644 14025 24708
rect 13511 24564 13575 24628
rect 13601 24564 13665 24628
rect 13691 24564 13755 24628
rect 13781 24564 13845 24628
rect 13871 24564 13935 24628
rect 13961 24564 14025 24628
rect 13511 24484 13575 24548
rect 13601 24484 13665 24548
rect 13691 24484 13755 24548
rect 13781 24484 13845 24548
rect 13871 24484 13935 24548
rect 13961 24484 14025 24548
rect 13511 24404 13575 24468
rect 13601 24404 13665 24468
rect 13691 24404 13755 24468
rect 13781 24404 13845 24468
rect 13871 24404 13935 24468
rect 13961 24404 14025 24468
rect 13511 24324 13575 24388
rect 13601 24324 13665 24388
rect 13691 24324 13755 24388
rect 13781 24324 13845 24388
rect 13871 24324 13935 24388
rect 13961 24324 14025 24388
rect 13511 24244 13575 24308
rect 13601 24244 13665 24308
rect 13691 24244 13755 24308
rect 13781 24244 13845 24308
rect 13871 24244 13935 24308
rect 13961 24244 14025 24308
rect 13511 24164 13575 24228
rect 13601 24164 13665 24228
rect 13691 24164 13755 24228
rect 13781 24164 13845 24228
rect 13871 24164 13935 24228
rect 13961 24164 14025 24228
rect 13511 24084 13575 24148
rect 13601 24084 13665 24148
rect 13691 24084 13755 24148
rect 13781 24084 13845 24148
rect 13871 24084 13935 24148
rect 13961 24084 14025 24148
rect 13511 24004 13575 24068
rect 13601 24004 13665 24068
rect 13691 24004 13755 24068
rect 13781 24004 13845 24068
rect 13871 24004 13935 24068
rect 13961 24004 14025 24068
rect 13511 23924 13575 23988
rect 13601 23924 13665 23988
rect 13691 23924 13755 23988
rect 13781 23924 13845 23988
rect 13871 23924 13935 23988
rect 13961 23924 14025 23988
rect 13511 23844 13575 23908
rect 13601 23844 13665 23908
rect 13691 23844 13755 23908
rect 13781 23844 13845 23908
rect 13871 23844 13935 23908
rect 13961 23844 14025 23908
rect 13511 23764 13575 23828
rect 13601 23764 13665 23828
rect 13691 23764 13755 23828
rect 13781 23764 13845 23828
rect 13871 23764 13935 23828
rect 13961 23764 14025 23828
rect 13511 23684 13575 23748
rect 13601 23684 13665 23748
rect 13691 23684 13755 23748
rect 13781 23684 13845 23748
rect 13871 23684 13935 23748
rect 13961 23684 14025 23748
rect 13511 23604 13575 23668
rect 13601 23604 13665 23668
rect 13691 23604 13755 23668
rect 13781 23604 13845 23668
rect 13871 23604 13935 23668
rect 13961 23604 14025 23668
rect 13511 23524 13575 23588
rect 13601 23524 13665 23588
rect 13691 23524 13755 23588
rect 13781 23524 13845 23588
rect 13871 23524 13935 23588
rect 13961 23524 14025 23588
rect 13511 23444 13575 23508
rect 13601 23444 13665 23508
rect 13691 23444 13755 23508
rect 13781 23444 13845 23508
rect 13871 23444 13935 23508
rect 13961 23444 14025 23508
rect 13511 23364 13575 23428
rect 13601 23364 13665 23428
rect 13691 23364 13755 23428
rect 13781 23364 13845 23428
rect 13871 23364 13935 23428
rect 13961 23364 14025 23428
rect 13511 23284 13575 23348
rect 13601 23284 13665 23348
rect 13691 23284 13755 23348
rect 13781 23284 13845 23348
rect 13871 23284 13935 23348
rect 13961 23284 14025 23348
rect 13511 23203 13575 23267
rect 13601 23203 13665 23267
rect 13691 23203 13755 23267
rect 13781 23203 13845 23267
rect 13871 23203 13935 23267
rect 13961 23203 14025 23267
rect 13511 23122 13575 23186
rect 13601 23122 13665 23186
rect 13691 23122 13755 23186
rect 13781 23122 13845 23186
rect 13871 23122 13935 23186
rect 13961 23122 14025 23186
rect 13511 23041 13575 23105
rect 13601 23041 13665 23105
rect 13691 23041 13755 23105
rect 13781 23041 13845 23105
rect 13871 23041 13935 23105
rect 13961 23041 14025 23105
rect 13511 22960 13575 23024
rect 13601 22960 13665 23024
rect 13691 22960 13755 23024
rect 13781 22960 13845 23024
rect 13871 22960 13935 23024
rect 13961 22960 14025 23024
rect 13511 22879 13575 22943
rect 13601 22879 13665 22943
rect 13691 22879 13755 22943
rect 13781 22879 13845 22943
rect 13871 22879 13935 22943
rect 13961 22879 14025 22943
rect 13511 22798 13575 22862
rect 13601 22798 13665 22862
rect 13691 22798 13755 22862
rect 13781 22798 13845 22862
rect 13871 22798 13935 22862
rect 13961 22798 14025 22862
rect 13511 22717 13575 22781
rect 13601 22717 13665 22781
rect 13691 22717 13755 22781
rect 13781 22717 13845 22781
rect 13871 22717 13935 22781
rect 13961 22717 14025 22781
rect 13511 22636 13575 22700
rect 13601 22636 13665 22700
rect 13691 22636 13755 22700
rect 13781 22636 13845 22700
rect 13871 22636 13935 22700
rect 13961 22636 14025 22700
rect 13511 22555 13575 22619
rect 13601 22555 13665 22619
rect 13691 22555 13755 22619
rect 13781 22555 13845 22619
rect 13871 22555 13935 22619
rect 13961 22555 14025 22619
rect 13511 22474 13575 22538
rect 13601 22474 13665 22538
rect 13691 22474 13755 22538
rect 13781 22474 13845 22538
rect 13871 22474 13935 22538
rect 13961 22474 14025 22538
rect 13511 22393 13575 22457
rect 13601 22393 13665 22457
rect 13691 22393 13755 22457
rect 13781 22393 13845 22457
rect 13871 22393 13935 22457
rect 13961 22393 14025 22457
rect 13511 22312 13575 22376
rect 13601 22312 13665 22376
rect 13691 22312 13755 22376
rect 13781 22312 13845 22376
rect 13871 22312 13935 22376
rect 13961 22312 14025 22376
rect 13511 22231 13575 22295
rect 13601 22231 13665 22295
rect 13691 22231 13755 22295
rect 13781 22231 13845 22295
rect 13871 22231 13935 22295
rect 13961 22231 14025 22295
rect 13511 22150 13575 22214
rect 13601 22150 13665 22214
rect 13691 22150 13755 22214
rect 13781 22150 13845 22214
rect 13871 22150 13935 22214
rect 13961 22150 14025 22214
rect 13511 22069 13575 22133
rect 13601 22069 13665 22133
rect 13691 22069 13755 22133
rect 13781 22069 13845 22133
rect 13871 22069 13935 22133
rect 13961 22069 14025 22133
rect 13511 21988 13575 22052
rect 13601 21988 13665 22052
rect 13691 21988 13755 22052
rect 13781 21988 13845 22052
rect 13871 21988 13935 22052
rect 13961 21988 14025 22052
rect 13511 21907 13575 21971
rect 13601 21907 13665 21971
rect 13691 21907 13755 21971
rect 13781 21907 13845 21971
rect 13871 21907 13935 21971
rect 13961 21907 14025 21971
rect 13511 21826 13575 21890
rect 13601 21826 13665 21890
rect 13691 21826 13755 21890
rect 13781 21826 13845 21890
rect 13871 21826 13935 21890
rect 13961 21826 14025 21890
rect 13511 21745 13575 21809
rect 13601 21745 13665 21809
rect 13691 21745 13755 21809
rect 13781 21745 13845 21809
rect 13871 21745 13935 21809
rect 13961 21745 14025 21809
rect 13511 21664 13575 21728
rect 13601 21664 13665 21728
rect 13691 21664 13755 21728
rect 13781 21664 13845 21728
rect 13871 21664 13935 21728
rect 13961 21664 14025 21728
rect 13511 21583 13575 21647
rect 13601 21583 13665 21647
rect 13691 21583 13755 21647
rect 13781 21583 13845 21647
rect 13871 21583 13935 21647
rect 13961 21583 14025 21647
rect 13511 21502 13575 21566
rect 13601 21502 13665 21566
rect 13691 21502 13755 21566
rect 13781 21502 13845 21566
rect 13871 21502 13935 21566
rect 13961 21502 14025 21566
rect 13511 21421 13575 21485
rect 13601 21421 13665 21485
rect 13691 21421 13755 21485
rect 13781 21421 13845 21485
rect 13871 21421 13935 21485
rect 13961 21421 14025 21485
rect 13511 21340 13575 21404
rect 13601 21340 13665 21404
rect 13691 21340 13755 21404
rect 13781 21340 13845 21404
rect 13871 21340 13935 21404
rect 13961 21340 14025 21404
rect 13511 21259 13575 21323
rect 13601 21259 13665 21323
rect 13691 21259 13755 21323
rect 13781 21259 13845 21323
rect 13871 21259 13935 21323
rect 13961 21259 14025 21323
rect 13511 21178 13575 21242
rect 13601 21178 13665 21242
rect 13691 21178 13755 21242
rect 13781 21178 13845 21242
rect 13871 21178 13935 21242
rect 13961 21178 14025 21242
rect 13511 21097 13575 21161
rect 13601 21097 13665 21161
rect 13691 21097 13755 21161
rect 13781 21097 13845 21161
rect 13871 21097 13935 21161
rect 13961 21097 14025 21161
rect 13511 21016 13575 21080
rect 13601 21016 13665 21080
rect 13691 21016 13755 21080
rect 13781 21016 13845 21080
rect 13871 21016 13935 21080
rect 13961 21016 14025 21080
rect 13412 20874 13476 20938
rect 13511 20935 13575 20999
rect 13601 20935 13665 20999
rect 13691 20935 13755 20999
rect 13781 20935 13845 20999
rect 13871 20935 13935 20999
rect 13961 20935 14025 20999
rect 13511 20854 13575 20918
rect 13601 20854 13665 20918
rect 13691 20854 13755 20918
rect 13781 20854 13845 20918
rect 13871 20854 13935 20918
rect 13961 20854 14025 20918
rect 13272 20760 13336 20824
rect 13362 20760 13426 20824
rect 13452 20760 13516 20824
rect 13542 20760 13606 20824
rect 13631 20760 13695 20824
rect 13740 20758 13804 20822
rect 13842 20751 13906 20815
rect 13272 20644 13336 20708
rect 13362 20644 13426 20708
rect 13452 20644 13516 20708
rect 13542 20644 13606 20708
rect 13631 20644 13695 20708
rect 13740 20647 13804 20711
rect 13131 20566 13195 20630
rect 13272 20528 13336 20592
rect 13362 20528 13426 20592
rect 13452 20528 13516 20592
rect 13542 20528 13606 20592
rect 13631 20528 13695 20592
rect 12952 20440 13016 20504
rect 13042 20440 13106 20504
rect 13132 20440 13196 20504
rect 13222 20440 13286 20504
rect 13311 20440 13375 20504
rect 13419 20404 13483 20468
rect 12952 20324 13016 20388
rect 13042 20324 13106 20388
rect 13132 20324 13196 20388
rect 13222 20324 13286 20388
rect 13311 20324 13375 20388
rect 1843 20076 1907 20140
rect 1947 20116 2011 20180
rect 2036 20116 2100 20180
rect 2126 20116 2190 20180
rect 2216 20116 2280 20180
rect 2306 20116 2370 20180
rect 1947 20000 2011 20064
rect 2036 20000 2100 20064
rect 2126 20000 2190 20064
rect 2216 20000 2280 20064
rect 2306 20000 2370 20064
rect 1947 19884 2011 19948
rect 2036 19884 2100 19948
rect 2126 19884 2190 19948
rect 2216 19884 2280 19948
rect 2306 19884 2370 19948
rect 2184 19735 2248 19799
rect 12806 20241 12870 20305
rect 12952 20208 13016 20272
rect 13042 20208 13106 20272
rect 13132 20208 13196 20272
rect 13222 20208 13286 20272
rect 13311 20208 13375 20272
rect 12628 20116 12692 20180
rect 12718 20116 12782 20180
rect 12808 20116 12872 20180
rect 12898 20116 12962 20180
rect 12987 20116 13051 20180
rect 13091 20076 13155 20140
rect 12141 20005 12205 20069
rect 12257 20005 12321 20069
rect 12372 20005 12436 20069
rect 12487 20005 12551 20069
rect 12628 20000 12692 20064
rect 12718 20000 12782 20064
rect 12808 20000 12872 20064
rect 12898 20000 12962 20064
rect 12987 20000 13051 20064
rect 12037 19890 12101 19954
rect 12141 19885 12205 19949
rect 12257 19885 12321 19949
rect 12372 19885 12436 19949
rect 12487 19885 12551 19949
rect 12628 19884 12692 19948
rect 12718 19884 12782 19948
rect 12808 19884 12872 19948
rect 12898 19884 12962 19948
rect 12987 19884 13051 19948
rect 11894 19779 11958 19843
rect 11978 19779 12042 19843
rect 12062 19779 12126 19843
rect 12146 19779 12210 19843
rect 12230 19779 12294 19843
rect 12314 19779 12378 19843
rect 12398 19779 12462 19843
rect 12482 19779 12546 19843
rect 12566 19779 12630 19843
rect 12650 19779 12714 19843
rect 12750 19735 12814 19799
rect 11790 19642 11854 19706
rect 11894 19663 11958 19727
rect 11978 19663 12042 19727
rect 12062 19663 12126 19727
rect 12146 19663 12210 19727
rect 12230 19663 12294 19727
rect 12314 19663 12378 19727
rect 12398 19663 12462 19727
rect 12482 19663 12546 19727
rect 12566 19663 12630 19727
rect 12650 19663 12714 19727
rect 11790 19549 11854 19613
rect 11894 19547 11958 19611
rect 11978 19547 12042 19611
rect 12062 19547 12126 19611
rect 12146 19547 12210 19611
rect 12230 19547 12294 19611
rect 12314 19547 12378 19611
rect 12398 19547 12462 19611
rect 12482 19547 12546 19611
rect 12566 19547 12630 19611
rect 12650 19547 12714 19611
rect 887 3022 2071 3646
rect 12887 3022 14071 3646
<< metal4 >>
rect 2266 34617 2667 34620
rect 2266 34553 2267 34617
rect 2331 34553 2350 34617
rect 2414 34553 2434 34617
rect 2498 34553 2518 34617
rect 2582 34553 2602 34617
rect 2666 34553 2667 34617
rect 2266 34523 2667 34553
rect 2122 34440 2204 34473
rect 2122 34376 2139 34440
rect 2203 34376 2204 34440
rect 2122 34343 2204 34376
rect 2266 34459 2267 34523
rect 2331 34459 2350 34523
rect 2414 34459 2434 34523
rect 2498 34459 2518 34523
rect 2582 34459 2602 34523
rect 2666 34459 2667 34523
rect 2266 34429 2667 34459
rect 2266 34365 2267 34429
rect 2331 34365 2350 34429
rect 2414 34365 2434 34429
rect 2498 34365 2518 34429
rect 2582 34365 2602 34429
rect 2666 34365 2667 34429
rect 2266 34335 2667 34365
rect 1993 34315 2221 34316
rect 1993 34251 1995 34315
rect 2059 34251 2075 34315
rect 2139 34251 2155 34315
rect 2219 34251 2221 34315
rect 1993 34219 2221 34251
rect 1864 34182 1946 34215
rect 1864 34118 1881 34182
rect 1945 34118 1946 34182
rect 1993 34155 1995 34219
rect 2059 34155 2075 34219
rect 2139 34155 2155 34219
rect 2219 34155 2221 34219
rect 1993 34154 2221 34155
rect 2266 34271 2267 34335
rect 2331 34271 2350 34335
rect 2414 34271 2434 34335
rect 2498 34271 2518 34335
rect 2582 34271 2602 34335
rect 2666 34271 2667 34335
rect 2266 34241 2667 34271
rect 2266 34177 2267 34241
rect 2331 34177 2350 34241
rect 2414 34177 2434 34241
rect 2498 34177 2518 34241
rect 2582 34177 2602 34241
rect 2666 34177 2667 34241
rect 1864 34085 1946 34118
rect 2266 34147 2667 34177
rect 2266 34083 2267 34147
rect 2331 34083 2350 34147
rect 2414 34083 2434 34147
rect 2498 34083 2518 34147
rect 2582 34083 2602 34147
rect 2666 34083 2667 34147
rect 2266 34080 2667 34083
rect 12331 34617 12733 34620
rect 12331 34553 12332 34617
rect 12396 34553 12416 34617
rect 12480 34553 12500 34617
rect 12564 34553 12584 34617
rect 12648 34553 12668 34617
rect 12732 34553 12733 34617
rect 12331 34523 12733 34553
rect 12331 34459 12332 34523
rect 12396 34459 12416 34523
rect 12480 34459 12500 34523
rect 12564 34459 12584 34523
rect 12648 34459 12668 34523
rect 12732 34459 12733 34523
rect 12331 34429 12733 34459
rect 12331 34365 12332 34429
rect 12396 34365 12416 34429
rect 12480 34365 12500 34429
rect 12564 34365 12584 34429
rect 12648 34365 12668 34429
rect 12732 34365 12733 34429
rect 12331 34335 12733 34365
rect 12794 34440 12876 34473
rect 12794 34376 12795 34440
rect 12859 34376 12876 34440
rect 12794 34343 12876 34376
rect 12331 34271 12332 34335
rect 12396 34271 12416 34335
rect 12480 34271 12500 34335
rect 12564 34271 12584 34335
rect 12648 34271 12668 34335
rect 12732 34271 12733 34335
rect 12331 34241 12733 34271
rect 12331 34177 12332 34241
rect 12396 34177 12416 34241
rect 12480 34177 12500 34241
rect 12564 34177 12584 34241
rect 12648 34177 12668 34241
rect 12732 34177 12733 34241
rect 12331 34147 12733 34177
rect 12777 34315 13005 34316
rect 12777 34251 12779 34315
rect 12843 34251 12859 34315
rect 12923 34251 12939 34315
rect 13003 34251 13005 34315
rect 12777 34219 13005 34251
rect 12777 34155 12779 34219
rect 12843 34155 12859 34219
rect 12923 34155 12939 34219
rect 13003 34155 13005 34219
rect 12777 34154 13005 34155
rect 13052 34182 13134 34215
rect 12331 34083 12332 34147
rect 12396 34083 12416 34147
rect 12480 34083 12500 34147
rect 12564 34083 12584 34147
rect 12648 34083 12668 34147
rect 12732 34083 12733 34147
rect 13052 34118 13053 34182
rect 13117 34118 13134 34182
rect 13052 34085 13134 34118
rect 12331 34080 12733 34083
rect 1738 34077 2163 34079
rect 1738 34013 1739 34077
rect 1803 34013 1828 34077
rect 1892 34013 1918 34077
rect 1982 34013 2008 34077
rect 2072 34013 2098 34077
rect 2162 34013 2163 34077
rect 12835 34077 13260 34079
rect 1738 33961 2163 34013
rect 1575 33885 1700 33918
rect 1575 33821 1635 33885
rect 1699 33821 1700 33885
rect 1575 33788 1700 33821
rect 1738 33897 1739 33961
rect 1803 33897 1828 33961
rect 1892 33897 1918 33961
rect 1982 33897 2008 33961
rect 2072 33897 2098 33961
rect 2162 33897 2163 33961
rect 2178 34008 2303 34041
rect 2178 33944 2238 34008
rect 2302 33944 2303 34008
rect 2178 33911 2303 33944
rect 12695 34008 12820 34041
rect 12695 33944 12696 34008
rect 12760 33944 12820 34008
rect 12695 33911 12820 33944
rect 12835 34013 12836 34077
rect 12900 34013 12926 34077
rect 12990 34013 13016 34077
rect 13080 34013 13106 34077
rect 13170 34013 13195 34077
rect 13259 34013 13260 34077
rect 12835 33961 13260 34013
rect 1738 33845 2163 33897
rect 1738 33781 1739 33845
rect 1803 33781 1828 33845
rect 1892 33781 1918 33845
rect 1982 33781 2008 33845
rect 2072 33781 2098 33845
rect 2162 33781 2163 33845
rect 1738 33779 2163 33781
rect 12835 33897 12836 33961
rect 12900 33897 12926 33961
rect 12990 33897 13016 33961
rect 13080 33897 13106 33961
rect 13170 33897 13195 33961
rect 13259 33897 13260 33961
rect 12835 33845 13260 33897
rect 12835 33781 12836 33845
rect 12900 33781 12926 33845
rect 12990 33781 13016 33845
rect 13080 33781 13106 33845
rect 13170 33781 13195 33845
rect 13259 33781 13260 33845
rect 13298 33885 13423 33918
rect 13298 33821 13299 33885
rect 13363 33821 13423 33885
rect 13298 33788 13423 33821
rect 12835 33779 13260 33781
rect 1414 33753 1839 33755
rect 13159 33753 13584 33755
rect 1414 33689 1415 33753
rect 1479 33689 1504 33753
rect 1568 33689 1594 33753
rect 1658 33689 1684 33753
rect 1748 33689 1774 33753
rect 1838 33689 1839 33753
rect 1414 33637 1839 33689
rect 1247 33557 1372 33590
rect 1247 33493 1307 33557
rect 1371 33493 1372 33557
rect 1247 33460 1372 33493
rect 1414 33573 1415 33637
rect 1479 33573 1504 33637
rect 1568 33573 1594 33637
rect 1658 33573 1684 33637
rect 1748 33573 1774 33637
rect 1838 33573 1839 33637
rect 1860 33720 1985 33753
rect 1860 33656 1920 33720
rect 1984 33656 1985 33720
rect 1860 33623 1985 33656
rect 13013 33720 13138 33753
rect 13013 33656 13014 33720
rect 13078 33656 13138 33720
rect 13013 33623 13138 33656
rect 13159 33689 13160 33753
rect 13224 33689 13250 33753
rect 13314 33689 13340 33753
rect 13404 33689 13430 33753
rect 13494 33689 13519 33753
rect 13583 33689 13584 33753
rect 13159 33637 13584 33689
rect 1414 33521 1839 33573
rect 1414 33457 1415 33521
rect 1479 33457 1504 33521
rect 1568 33457 1594 33521
rect 1658 33457 1684 33521
rect 1748 33457 1774 33521
rect 1838 33457 1839 33521
rect 1414 33455 1839 33457
rect 13159 33573 13160 33637
rect 13224 33573 13250 33637
rect 13314 33573 13340 33637
rect 13404 33573 13430 33637
rect 13494 33573 13519 33637
rect 13583 33573 13584 33637
rect 13159 33521 13584 33573
rect 13159 33457 13160 33521
rect 13224 33457 13250 33521
rect 13314 33457 13340 33521
rect 13404 33457 13430 33521
rect 13494 33457 13519 33521
rect 13583 33457 13584 33521
rect 13626 33557 13751 33590
rect 13626 33493 13627 33557
rect 13691 33493 13751 33557
rect 13626 33460 13751 33493
rect 13159 33455 13584 33457
rect 1094 33433 1519 33435
rect 1094 33369 1095 33433
rect 1159 33369 1184 33433
rect 1248 33369 1274 33433
rect 1338 33369 1364 33433
rect 1428 33369 1454 33433
rect 1518 33369 1519 33433
rect 13479 33433 13904 33435
rect 1094 33317 1519 33369
rect 1094 33253 1095 33317
rect 1159 33253 1184 33317
rect 1248 33253 1274 33317
rect 1338 33253 1364 33317
rect 1428 33253 1454 33317
rect 1518 33253 1519 33317
rect 1535 33395 1660 33428
rect 1535 33331 1595 33395
rect 1659 33331 1660 33395
rect 1535 33298 1660 33331
rect 13338 33395 13463 33428
rect 13338 33331 13339 33395
rect 13403 33331 13463 33395
rect 13338 33298 13463 33331
rect 13479 33369 13480 33433
rect 13544 33369 13570 33433
rect 13634 33369 13660 33433
rect 13724 33369 13750 33433
rect 13814 33369 13839 33433
rect 13903 33369 13904 33433
rect 13479 33317 13904 33369
rect 1094 33201 1519 33253
rect 1094 33137 1095 33201
rect 1159 33137 1184 33201
rect 1248 33137 1274 33201
rect 1338 33137 1364 33201
rect 1428 33137 1454 33201
rect 1518 33137 1519 33201
rect 1094 33135 1519 33137
rect 13479 33253 13480 33317
rect 13544 33253 13570 33317
rect 13634 33253 13660 33317
rect 13724 33253 13750 33317
rect 13814 33253 13839 33317
rect 13903 33253 13904 33317
rect 13479 33201 13904 33253
rect 13479 33137 13480 33201
rect 13544 33137 13570 33201
rect 13634 33137 13660 33201
rect 13724 33137 13750 33201
rect 13814 33137 13839 33201
rect 13903 33137 13904 33201
rect 13479 33135 13904 33137
rect 968 33108 1492 33109
rect 968 33044 973 33108
rect 1037 33044 1063 33108
rect 1127 33044 1153 33108
rect 1217 33044 1243 33108
rect 1307 33044 1333 33108
rect 1397 33044 1423 33108
rect 1487 33044 1492 33108
rect 968 33028 1492 33044
rect 968 32964 973 33028
rect 1037 32964 1063 33028
rect 1127 32964 1153 33028
rect 1217 32964 1243 33028
rect 1307 32964 1333 33028
rect 1397 32964 1423 33028
rect 1487 32964 1492 33028
rect 968 32948 1492 32964
rect 968 32884 973 32948
rect 1037 32884 1063 32948
rect 1127 32884 1153 32948
rect 1217 32884 1243 32948
rect 1307 32884 1333 32948
rect 1397 32884 1423 32948
rect 1487 32884 1492 32948
rect 968 32868 1492 32884
rect 968 32804 973 32868
rect 1037 32804 1063 32868
rect 1127 32804 1153 32868
rect 1217 32804 1243 32868
rect 1307 32804 1333 32868
rect 1397 32804 1423 32868
rect 1487 32804 1492 32868
rect 968 32788 1492 32804
rect 968 32724 973 32788
rect 1037 32724 1063 32788
rect 1127 32724 1153 32788
rect 1217 32724 1243 32788
rect 1307 32724 1333 32788
rect 1397 32724 1423 32788
rect 1487 32724 1492 32788
rect 968 32708 1492 32724
rect 968 32644 973 32708
rect 1037 32644 1063 32708
rect 1127 32644 1153 32708
rect 1217 32644 1243 32708
rect 1307 32644 1333 32708
rect 1397 32644 1423 32708
rect 1487 32644 1492 32708
rect 968 32628 1492 32644
rect 968 32564 973 32628
rect 1037 32564 1063 32628
rect 1127 32564 1153 32628
rect 1217 32564 1243 32628
rect 1307 32564 1333 32628
rect 1397 32564 1423 32628
rect 1487 32564 1492 32628
rect 968 32548 1492 32564
rect 968 32484 973 32548
rect 1037 32484 1063 32548
rect 1127 32484 1153 32548
rect 1217 32484 1243 32548
rect 1307 32484 1333 32548
rect 1397 32484 1423 32548
rect 1487 32484 1492 32548
rect 968 32468 1492 32484
rect 968 32404 973 32468
rect 1037 32404 1063 32468
rect 1127 32404 1153 32468
rect 1217 32404 1243 32468
rect 1307 32404 1333 32468
rect 1397 32404 1423 32468
rect 1487 32404 1492 32468
rect 968 32388 1492 32404
rect 968 32324 973 32388
rect 1037 32324 1063 32388
rect 1127 32324 1153 32388
rect 1217 32324 1243 32388
rect 1307 32324 1333 32388
rect 1397 32324 1423 32388
rect 1487 32324 1492 32388
rect 968 32308 1492 32324
rect 968 32244 973 32308
rect 1037 32244 1063 32308
rect 1127 32244 1153 32308
rect 1217 32244 1243 32308
rect 1307 32244 1333 32308
rect 1397 32244 1423 32308
rect 1487 32244 1492 32308
rect 968 32228 1492 32244
rect 968 32164 973 32228
rect 1037 32164 1063 32228
rect 1127 32164 1153 32228
rect 1217 32164 1243 32228
rect 1307 32164 1333 32228
rect 1397 32164 1423 32228
rect 1487 32164 1492 32228
rect 968 32148 1492 32164
rect 968 32084 973 32148
rect 1037 32084 1063 32148
rect 1127 32084 1153 32148
rect 1217 32084 1243 32148
rect 1307 32084 1333 32148
rect 1397 32084 1423 32148
rect 1487 32084 1492 32148
rect 968 32068 1492 32084
rect 968 32004 973 32068
rect 1037 32004 1063 32068
rect 1127 32004 1153 32068
rect 1217 32004 1243 32068
rect 1307 32004 1333 32068
rect 1397 32004 1423 32068
rect 1487 32004 1492 32068
rect 968 31988 1492 32004
rect 968 31924 973 31988
rect 1037 31924 1063 31988
rect 1127 31924 1153 31988
rect 1217 31924 1243 31988
rect 1307 31924 1333 31988
rect 1397 31924 1423 31988
rect 1487 31924 1492 31988
rect 968 31908 1492 31924
rect 968 31844 973 31908
rect 1037 31844 1063 31908
rect 1127 31844 1153 31908
rect 1217 31844 1243 31908
rect 1307 31844 1333 31908
rect 1397 31844 1423 31908
rect 1487 31844 1492 31908
rect 968 31828 1492 31844
rect 968 31764 973 31828
rect 1037 31764 1063 31828
rect 1127 31764 1153 31828
rect 1217 31764 1243 31828
rect 1307 31764 1333 31828
rect 1397 31764 1423 31828
rect 1487 31764 1492 31828
rect 968 31748 1492 31764
rect 968 31684 973 31748
rect 1037 31684 1063 31748
rect 1127 31684 1153 31748
rect 1217 31684 1243 31748
rect 1307 31684 1333 31748
rect 1397 31684 1423 31748
rect 1487 31684 1492 31748
rect 968 31668 1492 31684
rect 968 31604 973 31668
rect 1037 31604 1063 31668
rect 1127 31604 1153 31668
rect 1217 31604 1243 31668
rect 1307 31604 1333 31668
rect 1397 31604 1423 31668
rect 1487 31604 1492 31668
rect 968 31588 1492 31604
rect 968 31524 973 31588
rect 1037 31524 1063 31588
rect 1127 31524 1153 31588
rect 1217 31524 1243 31588
rect 1307 31524 1333 31588
rect 1397 31524 1423 31588
rect 1487 31524 1492 31588
rect 968 31508 1492 31524
rect 968 31444 973 31508
rect 1037 31444 1063 31508
rect 1127 31444 1153 31508
rect 1217 31444 1243 31508
rect 1307 31444 1333 31508
rect 1397 31444 1423 31508
rect 1487 31444 1492 31508
rect 968 31428 1492 31444
rect 968 31364 973 31428
rect 1037 31364 1063 31428
rect 1127 31364 1153 31428
rect 1217 31364 1243 31428
rect 1307 31364 1333 31428
rect 1397 31364 1423 31428
rect 1487 31364 1492 31428
rect 968 31348 1492 31364
rect 968 31284 973 31348
rect 1037 31284 1063 31348
rect 1127 31284 1153 31348
rect 1217 31284 1243 31348
rect 1307 31284 1333 31348
rect 1397 31284 1423 31348
rect 1487 31284 1492 31348
rect 968 31268 1492 31284
rect 968 31204 973 31268
rect 1037 31204 1063 31268
rect 1127 31204 1153 31268
rect 1217 31204 1243 31268
rect 1307 31204 1333 31268
rect 1397 31204 1423 31268
rect 1487 31204 1492 31268
rect 968 31188 1492 31204
rect 968 31124 973 31188
rect 1037 31124 1063 31188
rect 1127 31124 1153 31188
rect 1217 31124 1243 31188
rect 1307 31124 1333 31188
rect 1397 31124 1423 31188
rect 1487 31124 1492 31188
rect 968 31108 1492 31124
rect 968 31044 973 31108
rect 1037 31044 1063 31108
rect 1127 31044 1153 31108
rect 1217 31044 1243 31108
rect 1307 31044 1333 31108
rect 1397 31044 1423 31108
rect 1487 31044 1492 31108
rect 968 31028 1492 31044
rect 968 30964 973 31028
rect 1037 30964 1063 31028
rect 1127 30964 1153 31028
rect 1217 30964 1243 31028
rect 1307 30964 1333 31028
rect 1397 30964 1423 31028
rect 1487 30964 1492 31028
rect 968 30948 1492 30964
rect 968 30884 973 30948
rect 1037 30884 1063 30948
rect 1127 30884 1153 30948
rect 1217 30884 1243 30948
rect 1307 30884 1333 30948
rect 1397 30884 1423 30948
rect 1487 30884 1492 30948
rect 968 30868 1492 30884
rect 968 30804 973 30868
rect 1037 30804 1063 30868
rect 1127 30804 1153 30868
rect 1217 30804 1243 30868
rect 1307 30804 1333 30868
rect 1397 30804 1423 30868
rect 1487 30804 1492 30868
rect 968 30788 1492 30804
rect 968 30724 973 30788
rect 1037 30724 1063 30788
rect 1127 30724 1153 30788
rect 1217 30724 1243 30788
rect 1307 30724 1333 30788
rect 1397 30724 1423 30788
rect 1487 30724 1492 30788
rect 968 30708 1492 30724
rect 968 30644 973 30708
rect 1037 30644 1063 30708
rect 1127 30644 1153 30708
rect 1217 30644 1243 30708
rect 1307 30644 1333 30708
rect 1397 30644 1423 30708
rect 1487 30644 1492 30708
rect 968 30628 1492 30644
rect 968 30564 973 30628
rect 1037 30564 1063 30628
rect 1127 30564 1153 30628
rect 1217 30564 1243 30628
rect 1307 30564 1333 30628
rect 1397 30564 1423 30628
rect 1487 30564 1492 30628
rect 968 30548 1492 30564
rect 968 30484 973 30548
rect 1037 30484 1063 30548
rect 1127 30484 1153 30548
rect 1217 30484 1243 30548
rect 1307 30484 1333 30548
rect 1397 30484 1423 30548
rect 1487 30484 1492 30548
rect 968 30468 1492 30484
rect 968 30404 973 30468
rect 1037 30404 1063 30468
rect 1127 30404 1153 30468
rect 1217 30404 1243 30468
rect 1307 30404 1333 30468
rect 1397 30404 1423 30468
rect 1487 30404 1492 30468
rect 968 30388 1492 30404
rect 968 30324 973 30388
rect 1037 30324 1063 30388
rect 1127 30324 1153 30388
rect 1217 30324 1243 30388
rect 1307 30324 1333 30388
rect 1397 30324 1423 30388
rect 1487 30324 1492 30388
rect 968 30308 1492 30324
rect 968 30244 973 30308
rect 1037 30244 1063 30308
rect 1127 30244 1153 30308
rect 1217 30244 1243 30308
rect 1307 30244 1333 30308
rect 1397 30244 1423 30308
rect 1487 30244 1492 30308
rect 968 30228 1492 30244
rect 968 30164 973 30228
rect 1037 30164 1063 30228
rect 1127 30164 1153 30228
rect 1217 30164 1243 30228
rect 1307 30164 1333 30228
rect 1397 30164 1423 30228
rect 1487 30164 1492 30228
rect 968 30148 1492 30164
rect 968 30084 973 30148
rect 1037 30084 1063 30148
rect 1127 30084 1153 30148
rect 1217 30084 1243 30148
rect 1307 30084 1333 30148
rect 1397 30084 1423 30148
rect 1487 30084 1492 30148
rect 968 30068 1492 30084
rect 968 30004 973 30068
rect 1037 30004 1063 30068
rect 1127 30004 1153 30068
rect 1217 30004 1243 30068
rect 1307 30004 1333 30068
rect 1397 30004 1423 30068
rect 1487 30004 1492 30068
rect 968 29988 1492 30004
rect 968 29924 973 29988
rect 1037 29924 1063 29988
rect 1127 29924 1153 29988
rect 1217 29924 1243 29988
rect 1307 29924 1333 29988
rect 1397 29924 1423 29988
rect 1487 29924 1492 29988
rect 968 29908 1492 29924
rect 968 29844 973 29908
rect 1037 29844 1063 29908
rect 1127 29844 1153 29908
rect 1217 29844 1243 29908
rect 1307 29844 1333 29908
rect 1397 29844 1423 29908
rect 1487 29844 1492 29908
rect 968 29828 1492 29844
rect 968 29764 973 29828
rect 1037 29764 1063 29828
rect 1127 29764 1153 29828
rect 1217 29764 1243 29828
rect 1307 29764 1333 29828
rect 1397 29764 1423 29828
rect 1487 29764 1492 29828
rect 968 29748 1492 29764
rect 968 29684 973 29748
rect 1037 29684 1063 29748
rect 1127 29684 1153 29748
rect 1217 29684 1243 29748
rect 1307 29684 1333 29748
rect 1397 29684 1423 29748
rect 1487 29684 1492 29748
rect 968 29668 1492 29684
rect 968 29604 973 29668
rect 1037 29604 1063 29668
rect 1127 29604 1153 29668
rect 1217 29604 1243 29668
rect 1307 29604 1333 29668
rect 1397 29604 1423 29668
rect 1487 29604 1492 29668
rect 968 29588 1492 29604
rect 968 29524 973 29588
rect 1037 29524 1063 29588
rect 1127 29524 1153 29588
rect 1217 29524 1243 29588
rect 1307 29524 1333 29588
rect 1397 29524 1423 29588
rect 1487 29524 1492 29588
rect 968 29508 1492 29524
rect 968 29444 973 29508
rect 1037 29444 1063 29508
rect 1127 29444 1153 29508
rect 1217 29444 1243 29508
rect 1307 29444 1333 29508
rect 1397 29444 1423 29508
rect 1487 29444 1492 29508
rect 968 29428 1492 29444
rect 968 29364 973 29428
rect 1037 29364 1063 29428
rect 1127 29364 1153 29428
rect 1217 29364 1243 29428
rect 1307 29364 1333 29428
rect 1397 29364 1423 29428
rect 1487 29364 1492 29428
rect 968 29348 1492 29364
rect 968 29284 973 29348
rect 1037 29284 1063 29348
rect 1127 29284 1153 29348
rect 1217 29284 1243 29348
rect 1307 29284 1333 29348
rect 1397 29284 1423 29348
rect 1487 29284 1492 29348
rect 968 29268 1492 29284
rect 968 29204 973 29268
rect 1037 29204 1063 29268
rect 1127 29204 1153 29268
rect 1217 29204 1243 29268
rect 1307 29204 1333 29268
rect 1397 29204 1423 29268
rect 1487 29204 1492 29268
rect 968 29188 1492 29204
rect 968 29124 973 29188
rect 1037 29124 1063 29188
rect 1127 29124 1153 29188
rect 1217 29124 1243 29188
rect 1307 29124 1333 29188
rect 1397 29124 1423 29188
rect 1487 29124 1492 29188
rect 968 29108 1492 29124
rect 968 29044 973 29108
rect 1037 29044 1063 29108
rect 1127 29044 1153 29108
rect 1217 29044 1243 29108
rect 1307 29044 1333 29108
rect 1397 29044 1423 29108
rect 1487 29044 1492 29108
rect 968 29028 1492 29044
rect 968 28964 973 29028
rect 1037 28964 1063 29028
rect 1127 28964 1153 29028
rect 1217 28964 1243 29028
rect 1307 28964 1333 29028
rect 1397 28964 1423 29028
rect 1487 28964 1492 29028
rect 968 28948 1492 28964
rect 968 28884 973 28948
rect 1037 28884 1063 28948
rect 1127 28884 1153 28948
rect 1217 28884 1243 28948
rect 1307 28884 1333 28948
rect 1397 28884 1423 28948
rect 1487 28884 1492 28948
rect 968 28868 1492 28884
rect 968 28804 973 28868
rect 1037 28804 1063 28868
rect 1127 28804 1153 28868
rect 1217 28804 1243 28868
rect 1307 28804 1333 28868
rect 1397 28804 1423 28868
rect 1487 28804 1492 28868
rect 968 28788 1492 28804
rect 968 28724 973 28788
rect 1037 28724 1063 28788
rect 1127 28724 1153 28788
rect 1217 28724 1243 28788
rect 1307 28724 1333 28788
rect 1397 28724 1423 28788
rect 1487 28724 1492 28788
rect 968 28708 1492 28724
rect 968 28644 973 28708
rect 1037 28644 1063 28708
rect 1127 28644 1153 28708
rect 1217 28644 1243 28708
rect 1307 28644 1333 28708
rect 1397 28644 1423 28708
rect 1487 28644 1492 28708
rect 968 28628 1492 28644
rect 968 28564 973 28628
rect 1037 28564 1063 28628
rect 1127 28564 1153 28628
rect 1217 28564 1243 28628
rect 1307 28564 1333 28628
rect 1397 28564 1423 28628
rect 1487 28564 1492 28628
rect 968 28548 1492 28564
rect 968 28484 973 28548
rect 1037 28484 1063 28548
rect 1127 28484 1153 28548
rect 1217 28484 1243 28548
rect 1307 28484 1333 28548
rect 1397 28484 1423 28548
rect 1487 28484 1492 28548
rect 968 28468 1492 28484
rect 968 28404 973 28468
rect 1037 28404 1063 28468
rect 1127 28404 1153 28468
rect 1217 28404 1243 28468
rect 1307 28404 1333 28468
rect 1397 28404 1423 28468
rect 1487 28404 1492 28468
rect 968 28388 1492 28404
rect 968 28324 973 28388
rect 1037 28324 1063 28388
rect 1127 28324 1153 28388
rect 1217 28324 1243 28388
rect 1307 28324 1333 28388
rect 1397 28324 1423 28388
rect 1487 28324 1492 28388
rect 968 28308 1492 28324
rect 968 28244 973 28308
rect 1037 28244 1063 28308
rect 1127 28244 1153 28308
rect 1217 28244 1243 28308
rect 1307 28244 1333 28308
rect 1397 28244 1423 28308
rect 1487 28244 1492 28308
rect 968 28228 1492 28244
rect 968 28164 973 28228
rect 1037 28164 1063 28228
rect 1127 28164 1153 28228
rect 1217 28164 1243 28228
rect 1307 28164 1333 28228
rect 1397 28164 1423 28228
rect 1487 28164 1492 28228
rect 968 28148 1492 28164
rect 968 28084 973 28148
rect 1037 28084 1063 28148
rect 1127 28084 1153 28148
rect 1217 28084 1243 28148
rect 1307 28084 1333 28148
rect 1397 28084 1423 28148
rect 1487 28084 1492 28148
rect 968 28068 1492 28084
rect 968 28004 973 28068
rect 1037 28004 1063 28068
rect 1127 28004 1153 28068
rect 1217 28004 1243 28068
rect 1307 28004 1333 28068
rect 1397 28004 1423 28068
rect 1487 28004 1492 28068
rect 968 27988 1492 28004
rect 968 27924 973 27988
rect 1037 27924 1063 27988
rect 1127 27924 1153 27988
rect 1217 27924 1243 27988
rect 1307 27924 1333 27988
rect 1397 27924 1423 27988
rect 1487 27924 1492 27988
rect 968 27908 1492 27924
rect 968 27844 973 27908
rect 1037 27844 1063 27908
rect 1127 27844 1153 27908
rect 1217 27844 1243 27908
rect 1307 27844 1333 27908
rect 1397 27844 1423 27908
rect 1487 27844 1492 27908
rect 968 27828 1492 27844
rect 968 27764 973 27828
rect 1037 27764 1063 27828
rect 1127 27764 1153 27828
rect 1217 27764 1243 27828
rect 1307 27764 1333 27828
rect 1397 27764 1423 27828
rect 1487 27764 1492 27828
rect 968 27748 1492 27764
rect 968 27684 973 27748
rect 1037 27684 1063 27748
rect 1127 27684 1153 27748
rect 1217 27684 1243 27748
rect 1307 27684 1333 27748
rect 1397 27684 1423 27748
rect 1487 27684 1492 27748
rect 968 27668 1492 27684
rect 968 27604 973 27668
rect 1037 27604 1063 27668
rect 1127 27604 1153 27668
rect 1217 27604 1243 27668
rect 1307 27604 1333 27668
rect 1397 27604 1423 27668
rect 1487 27604 1492 27668
rect 968 27588 1492 27604
rect 968 27524 973 27588
rect 1037 27524 1063 27588
rect 1127 27524 1153 27588
rect 1217 27524 1243 27588
rect 1307 27524 1333 27588
rect 1397 27524 1423 27588
rect 1487 27524 1492 27588
rect 968 27508 1492 27524
rect 968 27444 973 27508
rect 1037 27444 1063 27508
rect 1127 27444 1153 27508
rect 1217 27444 1243 27508
rect 1307 27444 1333 27508
rect 1397 27444 1423 27508
rect 1487 27444 1492 27508
rect 968 27428 1492 27444
rect 968 27364 973 27428
rect 1037 27364 1063 27428
rect 1127 27364 1153 27428
rect 1217 27364 1243 27428
rect 1307 27364 1333 27428
rect 1397 27364 1423 27428
rect 1487 27364 1492 27428
rect 968 27348 1492 27364
rect 968 27284 973 27348
rect 1037 27284 1063 27348
rect 1127 27284 1153 27348
rect 1217 27284 1243 27348
rect 1307 27284 1333 27348
rect 1397 27284 1423 27348
rect 1487 27284 1492 27348
rect 968 27268 1492 27284
rect 968 27204 973 27268
rect 1037 27204 1063 27268
rect 1127 27204 1153 27268
rect 1217 27204 1243 27268
rect 1307 27204 1333 27268
rect 1397 27204 1423 27268
rect 1487 27204 1492 27268
rect 968 27188 1492 27204
rect 968 27124 973 27188
rect 1037 27124 1063 27188
rect 1127 27124 1153 27188
rect 1217 27124 1243 27188
rect 1307 27124 1333 27188
rect 1397 27124 1423 27188
rect 1487 27124 1492 27188
rect 968 27108 1492 27124
rect 968 27044 973 27108
rect 1037 27044 1063 27108
rect 1127 27044 1153 27108
rect 1217 27044 1243 27108
rect 1307 27044 1333 27108
rect 1397 27044 1423 27108
rect 1487 27044 1492 27108
rect 968 27028 1492 27044
rect 968 26964 973 27028
rect 1037 26964 1063 27028
rect 1127 26964 1153 27028
rect 1217 26964 1243 27028
rect 1307 26964 1333 27028
rect 1397 26964 1423 27028
rect 1487 26964 1492 27028
rect 968 26948 1492 26964
rect 968 26884 973 26948
rect 1037 26884 1063 26948
rect 1127 26884 1153 26948
rect 1217 26884 1243 26948
rect 1307 26884 1333 26948
rect 1397 26884 1423 26948
rect 1487 26884 1492 26948
rect 968 26868 1492 26884
rect 968 26804 973 26868
rect 1037 26804 1063 26868
rect 1127 26804 1153 26868
rect 1217 26804 1243 26868
rect 1307 26804 1333 26868
rect 1397 26804 1423 26868
rect 1487 26804 1492 26868
rect 968 26788 1492 26804
rect 968 26724 973 26788
rect 1037 26724 1063 26788
rect 1127 26724 1153 26788
rect 1217 26724 1243 26788
rect 1307 26724 1333 26788
rect 1397 26724 1423 26788
rect 1487 26724 1492 26788
rect 968 26708 1492 26724
rect 968 26644 973 26708
rect 1037 26644 1063 26708
rect 1127 26644 1153 26708
rect 1217 26644 1243 26708
rect 1307 26644 1333 26708
rect 1397 26644 1423 26708
rect 1487 26644 1492 26708
rect 968 26628 1492 26644
rect 968 26564 973 26628
rect 1037 26564 1063 26628
rect 1127 26564 1153 26628
rect 1217 26564 1243 26628
rect 1307 26564 1333 26628
rect 1397 26564 1423 26628
rect 1487 26564 1492 26628
rect 968 26548 1492 26564
rect 968 26484 973 26548
rect 1037 26484 1063 26548
rect 1127 26484 1153 26548
rect 1217 26484 1243 26548
rect 1307 26484 1333 26548
rect 1397 26484 1423 26548
rect 1487 26484 1492 26548
rect 968 26468 1492 26484
rect 968 26404 973 26468
rect 1037 26404 1063 26468
rect 1127 26404 1153 26468
rect 1217 26404 1243 26468
rect 1307 26404 1333 26468
rect 1397 26404 1423 26468
rect 1487 26404 1492 26468
rect 968 26388 1492 26404
rect 968 26324 973 26388
rect 1037 26324 1063 26388
rect 1127 26324 1153 26388
rect 1217 26324 1243 26388
rect 1307 26324 1333 26388
rect 1397 26324 1423 26388
rect 1487 26324 1492 26388
rect 968 26308 1492 26324
rect 968 26244 973 26308
rect 1037 26244 1063 26308
rect 1127 26244 1153 26308
rect 1217 26244 1243 26308
rect 1307 26244 1333 26308
rect 1397 26244 1423 26308
rect 1487 26244 1492 26308
rect 968 26228 1492 26244
rect 968 26164 973 26228
rect 1037 26164 1063 26228
rect 1127 26164 1153 26228
rect 1217 26164 1243 26228
rect 1307 26164 1333 26228
rect 1397 26164 1423 26228
rect 1487 26164 1492 26228
rect 968 26148 1492 26164
rect 968 26084 973 26148
rect 1037 26084 1063 26148
rect 1127 26084 1153 26148
rect 1217 26084 1243 26148
rect 1307 26084 1333 26148
rect 1397 26084 1423 26148
rect 1487 26084 1492 26148
rect 968 26068 1492 26084
rect 968 26004 973 26068
rect 1037 26004 1063 26068
rect 1127 26004 1153 26068
rect 1217 26004 1243 26068
rect 1307 26004 1333 26068
rect 1397 26004 1423 26068
rect 1487 26004 1492 26068
rect 968 25988 1492 26004
rect 968 25924 973 25988
rect 1037 25924 1063 25988
rect 1127 25924 1153 25988
rect 1217 25924 1243 25988
rect 1307 25924 1333 25988
rect 1397 25924 1423 25988
rect 1487 25924 1492 25988
rect 968 25908 1492 25924
rect 968 25844 973 25908
rect 1037 25844 1063 25908
rect 1127 25844 1153 25908
rect 1217 25844 1243 25908
rect 1307 25844 1333 25908
rect 1397 25844 1423 25908
rect 1487 25844 1492 25908
rect 968 25828 1492 25844
rect 968 25764 973 25828
rect 1037 25764 1063 25828
rect 1127 25764 1153 25828
rect 1217 25764 1243 25828
rect 1307 25764 1333 25828
rect 1397 25764 1423 25828
rect 1487 25764 1492 25828
rect 968 25748 1492 25764
rect 968 25684 973 25748
rect 1037 25684 1063 25748
rect 1127 25684 1153 25748
rect 1217 25684 1243 25748
rect 1307 25684 1333 25748
rect 1397 25684 1423 25748
rect 1487 25684 1492 25748
rect 968 25668 1492 25684
rect 968 25604 973 25668
rect 1037 25604 1063 25668
rect 1127 25604 1153 25668
rect 1217 25604 1243 25668
rect 1307 25604 1333 25668
rect 1397 25604 1423 25668
rect 1487 25604 1492 25668
rect 968 25588 1492 25604
rect 968 25524 973 25588
rect 1037 25524 1063 25588
rect 1127 25524 1153 25588
rect 1217 25524 1243 25588
rect 1307 25524 1333 25588
rect 1397 25524 1423 25588
rect 1487 25524 1492 25588
rect 968 25508 1492 25524
rect 968 25444 973 25508
rect 1037 25444 1063 25508
rect 1127 25444 1153 25508
rect 1217 25444 1243 25508
rect 1307 25444 1333 25508
rect 1397 25444 1423 25508
rect 1487 25444 1492 25508
rect 968 25428 1492 25444
rect 968 25364 973 25428
rect 1037 25364 1063 25428
rect 1127 25364 1153 25428
rect 1217 25364 1243 25428
rect 1307 25364 1333 25428
rect 1397 25364 1423 25428
rect 1487 25364 1492 25428
rect 968 25348 1492 25364
rect 968 25284 973 25348
rect 1037 25284 1063 25348
rect 1127 25284 1153 25348
rect 1217 25284 1243 25348
rect 1307 25284 1333 25348
rect 1397 25284 1423 25348
rect 1487 25284 1492 25348
rect 968 25268 1492 25284
rect 968 25204 973 25268
rect 1037 25204 1063 25268
rect 1127 25204 1153 25268
rect 1217 25204 1243 25268
rect 1307 25204 1333 25268
rect 1397 25204 1423 25268
rect 1487 25204 1492 25268
rect 968 25188 1492 25204
rect 968 25124 973 25188
rect 1037 25124 1063 25188
rect 1127 25124 1153 25188
rect 1217 25124 1243 25188
rect 1307 25124 1333 25188
rect 1397 25124 1423 25188
rect 1487 25124 1492 25188
rect 968 25108 1492 25124
rect 968 25044 973 25108
rect 1037 25044 1063 25108
rect 1127 25044 1153 25108
rect 1217 25044 1243 25108
rect 1307 25044 1333 25108
rect 1397 25044 1423 25108
rect 1487 25044 1492 25108
rect 968 25028 1492 25044
rect 968 24964 973 25028
rect 1037 24964 1063 25028
rect 1127 24964 1153 25028
rect 1217 24964 1243 25028
rect 1307 24964 1333 25028
rect 1397 24964 1423 25028
rect 1487 24964 1492 25028
rect 968 24948 1492 24964
rect 968 24884 973 24948
rect 1037 24884 1063 24948
rect 1127 24884 1153 24948
rect 1217 24884 1243 24948
rect 1307 24884 1333 24948
rect 1397 24884 1423 24948
rect 1487 24884 1492 24948
rect 968 24868 1492 24884
rect 968 24804 973 24868
rect 1037 24804 1063 24868
rect 1127 24804 1153 24868
rect 1217 24804 1243 24868
rect 1307 24804 1333 24868
rect 1397 24804 1423 24868
rect 1487 24804 1492 24868
rect 968 24788 1492 24804
rect 968 24724 973 24788
rect 1037 24724 1063 24788
rect 1127 24724 1153 24788
rect 1217 24724 1243 24788
rect 1307 24724 1333 24788
rect 1397 24724 1423 24788
rect 1487 24724 1492 24788
rect 968 24708 1492 24724
rect 968 24644 973 24708
rect 1037 24644 1063 24708
rect 1127 24644 1153 24708
rect 1217 24644 1243 24708
rect 1307 24644 1333 24708
rect 1397 24644 1423 24708
rect 1487 24644 1492 24708
rect 968 24628 1492 24644
rect 968 24564 973 24628
rect 1037 24564 1063 24628
rect 1127 24564 1153 24628
rect 1217 24564 1243 24628
rect 1307 24564 1333 24628
rect 1397 24564 1423 24628
rect 1487 24564 1492 24628
rect 968 24548 1492 24564
rect 968 24484 973 24548
rect 1037 24484 1063 24548
rect 1127 24484 1153 24548
rect 1217 24484 1243 24548
rect 1307 24484 1333 24548
rect 1397 24484 1423 24548
rect 1487 24484 1492 24548
rect 968 24468 1492 24484
rect 968 24404 973 24468
rect 1037 24404 1063 24468
rect 1127 24404 1153 24468
rect 1217 24404 1243 24468
rect 1307 24404 1333 24468
rect 1397 24404 1423 24468
rect 1487 24404 1492 24468
rect 968 24388 1492 24404
rect 968 24324 973 24388
rect 1037 24324 1063 24388
rect 1127 24324 1153 24388
rect 1217 24324 1243 24388
rect 1307 24324 1333 24388
rect 1397 24324 1423 24388
rect 1487 24324 1492 24388
rect 968 24308 1492 24324
rect 968 24244 973 24308
rect 1037 24244 1063 24308
rect 1127 24244 1153 24308
rect 1217 24244 1243 24308
rect 1307 24244 1333 24308
rect 1397 24244 1423 24308
rect 1487 24244 1492 24308
rect 968 24228 1492 24244
rect 968 24164 973 24228
rect 1037 24164 1063 24228
rect 1127 24164 1153 24228
rect 1217 24164 1243 24228
rect 1307 24164 1333 24228
rect 1397 24164 1423 24228
rect 1487 24164 1492 24228
rect 968 24148 1492 24164
rect 968 24084 973 24148
rect 1037 24084 1063 24148
rect 1127 24084 1153 24148
rect 1217 24084 1243 24148
rect 1307 24084 1333 24148
rect 1397 24084 1423 24148
rect 1487 24084 1492 24148
rect 968 24068 1492 24084
rect 968 24004 973 24068
rect 1037 24004 1063 24068
rect 1127 24004 1153 24068
rect 1217 24004 1243 24068
rect 1307 24004 1333 24068
rect 1397 24004 1423 24068
rect 1487 24004 1492 24068
rect 968 23988 1492 24004
rect 968 23924 973 23988
rect 1037 23924 1063 23988
rect 1127 23924 1153 23988
rect 1217 23924 1243 23988
rect 1307 23924 1333 23988
rect 1397 23924 1423 23988
rect 1487 23924 1492 23988
rect 968 23908 1492 23924
rect 968 23844 973 23908
rect 1037 23844 1063 23908
rect 1127 23844 1153 23908
rect 1217 23844 1243 23908
rect 1307 23844 1333 23908
rect 1397 23844 1423 23908
rect 1487 23844 1492 23908
rect 968 23828 1492 23844
rect 968 23764 973 23828
rect 1037 23764 1063 23828
rect 1127 23764 1153 23828
rect 1217 23764 1243 23828
rect 1307 23764 1333 23828
rect 1397 23764 1423 23828
rect 1487 23764 1492 23828
rect 968 23748 1492 23764
rect 968 23684 973 23748
rect 1037 23684 1063 23748
rect 1127 23684 1153 23748
rect 1217 23684 1243 23748
rect 1307 23684 1333 23748
rect 1397 23684 1423 23748
rect 1487 23684 1492 23748
rect 968 23668 1492 23684
rect 968 23604 973 23668
rect 1037 23604 1063 23668
rect 1127 23604 1153 23668
rect 1217 23604 1243 23668
rect 1307 23604 1333 23668
rect 1397 23604 1423 23668
rect 1487 23604 1492 23668
rect 968 23588 1492 23604
rect 968 23524 973 23588
rect 1037 23524 1063 23588
rect 1127 23524 1153 23588
rect 1217 23524 1243 23588
rect 1307 23524 1333 23588
rect 1397 23524 1423 23588
rect 1487 23524 1492 23588
rect 968 23508 1492 23524
rect 968 23444 973 23508
rect 1037 23444 1063 23508
rect 1127 23444 1153 23508
rect 1217 23444 1243 23508
rect 1307 23444 1333 23508
rect 1397 23444 1423 23508
rect 1487 23444 1492 23508
rect 968 23428 1492 23444
rect 968 23364 973 23428
rect 1037 23364 1063 23428
rect 1127 23364 1153 23428
rect 1217 23364 1243 23428
rect 1307 23364 1333 23428
rect 1397 23364 1423 23428
rect 1487 23364 1492 23428
rect 968 23348 1492 23364
rect 968 23284 973 23348
rect 1037 23284 1063 23348
rect 1127 23284 1153 23348
rect 1217 23284 1243 23348
rect 1307 23284 1333 23348
rect 1397 23284 1423 23348
rect 1487 23284 1492 23348
rect 968 23267 1492 23284
rect 968 23203 973 23267
rect 1037 23203 1063 23267
rect 1127 23203 1153 23267
rect 1217 23203 1243 23267
rect 1307 23203 1333 23267
rect 1397 23203 1423 23267
rect 1487 23203 1492 23267
rect 968 23186 1492 23203
rect 968 23122 973 23186
rect 1037 23122 1063 23186
rect 1127 23122 1153 23186
rect 1217 23122 1243 23186
rect 1307 23122 1333 23186
rect 1397 23122 1423 23186
rect 1487 23122 1492 23186
rect 968 23105 1492 23122
rect 968 23041 973 23105
rect 1037 23041 1063 23105
rect 1127 23041 1153 23105
rect 1217 23041 1243 23105
rect 1307 23041 1333 23105
rect 1397 23041 1423 23105
rect 1487 23041 1492 23105
rect 968 23024 1492 23041
rect 968 22960 973 23024
rect 1037 22960 1063 23024
rect 1127 22960 1153 23024
rect 1217 22960 1243 23024
rect 1307 22960 1333 23024
rect 1397 22960 1423 23024
rect 1487 22960 1492 23024
rect 968 22943 1492 22960
rect 968 22879 973 22943
rect 1037 22879 1063 22943
rect 1127 22879 1153 22943
rect 1217 22879 1243 22943
rect 1307 22879 1333 22943
rect 1397 22879 1423 22943
rect 1487 22879 1492 22943
rect 968 22862 1492 22879
rect 968 22798 973 22862
rect 1037 22798 1063 22862
rect 1127 22798 1153 22862
rect 1217 22798 1243 22862
rect 1307 22798 1333 22862
rect 1397 22798 1423 22862
rect 1487 22798 1492 22862
rect 968 22781 1492 22798
rect 968 22717 973 22781
rect 1037 22717 1063 22781
rect 1127 22717 1153 22781
rect 1217 22717 1243 22781
rect 1307 22717 1333 22781
rect 1397 22717 1423 22781
rect 1487 22717 1492 22781
rect 968 22700 1492 22717
rect 968 22636 973 22700
rect 1037 22636 1063 22700
rect 1127 22636 1153 22700
rect 1217 22636 1243 22700
rect 1307 22636 1333 22700
rect 1397 22636 1423 22700
rect 1487 22636 1492 22700
rect 968 22619 1492 22636
rect 968 22555 973 22619
rect 1037 22555 1063 22619
rect 1127 22555 1153 22619
rect 1217 22555 1243 22619
rect 1307 22555 1333 22619
rect 1397 22555 1423 22619
rect 1487 22555 1492 22619
rect 968 22538 1492 22555
rect 968 22474 973 22538
rect 1037 22474 1063 22538
rect 1127 22474 1153 22538
rect 1217 22474 1243 22538
rect 1307 22474 1333 22538
rect 1397 22474 1423 22538
rect 1487 22474 1492 22538
rect 968 22457 1492 22474
rect 968 22393 973 22457
rect 1037 22393 1063 22457
rect 1127 22393 1153 22457
rect 1217 22393 1243 22457
rect 1307 22393 1333 22457
rect 1397 22393 1423 22457
rect 1487 22393 1492 22457
rect 968 22376 1492 22393
rect 968 22312 973 22376
rect 1037 22312 1063 22376
rect 1127 22312 1153 22376
rect 1217 22312 1243 22376
rect 1307 22312 1333 22376
rect 1397 22312 1423 22376
rect 1487 22312 1492 22376
rect 968 22295 1492 22312
rect 968 22231 973 22295
rect 1037 22231 1063 22295
rect 1127 22231 1153 22295
rect 1217 22231 1243 22295
rect 1307 22231 1333 22295
rect 1397 22231 1423 22295
rect 1487 22231 1492 22295
rect 968 22214 1492 22231
rect 968 22150 973 22214
rect 1037 22150 1063 22214
rect 1127 22150 1153 22214
rect 1217 22150 1243 22214
rect 1307 22150 1333 22214
rect 1397 22150 1423 22214
rect 1487 22150 1492 22214
rect 968 22133 1492 22150
rect 968 22069 973 22133
rect 1037 22069 1063 22133
rect 1127 22069 1153 22133
rect 1217 22069 1243 22133
rect 1307 22069 1333 22133
rect 1397 22069 1423 22133
rect 1487 22069 1492 22133
rect 968 22052 1492 22069
rect 968 21988 973 22052
rect 1037 21988 1063 22052
rect 1127 21988 1153 22052
rect 1217 21988 1243 22052
rect 1307 21988 1333 22052
rect 1397 21988 1423 22052
rect 1487 21988 1492 22052
rect 968 21971 1492 21988
rect 968 21907 973 21971
rect 1037 21907 1063 21971
rect 1127 21907 1153 21971
rect 1217 21907 1243 21971
rect 1307 21907 1333 21971
rect 1397 21907 1423 21971
rect 1487 21907 1492 21971
rect 968 21890 1492 21907
rect 968 21826 973 21890
rect 1037 21826 1063 21890
rect 1127 21826 1153 21890
rect 1217 21826 1243 21890
rect 1307 21826 1333 21890
rect 1397 21826 1423 21890
rect 1487 21826 1492 21890
rect 968 21809 1492 21826
rect 968 21745 973 21809
rect 1037 21745 1063 21809
rect 1127 21745 1153 21809
rect 1217 21745 1243 21809
rect 1307 21745 1333 21809
rect 1397 21745 1423 21809
rect 1487 21745 1492 21809
rect 968 21728 1492 21745
rect 968 21664 973 21728
rect 1037 21664 1063 21728
rect 1127 21664 1153 21728
rect 1217 21664 1243 21728
rect 1307 21664 1333 21728
rect 1397 21664 1423 21728
rect 1487 21664 1492 21728
rect 968 21647 1492 21664
rect 968 21583 973 21647
rect 1037 21583 1063 21647
rect 1127 21583 1153 21647
rect 1217 21583 1243 21647
rect 1307 21583 1333 21647
rect 1397 21583 1423 21647
rect 1487 21583 1492 21647
rect 968 21566 1492 21583
rect 968 21502 973 21566
rect 1037 21502 1063 21566
rect 1127 21502 1153 21566
rect 1217 21502 1243 21566
rect 1307 21502 1333 21566
rect 1397 21502 1423 21566
rect 1487 21502 1492 21566
rect 968 21485 1492 21502
rect 968 21421 973 21485
rect 1037 21421 1063 21485
rect 1127 21421 1153 21485
rect 1217 21421 1243 21485
rect 1307 21421 1333 21485
rect 1397 21421 1423 21485
rect 1487 21421 1492 21485
rect 968 21404 1492 21421
rect 968 21340 973 21404
rect 1037 21340 1063 21404
rect 1127 21340 1153 21404
rect 1217 21340 1243 21404
rect 1307 21340 1333 21404
rect 1397 21340 1423 21404
rect 1487 21340 1492 21404
rect 968 21323 1492 21340
rect 968 21259 973 21323
rect 1037 21259 1063 21323
rect 1127 21259 1153 21323
rect 1217 21259 1243 21323
rect 1307 21259 1333 21323
rect 1397 21259 1423 21323
rect 1487 21259 1492 21323
rect 968 21242 1492 21259
rect 968 21178 973 21242
rect 1037 21178 1063 21242
rect 1127 21178 1153 21242
rect 1217 21178 1243 21242
rect 1307 21178 1333 21242
rect 1397 21178 1423 21242
rect 1487 21178 1492 21242
rect 968 21161 1492 21178
rect 968 21097 973 21161
rect 1037 21097 1063 21161
rect 1127 21097 1153 21161
rect 1217 21097 1243 21161
rect 1307 21097 1333 21161
rect 1397 21097 1423 21161
rect 1487 21097 1492 21161
rect 968 21080 1492 21097
rect 968 21016 973 21080
rect 1037 21016 1063 21080
rect 1127 21016 1153 21080
rect 1217 21016 1243 21080
rect 1307 21016 1333 21080
rect 1397 21016 1423 21080
rect 1487 21016 1492 21080
rect 968 20999 1492 21016
rect 968 20935 973 20999
rect 1037 20935 1063 20999
rect 1127 20935 1153 20999
rect 1217 20935 1243 20999
rect 1307 20935 1333 20999
rect 1397 20935 1423 20999
rect 1487 20971 1492 20999
rect 13506 33108 14030 33109
rect 13506 33044 13511 33108
rect 13575 33044 13601 33108
rect 13665 33044 13691 33108
rect 13755 33044 13781 33108
rect 13845 33044 13871 33108
rect 13935 33044 13961 33108
rect 14025 33044 14030 33108
rect 13506 33028 14030 33044
rect 13506 32964 13511 33028
rect 13575 32964 13601 33028
rect 13665 32964 13691 33028
rect 13755 32964 13781 33028
rect 13845 32964 13871 33028
rect 13935 32964 13961 33028
rect 14025 32964 14030 33028
rect 13506 32948 14030 32964
rect 13506 32884 13511 32948
rect 13575 32884 13601 32948
rect 13665 32884 13691 32948
rect 13755 32884 13781 32948
rect 13845 32884 13871 32948
rect 13935 32884 13961 32948
rect 14025 32884 14030 32948
rect 13506 32868 14030 32884
rect 13506 32804 13511 32868
rect 13575 32804 13601 32868
rect 13665 32804 13691 32868
rect 13755 32804 13781 32868
rect 13845 32804 13871 32868
rect 13935 32804 13961 32868
rect 14025 32804 14030 32868
rect 13506 32788 14030 32804
rect 13506 32724 13511 32788
rect 13575 32724 13601 32788
rect 13665 32724 13691 32788
rect 13755 32724 13781 32788
rect 13845 32724 13871 32788
rect 13935 32724 13961 32788
rect 14025 32724 14030 32788
rect 13506 32708 14030 32724
rect 13506 32644 13511 32708
rect 13575 32644 13601 32708
rect 13665 32644 13691 32708
rect 13755 32644 13781 32708
rect 13845 32644 13871 32708
rect 13935 32644 13961 32708
rect 14025 32644 14030 32708
rect 13506 32628 14030 32644
rect 13506 32564 13511 32628
rect 13575 32564 13601 32628
rect 13665 32564 13691 32628
rect 13755 32564 13781 32628
rect 13845 32564 13871 32628
rect 13935 32564 13961 32628
rect 14025 32564 14030 32628
rect 13506 32548 14030 32564
rect 13506 32484 13511 32548
rect 13575 32484 13601 32548
rect 13665 32484 13691 32548
rect 13755 32484 13781 32548
rect 13845 32484 13871 32548
rect 13935 32484 13961 32548
rect 14025 32484 14030 32548
rect 13506 32468 14030 32484
rect 13506 32404 13511 32468
rect 13575 32404 13601 32468
rect 13665 32404 13691 32468
rect 13755 32404 13781 32468
rect 13845 32404 13871 32468
rect 13935 32404 13961 32468
rect 14025 32404 14030 32468
rect 13506 32388 14030 32404
rect 13506 32324 13511 32388
rect 13575 32324 13601 32388
rect 13665 32324 13691 32388
rect 13755 32324 13781 32388
rect 13845 32324 13871 32388
rect 13935 32324 13961 32388
rect 14025 32324 14030 32388
rect 13506 32308 14030 32324
rect 13506 32244 13511 32308
rect 13575 32244 13601 32308
rect 13665 32244 13691 32308
rect 13755 32244 13781 32308
rect 13845 32244 13871 32308
rect 13935 32244 13961 32308
rect 14025 32244 14030 32308
rect 13506 32228 14030 32244
rect 13506 32164 13511 32228
rect 13575 32164 13601 32228
rect 13665 32164 13691 32228
rect 13755 32164 13781 32228
rect 13845 32164 13871 32228
rect 13935 32164 13961 32228
rect 14025 32164 14030 32228
rect 13506 32148 14030 32164
rect 13506 32084 13511 32148
rect 13575 32084 13601 32148
rect 13665 32084 13691 32148
rect 13755 32084 13781 32148
rect 13845 32084 13871 32148
rect 13935 32084 13961 32148
rect 14025 32084 14030 32148
rect 13506 32068 14030 32084
rect 13506 32004 13511 32068
rect 13575 32004 13601 32068
rect 13665 32004 13691 32068
rect 13755 32004 13781 32068
rect 13845 32004 13871 32068
rect 13935 32004 13961 32068
rect 14025 32004 14030 32068
rect 13506 31988 14030 32004
rect 13506 31924 13511 31988
rect 13575 31924 13601 31988
rect 13665 31924 13691 31988
rect 13755 31924 13781 31988
rect 13845 31924 13871 31988
rect 13935 31924 13961 31988
rect 14025 31924 14030 31988
rect 13506 31908 14030 31924
rect 13506 31844 13511 31908
rect 13575 31844 13601 31908
rect 13665 31844 13691 31908
rect 13755 31844 13781 31908
rect 13845 31844 13871 31908
rect 13935 31844 13961 31908
rect 14025 31844 14030 31908
rect 13506 31828 14030 31844
rect 13506 31764 13511 31828
rect 13575 31764 13601 31828
rect 13665 31764 13691 31828
rect 13755 31764 13781 31828
rect 13845 31764 13871 31828
rect 13935 31764 13961 31828
rect 14025 31764 14030 31828
rect 13506 31748 14030 31764
rect 13506 31684 13511 31748
rect 13575 31684 13601 31748
rect 13665 31684 13691 31748
rect 13755 31684 13781 31748
rect 13845 31684 13871 31748
rect 13935 31684 13961 31748
rect 14025 31684 14030 31748
rect 13506 31668 14030 31684
rect 13506 31604 13511 31668
rect 13575 31604 13601 31668
rect 13665 31604 13691 31668
rect 13755 31604 13781 31668
rect 13845 31604 13871 31668
rect 13935 31604 13961 31668
rect 14025 31604 14030 31668
rect 13506 31588 14030 31604
rect 13506 31524 13511 31588
rect 13575 31524 13601 31588
rect 13665 31524 13691 31588
rect 13755 31524 13781 31588
rect 13845 31524 13871 31588
rect 13935 31524 13961 31588
rect 14025 31524 14030 31588
rect 13506 31508 14030 31524
rect 13506 31444 13511 31508
rect 13575 31444 13601 31508
rect 13665 31444 13691 31508
rect 13755 31444 13781 31508
rect 13845 31444 13871 31508
rect 13935 31444 13961 31508
rect 14025 31444 14030 31508
rect 13506 31428 14030 31444
rect 13506 31364 13511 31428
rect 13575 31364 13601 31428
rect 13665 31364 13691 31428
rect 13755 31364 13781 31428
rect 13845 31364 13871 31428
rect 13935 31364 13961 31428
rect 14025 31364 14030 31428
rect 13506 31348 14030 31364
rect 13506 31284 13511 31348
rect 13575 31284 13601 31348
rect 13665 31284 13691 31348
rect 13755 31284 13781 31348
rect 13845 31284 13871 31348
rect 13935 31284 13961 31348
rect 14025 31284 14030 31348
rect 13506 31268 14030 31284
rect 13506 31204 13511 31268
rect 13575 31204 13601 31268
rect 13665 31204 13691 31268
rect 13755 31204 13781 31268
rect 13845 31204 13871 31268
rect 13935 31204 13961 31268
rect 14025 31204 14030 31268
rect 13506 31188 14030 31204
rect 13506 31124 13511 31188
rect 13575 31124 13601 31188
rect 13665 31124 13691 31188
rect 13755 31124 13781 31188
rect 13845 31124 13871 31188
rect 13935 31124 13961 31188
rect 14025 31124 14030 31188
rect 13506 31108 14030 31124
rect 13506 31044 13511 31108
rect 13575 31044 13601 31108
rect 13665 31044 13691 31108
rect 13755 31044 13781 31108
rect 13845 31044 13871 31108
rect 13935 31044 13961 31108
rect 14025 31044 14030 31108
rect 13506 31028 14030 31044
rect 13506 30964 13511 31028
rect 13575 30964 13601 31028
rect 13665 30964 13691 31028
rect 13755 30964 13781 31028
rect 13845 30964 13871 31028
rect 13935 30964 13961 31028
rect 14025 30964 14030 31028
rect 13506 30948 14030 30964
rect 13506 30884 13511 30948
rect 13575 30884 13601 30948
rect 13665 30884 13691 30948
rect 13755 30884 13781 30948
rect 13845 30884 13871 30948
rect 13935 30884 13961 30948
rect 14025 30884 14030 30948
rect 13506 30868 14030 30884
rect 13506 30804 13511 30868
rect 13575 30804 13601 30868
rect 13665 30804 13691 30868
rect 13755 30804 13781 30868
rect 13845 30804 13871 30868
rect 13935 30804 13961 30868
rect 14025 30804 14030 30868
rect 13506 30788 14030 30804
rect 13506 30724 13511 30788
rect 13575 30724 13601 30788
rect 13665 30724 13691 30788
rect 13755 30724 13781 30788
rect 13845 30724 13871 30788
rect 13935 30724 13961 30788
rect 14025 30724 14030 30788
rect 13506 30708 14030 30724
rect 13506 30644 13511 30708
rect 13575 30644 13601 30708
rect 13665 30644 13691 30708
rect 13755 30644 13781 30708
rect 13845 30644 13871 30708
rect 13935 30644 13961 30708
rect 14025 30644 14030 30708
rect 13506 30628 14030 30644
rect 13506 30564 13511 30628
rect 13575 30564 13601 30628
rect 13665 30564 13691 30628
rect 13755 30564 13781 30628
rect 13845 30564 13871 30628
rect 13935 30564 13961 30628
rect 14025 30564 14030 30628
rect 13506 30548 14030 30564
rect 13506 30484 13511 30548
rect 13575 30484 13601 30548
rect 13665 30484 13691 30548
rect 13755 30484 13781 30548
rect 13845 30484 13871 30548
rect 13935 30484 13961 30548
rect 14025 30484 14030 30548
rect 13506 30468 14030 30484
rect 13506 30404 13511 30468
rect 13575 30404 13601 30468
rect 13665 30404 13691 30468
rect 13755 30404 13781 30468
rect 13845 30404 13871 30468
rect 13935 30404 13961 30468
rect 14025 30404 14030 30468
rect 13506 30388 14030 30404
rect 13506 30324 13511 30388
rect 13575 30324 13601 30388
rect 13665 30324 13691 30388
rect 13755 30324 13781 30388
rect 13845 30324 13871 30388
rect 13935 30324 13961 30388
rect 14025 30324 14030 30388
rect 13506 30308 14030 30324
rect 13506 30244 13511 30308
rect 13575 30244 13601 30308
rect 13665 30244 13691 30308
rect 13755 30244 13781 30308
rect 13845 30244 13871 30308
rect 13935 30244 13961 30308
rect 14025 30244 14030 30308
rect 13506 30228 14030 30244
rect 13506 30164 13511 30228
rect 13575 30164 13601 30228
rect 13665 30164 13691 30228
rect 13755 30164 13781 30228
rect 13845 30164 13871 30228
rect 13935 30164 13961 30228
rect 14025 30164 14030 30228
rect 13506 30148 14030 30164
rect 13506 30084 13511 30148
rect 13575 30084 13601 30148
rect 13665 30084 13691 30148
rect 13755 30084 13781 30148
rect 13845 30084 13871 30148
rect 13935 30084 13961 30148
rect 14025 30084 14030 30148
rect 13506 30068 14030 30084
rect 13506 30004 13511 30068
rect 13575 30004 13601 30068
rect 13665 30004 13691 30068
rect 13755 30004 13781 30068
rect 13845 30004 13871 30068
rect 13935 30004 13961 30068
rect 14025 30004 14030 30068
rect 13506 29988 14030 30004
rect 13506 29924 13511 29988
rect 13575 29924 13601 29988
rect 13665 29924 13691 29988
rect 13755 29924 13781 29988
rect 13845 29924 13871 29988
rect 13935 29924 13961 29988
rect 14025 29924 14030 29988
rect 13506 29908 14030 29924
rect 13506 29844 13511 29908
rect 13575 29844 13601 29908
rect 13665 29844 13691 29908
rect 13755 29844 13781 29908
rect 13845 29844 13871 29908
rect 13935 29844 13961 29908
rect 14025 29844 14030 29908
rect 13506 29828 14030 29844
rect 13506 29764 13511 29828
rect 13575 29764 13601 29828
rect 13665 29764 13691 29828
rect 13755 29764 13781 29828
rect 13845 29764 13871 29828
rect 13935 29764 13961 29828
rect 14025 29764 14030 29828
rect 13506 29748 14030 29764
rect 13506 29684 13511 29748
rect 13575 29684 13601 29748
rect 13665 29684 13691 29748
rect 13755 29684 13781 29748
rect 13845 29684 13871 29748
rect 13935 29684 13961 29748
rect 14025 29684 14030 29748
rect 13506 29668 14030 29684
rect 13506 29604 13511 29668
rect 13575 29604 13601 29668
rect 13665 29604 13691 29668
rect 13755 29604 13781 29668
rect 13845 29604 13871 29668
rect 13935 29604 13961 29668
rect 14025 29604 14030 29668
rect 13506 29588 14030 29604
rect 13506 29524 13511 29588
rect 13575 29524 13601 29588
rect 13665 29524 13691 29588
rect 13755 29524 13781 29588
rect 13845 29524 13871 29588
rect 13935 29524 13961 29588
rect 14025 29524 14030 29588
rect 13506 29508 14030 29524
rect 13506 29444 13511 29508
rect 13575 29444 13601 29508
rect 13665 29444 13691 29508
rect 13755 29444 13781 29508
rect 13845 29444 13871 29508
rect 13935 29444 13961 29508
rect 14025 29444 14030 29508
rect 13506 29428 14030 29444
rect 13506 29364 13511 29428
rect 13575 29364 13601 29428
rect 13665 29364 13691 29428
rect 13755 29364 13781 29428
rect 13845 29364 13871 29428
rect 13935 29364 13961 29428
rect 14025 29364 14030 29428
rect 13506 29348 14030 29364
rect 13506 29284 13511 29348
rect 13575 29284 13601 29348
rect 13665 29284 13691 29348
rect 13755 29284 13781 29348
rect 13845 29284 13871 29348
rect 13935 29284 13961 29348
rect 14025 29284 14030 29348
rect 13506 29268 14030 29284
rect 13506 29204 13511 29268
rect 13575 29204 13601 29268
rect 13665 29204 13691 29268
rect 13755 29204 13781 29268
rect 13845 29204 13871 29268
rect 13935 29204 13961 29268
rect 14025 29204 14030 29268
rect 13506 29188 14030 29204
rect 13506 29124 13511 29188
rect 13575 29124 13601 29188
rect 13665 29124 13691 29188
rect 13755 29124 13781 29188
rect 13845 29124 13871 29188
rect 13935 29124 13961 29188
rect 14025 29124 14030 29188
rect 13506 29108 14030 29124
rect 13506 29044 13511 29108
rect 13575 29044 13601 29108
rect 13665 29044 13691 29108
rect 13755 29044 13781 29108
rect 13845 29044 13871 29108
rect 13935 29044 13961 29108
rect 14025 29044 14030 29108
rect 13506 29028 14030 29044
rect 13506 28964 13511 29028
rect 13575 28964 13601 29028
rect 13665 28964 13691 29028
rect 13755 28964 13781 29028
rect 13845 28964 13871 29028
rect 13935 28964 13961 29028
rect 14025 28964 14030 29028
rect 13506 28948 14030 28964
rect 13506 28884 13511 28948
rect 13575 28884 13601 28948
rect 13665 28884 13691 28948
rect 13755 28884 13781 28948
rect 13845 28884 13871 28948
rect 13935 28884 13961 28948
rect 14025 28884 14030 28948
rect 13506 28868 14030 28884
rect 13506 28804 13511 28868
rect 13575 28804 13601 28868
rect 13665 28804 13691 28868
rect 13755 28804 13781 28868
rect 13845 28804 13871 28868
rect 13935 28804 13961 28868
rect 14025 28804 14030 28868
rect 13506 28788 14030 28804
rect 13506 28724 13511 28788
rect 13575 28724 13601 28788
rect 13665 28724 13691 28788
rect 13755 28724 13781 28788
rect 13845 28724 13871 28788
rect 13935 28724 13961 28788
rect 14025 28724 14030 28788
rect 13506 28708 14030 28724
rect 13506 28644 13511 28708
rect 13575 28644 13601 28708
rect 13665 28644 13691 28708
rect 13755 28644 13781 28708
rect 13845 28644 13871 28708
rect 13935 28644 13961 28708
rect 14025 28644 14030 28708
rect 13506 28628 14030 28644
rect 13506 28564 13511 28628
rect 13575 28564 13601 28628
rect 13665 28564 13691 28628
rect 13755 28564 13781 28628
rect 13845 28564 13871 28628
rect 13935 28564 13961 28628
rect 14025 28564 14030 28628
rect 13506 28548 14030 28564
rect 13506 28484 13511 28548
rect 13575 28484 13601 28548
rect 13665 28484 13691 28548
rect 13755 28484 13781 28548
rect 13845 28484 13871 28548
rect 13935 28484 13961 28548
rect 14025 28484 14030 28548
rect 13506 28468 14030 28484
rect 13506 28404 13511 28468
rect 13575 28404 13601 28468
rect 13665 28404 13691 28468
rect 13755 28404 13781 28468
rect 13845 28404 13871 28468
rect 13935 28404 13961 28468
rect 14025 28404 14030 28468
rect 13506 28388 14030 28404
rect 13506 28324 13511 28388
rect 13575 28324 13601 28388
rect 13665 28324 13691 28388
rect 13755 28324 13781 28388
rect 13845 28324 13871 28388
rect 13935 28324 13961 28388
rect 14025 28324 14030 28388
rect 13506 28308 14030 28324
rect 13506 28244 13511 28308
rect 13575 28244 13601 28308
rect 13665 28244 13691 28308
rect 13755 28244 13781 28308
rect 13845 28244 13871 28308
rect 13935 28244 13961 28308
rect 14025 28244 14030 28308
rect 13506 28228 14030 28244
rect 13506 28164 13511 28228
rect 13575 28164 13601 28228
rect 13665 28164 13691 28228
rect 13755 28164 13781 28228
rect 13845 28164 13871 28228
rect 13935 28164 13961 28228
rect 14025 28164 14030 28228
rect 13506 28148 14030 28164
rect 13506 28084 13511 28148
rect 13575 28084 13601 28148
rect 13665 28084 13691 28148
rect 13755 28084 13781 28148
rect 13845 28084 13871 28148
rect 13935 28084 13961 28148
rect 14025 28084 14030 28148
rect 13506 28068 14030 28084
rect 13506 28004 13511 28068
rect 13575 28004 13601 28068
rect 13665 28004 13691 28068
rect 13755 28004 13781 28068
rect 13845 28004 13871 28068
rect 13935 28004 13961 28068
rect 14025 28004 14030 28068
rect 13506 27988 14030 28004
rect 13506 27924 13511 27988
rect 13575 27924 13601 27988
rect 13665 27924 13691 27988
rect 13755 27924 13781 27988
rect 13845 27924 13871 27988
rect 13935 27924 13961 27988
rect 14025 27924 14030 27988
rect 13506 27908 14030 27924
rect 13506 27844 13511 27908
rect 13575 27844 13601 27908
rect 13665 27844 13691 27908
rect 13755 27844 13781 27908
rect 13845 27844 13871 27908
rect 13935 27844 13961 27908
rect 14025 27844 14030 27908
rect 13506 27828 14030 27844
rect 13506 27764 13511 27828
rect 13575 27764 13601 27828
rect 13665 27764 13691 27828
rect 13755 27764 13781 27828
rect 13845 27764 13871 27828
rect 13935 27764 13961 27828
rect 14025 27764 14030 27828
rect 13506 27748 14030 27764
rect 13506 27684 13511 27748
rect 13575 27684 13601 27748
rect 13665 27684 13691 27748
rect 13755 27684 13781 27748
rect 13845 27684 13871 27748
rect 13935 27684 13961 27748
rect 14025 27684 14030 27748
rect 13506 27668 14030 27684
rect 13506 27604 13511 27668
rect 13575 27604 13601 27668
rect 13665 27604 13691 27668
rect 13755 27604 13781 27668
rect 13845 27604 13871 27668
rect 13935 27604 13961 27668
rect 14025 27604 14030 27668
rect 13506 27588 14030 27604
rect 13506 27524 13511 27588
rect 13575 27524 13601 27588
rect 13665 27524 13691 27588
rect 13755 27524 13781 27588
rect 13845 27524 13871 27588
rect 13935 27524 13961 27588
rect 14025 27524 14030 27588
rect 13506 27508 14030 27524
rect 13506 27444 13511 27508
rect 13575 27444 13601 27508
rect 13665 27444 13691 27508
rect 13755 27444 13781 27508
rect 13845 27444 13871 27508
rect 13935 27444 13961 27508
rect 14025 27444 14030 27508
rect 13506 27428 14030 27444
rect 13506 27364 13511 27428
rect 13575 27364 13601 27428
rect 13665 27364 13691 27428
rect 13755 27364 13781 27428
rect 13845 27364 13871 27428
rect 13935 27364 13961 27428
rect 14025 27364 14030 27428
rect 13506 27348 14030 27364
rect 13506 27284 13511 27348
rect 13575 27284 13601 27348
rect 13665 27284 13691 27348
rect 13755 27284 13781 27348
rect 13845 27284 13871 27348
rect 13935 27284 13961 27348
rect 14025 27284 14030 27348
rect 13506 27268 14030 27284
rect 13506 27204 13511 27268
rect 13575 27204 13601 27268
rect 13665 27204 13691 27268
rect 13755 27204 13781 27268
rect 13845 27204 13871 27268
rect 13935 27204 13961 27268
rect 14025 27204 14030 27268
rect 13506 27188 14030 27204
rect 13506 27124 13511 27188
rect 13575 27124 13601 27188
rect 13665 27124 13691 27188
rect 13755 27124 13781 27188
rect 13845 27124 13871 27188
rect 13935 27124 13961 27188
rect 14025 27124 14030 27188
rect 13506 27108 14030 27124
rect 13506 27044 13511 27108
rect 13575 27044 13601 27108
rect 13665 27044 13691 27108
rect 13755 27044 13781 27108
rect 13845 27044 13871 27108
rect 13935 27044 13961 27108
rect 14025 27044 14030 27108
rect 13506 27028 14030 27044
rect 13506 26964 13511 27028
rect 13575 26964 13601 27028
rect 13665 26964 13691 27028
rect 13755 26964 13781 27028
rect 13845 26964 13871 27028
rect 13935 26964 13961 27028
rect 14025 26964 14030 27028
rect 13506 26948 14030 26964
rect 13506 26884 13511 26948
rect 13575 26884 13601 26948
rect 13665 26884 13691 26948
rect 13755 26884 13781 26948
rect 13845 26884 13871 26948
rect 13935 26884 13961 26948
rect 14025 26884 14030 26948
rect 13506 26868 14030 26884
rect 13506 26804 13511 26868
rect 13575 26804 13601 26868
rect 13665 26804 13691 26868
rect 13755 26804 13781 26868
rect 13845 26804 13871 26868
rect 13935 26804 13961 26868
rect 14025 26804 14030 26868
rect 13506 26788 14030 26804
rect 13506 26724 13511 26788
rect 13575 26724 13601 26788
rect 13665 26724 13691 26788
rect 13755 26724 13781 26788
rect 13845 26724 13871 26788
rect 13935 26724 13961 26788
rect 14025 26724 14030 26788
rect 13506 26708 14030 26724
rect 13506 26644 13511 26708
rect 13575 26644 13601 26708
rect 13665 26644 13691 26708
rect 13755 26644 13781 26708
rect 13845 26644 13871 26708
rect 13935 26644 13961 26708
rect 14025 26644 14030 26708
rect 13506 26628 14030 26644
rect 13506 26564 13511 26628
rect 13575 26564 13601 26628
rect 13665 26564 13691 26628
rect 13755 26564 13781 26628
rect 13845 26564 13871 26628
rect 13935 26564 13961 26628
rect 14025 26564 14030 26628
rect 13506 26548 14030 26564
rect 13506 26484 13511 26548
rect 13575 26484 13601 26548
rect 13665 26484 13691 26548
rect 13755 26484 13781 26548
rect 13845 26484 13871 26548
rect 13935 26484 13961 26548
rect 14025 26484 14030 26548
rect 13506 26468 14030 26484
rect 13506 26404 13511 26468
rect 13575 26404 13601 26468
rect 13665 26404 13691 26468
rect 13755 26404 13781 26468
rect 13845 26404 13871 26468
rect 13935 26404 13961 26468
rect 14025 26404 14030 26468
rect 13506 26388 14030 26404
rect 13506 26324 13511 26388
rect 13575 26324 13601 26388
rect 13665 26324 13691 26388
rect 13755 26324 13781 26388
rect 13845 26324 13871 26388
rect 13935 26324 13961 26388
rect 14025 26324 14030 26388
rect 13506 26308 14030 26324
rect 13506 26244 13511 26308
rect 13575 26244 13601 26308
rect 13665 26244 13691 26308
rect 13755 26244 13781 26308
rect 13845 26244 13871 26308
rect 13935 26244 13961 26308
rect 14025 26244 14030 26308
rect 13506 26228 14030 26244
rect 13506 26164 13511 26228
rect 13575 26164 13601 26228
rect 13665 26164 13691 26228
rect 13755 26164 13781 26228
rect 13845 26164 13871 26228
rect 13935 26164 13961 26228
rect 14025 26164 14030 26228
rect 13506 26148 14030 26164
rect 13506 26084 13511 26148
rect 13575 26084 13601 26148
rect 13665 26084 13691 26148
rect 13755 26084 13781 26148
rect 13845 26084 13871 26148
rect 13935 26084 13961 26148
rect 14025 26084 14030 26148
rect 13506 26068 14030 26084
rect 13506 26004 13511 26068
rect 13575 26004 13601 26068
rect 13665 26004 13691 26068
rect 13755 26004 13781 26068
rect 13845 26004 13871 26068
rect 13935 26004 13961 26068
rect 14025 26004 14030 26068
rect 13506 25988 14030 26004
rect 13506 25924 13511 25988
rect 13575 25924 13601 25988
rect 13665 25924 13691 25988
rect 13755 25924 13781 25988
rect 13845 25924 13871 25988
rect 13935 25924 13961 25988
rect 14025 25924 14030 25988
rect 13506 25908 14030 25924
rect 13506 25844 13511 25908
rect 13575 25844 13601 25908
rect 13665 25844 13691 25908
rect 13755 25844 13781 25908
rect 13845 25844 13871 25908
rect 13935 25844 13961 25908
rect 14025 25844 14030 25908
rect 13506 25828 14030 25844
rect 13506 25764 13511 25828
rect 13575 25764 13601 25828
rect 13665 25764 13691 25828
rect 13755 25764 13781 25828
rect 13845 25764 13871 25828
rect 13935 25764 13961 25828
rect 14025 25764 14030 25828
rect 13506 25748 14030 25764
rect 13506 25684 13511 25748
rect 13575 25684 13601 25748
rect 13665 25684 13691 25748
rect 13755 25684 13781 25748
rect 13845 25684 13871 25748
rect 13935 25684 13961 25748
rect 14025 25684 14030 25748
rect 13506 25668 14030 25684
rect 13506 25604 13511 25668
rect 13575 25604 13601 25668
rect 13665 25604 13691 25668
rect 13755 25604 13781 25668
rect 13845 25604 13871 25668
rect 13935 25604 13961 25668
rect 14025 25604 14030 25668
rect 13506 25588 14030 25604
rect 13506 25524 13511 25588
rect 13575 25524 13601 25588
rect 13665 25524 13691 25588
rect 13755 25524 13781 25588
rect 13845 25524 13871 25588
rect 13935 25524 13961 25588
rect 14025 25524 14030 25588
rect 13506 25508 14030 25524
rect 13506 25444 13511 25508
rect 13575 25444 13601 25508
rect 13665 25444 13691 25508
rect 13755 25444 13781 25508
rect 13845 25444 13871 25508
rect 13935 25444 13961 25508
rect 14025 25444 14030 25508
rect 13506 25428 14030 25444
rect 13506 25364 13511 25428
rect 13575 25364 13601 25428
rect 13665 25364 13691 25428
rect 13755 25364 13781 25428
rect 13845 25364 13871 25428
rect 13935 25364 13961 25428
rect 14025 25364 14030 25428
rect 13506 25348 14030 25364
rect 13506 25284 13511 25348
rect 13575 25284 13601 25348
rect 13665 25284 13691 25348
rect 13755 25284 13781 25348
rect 13845 25284 13871 25348
rect 13935 25284 13961 25348
rect 14025 25284 14030 25348
rect 13506 25268 14030 25284
rect 13506 25204 13511 25268
rect 13575 25204 13601 25268
rect 13665 25204 13691 25268
rect 13755 25204 13781 25268
rect 13845 25204 13871 25268
rect 13935 25204 13961 25268
rect 14025 25204 14030 25268
rect 13506 25188 14030 25204
rect 13506 25124 13511 25188
rect 13575 25124 13601 25188
rect 13665 25124 13691 25188
rect 13755 25124 13781 25188
rect 13845 25124 13871 25188
rect 13935 25124 13961 25188
rect 14025 25124 14030 25188
rect 13506 25108 14030 25124
rect 13506 25044 13511 25108
rect 13575 25044 13601 25108
rect 13665 25044 13691 25108
rect 13755 25044 13781 25108
rect 13845 25044 13871 25108
rect 13935 25044 13961 25108
rect 14025 25044 14030 25108
rect 13506 25028 14030 25044
rect 13506 24964 13511 25028
rect 13575 24964 13601 25028
rect 13665 24964 13691 25028
rect 13755 24964 13781 25028
rect 13845 24964 13871 25028
rect 13935 24964 13961 25028
rect 14025 24964 14030 25028
rect 13506 24948 14030 24964
rect 13506 24884 13511 24948
rect 13575 24884 13601 24948
rect 13665 24884 13691 24948
rect 13755 24884 13781 24948
rect 13845 24884 13871 24948
rect 13935 24884 13961 24948
rect 14025 24884 14030 24948
rect 13506 24868 14030 24884
rect 13506 24804 13511 24868
rect 13575 24804 13601 24868
rect 13665 24804 13691 24868
rect 13755 24804 13781 24868
rect 13845 24804 13871 24868
rect 13935 24804 13961 24868
rect 14025 24804 14030 24868
rect 13506 24788 14030 24804
rect 13506 24724 13511 24788
rect 13575 24724 13601 24788
rect 13665 24724 13691 24788
rect 13755 24724 13781 24788
rect 13845 24724 13871 24788
rect 13935 24724 13961 24788
rect 14025 24724 14030 24788
rect 13506 24708 14030 24724
rect 13506 24644 13511 24708
rect 13575 24644 13601 24708
rect 13665 24644 13691 24708
rect 13755 24644 13781 24708
rect 13845 24644 13871 24708
rect 13935 24644 13961 24708
rect 14025 24644 14030 24708
rect 13506 24628 14030 24644
rect 13506 24564 13511 24628
rect 13575 24564 13601 24628
rect 13665 24564 13691 24628
rect 13755 24564 13781 24628
rect 13845 24564 13871 24628
rect 13935 24564 13961 24628
rect 14025 24564 14030 24628
rect 13506 24548 14030 24564
rect 13506 24484 13511 24548
rect 13575 24484 13601 24548
rect 13665 24484 13691 24548
rect 13755 24484 13781 24548
rect 13845 24484 13871 24548
rect 13935 24484 13961 24548
rect 14025 24484 14030 24548
rect 13506 24468 14030 24484
rect 13506 24404 13511 24468
rect 13575 24404 13601 24468
rect 13665 24404 13691 24468
rect 13755 24404 13781 24468
rect 13845 24404 13871 24468
rect 13935 24404 13961 24468
rect 14025 24404 14030 24468
rect 13506 24388 14030 24404
rect 13506 24324 13511 24388
rect 13575 24324 13601 24388
rect 13665 24324 13691 24388
rect 13755 24324 13781 24388
rect 13845 24324 13871 24388
rect 13935 24324 13961 24388
rect 14025 24324 14030 24388
rect 13506 24308 14030 24324
rect 13506 24244 13511 24308
rect 13575 24244 13601 24308
rect 13665 24244 13691 24308
rect 13755 24244 13781 24308
rect 13845 24244 13871 24308
rect 13935 24244 13961 24308
rect 14025 24244 14030 24308
rect 13506 24228 14030 24244
rect 13506 24164 13511 24228
rect 13575 24164 13601 24228
rect 13665 24164 13691 24228
rect 13755 24164 13781 24228
rect 13845 24164 13871 24228
rect 13935 24164 13961 24228
rect 14025 24164 14030 24228
rect 13506 24148 14030 24164
rect 13506 24084 13511 24148
rect 13575 24084 13601 24148
rect 13665 24084 13691 24148
rect 13755 24084 13781 24148
rect 13845 24084 13871 24148
rect 13935 24084 13961 24148
rect 14025 24084 14030 24148
rect 13506 24068 14030 24084
rect 13506 24004 13511 24068
rect 13575 24004 13601 24068
rect 13665 24004 13691 24068
rect 13755 24004 13781 24068
rect 13845 24004 13871 24068
rect 13935 24004 13961 24068
rect 14025 24004 14030 24068
rect 13506 23988 14030 24004
rect 13506 23924 13511 23988
rect 13575 23924 13601 23988
rect 13665 23924 13691 23988
rect 13755 23924 13781 23988
rect 13845 23924 13871 23988
rect 13935 23924 13961 23988
rect 14025 23924 14030 23988
rect 13506 23908 14030 23924
rect 13506 23844 13511 23908
rect 13575 23844 13601 23908
rect 13665 23844 13691 23908
rect 13755 23844 13781 23908
rect 13845 23844 13871 23908
rect 13935 23844 13961 23908
rect 14025 23844 14030 23908
rect 13506 23828 14030 23844
rect 13506 23764 13511 23828
rect 13575 23764 13601 23828
rect 13665 23764 13691 23828
rect 13755 23764 13781 23828
rect 13845 23764 13871 23828
rect 13935 23764 13961 23828
rect 14025 23764 14030 23828
rect 13506 23748 14030 23764
rect 13506 23684 13511 23748
rect 13575 23684 13601 23748
rect 13665 23684 13691 23748
rect 13755 23684 13781 23748
rect 13845 23684 13871 23748
rect 13935 23684 13961 23748
rect 14025 23684 14030 23748
rect 13506 23668 14030 23684
rect 13506 23604 13511 23668
rect 13575 23604 13601 23668
rect 13665 23604 13691 23668
rect 13755 23604 13781 23668
rect 13845 23604 13871 23668
rect 13935 23604 13961 23668
rect 14025 23604 14030 23668
rect 13506 23588 14030 23604
rect 13506 23524 13511 23588
rect 13575 23524 13601 23588
rect 13665 23524 13691 23588
rect 13755 23524 13781 23588
rect 13845 23524 13871 23588
rect 13935 23524 13961 23588
rect 14025 23524 14030 23588
rect 13506 23508 14030 23524
rect 13506 23444 13511 23508
rect 13575 23444 13601 23508
rect 13665 23444 13691 23508
rect 13755 23444 13781 23508
rect 13845 23444 13871 23508
rect 13935 23444 13961 23508
rect 14025 23444 14030 23508
rect 13506 23428 14030 23444
rect 13506 23364 13511 23428
rect 13575 23364 13601 23428
rect 13665 23364 13691 23428
rect 13755 23364 13781 23428
rect 13845 23364 13871 23428
rect 13935 23364 13961 23428
rect 14025 23364 14030 23428
rect 13506 23348 14030 23364
rect 13506 23284 13511 23348
rect 13575 23284 13601 23348
rect 13665 23284 13691 23348
rect 13755 23284 13781 23348
rect 13845 23284 13871 23348
rect 13935 23284 13961 23348
rect 14025 23284 14030 23348
rect 13506 23267 14030 23284
rect 13506 23203 13511 23267
rect 13575 23203 13601 23267
rect 13665 23203 13691 23267
rect 13755 23203 13781 23267
rect 13845 23203 13871 23267
rect 13935 23203 13961 23267
rect 14025 23203 14030 23267
rect 13506 23186 14030 23203
rect 13506 23122 13511 23186
rect 13575 23122 13601 23186
rect 13665 23122 13691 23186
rect 13755 23122 13781 23186
rect 13845 23122 13871 23186
rect 13935 23122 13961 23186
rect 14025 23122 14030 23186
rect 13506 23105 14030 23122
rect 13506 23041 13511 23105
rect 13575 23041 13601 23105
rect 13665 23041 13691 23105
rect 13755 23041 13781 23105
rect 13845 23041 13871 23105
rect 13935 23041 13961 23105
rect 14025 23041 14030 23105
rect 13506 23024 14030 23041
rect 13506 22960 13511 23024
rect 13575 22960 13601 23024
rect 13665 22960 13691 23024
rect 13755 22960 13781 23024
rect 13845 22960 13871 23024
rect 13935 22960 13961 23024
rect 14025 22960 14030 23024
rect 13506 22943 14030 22960
rect 13506 22879 13511 22943
rect 13575 22879 13601 22943
rect 13665 22879 13691 22943
rect 13755 22879 13781 22943
rect 13845 22879 13871 22943
rect 13935 22879 13961 22943
rect 14025 22879 14030 22943
rect 13506 22862 14030 22879
rect 13506 22798 13511 22862
rect 13575 22798 13601 22862
rect 13665 22798 13691 22862
rect 13755 22798 13781 22862
rect 13845 22798 13871 22862
rect 13935 22798 13961 22862
rect 14025 22798 14030 22862
rect 13506 22781 14030 22798
rect 13506 22717 13511 22781
rect 13575 22717 13601 22781
rect 13665 22717 13691 22781
rect 13755 22717 13781 22781
rect 13845 22717 13871 22781
rect 13935 22717 13961 22781
rect 14025 22717 14030 22781
rect 13506 22700 14030 22717
rect 13506 22636 13511 22700
rect 13575 22636 13601 22700
rect 13665 22636 13691 22700
rect 13755 22636 13781 22700
rect 13845 22636 13871 22700
rect 13935 22636 13961 22700
rect 14025 22636 14030 22700
rect 13506 22619 14030 22636
rect 13506 22555 13511 22619
rect 13575 22555 13601 22619
rect 13665 22555 13691 22619
rect 13755 22555 13781 22619
rect 13845 22555 13871 22619
rect 13935 22555 13961 22619
rect 14025 22555 14030 22619
rect 13506 22538 14030 22555
rect 13506 22474 13511 22538
rect 13575 22474 13601 22538
rect 13665 22474 13691 22538
rect 13755 22474 13781 22538
rect 13845 22474 13871 22538
rect 13935 22474 13961 22538
rect 14025 22474 14030 22538
rect 13506 22457 14030 22474
rect 13506 22393 13511 22457
rect 13575 22393 13601 22457
rect 13665 22393 13691 22457
rect 13755 22393 13781 22457
rect 13845 22393 13871 22457
rect 13935 22393 13961 22457
rect 14025 22393 14030 22457
rect 13506 22376 14030 22393
rect 13506 22312 13511 22376
rect 13575 22312 13601 22376
rect 13665 22312 13691 22376
rect 13755 22312 13781 22376
rect 13845 22312 13871 22376
rect 13935 22312 13961 22376
rect 14025 22312 14030 22376
rect 13506 22295 14030 22312
rect 13506 22231 13511 22295
rect 13575 22231 13601 22295
rect 13665 22231 13691 22295
rect 13755 22231 13781 22295
rect 13845 22231 13871 22295
rect 13935 22231 13961 22295
rect 14025 22231 14030 22295
rect 13506 22214 14030 22231
rect 13506 22150 13511 22214
rect 13575 22150 13601 22214
rect 13665 22150 13691 22214
rect 13755 22150 13781 22214
rect 13845 22150 13871 22214
rect 13935 22150 13961 22214
rect 14025 22150 14030 22214
rect 13506 22133 14030 22150
rect 13506 22069 13511 22133
rect 13575 22069 13601 22133
rect 13665 22069 13691 22133
rect 13755 22069 13781 22133
rect 13845 22069 13871 22133
rect 13935 22069 13961 22133
rect 14025 22069 14030 22133
rect 13506 22052 14030 22069
rect 13506 21988 13511 22052
rect 13575 21988 13601 22052
rect 13665 21988 13691 22052
rect 13755 21988 13781 22052
rect 13845 21988 13871 22052
rect 13935 21988 13961 22052
rect 14025 21988 14030 22052
rect 13506 21971 14030 21988
rect 13506 21907 13511 21971
rect 13575 21907 13601 21971
rect 13665 21907 13691 21971
rect 13755 21907 13781 21971
rect 13845 21907 13871 21971
rect 13935 21907 13961 21971
rect 14025 21907 14030 21971
rect 13506 21890 14030 21907
rect 13506 21826 13511 21890
rect 13575 21826 13601 21890
rect 13665 21826 13691 21890
rect 13755 21826 13781 21890
rect 13845 21826 13871 21890
rect 13935 21826 13961 21890
rect 14025 21826 14030 21890
rect 13506 21809 14030 21826
rect 13506 21745 13511 21809
rect 13575 21745 13601 21809
rect 13665 21745 13691 21809
rect 13755 21745 13781 21809
rect 13845 21745 13871 21809
rect 13935 21745 13961 21809
rect 14025 21745 14030 21809
rect 13506 21728 14030 21745
rect 13506 21664 13511 21728
rect 13575 21664 13601 21728
rect 13665 21664 13691 21728
rect 13755 21664 13781 21728
rect 13845 21664 13871 21728
rect 13935 21664 13961 21728
rect 14025 21664 14030 21728
rect 13506 21647 14030 21664
rect 13506 21583 13511 21647
rect 13575 21583 13601 21647
rect 13665 21583 13691 21647
rect 13755 21583 13781 21647
rect 13845 21583 13871 21647
rect 13935 21583 13961 21647
rect 14025 21583 14030 21647
rect 13506 21566 14030 21583
rect 13506 21502 13511 21566
rect 13575 21502 13601 21566
rect 13665 21502 13691 21566
rect 13755 21502 13781 21566
rect 13845 21502 13871 21566
rect 13935 21502 13961 21566
rect 14025 21502 14030 21566
rect 13506 21485 14030 21502
rect 13506 21421 13511 21485
rect 13575 21421 13601 21485
rect 13665 21421 13691 21485
rect 13755 21421 13781 21485
rect 13845 21421 13871 21485
rect 13935 21421 13961 21485
rect 14025 21421 14030 21485
rect 13506 21404 14030 21421
rect 13506 21340 13511 21404
rect 13575 21340 13601 21404
rect 13665 21340 13691 21404
rect 13755 21340 13781 21404
rect 13845 21340 13871 21404
rect 13935 21340 13961 21404
rect 14025 21340 14030 21404
rect 13506 21323 14030 21340
rect 13506 21259 13511 21323
rect 13575 21259 13601 21323
rect 13665 21259 13691 21323
rect 13755 21259 13781 21323
rect 13845 21259 13871 21323
rect 13935 21259 13961 21323
rect 14025 21259 14030 21323
rect 13506 21242 14030 21259
rect 13506 21178 13511 21242
rect 13575 21178 13601 21242
rect 13665 21178 13691 21242
rect 13755 21178 13781 21242
rect 13845 21178 13871 21242
rect 13935 21178 13961 21242
rect 14025 21178 14030 21242
rect 13506 21161 14030 21178
rect 13506 21097 13511 21161
rect 13575 21097 13601 21161
rect 13665 21097 13691 21161
rect 13755 21097 13781 21161
rect 13845 21097 13871 21161
rect 13935 21097 13961 21161
rect 14025 21097 14030 21161
rect 13506 21080 14030 21097
rect 13506 21016 13511 21080
rect 13575 21016 13601 21080
rect 13665 21016 13691 21080
rect 13755 21016 13781 21080
rect 13845 21016 13871 21080
rect 13935 21016 13961 21080
rect 14025 21016 14030 21080
rect 13506 20999 14030 21016
rect 13506 20971 13511 20999
rect 1487 20938 1587 20971
rect 1487 20935 1522 20938
rect 968 20918 1522 20935
rect 968 20854 973 20918
rect 1037 20854 1063 20918
rect 1127 20854 1153 20918
rect 1217 20854 1243 20918
rect 1307 20854 1333 20918
rect 1397 20854 1423 20918
rect 1487 20874 1522 20918
rect 1586 20874 1587 20938
rect 1487 20854 1587 20874
rect 968 20853 1587 20854
rect 1462 20841 1587 20853
rect 13411 20938 13511 20971
rect 13411 20874 13412 20938
rect 13476 20935 13511 20938
rect 13575 20935 13601 20999
rect 13665 20935 13691 20999
rect 13755 20935 13781 20999
rect 13845 20935 13871 20999
rect 13935 20935 13961 20999
rect 14025 20935 14030 20999
rect 13476 20918 14030 20935
rect 13476 20874 13511 20918
rect 13411 20854 13511 20874
rect 13575 20854 13601 20918
rect 13665 20854 13691 20918
rect 13755 20854 13781 20918
rect 13845 20854 13871 20918
rect 13935 20854 13961 20918
rect 14025 20854 14030 20918
rect 13411 20853 14030 20854
rect 13411 20841 13536 20853
rect 1302 20824 1727 20826
rect 1131 20782 1256 20815
rect 1131 20718 1132 20782
rect 1196 20718 1256 20782
rect 1131 20685 1256 20718
rect 1302 20760 1303 20824
rect 1367 20760 1392 20824
rect 1456 20760 1482 20824
rect 1546 20760 1572 20824
rect 1636 20760 1662 20824
rect 1726 20760 1727 20824
rect 1302 20708 1727 20760
rect 1302 20644 1303 20708
rect 1367 20644 1392 20708
rect 1456 20644 1482 20708
rect 1546 20644 1572 20708
rect 1636 20644 1662 20708
rect 1726 20644 1727 20708
rect 13271 20824 13696 20826
rect 13271 20760 13272 20824
rect 13336 20760 13362 20824
rect 13426 20760 13452 20824
rect 13516 20760 13542 20824
rect 13606 20760 13631 20824
rect 13695 20760 13696 20824
rect 13271 20708 13696 20760
rect 1302 20592 1727 20644
rect 1302 20528 1303 20592
rect 1367 20528 1392 20592
rect 1456 20528 1482 20592
rect 1546 20528 1572 20592
rect 1636 20528 1662 20592
rect 1726 20528 1727 20592
rect 1743 20630 1868 20663
rect 1743 20566 1803 20630
rect 1867 20566 1868 20630
rect 1743 20533 1868 20566
rect 13130 20630 13255 20663
rect 13130 20566 13131 20630
rect 13195 20566 13255 20630
rect 13130 20533 13255 20566
rect 13271 20644 13272 20708
rect 13336 20644 13362 20708
rect 13426 20644 13452 20708
rect 13516 20644 13542 20708
rect 13606 20644 13631 20708
rect 13695 20644 13696 20708
rect 13710 20822 13834 20823
rect 13710 20758 13740 20822
rect 13804 20758 13834 20822
rect 13710 20711 13834 20758
rect 13840 20815 13907 20848
rect 13840 20751 13842 20815
rect 13906 20751 13907 20815
rect 13840 20718 13907 20751
rect 13710 20647 13740 20711
rect 13804 20647 13834 20711
rect 13710 20646 13834 20647
rect 13271 20592 13696 20644
rect 1302 20526 1727 20528
rect 13271 20528 13272 20592
rect 13336 20528 13362 20592
rect 13426 20528 13452 20592
rect 13516 20528 13542 20592
rect 13606 20528 13631 20592
rect 13695 20528 13696 20592
rect 13271 20526 13696 20528
rect 1622 20504 2047 20506
rect 1455 20468 1580 20501
rect 1455 20404 1515 20468
rect 1579 20404 1580 20468
rect 1455 20371 1580 20404
rect 1622 20440 1623 20504
rect 1687 20440 1712 20504
rect 1776 20440 1802 20504
rect 1866 20440 1892 20504
rect 1956 20440 1982 20504
rect 2046 20440 2047 20504
rect 1622 20388 2047 20440
rect 1622 20324 1623 20388
rect 1687 20324 1712 20388
rect 1776 20324 1802 20388
rect 1866 20324 1892 20388
rect 1956 20324 1982 20388
rect 2046 20324 2047 20388
rect 12951 20504 13376 20506
rect 12951 20440 12952 20504
rect 13016 20440 13042 20504
rect 13106 20440 13132 20504
rect 13196 20440 13222 20504
rect 13286 20440 13311 20504
rect 13375 20440 13376 20504
rect 12951 20388 13376 20440
rect 1622 20272 2047 20324
rect 1622 20208 1623 20272
rect 1687 20208 1712 20272
rect 1776 20208 1802 20272
rect 1866 20208 1892 20272
rect 1956 20208 1982 20272
rect 2046 20208 2047 20272
rect 2068 20305 2193 20338
rect 2068 20241 2128 20305
rect 2192 20241 2193 20305
rect 2068 20208 2193 20241
rect 12805 20305 12930 20338
rect 12805 20241 12806 20305
rect 12870 20241 12930 20305
rect 12805 20208 12930 20241
rect 12951 20324 12952 20388
rect 13016 20324 13042 20388
rect 13106 20324 13132 20388
rect 13196 20324 13222 20388
rect 13286 20324 13311 20388
rect 13375 20324 13376 20388
rect 13418 20468 13543 20501
rect 13418 20404 13419 20468
rect 13483 20404 13543 20468
rect 13418 20371 13543 20404
rect 12951 20272 13376 20324
rect 12951 20208 12952 20272
rect 13016 20208 13042 20272
rect 13106 20208 13132 20272
rect 13196 20208 13222 20272
rect 13286 20208 13311 20272
rect 13375 20208 13376 20272
rect 1622 20206 2047 20208
rect 12951 20206 13376 20208
rect 1946 20180 2371 20182
rect 1783 20140 1908 20173
rect 1783 20076 1843 20140
rect 1907 20076 1908 20140
rect 1783 20043 1908 20076
rect 1946 20116 1947 20180
rect 2011 20116 2036 20180
rect 2100 20116 2126 20180
rect 2190 20116 2216 20180
rect 2280 20116 2306 20180
rect 2370 20116 2371 20180
rect 1946 20064 2371 20116
rect 12627 20180 13052 20182
rect 12627 20116 12628 20180
rect 12692 20116 12718 20180
rect 12782 20116 12808 20180
rect 12872 20116 12898 20180
rect 12962 20116 12987 20180
rect 13051 20116 13052 20180
rect 1946 20000 1947 20064
rect 2011 20000 2036 20064
rect 2100 20000 2126 20064
rect 2190 20000 2216 20064
rect 2280 20000 2306 20064
rect 2370 20000 2371 20064
rect 1946 19948 2371 20000
rect 12140 20069 12552 20070
rect 12140 20005 12141 20069
rect 12205 20005 12257 20069
rect 12321 20005 12372 20069
rect 12436 20005 12487 20069
rect 12551 20005 12552 20069
rect 1946 19884 1947 19948
rect 2011 19884 2036 19948
rect 2100 19884 2126 19948
rect 2190 19884 2216 19948
rect 2280 19884 2306 19948
rect 2370 19884 2371 19948
rect 1946 19882 2371 19884
rect 12036 19954 12126 19987
rect 12036 19890 12037 19954
rect 12101 19890 12126 19954
rect 12036 19857 12126 19890
rect 12140 19949 12552 20005
rect 12140 19885 12141 19949
rect 12205 19885 12257 19949
rect 12321 19885 12372 19949
rect 12436 19885 12487 19949
rect 12551 19885 12552 19949
rect 12140 19884 12552 19885
rect 12627 20064 13052 20116
rect 12627 20000 12628 20064
rect 12692 20000 12718 20064
rect 12782 20000 12808 20064
rect 12872 20000 12898 20064
rect 12962 20000 12987 20064
rect 13051 20000 13052 20064
rect 13090 20140 13215 20173
rect 13090 20076 13091 20140
rect 13155 20076 13215 20140
rect 13090 20043 13215 20076
rect 12627 19948 13052 20000
rect 12627 19884 12628 19948
rect 12692 19884 12718 19948
rect 12782 19884 12808 19948
rect 12872 19884 12898 19948
rect 12962 19884 12987 19948
rect 13051 19884 13052 19948
rect 12627 19882 13052 19884
rect 11893 19843 12715 19845
rect 2124 19799 2249 19832
rect 2124 19735 2184 19799
rect 2248 19735 2249 19799
rect 2124 19702 2249 19735
rect 11893 19779 11894 19843
rect 11958 19779 11978 19843
rect 12042 19779 12062 19843
rect 12126 19779 12146 19843
rect 12210 19779 12230 19843
rect 12294 19779 12314 19843
rect 12378 19779 12398 19843
rect 12462 19779 12482 19843
rect 12546 19779 12566 19843
rect 12630 19779 12650 19843
rect 12714 19779 12715 19843
rect 11893 19727 12715 19779
rect 11760 19706 11884 19707
rect 11760 19642 11790 19706
rect 11854 19642 11884 19706
rect 11760 19613 11884 19642
rect 11760 19549 11790 19613
rect 11854 19549 11884 19613
rect 11760 19548 11884 19549
rect 11893 19663 11894 19727
rect 11958 19663 11978 19727
rect 12042 19663 12062 19727
rect 12126 19663 12146 19727
rect 12210 19663 12230 19727
rect 12294 19663 12314 19727
rect 12378 19663 12398 19727
rect 12462 19663 12482 19727
rect 12546 19663 12566 19727
rect 12630 19663 12650 19727
rect 12714 19663 12715 19727
rect 12749 19799 12874 19832
rect 12749 19735 12750 19799
rect 12814 19735 12874 19799
rect 12749 19702 12874 19735
rect 11893 19611 12715 19663
rect 11893 19547 11894 19611
rect 11958 19547 11978 19611
rect 12042 19547 12062 19611
rect 12126 19547 12146 19611
rect 12210 19547 12230 19611
rect 12294 19547 12314 19611
rect 12378 19547 12398 19611
rect 12462 19547 12482 19611
rect 12546 19547 12566 19611
rect 12630 19547 12650 19611
rect 12714 19547 12715 19611
rect 11893 19545 12715 19547
rect 886 3646 2072 3658
rect 886 3022 887 3646
rect 2071 3022 2072 3646
rect 886 3010 2072 3022
rect 6886 3010 8072 3658
rect 12886 3646 14072 3658
rect 12886 3022 12887 3646
rect 14071 3022 14072 3646
rect 12886 3010 14072 3022
use sky130_fd_io__com_busses_esd  sky130_fd_io__com_busses_esd_0
timestamp 1644511149
transform 1 0 8 0 1 550
box 0 -142 15000 39451
<< properties >>
string GDS_END 265690
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io__analog.gds
string GDS_START 148
<< end >>
