magic
tech sky130B
timestamp 1644511149
<< properties >>
string GDS_END 49972
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 49648
<< end >>
