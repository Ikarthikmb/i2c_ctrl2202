magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 26 21 612 203
rect 29 -17 63 21
<< locali >>
rect 17 199 156 265
rect 190 199 252 493
rect 286 333 396 493
rect 530 333 627 493
rect 286 299 627 333
rect 286 199 356 265
rect 397 64 440 265
rect 489 165 532 299
rect 566 199 627 265
rect 489 51 627 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 299 156 527
rect 430 367 496 527
rect 17 17 114 165
rect 148 131 350 165
rect 148 51 182 131
rect 216 17 282 97
rect 316 51 350 131
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
rlabel locali s 17 199 156 265 6 A1
port 1 nsew signal input
rlabel locali s 190 199 252 493 6 A2
port 2 nsew signal input
rlabel locali s 286 199 356 265 6 A3
port 3 nsew signal input
rlabel locali s 397 64 440 265 6 B1
port 4 nsew signal input
rlabel locali s 566 199 627 265 6 C1
port 5 nsew signal input
rlabel metal1 s 0 -48 644 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 26 21 612 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 682 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 644 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 489 51 627 165 6 Y
port 10 nsew signal output
rlabel locali s 489 165 532 299 6 Y
port 10 nsew signal output
rlabel locali s 286 299 627 333 6 Y
port 10 nsew signal output
rlabel locali s 530 333 627 493 6 Y
port 10 nsew signal output
rlabel locali s 286 333 396 493 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 644 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 886694
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 879846
<< end >>
