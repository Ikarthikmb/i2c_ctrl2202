magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 26 21 612 157
rect 29 -17 63 21
<< scnmos >>
rect 108 47 138 131
rect 192 47 222 131
rect 276 47 306 131
rect 428 47 458 131
rect 500 47 530 131
<< scpmoshvt >>
rect 108 369 138 497
rect 192 369 222 497
rect 276 369 306 497
rect 396 369 426 497
rect 500 369 530 497
<< ndiff >>
rect 52 106 108 131
rect 52 72 64 106
rect 98 72 108 106
rect 52 47 108 72
rect 138 106 192 131
rect 138 72 148 106
rect 182 72 192 106
rect 138 47 192 72
rect 222 89 276 131
rect 222 55 232 89
rect 266 55 276 89
rect 222 47 276 55
rect 306 106 428 131
rect 306 72 316 106
rect 350 72 428 106
rect 306 47 428 72
rect 458 47 500 131
rect 530 106 586 131
rect 530 72 540 106
rect 574 72 586 106
rect 530 47 586 72
<< pdiff >>
rect 52 484 108 497
rect 52 450 64 484
rect 98 450 108 484
rect 52 416 108 450
rect 52 382 64 416
rect 98 382 108 416
rect 52 369 108 382
rect 138 369 192 497
rect 222 369 276 497
rect 306 484 396 497
rect 306 450 334 484
rect 368 450 396 484
rect 306 416 396 450
rect 306 382 334 416
rect 368 382 396 416
rect 306 369 396 382
rect 426 484 500 497
rect 426 450 446 484
rect 480 450 500 484
rect 426 416 500 450
rect 426 382 446 416
rect 480 382 500 416
rect 426 369 500 382
rect 530 484 592 497
rect 530 450 546 484
rect 580 450 592 484
rect 530 416 592 450
rect 530 382 546 416
rect 580 382 592 416
rect 530 369 592 382
<< ndiffc >>
rect 64 72 98 106
rect 148 72 182 106
rect 232 55 266 89
rect 316 72 350 106
rect 540 72 574 106
<< pdiffc >>
rect 64 450 98 484
rect 64 382 98 416
rect 334 450 368 484
rect 334 382 368 416
rect 446 450 480 484
rect 446 382 480 416
rect 546 450 580 484
rect 546 382 580 416
<< poly >>
rect 108 497 138 523
rect 192 497 222 523
rect 276 497 306 523
rect 396 497 426 523
rect 500 497 530 523
rect 108 265 138 369
rect 192 265 222 369
rect 276 265 306 369
rect 396 265 426 369
rect 500 265 530 369
rect 54 249 138 265
rect 54 215 64 249
rect 98 215 138 249
rect 54 199 138 215
rect 180 249 234 265
rect 180 215 190 249
rect 224 215 234 249
rect 180 199 234 215
rect 276 249 330 265
rect 276 215 286 249
rect 320 215 330 249
rect 276 199 330 215
rect 396 249 458 265
rect 396 215 406 249
rect 440 215 458 249
rect 396 199 458 215
rect 108 131 138 199
rect 192 131 222 199
rect 276 131 306 199
rect 428 131 458 199
rect 500 249 610 265
rect 500 215 566 249
rect 600 215 610 249
rect 500 199 610 215
rect 500 131 530 199
rect 108 21 138 47
rect 192 21 222 47
rect 276 21 306 47
rect 428 21 458 47
rect 500 21 530 47
<< polycont >>
rect 64 215 98 249
rect 190 215 224 249
rect 286 215 320 249
rect 406 215 440 249
rect 566 215 600 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 17 484 156 527
rect 17 450 64 484
rect 98 450 156 484
rect 17 416 156 450
rect 17 382 64 416
rect 98 382 156 416
rect 17 359 156 382
rect 17 249 156 325
rect 17 215 64 249
rect 98 215 156 249
rect 17 199 156 215
rect 190 249 252 493
rect 286 484 396 493
rect 286 450 334 484
rect 368 450 396 484
rect 286 416 396 450
rect 286 382 334 416
rect 368 382 396 416
rect 286 333 396 382
rect 430 484 496 527
rect 430 450 446 484
rect 480 450 496 484
rect 430 416 496 450
rect 430 382 446 416
rect 480 382 496 416
rect 430 367 496 382
rect 530 484 627 493
rect 530 450 546 484
rect 580 450 627 484
rect 530 416 627 450
rect 530 382 546 416
rect 580 382 627 416
rect 530 333 627 382
rect 286 299 627 333
rect 224 215 252 249
rect 190 199 252 215
rect 286 249 356 265
rect 320 215 356 249
rect 286 199 356 215
rect 397 249 440 265
rect 397 215 406 249
rect 17 153 114 199
rect 148 131 350 165
rect 17 106 114 119
rect 17 72 64 106
rect 98 72 114 106
rect 17 17 114 72
rect 148 106 182 131
rect 316 106 350 131
rect 148 51 182 72
rect 216 89 282 97
rect 216 55 232 89
rect 266 55 282 89
rect 216 17 282 55
rect 316 51 350 72
rect 397 52 440 215
rect 489 119 532 299
rect 566 249 627 265
rect 600 215 627 249
rect 566 153 627 215
rect 489 106 627 119
rect 489 72 540 106
rect 574 72 627 106
rect 489 51 627 72
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 213 425 247 459 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 581 153 615 187 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 357 247 391 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 121 289 155 323 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 581 85 615 119 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 A3
port 3 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 B1
port 4 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 121 221 155 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 153 523 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 489 85 523 119 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 489 289 523 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 305 357 339 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 305 425 339 459 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 581 425 615 459 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 581 357 615 391 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o311ai_0
rlabel metal1 s 0 -48 644 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 879788
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 872362
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 3.220 0.000 
<< end >>
