magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 458 163 735 203
rect 1 27 735 163
rect 29 -17 63 27
rect 461 21 735 27
<< locali >>
rect 29 149 82 265
rect 363 425 458 493
rect 575 359 632 493
rect 402 153 484 249
rect 598 289 632 359
rect 598 185 719 289
rect 402 61 444 153
rect 598 143 632 185
rect 583 51 632 143
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 17 315 80 527
rect 206 426 329 527
rect 116 249 171 381
rect 210 319 257 392
rect 291 391 329 426
rect 291 353 357 391
rect 402 319 440 378
rect 492 358 535 527
rect 210 285 564 319
rect 116 203 283 249
rect 17 17 71 115
rect 116 61 171 203
rect 317 114 368 285
rect 211 61 368 114
rect 518 199 564 285
rect 666 325 719 527
rect 482 17 548 116
rect 666 17 719 149
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
<< metal1 >>
rect 0 561 736 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 736 561
rect 0 496 736 527
rect 0 17 736 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 736 17
rect 0 -48 736 -17
<< labels >>
rlabel locali s 29 149 82 265 6 A_N
port 1 nsew signal input
rlabel locali s 363 425 458 493 6 B
port 2 nsew signal input
rlabel locali s 402 61 444 153 6 C
port 3 nsew signal input
rlabel locali s 402 153 484 249 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 736 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 461 21 735 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 29 -17 63 27 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 27 735 163 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 458 163 735 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 583 51 632 143 6 X
port 8 nsew signal output
rlabel locali s 598 143 632 185 6 X
port 8 nsew signal output
rlabel locali s 598 185 719 289 6 X
port 8 nsew signal output
rlabel locali s 598 289 632 359 6 X
port 8 nsew signal output
rlabel locali s 575 359 632 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3884062
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3877514
<< end >>
