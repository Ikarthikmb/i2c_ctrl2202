magic
tech sky130B
timestamp 1644511149
<< properties >>
string GDS_END 15433544
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15432068
<< end >>
