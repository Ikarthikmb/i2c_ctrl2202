/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/sky130A/libs.tech/ngspice/sonos_see_e/end_of_life.spice