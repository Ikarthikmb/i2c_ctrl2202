magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 157 157 549 203
rect 59 21 549 157
rect 59 17 63 21
rect 29 -17 63 17
<< scnmos >>
rect 138 47 168 131
rect 236 47 266 177
rect 354 47 384 177
rect 440 47 470 177
<< scpmoshvt >>
rect 80 413 110 497
rect 270 297 300 497
rect 356 297 386 497
rect 442 297 472 497
<< ndiff >>
rect 183 157 236 177
rect 183 131 191 157
rect 85 107 138 131
rect 85 73 93 107
rect 127 73 138 107
rect 85 47 138 73
rect 168 123 191 131
rect 225 123 236 157
rect 168 89 236 123
rect 168 55 191 89
rect 225 55 236 89
rect 168 47 236 55
rect 266 129 354 177
rect 266 95 293 129
rect 327 95 354 129
rect 266 47 354 95
rect 384 47 440 177
rect 470 161 523 177
rect 470 127 481 161
rect 515 127 523 161
rect 470 93 523 127
rect 470 59 481 93
rect 515 59 523 93
rect 470 47 523 59
<< pdiff >>
rect 27 471 80 497
rect 27 437 35 471
rect 69 437 80 471
rect 27 413 80 437
rect 110 485 163 497
rect 110 451 121 485
rect 155 451 163 485
rect 110 413 163 451
rect 217 479 270 497
rect 217 445 225 479
rect 259 445 270 479
rect 217 411 270 445
rect 217 377 225 411
rect 259 377 270 411
rect 217 343 270 377
rect 217 309 225 343
rect 259 309 270 343
rect 217 297 270 309
rect 300 475 356 497
rect 300 441 311 475
rect 345 441 356 475
rect 300 407 356 441
rect 300 373 311 407
rect 345 373 356 407
rect 300 297 356 373
rect 386 489 442 497
rect 386 455 397 489
rect 431 455 442 489
rect 386 421 442 455
rect 386 387 397 421
rect 431 387 442 421
rect 386 297 442 387
rect 472 475 525 497
rect 472 441 483 475
rect 517 441 525 475
rect 472 407 525 441
rect 472 373 483 407
rect 517 373 525 407
rect 472 297 525 373
<< ndiffc >>
rect 93 73 127 107
rect 191 123 225 157
rect 191 55 225 89
rect 293 95 327 129
rect 481 127 515 161
rect 481 59 515 93
<< pdiffc >>
rect 35 437 69 471
rect 121 451 155 485
rect 225 445 259 479
rect 225 377 259 411
rect 225 309 259 343
rect 311 441 345 475
rect 311 373 345 407
rect 397 455 431 489
rect 397 387 431 421
rect 483 441 517 475
rect 483 373 517 407
<< poly >>
rect 80 497 110 523
rect 270 497 300 523
rect 356 497 386 523
rect 442 497 472 523
rect 80 393 110 413
rect 21 363 110 393
rect 21 317 75 363
rect 21 283 31 317
rect 65 283 75 317
rect 21 249 75 283
rect 21 215 31 249
rect 65 215 75 249
rect 117 305 171 321
rect 117 271 127 305
rect 161 277 171 305
rect 270 277 300 297
rect 161 271 300 277
rect 117 237 300 271
rect 356 265 386 297
rect 442 265 472 297
rect 344 249 398 265
rect 21 181 75 215
rect 21 151 168 181
rect 236 177 266 237
rect 344 215 354 249
rect 388 215 398 249
rect 344 199 398 215
rect 440 249 524 265
rect 440 215 480 249
rect 514 215 524 249
rect 440 199 524 215
rect 354 177 384 199
rect 440 177 470 199
rect 138 131 168 151
rect 138 21 168 47
rect 236 21 266 47
rect 354 21 384 47
rect 440 21 470 47
<< polycont >>
rect 31 283 65 317
rect 31 215 65 249
rect 127 271 161 305
rect 354 215 388 249
rect 480 215 514 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 19 471 71 487
rect 19 437 35 471
rect 69 437 71 471
rect 105 485 171 527
rect 105 451 121 485
rect 155 451 171 485
rect 105 445 171 451
rect 209 479 275 491
rect 209 445 225 479
rect 259 445 275 479
rect 19 409 71 437
rect 209 411 275 445
rect 19 369 171 409
rect 21 317 67 333
rect 21 283 31 317
rect 65 283 67 317
rect 21 249 67 283
rect 21 215 31 249
rect 65 215 67 249
rect 21 195 67 215
rect 103 305 171 369
rect 103 271 127 305
rect 161 271 171 305
rect 103 233 171 271
rect 209 377 225 411
rect 259 377 275 411
rect 209 343 275 377
rect 209 309 225 343
rect 259 309 275 343
rect 209 269 275 309
rect 309 475 347 491
rect 309 441 311 475
rect 345 441 347 475
rect 309 407 347 441
rect 309 373 311 407
rect 345 373 347 407
rect 381 489 447 527
rect 381 455 397 489
rect 431 455 447 489
rect 381 421 447 455
rect 381 387 397 421
rect 431 387 447 421
rect 381 381 447 387
rect 483 475 517 491
rect 483 407 517 441
rect 309 345 347 373
rect 483 345 517 373
rect 309 305 517 345
rect 103 143 149 233
rect 209 209 316 269
rect 73 107 149 143
rect 73 73 93 107
rect 127 73 149 107
rect 73 53 149 73
rect 185 157 231 173
rect 185 123 191 157
rect 225 123 231 157
rect 185 89 231 123
rect 185 55 191 89
rect 225 55 231 89
rect 185 17 231 55
rect 267 159 316 209
rect 352 249 431 269
rect 352 215 354 249
rect 388 215 431 249
rect 352 199 431 215
rect 470 249 528 269
rect 470 215 480 249
rect 514 215 528 249
rect 470 199 528 215
rect 267 129 353 159
rect 267 95 293 129
rect 327 95 353 129
rect 267 53 353 95
rect 389 75 431 199
rect 465 161 531 163
rect 465 127 481 161
rect 515 127 531 161
rect 465 93 531 127
rect 465 59 481 93
rect 515 59 531 93
rect 465 17 531 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
<< metal1 >>
rect 0 561 552 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 552 561
rect 0 496 552 527
rect 0 17 552 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 552 17
rect 0 -48 552 -17
<< labels >>
flabel locali s 305 85 339 119 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 213 221 247 255 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 215 425 249 459 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 215 289 249 323 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 215 357 249 391 0 FreeSans 200 0 0 0 Y
port 8 nsew signal output
flabel locali s 397 85 431 119 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 489 221 523 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 29 289 63 323 0 FreeSans 200 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 397 153 431 187 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a21boi_1
rlabel metal1 s 0 -48 552 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 552 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 552 544
string GDS_END 4006180
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3999944
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 13.800 0.000 
<< end >>
