magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< locali >>
rect 60243 77697 60277 77713
rect 60243 77647 60277 77663
rect 60243 76207 60277 76223
rect 60243 76157 60277 76173
rect 60243 74869 60277 74885
rect 60243 74819 60277 74835
rect 60243 73379 60277 73395
rect 60243 73329 60277 73345
rect 60243 72041 60277 72057
rect 60243 71991 60277 72007
rect 60243 70551 60277 70567
rect 60243 70501 60277 70517
rect 60243 69213 60277 69229
rect 60243 69163 60277 69179
rect 60243 67723 60277 67739
rect 60243 67673 60277 67689
rect 55077 64616 55111 64632
rect 55111 64582 55257 64616
rect 55077 64566 55111 64582
rect 12139 64376 12173 64392
rect 11993 64342 12139 64376
rect 12139 64326 12173 64342
rect 55077 64376 55111 64392
rect 55111 64342 55257 64376
rect 55077 64326 55111 64342
rect 12139 63826 12173 63842
rect 11993 63792 12139 63826
rect 12139 63776 12173 63792
rect 55077 63826 55111 63842
rect 55111 63792 55257 63826
rect 55077 63776 55111 63792
rect 12139 63586 12173 63602
rect 11993 63552 12139 63586
rect 12139 63536 12173 63552
rect 55077 63586 55111 63602
rect 55111 63552 55257 63586
rect 55077 63536 55111 63552
rect 12139 63036 12173 63052
rect 11993 63002 12139 63036
rect 12139 62986 12173 63002
rect 55077 63036 55111 63052
rect 55111 63002 55257 63036
rect 55077 62986 55111 63002
rect 12139 62796 12173 62812
rect 11993 62762 12139 62796
rect 12139 62746 12173 62762
rect 55077 62796 55111 62812
rect 55111 62762 55257 62796
rect 55077 62746 55111 62762
rect 12139 62246 12173 62262
rect 11993 62212 12139 62246
rect 12139 62196 12173 62212
rect 55077 62246 55111 62262
rect 55111 62212 55257 62246
rect 55077 62196 55111 62212
rect 12139 62006 12173 62022
rect 11993 61972 12139 62006
rect 12139 61956 12173 61972
rect 55077 62006 55111 62022
rect 55111 61972 55257 62006
rect 55077 61956 55111 61972
rect 12139 61456 12173 61472
rect 11993 61422 12139 61456
rect 12139 61406 12173 61422
rect 55077 61456 55111 61472
rect 55111 61422 55257 61456
rect 55077 61406 55111 61422
rect 12139 61216 12173 61232
rect 11993 61182 12139 61216
rect 12139 61166 12173 61182
rect 55077 61216 55111 61232
rect 55111 61182 55257 61216
rect 55077 61166 55111 61182
rect 12139 60666 12173 60682
rect 11993 60632 12139 60666
rect 12139 60616 12173 60632
rect 55077 60666 55111 60682
rect 55111 60632 55257 60666
rect 55077 60616 55111 60632
rect 12139 60426 12173 60442
rect 11993 60392 12139 60426
rect 12139 60376 12173 60392
rect 55077 60426 55111 60442
rect 55111 60392 55257 60426
rect 55077 60376 55111 60392
rect 12139 59876 12173 59892
rect 11993 59842 12139 59876
rect 12139 59826 12173 59842
rect 55077 59876 55111 59892
rect 55111 59842 55257 59876
rect 55077 59826 55111 59842
rect 12139 59636 12173 59652
rect 11993 59602 12139 59636
rect 12139 59586 12173 59602
rect 55077 59636 55111 59652
rect 55111 59602 55257 59636
rect 55077 59586 55111 59602
rect 12139 59086 12173 59102
rect 11993 59052 12139 59086
rect 12139 59036 12173 59052
rect 55077 59086 55111 59102
rect 55111 59052 55257 59086
rect 55077 59036 55111 59052
rect 12139 58846 12173 58862
rect 11993 58812 12139 58846
rect 12139 58796 12173 58812
rect 55077 58846 55111 58862
rect 55111 58812 55257 58846
rect 55077 58796 55111 58812
rect 12139 58296 12173 58312
rect 11993 58262 12139 58296
rect 12139 58246 12173 58262
rect 55077 58296 55111 58312
rect 55111 58262 55257 58296
rect 55077 58246 55111 58262
rect 12139 58056 12173 58072
rect 11993 58022 12139 58056
rect 12139 58006 12173 58022
rect 55077 58056 55111 58072
rect 55111 58022 55257 58056
rect 55077 58006 55111 58022
rect 12139 57506 12173 57522
rect 11993 57472 12139 57506
rect 12139 57456 12173 57472
rect 55077 57506 55111 57522
rect 55111 57472 55257 57506
rect 55077 57456 55111 57472
rect 12139 57266 12173 57282
rect 11993 57232 12139 57266
rect 12139 57216 12173 57232
rect 55077 57266 55111 57282
rect 55111 57232 55257 57266
rect 55077 57216 55111 57232
rect 12139 56716 12173 56732
rect 11993 56682 12139 56716
rect 12139 56666 12173 56682
rect 55077 56716 55111 56732
rect 55111 56682 55257 56716
rect 55077 56666 55111 56682
rect 12139 56476 12173 56492
rect 11993 56442 12139 56476
rect 12139 56426 12173 56442
rect 55077 56476 55111 56492
rect 55111 56442 55257 56476
rect 55077 56426 55111 56442
rect 12139 55926 12173 55942
rect 11993 55892 12139 55926
rect 12139 55876 12173 55892
rect 55077 55926 55111 55942
rect 55111 55892 55257 55926
rect 55077 55876 55111 55892
rect 12139 55686 12173 55702
rect 11993 55652 12139 55686
rect 12139 55636 12173 55652
rect 55077 55686 55111 55702
rect 55111 55652 55257 55686
rect 55077 55636 55111 55652
rect 12139 55136 12173 55152
rect 11993 55102 12139 55136
rect 12139 55086 12173 55102
rect 55077 55136 55111 55152
rect 55111 55102 55257 55136
rect 55077 55086 55111 55102
rect 12139 54896 12173 54912
rect 11993 54862 12139 54896
rect 12139 54846 12173 54862
rect 55077 54896 55111 54912
rect 55111 54862 55257 54896
rect 55077 54846 55111 54862
rect 12139 54346 12173 54362
rect 11993 54312 12139 54346
rect 12139 54296 12173 54312
rect 55077 54346 55111 54362
rect 55111 54312 55257 54346
rect 55077 54296 55111 54312
rect 12139 54106 12173 54122
rect 11993 54072 12139 54106
rect 12139 54056 12173 54072
rect 55077 54106 55111 54122
rect 55111 54072 55257 54106
rect 55077 54056 55111 54072
rect 12139 53556 12173 53572
rect 11993 53522 12139 53556
rect 12139 53506 12173 53522
rect 55077 53556 55111 53572
rect 55111 53522 55257 53556
rect 55077 53506 55111 53522
rect 12139 53316 12173 53332
rect 11993 53282 12139 53316
rect 12139 53266 12173 53282
rect 55077 53316 55111 53332
rect 55111 53282 55257 53316
rect 55077 53266 55111 53282
rect 12139 52766 12173 52782
rect 11993 52732 12139 52766
rect 12139 52716 12173 52732
rect 55077 52766 55111 52782
rect 55111 52732 55257 52766
rect 55077 52716 55111 52732
rect 12139 52526 12173 52542
rect 11993 52492 12139 52526
rect 12139 52476 12173 52492
rect 55077 52526 55111 52542
rect 55111 52492 55257 52526
rect 55077 52476 55111 52492
rect 12139 51976 12173 51992
rect 11993 51942 12139 51976
rect 12139 51926 12173 51942
rect 55077 51976 55111 51992
rect 55111 51942 55257 51976
rect 55077 51926 55111 51942
rect 12139 51736 12173 51752
rect 11993 51702 12139 51736
rect 12139 51686 12173 51702
rect 55077 51736 55111 51752
rect 55111 51702 55257 51736
rect 55077 51686 55111 51702
rect 12139 51186 12173 51202
rect 11993 51152 12139 51186
rect 12139 51136 12173 51152
rect 55077 51186 55111 51202
rect 55111 51152 55257 51186
rect 55077 51136 55111 51152
rect 12139 50946 12173 50962
rect 11993 50912 12139 50946
rect 12139 50896 12173 50912
rect 55077 50946 55111 50962
rect 55111 50912 55257 50946
rect 55077 50896 55111 50912
rect 12139 50396 12173 50412
rect 11993 50362 12139 50396
rect 12139 50346 12173 50362
rect 55077 50396 55111 50412
rect 55111 50362 55257 50396
rect 55077 50346 55111 50362
rect 12139 50156 12173 50172
rect 11993 50122 12139 50156
rect 12139 50106 12173 50122
rect 55077 50156 55111 50172
rect 55111 50122 55257 50156
rect 55077 50106 55111 50122
rect 12139 49606 12173 49622
rect 11993 49572 12139 49606
rect 12139 49556 12173 49572
rect 55077 49606 55111 49622
rect 55111 49572 55257 49606
rect 55077 49556 55111 49572
rect 12139 49366 12173 49382
rect 11993 49332 12139 49366
rect 12139 49316 12173 49332
rect 55077 49366 55111 49382
rect 55111 49332 55257 49366
rect 55077 49316 55111 49332
rect 12139 48816 12173 48832
rect 11993 48782 12139 48816
rect 12139 48766 12173 48782
rect 55077 48816 55111 48832
rect 55111 48782 55257 48816
rect 55077 48766 55111 48782
rect 12139 48576 12173 48592
rect 11993 48542 12139 48576
rect 12139 48526 12173 48542
rect 55077 48576 55111 48592
rect 55111 48542 55257 48576
rect 55077 48526 55111 48542
rect 12139 48026 12173 48042
rect 11993 47992 12139 48026
rect 12139 47976 12173 47992
rect 55077 48026 55111 48042
rect 55111 47992 55257 48026
rect 55077 47976 55111 47992
rect 12139 47786 12173 47802
rect 11993 47752 12139 47786
rect 12139 47736 12173 47752
rect 55077 47786 55111 47802
rect 55111 47752 55257 47786
rect 55077 47736 55111 47752
rect 12139 47236 12173 47252
rect 11993 47202 12139 47236
rect 12139 47186 12173 47202
rect 55077 47236 55111 47252
rect 55111 47202 55257 47236
rect 55077 47186 55111 47202
rect 12139 46996 12173 47012
rect 11993 46962 12139 46996
rect 12139 46946 12173 46962
rect 55077 46996 55111 47012
rect 55111 46962 55257 46996
rect 55077 46946 55111 46962
rect 12139 46446 12173 46462
rect 11993 46412 12139 46446
rect 12139 46396 12173 46412
rect 55077 46446 55111 46462
rect 55111 46412 55257 46446
rect 55077 46396 55111 46412
rect 12139 46206 12173 46222
rect 11993 46172 12139 46206
rect 12139 46156 12173 46172
rect 55077 46206 55111 46222
rect 55111 46172 55257 46206
rect 55077 46156 55111 46172
rect 12139 45656 12173 45672
rect 11993 45622 12139 45656
rect 12139 45606 12173 45622
rect 55077 45656 55111 45672
rect 55111 45622 55257 45656
rect 55077 45606 55111 45622
rect 12139 45416 12173 45432
rect 11993 45382 12139 45416
rect 12139 45366 12173 45382
rect 55077 45416 55111 45432
rect 55111 45382 55257 45416
rect 55077 45366 55111 45382
rect 12139 44866 12173 44882
rect 11993 44832 12139 44866
rect 12139 44816 12173 44832
rect 55077 44866 55111 44882
rect 55111 44832 55257 44866
rect 55077 44816 55111 44832
rect 12139 44626 12173 44642
rect 11993 44592 12139 44626
rect 12139 44576 12173 44592
rect 55077 44626 55111 44642
rect 55111 44592 55257 44626
rect 55077 44576 55111 44592
rect 12139 44076 12173 44092
rect 11993 44042 12139 44076
rect 12139 44026 12173 44042
rect 55077 44076 55111 44092
rect 55111 44042 55257 44076
rect 55077 44026 55111 44042
rect 12139 43836 12173 43852
rect 11993 43802 12139 43836
rect 12139 43786 12173 43802
rect 55077 43836 55111 43852
rect 55111 43802 55257 43836
rect 55077 43786 55111 43802
rect 12139 43286 12173 43302
rect 11993 43252 12139 43286
rect 12139 43236 12173 43252
rect 55077 43286 55111 43302
rect 55111 43252 55257 43286
rect 55077 43236 55111 43252
rect 12139 43046 12173 43062
rect 11993 43012 12139 43046
rect 12139 42996 12173 43012
rect 55077 43046 55111 43062
rect 55111 43012 55257 43046
rect 55077 42996 55111 43012
rect 12139 42496 12173 42512
rect 11993 42462 12139 42496
rect 12139 42446 12173 42462
rect 55077 42496 55111 42512
rect 55111 42462 55257 42496
rect 55077 42446 55111 42462
rect 12139 42256 12173 42272
rect 11993 42222 12139 42256
rect 12139 42206 12173 42222
rect 55077 42256 55111 42272
rect 55111 42222 55257 42256
rect 55077 42206 55111 42222
rect 12139 41706 12173 41722
rect 11993 41672 12139 41706
rect 12139 41656 12173 41672
rect 55077 41706 55111 41722
rect 55111 41672 55257 41706
rect 55077 41656 55111 41672
rect 12139 41466 12173 41482
rect 11993 41432 12139 41466
rect 12139 41416 12173 41432
rect 55077 41466 55111 41482
rect 55111 41432 55257 41466
rect 55077 41416 55111 41432
rect 12139 40916 12173 40932
rect 11993 40882 12139 40916
rect 12139 40866 12173 40882
rect 55077 40916 55111 40932
rect 55111 40882 55257 40916
rect 55077 40866 55111 40882
rect 12139 40676 12173 40692
rect 11993 40642 12139 40676
rect 12139 40626 12173 40642
rect 55077 40676 55111 40692
rect 55111 40642 55257 40676
rect 55077 40626 55111 40642
rect 12139 40126 12173 40142
rect 11993 40092 12139 40126
rect 12139 40076 12173 40092
rect 55077 40126 55111 40142
rect 55111 40092 55257 40126
rect 55077 40076 55111 40092
rect 12139 39886 12173 39902
rect 11993 39852 12139 39886
rect 12139 39836 12173 39852
rect 55077 39886 55111 39902
rect 55111 39852 55257 39886
rect 55077 39836 55111 39852
rect 12139 39336 12173 39352
rect 11993 39302 12139 39336
rect 12139 39286 12173 39302
rect 55077 39336 55111 39352
rect 55111 39302 55257 39336
rect 55077 39286 55111 39302
rect 12139 39096 12173 39112
rect 11993 39062 12139 39096
rect 12139 39046 12173 39062
rect 55077 39096 55111 39112
rect 55111 39062 55257 39096
rect 55077 39046 55111 39062
rect 12139 38546 12173 38562
rect 11993 38512 12139 38546
rect 12139 38496 12173 38512
rect 55077 38546 55111 38562
rect 55111 38512 55257 38546
rect 55077 38496 55111 38512
rect 12139 38306 12173 38322
rect 11993 38272 12139 38306
rect 12139 38256 12173 38272
rect 55077 38306 55111 38322
rect 55111 38272 55257 38306
rect 55077 38256 55111 38272
rect 12139 37756 12173 37772
rect 11993 37722 12139 37756
rect 12139 37706 12173 37722
rect 55077 37756 55111 37772
rect 55111 37722 55257 37756
rect 55077 37706 55111 37722
rect 12139 37516 12173 37532
rect 11993 37482 12139 37516
rect 12139 37466 12173 37482
rect 55077 37516 55111 37532
rect 55111 37482 55257 37516
rect 55077 37466 55111 37482
rect 12139 36966 12173 36982
rect 11993 36932 12139 36966
rect 12139 36916 12173 36932
rect 55077 36966 55111 36982
rect 55111 36932 55257 36966
rect 55077 36916 55111 36932
rect 12139 36726 12173 36742
rect 11993 36692 12139 36726
rect 12139 36676 12173 36692
rect 55077 36726 55111 36742
rect 55111 36692 55257 36726
rect 55077 36676 55111 36692
rect 12139 36176 12173 36192
rect 11993 36142 12139 36176
rect 12139 36126 12173 36142
rect 55077 36176 55111 36192
rect 55111 36142 55257 36176
rect 55077 36126 55111 36142
rect 12139 35936 12173 35952
rect 11993 35902 12139 35936
rect 12139 35886 12173 35902
rect 55077 35936 55111 35952
rect 55111 35902 55257 35936
rect 55077 35886 55111 35902
rect 12139 35386 12173 35402
rect 11993 35352 12139 35386
rect 12139 35336 12173 35352
rect 55077 35386 55111 35402
rect 55111 35352 55257 35386
rect 55077 35336 55111 35352
rect 12139 35146 12173 35162
rect 11993 35112 12139 35146
rect 12139 35096 12173 35112
rect 55077 35146 55111 35162
rect 55111 35112 55257 35146
rect 55077 35096 55111 35112
rect 12139 34596 12173 34612
rect 11993 34562 12139 34596
rect 12139 34546 12173 34562
rect 55077 34596 55111 34612
rect 55111 34562 55257 34596
rect 55077 34546 55111 34562
rect 12139 34356 12173 34372
rect 11993 34322 12139 34356
rect 12139 34306 12173 34322
rect 55077 34356 55111 34372
rect 55111 34322 55257 34356
rect 55077 34306 55111 34322
rect 12139 33806 12173 33822
rect 11993 33772 12139 33806
rect 12139 33756 12173 33772
rect 55077 33806 55111 33822
rect 55111 33772 55257 33806
rect 55077 33756 55111 33772
rect 12139 33566 12173 33582
rect 11993 33532 12139 33566
rect 12139 33516 12173 33532
rect 55077 33566 55111 33582
rect 55111 33532 55257 33566
rect 55077 33516 55111 33532
rect 12139 33016 12173 33032
rect 11993 32982 12139 33016
rect 12139 32966 12173 32982
rect 55077 33016 55111 33032
rect 55111 32982 55257 33016
rect 55077 32966 55111 32982
rect 12139 32776 12173 32792
rect 11993 32742 12139 32776
rect 12139 32726 12173 32742
rect 55077 32776 55111 32792
rect 55111 32742 55257 32776
rect 55077 32726 55111 32742
rect 12139 32226 12173 32242
rect 11993 32192 12139 32226
rect 12139 32176 12173 32192
rect 55077 32226 55111 32242
rect 55111 32192 55257 32226
rect 55077 32176 55111 32192
rect 12139 31986 12173 32002
rect 11993 31952 12139 31986
rect 12139 31936 12173 31952
rect 55077 31986 55111 32002
rect 55111 31952 55257 31986
rect 55077 31936 55111 31952
rect 12139 31436 12173 31452
rect 11993 31402 12139 31436
rect 12139 31386 12173 31402
rect 55077 31436 55111 31452
rect 55111 31402 55257 31436
rect 55077 31386 55111 31402
rect 12139 31196 12173 31212
rect 11993 31162 12139 31196
rect 12139 31146 12173 31162
rect 55077 31196 55111 31212
rect 55111 31162 55257 31196
rect 55077 31146 55111 31162
rect 12139 30646 12173 30662
rect 11993 30612 12139 30646
rect 12139 30596 12173 30612
rect 55077 30646 55111 30662
rect 55111 30612 55257 30646
rect 55077 30596 55111 30612
rect 12139 30406 12173 30422
rect 11993 30372 12139 30406
rect 12139 30356 12173 30372
rect 55077 30406 55111 30422
rect 55111 30372 55257 30406
rect 55077 30356 55111 30372
rect 12139 29856 12173 29872
rect 11993 29822 12139 29856
rect 12139 29806 12173 29822
rect 55077 29856 55111 29872
rect 55111 29822 55257 29856
rect 55077 29806 55111 29822
rect 12139 29616 12173 29632
rect 11993 29582 12139 29616
rect 12139 29566 12173 29582
rect 55077 29616 55111 29632
rect 55111 29582 55257 29616
rect 55077 29566 55111 29582
rect 12139 29066 12173 29082
rect 11993 29032 12139 29066
rect 12139 29016 12173 29032
rect 55077 29066 55111 29082
rect 55111 29032 55257 29066
rect 55077 29016 55111 29032
rect 12139 28826 12173 28842
rect 11993 28792 12139 28826
rect 12139 28776 12173 28792
rect 55077 28826 55111 28842
rect 55111 28792 55257 28826
rect 55077 28776 55111 28792
rect 12139 28276 12173 28292
rect 11993 28242 12139 28276
rect 12139 28226 12173 28242
rect 55077 28276 55111 28292
rect 55111 28242 55257 28276
rect 55077 28226 55111 28242
rect 12139 28036 12173 28052
rect 11993 28002 12139 28036
rect 12139 27986 12173 28002
rect 55077 28036 55111 28052
rect 55111 28002 55257 28036
rect 55077 27986 55111 28002
rect 12139 27486 12173 27502
rect 11993 27452 12139 27486
rect 12139 27436 12173 27452
rect 55077 27486 55111 27502
rect 55111 27452 55257 27486
rect 55077 27436 55111 27452
rect 12139 27246 12173 27262
rect 11993 27212 12139 27246
rect 12139 27196 12173 27212
rect 55077 27246 55111 27262
rect 55111 27212 55257 27246
rect 55077 27196 55111 27212
rect 12139 26696 12173 26712
rect 11993 26662 12139 26696
rect 12139 26646 12173 26662
rect 55077 26696 55111 26712
rect 55111 26662 55257 26696
rect 55077 26646 55111 26662
rect 12139 26456 12173 26472
rect 11993 26422 12139 26456
rect 12139 26406 12173 26422
rect 55077 26456 55111 26472
rect 55111 26422 55257 26456
rect 55077 26406 55111 26422
rect 12139 25906 12173 25922
rect 11993 25872 12139 25906
rect 12139 25856 12173 25872
rect 55077 25906 55111 25922
rect 55111 25872 55257 25906
rect 55077 25856 55111 25872
rect 12139 25666 12173 25682
rect 11993 25632 12139 25666
rect 12139 25616 12173 25632
rect 55077 25666 55111 25682
rect 55111 25632 55257 25666
rect 55077 25616 55111 25632
rect 12139 25116 12173 25132
rect 11993 25082 12139 25116
rect 12139 25066 12173 25082
rect 55077 25116 55111 25132
rect 55111 25082 55257 25116
rect 55077 25066 55111 25082
rect 12139 24876 12173 24892
rect 11993 24842 12139 24876
rect 12139 24826 12173 24842
rect 55077 24876 55111 24892
rect 55111 24842 55257 24876
rect 55077 24826 55111 24842
rect 12139 24326 12173 24342
rect 11993 24292 12139 24326
rect 12139 24276 12173 24292
rect 55077 24326 55111 24342
rect 55111 24292 55257 24326
rect 55077 24276 55111 24292
rect 12139 24086 12173 24102
rect 11993 24052 12139 24086
rect 12139 24036 12173 24052
rect 55077 24086 55111 24102
rect 55111 24052 55257 24086
rect 55077 24036 55111 24052
rect 12139 23536 12173 23552
rect 11993 23502 12139 23536
rect 12139 23486 12173 23502
rect 55077 23536 55111 23552
rect 55111 23502 55257 23536
rect 55077 23486 55111 23502
rect 12139 23296 12173 23312
rect 11993 23262 12139 23296
rect 12139 23246 12173 23262
rect 55077 23296 55111 23312
rect 55111 23262 55257 23296
rect 55077 23246 55111 23262
rect 12139 22746 12173 22762
rect 11993 22712 12139 22746
rect 12139 22696 12173 22712
rect 55077 22746 55111 22762
rect 55111 22712 55257 22746
rect 55077 22696 55111 22712
rect 12139 22506 12173 22522
rect 11993 22472 12139 22506
rect 12139 22456 12173 22472
rect 55077 22506 55111 22522
rect 55111 22472 55257 22506
rect 55077 22456 55111 22472
rect 12139 21956 12173 21972
rect 11993 21922 12139 21956
rect 12139 21906 12173 21922
rect 55077 21956 55111 21972
rect 55111 21922 55257 21956
rect 55077 21906 55111 21922
rect 12139 21716 12173 21732
rect 11993 21682 12139 21716
rect 12139 21666 12173 21682
rect 55077 21716 55111 21732
rect 55111 21682 55257 21716
rect 55077 21666 55111 21682
rect 12139 21166 12173 21182
rect 11993 21132 12139 21166
rect 12139 21116 12173 21132
rect 55077 21166 55111 21182
rect 55111 21132 55257 21166
rect 55077 21116 55111 21132
rect 12139 20926 12173 20942
rect 11993 20892 12139 20926
rect 12139 20876 12173 20892
rect 55077 20926 55111 20942
rect 55111 20892 55257 20926
rect 55077 20876 55111 20892
rect 12139 20376 12173 20392
rect 11993 20342 12139 20376
rect 12139 20326 12173 20342
rect 55077 20376 55111 20392
rect 55111 20342 55257 20376
rect 55077 20326 55111 20342
rect 12139 20136 12173 20152
rect 11993 20102 12139 20136
rect 12139 20086 12173 20102
rect 55077 20136 55111 20152
rect 55111 20102 55257 20136
rect 55077 20086 55111 20102
rect 12139 19586 12173 19602
rect 11993 19552 12139 19586
rect 12139 19536 12173 19552
rect 55077 19586 55111 19602
rect 55111 19552 55257 19586
rect 55077 19536 55111 19552
rect 12139 19346 12173 19362
rect 11993 19312 12139 19346
rect 12139 19296 12173 19312
rect 55077 19346 55111 19362
rect 55111 19312 55257 19346
rect 55077 19296 55111 19312
rect 12139 18796 12173 18812
rect 11993 18762 12139 18796
rect 12139 18746 12173 18762
rect 55077 18796 55111 18812
rect 55111 18762 55257 18796
rect 55077 18746 55111 18762
rect 12139 18556 12173 18572
rect 11993 18522 12139 18556
rect 12139 18506 12173 18522
rect 55077 18556 55111 18572
rect 55111 18522 55257 18556
rect 55077 18506 55111 18522
rect 12139 18006 12173 18022
rect 11993 17972 12139 18006
rect 12139 17956 12173 17972
rect 55077 18006 55111 18022
rect 55111 17972 55257 18006
rect 55077 17956 55111 17972
rect 12139 17766 12173 17782
rect 11993 17732 12139 17766
rect 12139 17716 12173 17732
rect 55077 17766 55111 17782
rect 55111 17732 55257 17766
rect 55077 17716 55111 17732
rect 12139 17216 12173 17232
rect 11993 17182 12139 17216
rect 12139 17166 12173 17182
rect 55077 17216 55111 17232
rect 55111 17182 55257 17216
rect 55077 17166 55111 17182
rect 12139 16976 12173 16992
rect 11993 16942 12139 16976
rect 12139 16926 12173 16942
rect 55077 16976 55111 16992
rect 55111 16942 55257 16976
rect 55077 16926 55111 16942
rect 12139 16426 12173 16442
rect 11993 16392 12139 16426
rect 12139 16376 12173 16392
rect 55077 16426 55111 16442
rect 55111 16392 55257 16426
rect 55077 16376 55111 16392
rect 12139 16186 12173 16202
rect 11993 16152 12139 16186
rect 12139 16136 12173 16152
rect 55077 16186 55111 16202
rect 55111 16152 55257 16186
rect 55077 16136 55111 16152
rect 12139 15636 12173 15652
rect 11993 15602 12139 15636
rect 12139 15586 12173 15602
rect 55077 15636 55111 15652
rect 55111 15602 55257 15636
rect 55077 15586 55111 15602
rect 12139 15396 12173 15412
rect 11993 15362 12139 15396
rect 12139 15346 12173 15362
rect 55077 15396 55111 15412
rect 55111 15362 55257 15396
rect 55077 15346 55111 15362
rect 12139 14846 12173 14862
rect 11993 14812 12139 14846
rect 12139 14796 12173 14812
rect 55077 14846 55111 14862
rect 55111 14812 55257 14846
rect 55077 14796 55111 14812
rect 12139 14606 12173 14622
rect 11993 14572 12139 14606
rect 12139 14556 12173 14572
rect 55077 14606 55111 14622
rect 55111 14572 55257 14606
rect 55077 14556 55111 14572
rect 12139 14056 12173 14072
rect 11993 14022 12139 14056
rect 12139 14006 12173 14022
rect 55077 14056 55111 14072
rect 55111 14022 55257 14056
rect 55077 14006 55111 14022
rect 12139 13816 12173 13832
rect 11993 13782 12139 13816
rect 12139 13766 12173 13782
rect 6849 10709 6883 10725
rect 6849 10659 6883 10675
rect 6849 9219 6883 9235
rect 6849 9169 6883 9185
rect 6849 7881 6883 7897
rect 6849 7831 6883 7847
rect 6849 6391 6883 6407
rect 6849 6341 6883 6357
rect 6849 5053 6883 5069
rect 6849 5003 6883 5019
rect 6849 3563 6883 3579
rect 6849 3513 6883 3529
rect 6849 2225 6883 2241
rect 6849 2175 6883 2191
rect 6849 735 6883 751
rect 6849 685 6883 701
<< viali >>
rect 60243 77663 60277 77697
rect 60243 76173 60277 76207
rect 60243 74835 60277 74869
rect 60243 73345 60277 73379
rect 60243 72007 60277 72041
rect 60243 70517 60277 70551
rect 60243 69179 60277 69213
rect 60243 67689 60277 67723
rect 55077 64582 55111 64616
rect 12139 64342 12173 64376
rect 55077 64342 55111 64376
rect 12139 63792 12173 63826
rect 55077 63792 55111 63826
rect 12139 63552 12173 63586
rect 55077 63552 55111 63586
rect 12139 63002 12173 63036
rect 55077 63002 55111 63036
rect 12139 62762 12173 62796
rect 55077 62762 55111 62796
rect 12139 62212 12173 62246
rect 55077 62212 55111 62246
rect 12139 61972 12173 62006
rect 55077 61972 55111 62006
rect 12139 61422 12173 61456
rect 55077 61422 55111 61456
rect 12139 61182 12173 61216
rect 55077 61182 55111 61216
rect 12139 60632 12173 60666
rect 55077 60632 55111 60666
rect 12139 60392 12173 60426
rect 55077 60392 55111 60426
rect 12139 59842 12173 59876
rect 55077 59842 55111 59876
rect 12139 59602 12173 59636
rect 55077 59602 55111 59636
rect 12139 59052 12173 59086
rect 55077 59052 55111 59086
rect 12139 58812 12173 58846
rect 55077 58812 55111 58846
rect 12139 58262 12173 58296
rect 55077 58262 55111 58296
rect 12139 58022 12173 58056
rect 55077 58022 55111 58056
rect 12139 57472 12173 57506
rect 55077 57472 55111 57506
rect 12139 57232 12173 57266
rect 55077 57232 55111 57266
rect 12139 56682 12173 56716
rect 55077 56682 55111 56716
rect 12139 56442 12173 56476
rect 55077 56442 55111 56476
rect 12139 55892 12173 55926
rect 55077 55892 55111 55926
rect 12139 55652 12173 55686
rect 55077 55652 55111 55686
rect 12139 55102 12173 55136
rect 55077 55102 55111 55136
rect 12139 54862 12173 54896
rect 55077 54862 55111 54896
rect 12139 54312 12173 54346
rect 55077 54312 55111 54346
rect 12139 54072 12173 54106
rect 55077 54072 55111 54106
rect 12139 53522 12173 53556
rect 55077 53522 55111 53556
rect 12139 53282 12173 53316
rect 55077 53282 55111 53316
rect 12139 52732 12173 52766
rect 55077 52732 55111 52766
rect 12139 52492 12173 52526
rect 55077 52492 55111 52526
rect 12139 51942 12173 51976
rect 55077 51942 55111 51976
rect 12139 51702 12173 51736
rect 55077 51702 55111 51736
rect 12139 51152 12173 51186
rect 55077 51152 55111 51186
rect 12139 50912 12173 50946
rect 55077 50912 55111 50946
rect 12139 50362 12173 50396
rect 55077 50362 55111 50396
rect 12139 50122 12173 50156
rect 55077 50122 55111 50156
rect 12139 49572 12173 49606
rect 55077 49572 55111 49606
rect 12139 49332 12173 49366
rect 55077 49332 55111 49366
rect 12139 48782 12173 48816
rect 55077 48782 55111 48816
rect 12139 48542 12173 48576
rect 55077 48542 55111 48576
rect 12139 47992 12173 48026
rect 55077 47992 55111 48026
rect 12139 47752 12173 47786
rect 55077 47752 55111 47786
rect 12139 47202 12173 47236
rect 55077 47202 55111 47236
rect 12139 46962 12173 46996
rect 55077 46962 55111 46996
rect 12139 46412 12173 46446
rect 55077 46412 55111 46446
rect 12139 46172 12173 46206
rect 55077 46172 55111 46206
rect 12139 45622 12173 45656
rect 55077 45622 55111 45656
rect 12139 45382 12173 45416
rect 55077 45382 55111 45416
rect 12139 44832 12173 44866
rect 55077 44832 55111 44866
rect 12139 44592 12173 44626
rect 55077 44592 55111 44626
rect 12139 44042 12173 44076
rect 55077 44042 55111 44076
rect 12139 43802 12173 43836
rect 55077 43802 55111 43836
rect 12139 43252 12173 43286
rect 55077 43252 55111 43286
rect 12139 43012 12173 43046
rect 55077 43012 55111 43046
rect 12139 42462 12173 42496
rect 55077 42462 55111 42496
rect 12139 42222 12173 42256
rect 55077 42222 55111 42256
rect 12139 41672 12173 41706
rect 55077 41672 55111 41706
rect 12139 41432 12173 41466
rect 55077 41432 55111 41466
rect 12139 40882 12173 40916
rect 55077 40882 55111 40916
rect 12139 40642 12173 40676
rect 55077 40642 55111 40676
rect 12139 40092 12173 40126
rect 55077 40092 55111 40126
rect 12139 39852 12173 39886
rect 55077 39852 55111 39886
rect 12139 39302 12173 39336
rect 55077 39302 55111 39336
rect 12139 39062 12173 39096
rect 55077 39062 55111 39096
rect 12139 38512 12173 38546
rect 55077 38512 55111 38546
rect 12139 38272 12173 38306
rect 55077 38272 55111 38306
rect 12139 37722 12173 37756
rect 55077 37722 55111 37756
rect 12139 37482 12173 37516
rect 55077 37482 55111 37516
rect 12139 36932 12173 36966
rect 55077 36932 55111 36966
rect 12139 36692 12173 36726
rect 55077 36692 55111 36726
rect 12139 36142 12173 36176
rect 55077 36142 55111 36176
rect 12139 35902 12173 35936
rect 55077 35902 55111 35936
rect 12139 35352 12173 35386
rect 55077 35352 55111 35386
rect 12139 35112 12173 35146
rect 55077 35112 55111 35146
rect 12139 34562 12173 34596
rect 55077 34562 55111 34596
rect 12139 34322 12173 34356
rect 55077 34322 55111 34356
rect 12139 33772 12173 33806
rect 55077 33772 55111 33806
rect 12139 33532 12173 33566
rect 55077 33532 55111 33566
rect 12139 32982 12173 33016
rect 55077 32982 55111 33016
rect 12139 32742 12173 32776
rect 55077 32742 55111 32776
rect 12139 32192 12173 32226
rect 55077 32192 55111 32226
rect 12139 31952 12173 31986
rect 55077 31952 55111 31986
rect 12139 31402 12173 31436
rect 55077 31402 55111 31436
rect 12139 31162 12173 31196
rect 55077 31162 55111 31196
rect 12139 30612 12173 30646
rect 55077 30612 55111 30646
rect 12139 30372 12173 30406
rect 55077 30372 55111 30406
rect 12139 29822 12173 29856
rect 55077 29822 55111 29856
rect 12139 29582 12173 29616
rect 55077 29582 55111 29616
rect 12139 29032 12173 29066
rect 55077 29032 55111 29066
rect 12139 28792 12173 28826
rect 55077 28792 55111 28826
rect 12139 28242 12173 28276
rect 55077 28242 55111 28276
rect 12139 28002 12173 28036
rect 55077 28002 55111 28036
rect 12139 27452 12173 27486
rect 55077 27452 55111 27486
rect 12139 27212 12173 27246
rect 55077 27212 55111 27246
rect 12139 26662 12173 26696
rect 55077 26662 55111 26696
rect 12139 26422 12173 26456
rect 55077 26422 55111 26456
rect 12139 25872 12173 25906
rect 55077 25872 55111 25906
rect 12139 25632 12173 25666
rect 55077 25632 55111 25666
rect 12139 25082 12173 25116
rect 55077 25082 55111 25116
rect 12139 24842 12173 24876
rect 55077 24842 55111 24876
rect 12139 24292 12173 24326
rect 55077 24292 55111 24326
rect 12139 24052 12173 24086
rect 55077 24052 55111 24086
rect 12139 23502 12173 23536
rect 55077 23502 55111 23536
rect 12139 23262 12173 23296
rect 55077 23262 55111 23296
rect 12139 22712 12173 22746
rect 55077 22712 55111 22746
rect 12139 22472 12173 22506
rect 55077 22472 55111 22506
rect 12139 21922 12173 21956
rect 55077 21922 55111 21956
rect 12139 21682 12173 21716
rect 55077 21682 55111 21716
rect 12139 21132 12173 21166
rect 55077 21132 55111 21166
rect 12139 20892 12173 20926
rect 55077 20892 55111 20926
rect 12139 20342 12173 20376
rect 55077 20342 55111 20376
rect 12139 20102 12173 20136
rect 55077 20102 55111 20136
rect 12139 19552 12173 19586
rect 55077 19552 55111 19586
rect 12139 19312 12173 19346
rect 55077 19312 55111 19346
rect 12139 18762 12173 18796
rect 55077 18762 55111 18796
rect 12139 18522 12173 18556
rect 55077 18522 55111 18556
rect 12139 17972 12173 18006
rect 55077 17972 55111 18006
rect 12139 17732 12173 17766
rect 55077 17732 55111 17766
rect 12139 17182 12173 17216
rect 55077 17182 55111 17216
rect 12139 16942 12173 16976
rect 55077 16942 55111 16976
rect 12139 16392 12173 16426
rect 55077 16392 55111 16426
rect 12139 16152 12173 16186
rect 55077 16152 55111 16186
rect 12139 15602 12173 15636
rect 55077 15602 55111 15636
rect 12139 15362 12173 15396
rect 55077 15362 55111 15396
rect 12139 14812 12173 14846
rect 55077 14812 55111 14846
rect 12139 14572 12173 14606
rect 55077 14572 55111 14606
rect 12139 14022 12173 14056
rect 55077 14022 55111 14056
rect 12139 13782 12173 13816
rect 6849 10675 6883 10709
rect 6849 9185 6883 9219
rect 6849 7847 6883 7881
rect 6849 6357 6883 6391
rect 6849 5019 6883 5053
rect 6849 3529 6883 3563
rect 6849 2191 6883 2225
rect 6849 701 6883 735
<< metal1 >>
rect 60228 77654 60234 77706
rect 60286 77654 60292 77706
rect 62770 77651 62816 77709
rect 60228 76164 60234 76216
rect 60286 76164 60292 76216
rect 62646 76161 62692 76219
rect 60228 74826 60234 74878
rect 60286 74826 60292 74878
rect 62522 74823 62568 74881
rect 60228 73336 60234 73388
rect 60286 73336 60292 73388
rect 60228 71998 60234 72050
rect 60286 71998 60292 72050
rect 13761 71461 13807 71715
rect 18753 71461 18799 71715
rect 23745 71461 23791 71715
rect 28737 71461 28783 71715
rect 33729 71461 33775 71715
rect 38721 71461 38767 71715
rect 43713 71461 43759 71715
rect 48705 71461 48751 71715
rect 60228 70508 60234 70560
rect 60286 70508 60292 70560
rect 60228 69170 60234 69222
rect 60286 69170 60292 69222
rect 60228 67680 60234 67732
rect 60286 67680 60292 67732
rect 53641 66373 53647 66425
rect 53699 66373 53705 66425
rect 53659 66275 53687 66373
rect 13723 65409 13751 65521
rect 14187 65409 14215 65521
rect 13723 65381 13983 65409
rect 13955 65269 13983 65381
rect 14027 65381 14215 65409
rect 14347 65409 14375 65521
rect 14811 65409 14839 65521
rect 14347 65381 14535 65409
rect 14027 65269 14055 65381
rect 14507 65269 14535 65381
rect 14579 65381 14839 65409
rect 14971 65409 14999 65521
rect 15435 65409 15463 65521
rect 14971 65381 15231 65409
rect 14579 65269 14607 65381
rect 15203 65269 15231 65381
rect 15275 65381 15463 65409
rect 15595 65409 15623 65521
rect 16059 65409 16087 65521
rect 15595 65381 15783 65409
rect 15275 65269 15303 65381
rect 15755 65269 15783 65381
rect 15827 65381 16087 65409
rect 16219 65409 16247 65521
rect 16683 65409 16711 65521
rect 16219 65381 16479 65409
rect 15827 65269 15855 65381
rect 16451 65269 16479 65381
rect 16523 65381 16711 65409
rect 16843 65409 16871 65521
rect 17307 65409 17335 65521
rect 16843 65381 17031 65409
rect 16523 65269 16551 65381
rect 17003 65269 17031 65381
rect 17075 65381 17335 65409
rect 17467 65409 17495 65521
rect 17931 65409 17959 65521
rect 17467 65381 17727 65409
rect 17075 65269 17103 65381
rect 17699 65269 17727 65381
rect 17771 65381 17959 65409
rect 18091 65409 18119 65521
rect 18555 65409 18583 65521
rect 18091 65381 18279 65409
rect 17771 65269 17799 65381
rect 18251 65269 18279 65381
rect 18323 65381 18583 65409
rect 18715 65409 18743 65521
rect 19179 65409 19207 65521
rect 18715 65381 18975 65409
rect 18323 65269 18351 65381
rect 18947 65269 18975 65381
rect 19019 65381 19207 65409
rect 19339 65409 19367 65521
rect 19803 65409 19831 65521
rect 19339 65381 19527 65409
rect 19019 65269 19047 65381
rect 19499 65269 19527 65381
rect 19571 65381 19831 65409
rect 19963 65409 19991 65521
rect 20427 65409 20455 65521
rect 19963 65381 20223 65409
rect 19571 65269 19599 65381
rect 20195 65269 20223 65381
rect 20267 65381 20455 65409
rect 20587 65409 20615 65521
rect 21051 65409 21079 65521
rect 20587 65381 20775 65409
rect 20267 65269 20295 65381
rect 20747 65269 20775 65381
rect 20819 65381 21079 65409
rect 21211 65409 21239 65521
rect 21675 65409 21703 65521
rect 21211 65381 21471 65409
rect 20819 65269 20847 65381
rect 21443 65269 21471 65381
rect 21515 65381 21703 65409
rect 21835 65409 21863 65521
rect 22299 65409 22327 65521
rect 21835 65381 22023 65409
rect 21515 65269 21543 65381
rect 21995 65269 22023 65381
rect 22067 65381 22327 65409
rect 22459 65409 22487 65521
rect 22923 65409 22951 65521
rect 22459 65381 22719 65409
rect 22067 65269 22095 65381
rect 22691 65269 22719 65381
rect 22763 65381 22951 65409
rect 23083 65409 23111 65521
rect 23547 65409 23575 65521
rect 23083 65381 23271 65409
rect 22763 65269 22791 65381
rect 23243 65269 23271 65381
rect 23315 65381 23575 65409
rect 23707 65409 23735 65521
rect 24171 65409 24199 65521
rect 23707 65381 23967 65409
rect 23315 65269 23343 65381
rect 23939 65269 23967 65381
rect 24011 65381 24199 65409
rect 24331 65409 24359 65521
rect 24795 65409 24823 65521
rect 24331 65381 24519 65409
rect 24011 65269 24039 65381
rect 24491 65269 24519 65381
rect 24563 65381 24823 65409
rect 24955 65409 24983 65521
rect 25419 65409 25447 65521
rect 24955 65381 25215 65409
rect 24563 65269 24591 65381
rect 25187 65269 25215 65381
rect 25259 65381 25447 65409
rect 25579 65409 25607 65521
rect 26043 65409 26071 65521
rect 25579 65381 25767 65409
rect 25259 65269 25287 65381
rect 25739 65269 25767 65381
rect 25811 65381 26071 65409
rect 26203 65409 26231 65521
rect 26667 65409 26695 65521
rect 26203 65381 26463 65409
rect 25811 65269 25839 65381
rect 26435 65269 26463 65381
rect 26507 65381 26695 65409
rect 26827 65409 26855 65521
rect 27291 65409 27319 65521
rect 26827 65381 27015 65409
rect 26507 65269 26535 65381
rect 26987 65269 27015 65381
rect 27059 65381 27319 65409
rect 27451 65409 27479 65521
rect 27915 65409 27943 65521
rect 27451 65381 27711 65409
rect 27059 65269 27087 65381
rect 27683 65269 27711 65381
rect 27755 65381 27943 65409
rect 28075 65409 28103 65521
rect 28539 65409 28567 65521
rect 28075 65381 28263 65409
rect 27755 65269 27783 65381
rect 28235 65269 28263 65381
rect 28307 65381 28567 65409
rect 28699 65409 28727 65521
rect 29163 65409 29191 65521
rect 28699 65381 28959 65409
rect 28307 65269 28335 65381
rect 28931 65269 28959 65381
rect 29003 65381 29191 65409
rect 29323 65409 29351 65521
rect 29787 65409 29815 65521
rect 29323 65381 29511 65409
rect 29003 65269 29031 65381
rect 29483 65269 29511 65381
rect 29555 65381 29815 65409
rect 29947 65409 29975 65521
rect 30411 65409 30439 65521
rect 29947 65381 30207 65409
rect 29555 65269 29583 65381
rect 30179 65269 30207 65381
rect 30251 65381 30439 65409
rect 30571 65409 30599 65521
rect 31035 65409 31063 65521
rect 30571 65381 30759 65409
rect 30251 65269 30279 65381
rect 30731 65269 30759 65381
rect 30803 65381 31063 65409
rect 31195 65409 31223 65521
rect 31659 65409 31687 65521
rect 31195 65381 31455 65409
rect 30803 65269 30831 65381
rect 31427 65269 31455 65381
rect 31499 65381 31687 65409
rect 31819 65409 31847 65521
rect 32283 65409 32311 65521
rect 31819 65381 32007 65409
rect 31499 65269 31527 65381
rect 31979 65269 32007 65381
rect 32051 65381 32311 65409
rect 32443 65409 32471 65521
rect 32907 65409 32935 65521
rect 32443 65381 32703 65409
rect 32051 65269 32079 65381
rect 32675 65269 32703 65381
rect 32747 65381 32935 65409
rect 33067 65409 33095 65521
rect 33531 65409 33559 65521
rect 33067 65381 33255 65409
rect 32747 65269 32775 65381
rect 33227 65269 33255 65381
rect 33299 65381 33559 65409
rect 33691 65409 33719 65521
rect 34155 65409 34183 65521
rect 33691 65381 33951 65409
rect 33299 65269 33327 65381
rect 33923 65269 33951 65381
rect 33995 65381 34183 65409
rect 34315 65409 34343 65521
rect 34779 65409 34807 65521
rect 34315 65381 34503 65409
rect 33995 65269 34023 65381
rect 34475 65269 34503 65381
rect 34547 65381 34807 65409
rect 34939 65409 34967 65521
rect 35403 65409 35431 65521
rect 34939 65381 35199 65409
rect 34547 65269 34575 65381
rect 35171 65269 35199 65381
rect 35243 65381 35431 65409
rect 35563 65409 35591 65521
rect 36027 65409 36055 65521
rect 35563 65381 35751 65409
rect 35243 65269 35271 65381
rect 35723 65269 35751 65381
rect 35795 65381 36055 65409
rect 36187 65409 36215 65521
rect 36651 65409 36679 65521
rect 36187 65381 36447 65409
rect 35795 65269 35823 65381
rect 36419 65269 36447 65381
rect 36491 65381 36679 65409
rect 36811 65409 36839 65521
rect 37275 65409 37303 65521
rect 36811 65381 36999 65409
rect 36491 65269 36519 65381
rect 36971 65269 36999 65381
rect 37043 65381 37303 65409
rect 37435 65409 37463 65521
rect 37899 65409 37927 65521
rect 37435 65381 37695 65409
rect 37043 65269 37071 65381
rect 37667 65269 37695 65381
rect 37739 65381 37927 65409
rect 38059 65409 38087 65521
rect 38523 65409 38551 65521
rect 38059 65381 38247 65409
rect 37739 65269 37767 65381
rect 38219 65269 38247 65381
rect 38291 65381 38551 65409
rect 38683 65409 38711 65521
rect 39147 65409 39175 65521
rect 38683 65381 38943 65409
rect 38291 65269 38319 65381
rect 38915 65269 38943 65381
rect 38987 65381 39175 65409
rect 39307 65409 39335 65521
rect 39771 65409 39799 65521
rect 39307 65381 39495 65409
rect 38987 65269 39015 65381
rect 39467 65269 39495 65381
rect 39539 65381 39799 65409
rect 39931 65409 39959 65521
rect 40395 65409 40423 65521
rect 39931 65381 40191 65409
rect 39539 65269 39567 65381
rect 40163 65269 40191 65381
rect 40235 65381 40423 65409
rect 40555 65409 40583 65521
rect 41019 65409 41047 65521
rect 40555 65381 40743 65409
rect 40235 65269 40263 65381
rect 40715 65269 40743 65381
rect 40787 65381 41047 65409
rect 41179 65409 41207 65521
rect 41643 65409 41671 65521
rect 41179 65381 41439 65409
rect 40787 65269 40815 65381
rect 41411 65269 41439 65381
rect 41483 65381 41671 65409
rect 41803 65409 41831 65521
rect 42267 65409 42295 65521
rect 41803 65381 41991 65409
rect 41483 65269 41511 65381
rect 41963 65269 41991 65381
rect 42035 65381 42295 65409
rect 42427 65409 42455 65521
rect 42891 65409 42919 65521
rect 42427 65381 42687 65409
rect 42035 65269 42063 65381
rect 42659 65269 42687 65381
rect 42731 65381 42919 65409
rect 43051 65409 43079 65521
rect 43515 65409 43543 65521
rect 43051 65381 43239 65409
rect 42731 65269 42759 65381
rect 43211 65269 43239 65381
rect 43283 65381 43543 65409
rect 43675 65409 43703 65521
rect 44139 65409 44167 65521
rect 43675 65381 43935 65409
rect 43283 65269 43311 65381
rect 43907 65269 43935 65381
rect 43979 65381 44167 65409
rect 44299 65409 44327 65521
rect 44763 65409 44791 65521
rect 44299 65381 44487 65409
rect 43979 65269 44007 65381
rect 44459 65269 44487 65381
rect 44531 65381 44791 65409
rect 44923 65409 44951 65521
rect 45387 65409 45415 65521
rect 44923 65381 45183 65409
rect 44531 65269 44559 65381
rect 45155 65269 45183 65381
rect 45227 65381 45415 65409
rect 45547 65409 45575 65521
rect 46011 65409 46039 65521
rect 45547 65381 45735 65409
rect 45227 65269 45255 65381
rect 45707 65269 45735 65381
rect 45779 65381 46039 65409
rect 46171 65409 46199 65521
rect 46635 65409 46663 65521
rect 46171 65381 46431 65409
rect 45779 65269 45807 65381
rect 46403 65269 46431 65381
rect 46475 65381 46663 65409
rect 46795 65409 46823 65521
rect 47259 65409 47287 65521
rect 46795 65381 46983 65409
rect 46475 65269 46503 65381
rect 46955 65269 46983 65381
rect 47027 65381 47287 65409
rect 47419 65409 47447 65521
rect 47883 65409 47911 65521
rect 47419 65381 47679 65409
rect 47027 65269 47055 65381
rect 47651 65269 47679 65381
rect 47723 65381 47911 65409
rect 48043 65409 48071 65521
rect 48507 65409 48535 65521
rect 48043 65381 48231 65409
rect 47723 65269 47751 65381
rect 48203 65269 48231 65381
rect 48275 65381 48535 65409
rect 48667 65409 48695 65521
rect 49131 65409 49159 65521
rect 48667 65381 48927 65409
rect 48275 65269 48303 65381
rect 48899 65269 48927 65381
rect 48971 65381 49159 65409
rect 49291 65409 49319 65521
rect 49755 65409 49783 65521
rect 49291 65381 49479 65409
rect 48971 65269 48999 65381
rect 49451 65269 49479 65381
rect 49523 65381 49783 65409
rect 49915 65409 49943 65521
rect 50379 65409 50407 65521
rect 49915 65381 50175 65409
rect 49523 65269 49551 65381
rect 50147 65269 50175 65381
rect 50219 65381 50407 65409
rect 50539 65409 50567 65521
rect 51003 65409 51031 65521
rect 50539 65381 50727 65409
rect 50219 65269 50247 65381
rect 50699 65269 50727 65381
rect 50771 65381 51031 65409
rect 51163 65409 51191 65521
rect 51627 65409 51655 65521
rect 51163 65381 51423 65409
rect 50771 65269 50799 65381
rect 51395 65269 51423 65381
rect 51467 65381 51655 65409
rect 51787 65409 51815 65521
rect 52251 65409 52279 65521
rect 51787 65381 51975 65409
rect 51467 65269 51495 65381
rect 51947 65269 51975 65381
rect 52019 65381 52279 65409
rect 52411 65409 52439 65521
rect 52875 65409 52903 65521
rect 52411 65381 52671 65409
rect 52019 65269 52047 65381
rect 52643 65269 52671 65381
rect 52715 65381 52903 65409
rect 53035 65409 53063 65521
rect 53499 65409 53527 65521
rect 53035 65381 53223 65409
rect 52715 65269 52743 65381
rect 53195 65269 53223 65381
rect 53267 65381 53527 65409
rect 53659 65409 53687 65521
rect 54123 65409 54151 65521
rect 53659 65381 53919 65409
rect 53267 65269 53295 65381
rect 53891 65269 53919 65381
rect 53963 65381 54151 65409
rect 53963 65269 53991 65381
rect 55062 64573 55068 64625
rect 55120 64573 55126 64625
rect 12124 64333 12130 64385
rect 12182 64333 12188 64385
rect 55062 64333 55068 64385
rect 55120 64333 55126 64385
rect 12124 63783 12130 63835
rect 12182 63783 12188 63835
rect 55062 63783 55068 63835
rect 55120 63783 55126 63835
rect 12124 63543 12130 63595
rect 12182 63543 12188 63595
rect 55062 63543 55068 63595
rect 55120 63543 55126 63595
rect 12124 62993 12130 63045
rect 12182 62993 12188 63045
rect 55062 62993 55068 63045
rect 55120 62993 55126 63045
rect 12124 62753 12130 62805
rect 12182 62753 12188 62805
rect 55062 62753 55068 62805
rect 55120 62753 55126 62805
rect 12124 62203 12130 62255
rect 12182 62203 12188 62255
rect 55062 62203 55068 62255
rect 55120 62203 55126 62255
rect 12124 61963 12130 62015
rect 12182 61963 12188 62015
rect 55062 61963 55068 62015
rect 55120 61963 55126 62015
rect 12124 61413 12130 61465
rect 12182 61413 12188 61465
rect 55062 61413 55068 61465
rect 55120 61413 55126 61465
rect 12124 61173 12130 61225
rect 12182 61173 12188 61225
rect 55062 61173 55068 61225
rect 55120 61173 55126 61225
rect 12124 60623 12130 60675
rect 12182 60623 12188 60675
rect 55062 60623 55068 60675
rect 55120 60623 55126 60675
rect 12124 60383 12130 60435
rect 12182 60383 12188 60435
rect 55062 60383 55068 60435
rect 55120 60383 55126 60435
rect 12124 59833 12130 59885
rect 12182 59833 12188 59885
rect 55062 59833 55068 59885
rect 55120 59833 55126 59885
rect 12124 59593 12130 59645
rect 12182 59593 12188 59645
rect 55062 59593 55068 59645
rect 55120 59593 55126 59645
rect 12124 59043 12130 59095
rect 12182 59043 12188 59095
rect 55062 59043 55068 59095
rect 55120 59043 55126 59095
rect 12124 58803 12130 58855
rect 12182 58803 12188 58855
rect 55062 58803 55068 58855
rect 55120 58803 55126 58855
rect 12124 58253 12130 58305
rect 12182 58253 12188 58305
rect 55062 58253 55068 58305
rect 55120 58253 55126 58305
rect 12124 58013 12130 58065
rect 12182 58013 12188 58065
rect 55062 58013 55068 58065
rect 55120 58013 55126 58065
rect 12124 57463 12130 57515
rect 12182 57463 12188 57515
rect 55062 57463 55068 57515
rect 55120 57463 55126 57515
rect 12124 57223 12130 57275
rect 12182 57223 12188 57275
rect 55062 57223 55068 57275
rect 55120 57223 55126 57275
rect 12124 56673 12130 56725
rect 12182 56673 12188 56725
rect 55062 56673 55068 56725
rect 55120 56673 55126 56725
rect 12124 56433 12130 56485
rect 12182 56433 12188 56485
rect 55062 56433 55068 56485
rect 55120 56433 55126 56485
rect 12124 55883 12130 55935
rect 12182 55883 12188 55935
rect 55062 55883 55068 55935
rect 55120 55883 55126 55935
rect 12124 55643 12130 55695
rect 12182 55643 12188 55695
rect 55062 55643 55068 55695
rect 55120 55643 55126 55695
rect 12124 55093 12130 55145
rect 12182 55093 12188 55145
rect 55062 55093 55068 55145
rect 55120 55093 55126 55145
rect 12124 54853 12130 54905
rect 12182 54853 12188 54905
rect 55062 54853 55068 54905
rect 55120 54853 55126 54905
rect 12124 54303 12130 54355
rect 12182 54303 12188 54355
rect 55062 54303 55068 54355
rect 55120 54303 55126 54355
rect 12124 54063 12130 54115
rect 12182 54063 12188 54115
rect 55062 54063 55068 54115
rect 55120 54063 55126 54115
rect 12124 53513 12130 53565
rect 12182 53513 12188 53565
rect 55062 53513 55068 53565
rect 55120 53513 55126 53565
rect 12124 53273 12130 53325
rect 12182 53273 12188 53325
rect 55062 53273 55068 53325
rect 55120 53273 55126 53325
rect 12124 52723 12130 52775
rect 12182 52723 12188 52775
rect 55062 52723 55068 52775
rect 55120 52723 55126 52775
rect 12124 52483 12130 52535
rect 12182 52483 12188 52535
rect 55062 52483 55068 52535
rect 55120 52483 55126 52535
rect 12124 51933 12130 51985
rect 12182 51933 12188 51985
rect 55062 51933 55068 51985
rect 55120 51933 55126 51985
rect 12124 51693 12130 51745
rect 12182 51693 12188 51745
rect 55062 51693 55068 51745
rect 55120 51693 55126 51745
rect 12124 51143 12130 51195
rect 12182 51143 12188 51195
rect 55062 51143 55068 51195
rect 55120 51143 55126 51195
rect 12124 50903 12130 50955
rect 12182 50903 12188 50955
rect 55062 50903 55068 50955
rect 55120 50903 55126 50955
rect 12124 50353 12130 50405
rect 12182 50353 12188 50405
rect 55062 50353 55068 50405
rect 55120 50353 55126 50405
rect 12124 50113 12130 50165
rect 12182 50113 12188 50165
rect 55062 50113 55068 50165
rect 55120 50113 55126 50165
rect 12124 49563 12130 49615
rect 12182 49563 12188 49615
rect 55062 49563 55068 49615
rect 55120 49563 55126 49615
rect 12124 49323 12130 49375
rect 12182 49323 12188 49375
rect 55062 49323 55068 49375
rect 55120 49323 55126 49375
rect 12124 48773 12130 48825
rect 12182 48773 12188 48825
rect 55062 48773 55068 48825
rect 55120 48773 55126 48825
rect 12124 48533 12130 48585
rect 12182 48533 12188 48585
rect 55062 48533 55068 48585
rect 55120 48533 55126 48585
rect 12124 47983 12130 48035
rect 12182 47983 12188 48035
rect 55062 47983 55068 48035
rect 55120 47983 55126 48035
rect 12124 47743 12130 47795
rect 12182 47743 12188 47795
rect 55062 47743 55068 47795
rect 55120 47743 55126 47795
rect 12124 47193 12130 47245
rect 12182 47193 12188 47245
rect 55062 47193 55068 47245
rect 55120 47193 55126 47245
rect 12124 46953 12130 47005
rect 12182 46953 12188 47005
rect 55062 46953 55068 47005
rect 55120 46953 55126 47005
rect 12124 46403 12130 46455
rect 12182 46403 12188 46455
rect 55062 46403 55068 46455
rect 55120 46403 55126 46455
rect 12124 46163 12130 46215
rect 12182 46163 12188 46215
rect 55062 46163 55068 46215
rect 55120 46163 55126 46215
rect 12124 45613 12130 45665
rect 12182 45613 12188 45665
rect 55062 45613 55068 45665
rect 55120 45613 55126 45665
rect 12124 45373 12130 45425
rect 12182 45373 12188 45425
rect 55062 45373 55068 45425
rect 55120 45373 55126 45425
rect 12124 44823 12130 44875
rect 12182 44823 12188 44875
rect 55062 44823 55068 44875
rect 55120 44823 55126 44875
rect 12124 44583 12130 44635
rect 12182 44583 12188 44635
rect 55062 44583 55068 44635
rect 55120 44583 55126 44635
rect 12124 44033 12130 44085
rect 12182 44033 12188 44085
rect 55062 44033 55068 44085
rect 55120 44033 55126 44085
rect 12124 43793 12130 43845
rect 12182 43793 12188 43845
rect 55062 43793 55068 43845
rect 55120 43793 55126 43845
rect 12124 43243 12130 43295
rect 12182 43243 12188 43295
rect 55062 43243 55068 43295
rect 55120 43243 55126 43295
rect 12124 43003 12130 43055
rect 12182 43003 12188 43055
rect 55062 43003 55068 43055
rect 55120 43003 55126 43055
rect 12124 42453 12130 42505
rect 12182 42453 12188 42505
rect 55062 42453 55068 42505
rect 55120 42453 55126 42505
rect 12124 42213 12130 42265
rect 12182 42213 12188 42265
rect 55062 42213 55068 42265
rect 55120 42213 55126 42265
rect 12124 41663 12130 41715
rect 12182 41663 12188 41715
rect 55062 41663 55068 41715
rect 55120 41663 55126 41715
rect 12124 41423 12130 41475
rect 12182 41423 12188 41475
rect 55062 41423 55068 41475
rect 55120 41423 55126 41475
rect 12124 40873 12130 40925
rect 12182 40873 12188 40925
rect 55062 40873 55068 40925
rect 55120 40873 55126 40925
rect 12124 40633 12130 40685
rect 12182 40633 12188 40685
rect 55062 40633 55068 40685
rect 55120 40633 55126 40685
rect 12124 40083 12130 40135
rect 12182 40083 12188 40135
rect 55062 40083 55068 40135
rect 55120 40083 55126 40135
rect 12124 39843 12130 39895
rect 12182 39843 12188 39895
rect 55062 39843 55068 39895
rect 55120 39843 55126 39895
rect 12124 39293 12130 39345
rect 12182 39293 12188 39345
rect 55062 39293 55068 39345
rect 55120 39293 55126 39345
rect 12124 39053 12130 39105
rect 12182 39053 12188 39105
rect 55062 39053 55068 39105
rect 55120 39053 55126 39105
rect 12124 38503 12130 38555
rect 12182 38503 12188 38555
rect 55062 38503 55068 38555
rect 55120 38503 55126 38555
rect 12124 38263 12130 38315
rect 12182 38263 12188 38315
rect 55062 38263 55068 38315
rect 55120 38263 55126 38315
rect 12124 37713 12130 37765
rect 12182 37713 12188 37765
rect 55062 37713 55068 37765
rect 55120 37713 55126 37765
rect 12124 37473 12130 37525
rect 12182 37473 12188 37525
rect 55062 37473 55068 37525
rect 55120 37473 55126 37525
rect 12124 36923 12130 36975
rect 12182 36923 12188 36975
rect 55062 36923 55068 36975
rect 55120 36923 55126 36975
rect 12124 36683 12130 36735
rect 12182 36683 12188 36735
rect 55062 36683 55068 36735
rect 55120 36683 55126 36735
rect 12124 36133 12130 36185
rect 12182 36133 12188 36185
rect 55062 36133 55068 36185
rect 55120 36133 55126 36185
rect 12124 35893 12130 35945
rect 12182 35893 12188 35945
rect 55062 35893 55068 35945
rect 55120 35893 55126 35945
rect 12124 35343 12130 35395
rect 12182 35343 12188 35395
rect 55062 35343 55068 35395
rect 55120 35343 55126 35395
rect 12124 35103 12130 35155
rect 12182 35103 12188 35155
rect 55062 35103 55068 35155
rect 55120 35103 55126 35155
rect 12124 34553 12130 34605
rect 12182 34553 12188 34605
rect 55062 34553 55068 34605
rect 55120 34553 55126 34605
rect 12124 34313 12130 34365
rect 12182 34313 12188 34365
rect 55062 34313 55068 34365
rect 55120 34313 55126 34365
rect 12124 33763 12130 33815
rect 12182 33763 12188 33815
rect 55062 33763 55068 33815
rect 55120 33763 55126 33815
rect 12124 33523 12130 33575
rect 12182 33523 12188 33575
rect 55062 33523 55068 33575
rect 55120 33523 55126 33575
rect 12124 32973 12130 33025
rect 12182 32973 12188 33025
rect 55062 32973 55068 33025
rect 55120 32973 55126 33025
rect 12124 32733 12130 32785
rect 12182 32733 12188 32785
rect 55062 32733 55068 32785
rect 55120 32733 55126 32785
rect 12124 32183 12130 32235
rect 12182 32183 12188 32235
rect 55062 32183 55068 32235
rect 55120 32183 55126 32235
rect 12124 31943 12130 31995
rect 12182 31943 12188 31995
rect 55062 31943 55068 31995
rect 55120 31943 55126 31995
rect 12124 31393 12130 31445
rect 12182 31393 12188 31445
rect 55062 31393 55068 31445
rect 55120 31393 55126 31445
rect 12124 31153 12130 31205
rect 12182 31153 12188 31205
rect 55062 31153 55068 31205
rect 55120 31153 55126 31205
rect 12124 30603 12130 30655
rect 12182 30603 12188 30655
rect 55062 30603 55068 30655
rect 55120 30603 55126 30655
rect 12124 30363 12130 30415
rect 12182 30363 12188 30415
rect 55062 30363 55068 30415
rect 55120 30363 55126 30415
rect 12124 29813 12130 29865
rect 12182 29813 12188 29865
rect 55062 29813 55068 29865
rect 55120 29813 55126 29865
rect 12124 29573 12130 29625
rect 12182 29573 12188 29625
rect 55062 29573 55068 29625
rect 55120 29573 55126 29625
rect 12124 29023 12130 29075
rect 12182 29023 12188 29075
rect 55062 29023 55068 29075
rect 55120 29023 55126 29075
rect 12124 28783 12130 28835
rect 12182 28783 12188 28835
rect 55062 28783 55068 28835
rect 55120 28783 55126 28835
rect 12124 28233 12130 28285
rect 12182 28233 12188 28285
rect 55062 28233 55068 28285
rect 55120 28233 55126 28285
rect 12124 27993 12130 28045
rect 12182 27993 12188 28045
rect 55062 27993 55068 28045
rect 55120 27993 55126 28045
rect 12124 27443 12130 27495
rect 12182 27443 12188 27495
rect 55062 27443 55068 27495
rect 55120 27443 55126 27495
rect 12124 27203 12130 27255
rect 12182 27203 12188 27255
rect 55062 27203 55068 27255
rect 55120 27203 55126 27255
rect 12124 26653 12130 26705
rect 12182 26653 12188 26705
rect 55062 26653 55068 26705
rect 55120 26653 55126 26705
rect 12124 26413 12130 26465
rect 12182 26413 12188 26465
rect 55062 26413 55068 26465
rect 55120 26413 55126 26465
rect 12124 25863 12130 25915
rect 12182 25863 12188 25915
rect 55062 25863 55068 25915
rect 55120 25863 55126 25915
rect 12124 25623 12130 25675
rect 12182 25623 12188 25675
rect 55062 25623 55068 25675
rect 55120 25623 55126 25675
rect 12124 25073 12130 25125
rect 12182 25073 12188 25125
rect 55062 25073 55068 25125
rect 55120 25073 55126 25125
rect 12124 24833 12130 24885
rect 12182 24833 12188 24885
rect 55062 24833 55068 24885
rect 55120 24833 55126 24885
rect 12124 24283 12130 24335
rect 12182 24283 12188 24335
rect 55062 24283 55068 24335
rect 55120 24283 55126 24335
rect 12124 24043 12130 24095
rect 12182 24043 12188 24095
rect 55062 24043 55068 24095
rect 55120 24043 55126 24095
rect 12124 23493 12130 23545
rect 12182 23493 12188 23545
rect 55062 23493 55068 23545
rect 55120 23493 55126 23545
rect 12124 23253 12130 23305
rect 12182 23253 12188 23305
rect 55062 23253 55068 23305
rect 55120 23253 55126 23305
rect 12124 22703 12130 22755
rect 12182 22703 12188 22755
rect 55062 22703 55068 22755
rect 55120 22703 55126 22755
rect 12124 22463 12130 22515
rect 12182 22463 12188 22515
rect 55062 22463 55068 22515
rect 55120 22463 55126 22515
rect 12124 21913 12130 21965
rect 12182 21913 12188 21965
rect 55062 21913 55068 21965
rect 55120 21913 55126 21965
rect 19 13919 47 21819
rect 99 13919 127 21819
rect 179 13919 207 21819
rect 259 13919 287 21819
rect 339 13919 367 21819
rect 419 13919 447 21819
rect 499 13919 527 21819
rect 12124 21673 12130 21725
rect 12182 21673 12188 21725
rect 55062 21673 55068 21725
rect 55120 21673 55126 21725
rect 12124 21123 12130 21175
rect 12182 21123 12188 21175
rect 55062 21123 55068 21175
rect 55120 21123 55126 21175
rect 12124 20883 12130 20935
rect 12182 20883 12188 20935
rect 55062 20883 55068 20935
rect 55120 20883 55126 20935
rect 12124 20333 12130 20385
rect 12182 20333 12188 20385
rect 55062 20333 55068 20385
rect 55120 20333 55126 20385
rect 12124 20093 12130 20145
rect 12182 20093 12188 20145
rect 55062 20093 55068 20145
rect 55120 20093 55126 20145
rect 12124 19543 12130 19595
rect 12182 19543 12188 19595
rect 55062 19543 55068 19595
rect 55120 19543 55126 19595
rect 12124 19303 12130 19355
rect 12182 19303 12188 19355
rect 55062 19303 55068 19355
rect 55120 19303 55126 19355
rect 12124 18753 12130 18805
rect 12182 18753 12188 18805
rect 55062 18753 55068 18805
rect 55120 18753 55126 18805
rect 12124 18513 12130 18565
rect 12182 18513 12188 18565
rect 55062 18513 55068 18565
rect 55120 18513 55126 18565
rect 12124 17963 12130 18015
rect 12182 17963 12188 18015
rect 55062 17963 55068 18015
rect 55120 17963 55126 18015
rect 12124 17723 12130 17775
rect 12182 17723 12188 17775
rect 55062 17723 55068 17775
rect 55120 17723 55126 17775
rect 12124 17173 12130 17225
rect 12182 17173 12188 17225
rect 55062 17173 55068 17225
rect 55120 17173 55126 17225
rect 12124 16933 12130 16985
rect 12182 16933 12188 16985
rect 55062 16933 55068 16985
rect 55120 16933 55126 16985
rect 12124 16383 12130 16435
rect 12182 16383 12188 16435
rect 55062 16383 55068 16435
rect 55120 16383 55126 16435
rect 12124 16143 12130 16195
rect 12182 16143 12188 16195
rect 55062 16143 55068 16195
rect 55120 16143 55126 16195
rect 12124 15593 12130 15645
rect 12182 15593 12188 15645
rect 55062 15593 55068 15645
rect 55120 15593 55126 15645
rect 12124 15353 12130 15405
rect 12182 15353 12188 15405
rect 55062 15353 55068 15405
rect 55120 15353 55126 15405
rect 12124 14803 12130 14855
rect 12182 14803 12188 14855
rect 55062 14803 55068 14855
rect 55120 14803 55126 14855
rect 12124 14563 12130 14615
rect 12182 14563 12188 14615
rect 55062 14563 55068 14615
rect 55120 14563 55126 14615
rect 12124 14013 12130 14065
rect 12182 14013 12188 14065
rect 55062 14013 55068 14065
rect 55120 14013 55126 14065
rect 66723 13919 66751 21819
rect 66803 13919 66831 21819
rect 66883 13919 66911 21819
rect 66963 13919 66991 21819
rect 67043 13919 67071 21819
rect 67123 13919 67151 21819
rect 67203 13919 67231 21819
rect 12124 13773 12130 13825
rect 12182 13773 12188 13825
rect 13475 13017 13503 13129
rect 13099 12989 13503 13017
rect 13547 13017 13575 13129
rect 13739 13017 13767 13129
rect 13547 12989 13591 13017
rect 13099 12877 13127 12989
rect 13563 12877 13591 12989
rect 13723 12989 13767 13017
rect 13811 13017 13839 13129
rect 14723 13017 14751 13129
rect 13811 12989 14215 13017
rect 13723 12877 13751 12989
rect 14187 12877 14215 12989
rect 14347 12989 14751 13017
rect 14795 13017 14823 13129
rect 14987 13017 15015 13129
rect 14795 12989 14839 13017
rect 14347 12877 14375 12989
rect 14811 12877 14839 12989
rect 14971 12989 15015 13017
rect 15059 13017 15087 13129
rect 15971 13017 15999 13129
rect 15059 12989 15463 13017
rect 14971 12877 14999 12989
rect 15435 12877 15463 12989
rect 15595 12989 15999 13017
rect 16043 13017 16071 13129
rect 16235 13017 16263 13129
rect 16043 12989 16087 13017
rect 15595 12877 15623 12989
rect 16059 12877 16087 12989
rect 16219 12989 16263 13017
rect 16307 13017 16335 13129
rect 17219 13017 17247 13129
rect 16307 12989 16711 13017
rect 16219 12877 16247 12989
rect 16683 12877 16711 12989
rect 16843 12989 17247 13017
rect 17291 13017 17319 13129
rect 17483 13017 17511 13129
rect 17291 12989 17335 13017
rect 16843 12877 16871 12989
rect 17307 12877 17335 12989
rect 17467 12989 17511 13017
rect 17555 13017 17583 13129
rect 18467 13017 18495 13129
rect 17555 12989 17959 13017
rect 17467 12877 17495 12989
rect 17931 12877 17959 12989
rect 18091 12989 18495 13017
rect 18539 13017 18567 13129
rect 18731 13017 18759 13129
rect 18539 12989 18583 13017
rect 18091 12877 18119 12989
rect 18555 12877 18583 12989
rect 18715 12989 18759 13017
rect 18803 13017 18831 13129
rect 19715 13017 19743 13129
rect 18803 12989 19207 13017
rect 18715 12877 18743 12989
rect 19179 12877 19207 12989
rect 19339 12989 19743 13017
rect 19787 13017 19815 13129
rect 19979 13017 20007 13129
rect 19787 12989 19831 13017
rect 19339 12877 19367 12989
rect 19803 12877 19831 12989
rect 19963 12989 20007 13017
rect 20051 13017 20079 13129
rect 20963 13017 20991 13129
rect 20051 12989 20455 13017
rect 19963 12877 19991 12989
rect 20427 12877 20455 12989
rect 20587 12989 20991 13017
rect 21035 13017 21063 13129
rect 21227 13017 21255 13129
rect 21035 12989 21079 13017
rect 20587 12877 20615 12989
rect 21051 12877 21079 12989
rect 21211 12989 21255 13017
rect 21299 13017 21327 13129
rect 22211 13017 22239 13129
rect 21299 12989 21703 13017
rect 21211 12877 21239 12989
rect 21675 12877 21703 12989
rect 21835 12989 22239 13017
rect 22283 13017 22311 13129
rect 22475 13017 22503 13129
rect 22283 12989 22327 13017
rect 21835 12877 21863 12989
rect 22299 12877 22327 12989
rect 22459 12989 22503 13017
rect 22547 13017 22575 13129
rect 23459 13017 23487 13129
rect 22547 12989 22951 13017
rect 22459 12877 22487 12989
rect 22923 12877 22951 12989
rect 23083 12989 23487 13017
rect 23531 13017 23559 13129
rect 23723 13017 23751 13129
rect 23531 12989 23575 13017
rect 23083 12877 23111 12989
rect 23547 12877 23575 12989
rect 23707 12989 23751 13017
rect 23795 13017 23823 13129
rect 24707 13017 24735 13129
rect 23795 12989 24199 13017
rect 23707 12877 23735 12989
rect 24171 12877 24199 12989
rect 24331 12989 24735 13017
rect 24779 13017 24807 13129
rect 24971 13017 24999 13129
rect 24779 12989 24823 13017
rect 24331 12877 24359 12989
rect 24795 12877 24823 12989
rect 24955 12989 24999 13017
rect 25043 13017 25071 13129
rect 25955 13017 25983 13129
rect 25043 12989 25447 13017
rect 24955 12877 24983 12989
rect 25419 12877 25447 12989
rect 25579 12989 25983 13017
rect 26027 13017 26055 13129
rect 26219 13017 26247 13129
rect 26027 12989 26071 13017
rect 25579 12877 25607 12989
rect 26043 12877 26071 12989
rect 26203 12989 26247 13017
rect 26291 13017 26319 13129
rect 27203 13017 27231 13129
rect 26291 12989 26695 13017
rect 26203 12877 26231 12989
rect 26667 12877 26695 12989
rect 26827 12989 27231 13017
rect 27275 13017 27303 13129
rect 27467 13017 27495 13129
rect 27275 12989 27319 13017
rect 26827 12877 26855 12989
rect 27291 12877 27319 12989
rect 27451 12989 27495 13017
rect 27539 13017 27567 13129
rect 28451 13017 28479 13129
rect 27539 12989 27943 13017
rect 27451 12877 27479 12989
rect 27915 12877 27943 12989
rect 28075 12989 28479 13017
rect 28523 13017 28551 13129
rect 28715 13017 28743 13129
rect 28523 12989 28567 13017
rect 28075 12877 28103 12989
rect 28539 12877 28567 12989
rect 28699 12989 28743 13017
rect 28787 13017 28815 13129
rect 29699 13017 29727 13129
rect 28787 12989 29191 13017
rect 28699 12877 28727 12989
rect 29163 12877 29191 12989
rect 29323 12989 29727 13017
rect 29771 13017 29799 13129
rect 29963 13017 29991 13129
rect 29771 12989 29815 13017
rect 29323 12877 29351 12989
rect 29787 12877 29815 12989
rect 29947 12989 29991 13017
rect 30035 13017 30063 13129
rect 30947 13017 30975 13129
rect 30035 12989 30439 13017
rect 29947 12877 29975 12989
rect 30411 12877 30439 12989
rect 30571 12989 30975 13017
rect 31019 13017 31047 13129
rect 31211 13017 31239 13129
rect 31019 12989 31063 13017
rect 30571 12877 30599 12989
rect 31035 12877 31063 12989
rect 31195 12989 31239 13017
rect 31283 13017 31311 13129
rect 32195 13017 32223 13129
rect 31283 12989 31687 13017
rect 31195 12877 31223 12989
rect 31659 12877 31687 12989
rect 31819 12989 32223 13017
rect 32267 13017 32295 13129
rect 32459 13017 32487 13129
rect 32267 12989 32311 13017
rect 31819 12877 31847 12989
rect 32283 12877 32311 12989
rect 32443 12989 32487 13017
rect 32531 13017 32559 13129
rect 33443 13017 33471 13129
rect 32531 12989 32935 13017
rect 32443 12877 32471 12989
rect 32907 12877 32935 12989
rect 33067 12989 33471 13017
rect 33515 13017 33543 13129
rect 33707 13017 33735 13129
rect 33515 12989 33559 13017
rect 33067 12877 33095 12989
rect 33531 12877 33559 12989
rect 33691 12989 33735 13017
rect 33779 13017 33807 13129
rect 34691 13017 34719 13129
rect 33779 12989 34183 13017
rect 33691 12877 33719 12989
rect 34155 12877 34183 12989
rect 34315 12989 34719 13017
rect 34763 13017 34791 13129
rect 34955 13017 34983 13129
rect 34763 12989 34807 13017
rect 34315 12877 34343 12989
rect 34779 12877 34807 12989
rect 34939 12989 34983 13017
rect 35027 13017 35055 13129
rect 35939 13017 35967 13129
rect 35027 12989 35431 13017
rect 34939 12877 34967 12989
rect 35403 12877 35431 12989
rect 35563 12989 35967 13017
rect 36011 13017 36039 13129
rect 36203 13017 36231 13129
rect 36011 12989 36055 13017
rect 35563 12877 35591 12989
rect 36027 12877 36055 12989
rect 36187 12989 36231 13017
rect 36275 13017 36303 13129
rect 37187 13017 37215 13129
rect 36275 12989 36679 13017
rect 36187 12877 36215 12989
rect 36651 12877 36679 12989
rect 36811 12989 37215 13017
rect 37259 13017 37287 13129
rect 37451 13017 37479 13129
rect 37259 12989 37303 13017
rect 36811 12877 36839 12989
rect 37275 12877 37303 12989
rect 37435 12989 37479 13017
rect 37523 13017 37551 13129
rect 38435 13017 38463 13129
rect 37523 12989 37927 13017
rect 37435 12877 37463 12989
rect 37899 12877 37927 12989
rect 38059 12989 38463 13017
rect 38507 13017 38535 13129
rect 38699 13017 38727 13129
rect 38507 12989 38551 13017
rect 38059 12877 38087 12989
rect 38523 12877 38551 12989
rect 38683 12989 38727 13017
rect 38771 13017 38799 13129
rect 39683 13017 39711 13129
rect 38771 12989 39175 13017
rect 38683 12877 38711 12989
rect 39147 12877 39175 12989
rect 39307 12989 39711 13017
rect 39755 13017 39783 13129
rect 39947 13017 39975 13129
rect 39755 12989 39799 13017
rect 39307 12877 39335 12989
rect 39771 12877 39799 12989
rect 39931 12989 39975 13017
rect 40019 13017 40047 13129
rect 40931 13017 40959 13129
rect 40019 12989 40423 13017
rect 39931 12877 39959 12989
rect 40395 12877 40423 12989
rect 40555 12989 40959 13017
rect 41003 13017 41031 13129
rect 41195 13017 41223 13129
rect 41003 12989 41047 13017
rect 40555 12877 40583 12989
rect 41019 12877 41047 12989
rect 41179 12989 41223 13017
rect 41267 13017 41295 13129
rect 42179 13017 42207 13129
rect 41267 12989 41671 13017
rect 41179 12877 41207 12989
rect 41643 12877 41671 12989
rect 41803 12989 42207 13017
rect 42251 13017 42279 13129
rect 42443 13017 42471 13129
rect 42251 12989 42295 13017
rect 41803 12877 41831 12989
rect 42267 12877 42295 12989
rect 42427 12989 42471 13017
rect 42515 13017 42543 13129
rect 43427 13017 43455 13129
rect 42515 12989 42919 13017
rect 42427 12877 42455 12989
rect 42891 12877 42919 12989
rect 43051 12989 43455 13017
rect 43499 13017 43527 13129
rect 43691 13017 43719 13129
rect 43499 12989 43543 13017
rect 43051 12877 43079 12989
rect 43515 12877 43543 12989
rect 43675 12989 43719 13017
rect 43763 13017 43791 13129
rect 44675 13017 44703 13129
rect 43763 12989 44167 13017
rect 43675 12877 43703 12989
rect 44139 12877 44167 12989
rect 44299 12989 44703 13017
rect 44747 13017 44775 13129
rect 44939 13017 44967 13129
rect 44747 12989 44791 13017
rect 44299 12877 44327 12989
rect 44763 12877 44791 12989
rect 44923 12989 44967 13017
rect 45011 13017 45039 13129
rect 45923 13017 45951 13129
rect 45011 12989 45415 13017
rect 44923 12877 44951 12989
rect 45387 12877 45415 12989
rect 45547 12989 45951 13017
rect 45995 13017 46023 13129
rect 46187 13017 46215 13129
rect 45995 12989 46039 13017
rect 45547 12877 45575 12989
rect 46011 12877 46039 12989
rect 46171 12989 46215 13017
rect 46259 13017 46287 13129
rect 47171 13017 47199 13129
rect 46259 12989 46663 13017
rect 46171 12877 46199 12989
rect 46635 12877 46663 12989
rect 46795 12989 47199 13017
rect 47243 13017 47271 13129
rect 47435 13017 47463 13129
rect 47243 12989 47287 13017
rect 46795 12877 46823 12989
rect 47259 12877 47287 12989
rect 47419 12989 47463 13017
rect 47507 13017 47535 13129
rect 48419 13017 48447 13129
rect 47507 12989 47911 13017
rect 47419 12877 47447 12989
rect 47883 12877 47911 12989
rect 48043 12989 48447 13017
rect 48491 13017 48519 13129
rect 48683 13017 48711 13129
rect 48491 12989 48535 13017
rect 48043 12877 48071 12989
rect 48507 12877 48535 12989
rect 48667 12989 48711 13017
rect 48755 13017 48783 13129
rect 49667 13017 49695 13129
rect 48755 12989 49159 13017
rect 48667 12877 48695 12989
rect 49131 12877 49159 12989
rect 49291 12989 49695 13017
rect 49739 13017 49767 13129
rect 49931 13017 49959 13129
rect 49739 12989 49783 13017
rect 49291 12877 49319 12989
rect 49755 12877 49783 12989
rect 49915 12989 49959 13017
rect 50003 13017 50031 13129
rect 50915 13017 50943 13129
rect 50003 12989 50407 13017
rect 49915 12877 49943 12989
rect 50379 12877 50407 12989
rect 50539 12989 50943 13017
rect 50987 13017 51015 13129
rect 51179 13017 51207 13129
rect 50987 12989 51031 13017
rect 50539 12877 50567 12989
rect 51003 12877 51031 12989
rect 51163 12989 51207 13017
rect 51251 13017 51279 13129
rect 52163 13017 52191 13129
rect 51251 12989 51655 13017
rect 51163 12877 51191 12989
rect 51627 12877 51655 12989
rect 51787 12989 52191 13017
rect 52235 13017 52263 13129
rect 52427 13017 52455 13129
rect 52235 12989 52279 13017
rect 51787 12877 51815 12989
rect 52251 12877 52279 12989
rect 52411 12989 52455 13017
rect 52499 13017 52527 13129
rect 53411 13017 53439 13129
rect 52499 12989 52903 13017
rect 52411 12877 52439 12989
rect 52875 12877 52903 12989
rect 53035 12989 53439 13017
rect 53483 13017 53511 13129
rect 53483 12989 53527 13017
rect 53035 12877 53063 12989
rect 53499 12877 53527 12989
rect 13563 12025 13591 12123
rect 13545 11973 13551 12025
rect 13603 11973 13609 12025
rect 6834 10666 6840 10718
rect 6892 10666 6898 10718
rect 6834 9176 6840 9228
rect 6892 9176 6898 9228
rect 6834 7838 6840 7890
rect 6892 7838 6898 7890
rect 13761 6683 13807 6937
rect 18753 6683 18799 6937
rect 23745 6683 23791 6937
rect 28737 6683 28783 6937
rect 33729 6683 33775 6937
rect 38721 6683 38767 6937
rect 43713 6683 43759 6937
rect 48705 6683 48751 6937
rect 6834 6348 6840 6400
rect 6892 6348 6898 6400
rect 6834 5010 6840 5062
rect 6892 5010 6898 5062
rect 13912 4424 13972 4480
rect 18904 4424 18964 4480
rect 23896 4424 23956 4480
rect 28888 4424 28948 4480
rect 33880 4424 33940 4480
rect 38872 4424 38932 4480
rect 43864 4424 43924 4480
rect 48856 4424 48916 4480
rect 4558 3517 4604 3575
rect 6834 3520 6840 3572
rect 6892 3520 6898 3572
rect 4434 2179 4480 2237
rect 6834 2182 6840 2234
rect 6892 2182 6898 2234
rect 4310 689 4356 747
rect 6834 692 6840 744
rect 6892 692 6898 744
<< via1 >>
rect 60234 77697 60286 77706
rect 60234 77663 60243 77697
rect 60243 77663 60277 77697
rect 60277 77663 60286 77697
rect 60234 77654 60286 77663
rect 60234 76207 60286 76216
rect 60234 76173 60243 76207
rect 60243 76173 60277 76207
rect 60277 76173 60286 76207
rect 60234 76164 60286 76173
rect 60234 74869 60286 74878
rect 60234 74835 60243 74869
rect 60243 74835 60277 74869
rect 60277 74835 60286 74869
rect 60234 74826 60286 74835
rect 60234 73379 60286 73388
rect 60234 73345 60243 73379
rect 60243 73345 60277 73379
rect 60277 73345 60286 73379
rect 60234 73336 60286 73345
rect 60234 72041 60286 72050
rect 60234 72007 60243 72041
rect 60243 72007 60277 72041
rect 60277 72007 60286 72041
rect 60234 71998 60286 72007
rect 60234 70551 60286 70560
rect 60234 70517 60243 70551
rect 60243 70517 60277 70551
rect 60277 70517 60286 70551
rect 60234 70508 60286 70517
rect 60234 69213 60286 69222
rect 60234 69179 60243 69213
rect 60243 69179 60277 69213
rect 60277 69179 60286 69213
rect 60234 69170 60286 69179
rect 60234 67723 60286 67732
rect 60234 67689 60243 67723
rect 60243 67689 60277 67723
rect 60277 67689 60286 67723
rect 60234 67680 60286 67689
rect 53647 66373 53699 66425
rect 55068 64616 55120 64625
rect 55068 64582 55077 64616
rect 55077 64582 55111 64616
rect 55111 64582 55120 64616
rect 55068 64573 55120 64582
rect 12130 64376 12182 64385
rect 12130 64342 12139 64376
rect 12139 64342 12173 64376
rect 12173 64342 12182 64376
rect 12130 64333 12182 64342
rect 55068 64376 55120 64385
rect 55068 64342 55077 64376
rect 55077 64342 55111 64376
rect 55111 64342 55120 64376
rect 55068 64333 55120 64342
rect 12130 63826 12182 63835
rect 12130 63792 12139 63826
rect 12139 63792 12173 63826
rect 12173 63792 12182 63826
rect 12130 63783 12182 63792
rect 55068 63826 55120 63835
rect 55068 63792 55077 63826
rect 55077 63792 55111 63826
rect 55111 63792 55120 63826
rect 55068 63783 55120 63792
rect 12130 63586 12182 63595
rect 12130 63552 12139 63586
rect 12139 63552 12173 63586
rect 12173 63552 12182 63586
rect 12130 63543 12182 63552
rect 55068 63586 55120 63595
rect 55068 63552 55077 63586
rect 55077 63552 55111 63586
rect 55111 63552 55120 63586
rect 55068 63543 55120 63552
rect 12130 63036 12182 63045
rect 12130 63002 12139 63036
rect 12139 63002 12173 63036
rect 12173 63002 12182 63036
rect 12130 62993 12182 63002
rect 55068 63036 55120 63045
rect 55068 63002 55077 63036
rect 55077 63002 55111 63036
rect 55111 63002 55120 63036
rect 55068 62993 55120 63002
rect 12130 62796 12182 62805
rect 12130 62762 12139 62796
rect 12139 62762 12173 62796
rect 12173 62762 12182 62796
rect 12130 62753 12182 62762
rect 55068 62796 55120 62805
rect 55068 62762 55077 62796
rect 55077 62762 55111 62796
rect 55111 62762 55120 62796
rect 55068 62753 55120 62762
rect 12130 62246 12182 62255
rect 12130 62212 12139 62246
rect 12139 62212 12173 62246
rect 12173 62212 12182 62246
rect 12130 62203 12182 62212
rect 55068 62246 55120 62255
rect 55068 62212 55077 62246
rect 55077 62212 55111 62246
rect 55111 62212 55120 62246
rect 55068 62203 55120 62212
rect 12130 62006 12182 62015
rect 12130 61972 12139 62006
rect 12139 61972 12173 62006
rect 12173 61972 12182 62006
rect 12130 61963 12182 61972
rect 55068 62006 55120 62015
rect 55068 61972 55077 62006
rect 55077 61972 55111 62006
rect 55111 61972 55120 62006
rect 55068 61963 55120 61972
rect 12130 61456 12182 61465
rect 12130 61422 12139 61456
rect 12139 61422 12173 61456
rect 12173 61422 12182 61456
rect 12130 61413 12182 61422
rect 55068 61456 55120 61465
rect 55068 61422 55077 61456
rect 55077 61422 55111 61456
rect 55111 61422 55120 61456
rect 55068 61413 55120 61422
rect 12130 61216 12182 61225
rect 12130 61182 12139 61216
rect 12139 61182 12173 61216
rect 12173 61182 12182 61216
rect 12130 61173 12182 61182
rect 55068 61216 55120 61225
rect 55068 61182 55077 61216
rect 55077 61182 55111 61216
rect 55111 61182 55120 61216
rect 55068 61173 55120 61182
rect 12130 60666 12182 60675
rect 12130 60632 12139 60666
rect 12139 60632 12173 60666
rect 12173 60632 12182 60666
rect 12130 60623 12182 60632
rect 55068 60666 55120 60675
rect 55068 60632 55077 60666
rect 55077 60632 55111 60666
rect 55111 60632 55120 60666
rect 55068 60623 55120 60632
rect 12130 60426 12182 60435
rect 12130 60392 12139 60426
rect 12139 60392 12173 60426
rect 12173 60392 12182 60426
rect 12130 60383 12182 60392
rect 55068 60426 55120 60435
rect 55068 60392 55077 60426
rect 55077 60392 55111 60426
rect 55111 60392 55120 60426
rect 55068 60383 55120 60392
rect 12130 59876 12182 59885
rect 12130 59842 12139 59876
rect 12139 59842 12173 59876
rect 12173 59842 12182 59876
rect 12130 59833 12182 59842
rect 55068 59876 55120 59885
rect 55068 59842 55077 59876
rect 55077 59842 55111 59876
rect 55111 59842 55120 59876
rect 55068 59833 55120 59842
rect 12130 59636 12182 59645
rect 12130 59602 12139 59636
rect 12139 59602 12173 59636
rect 12173 59602 12182 59636
rect 12130 59593 12182 59602
rect 55068 59636 55120 59645
rect 55068 59602 55077 59636
rect 55077 59602 55111 59636
rect 55111 59602 55120 59636
rect 55068 59593 55120 59602
rect 12130 59086 12182 59095
rect 12130 59052 12139 59086
rect 12139 59052 12173 59086
rect 12173 59052 12182 59086
rect 12130 59043 12182 59052
rect 55068 59086 55120 59095
rect 55068 59052 55077 59086
rect 55077 59052 55111 59086
rect 55111 59052 55120 59086
rect 55068 59043 55120 59052
rect 12130 58846 12182 58855
rect 12130 58812 12139 58846
rect 12139 58812 12173 58846
rect 12173 58812 12182 58846
rect 12130 58803 12182 58812
rect 55068 58846 55120 58855
rect 55068 58812 55077 58846
rect 55077 58812 55111 58846
rect 55111 58812 55120 58846
rect 55068 58803 55120 58812
rect 12130 58296 12182 58305
rect 12130 58262 12139 58296
rect 12139 58262 12173 58296
rect 12173 58262 12182 58296
rect 12130 58253 12182 58262
rect 55068 58296 55120 58305
rect 55068 58262 55077 58296
rect 55077 58262 55111 58296
rect 55111 58262 55120 58296
rect 55068 58253 55120 58262
rect 12130 58056 12182 58065
rect 12130 58022 12139 58056
rect 12139 58022 12173 58056
rect 12173 58022 12182 58056
rect 12130 58013 12182 58022
rect 55068 58056 55120 58065
rect 55068 58022 55077 58056
rect 55077 58022 55111 58056
rect 55111 58022 55120 58056
rect 55068 58013 55120 58022
rect 12130 57506 12182 57515
rect 12130 57472 12139 57506
rect 12139 57472 12173 57506
rect 12173 57472 12182 57506
rect 12130 57463 12182 57472
rect 55068 57506 55120 57515
rect 55068 57472 55077 57506
rect 55077 57472 55111 57506
rect 55111 57472 55120 57506
rect 55068 57463 55120 57472
rect 12130 57266 12182 57275
rect 12130 57232 12139 57266
rect 12139 57232 12173 57266
rect 12173 57232 12182 57266
rect 12130 57223 12182 57232
rect 55068 57266 55120 57275
rect 55068 57232 55077 57266
rect 55077 57232 55111 57266
rect 55111 57232 55120 57266
rect 55068 57223 55120 57232
rect 12130 56716 12182 56725
rect 12130 56682 12139 56716
rect 12139 56682 12173 56716
rect 12173 56682 12182 56716
rect 12130 56673 12182 56682
rect 55068 56716 55120 56725
rect 55068 56682 55077 56716
rect 55077 56682 55111 56716
rect 55111 56682 55120 56716
rect 55068 56673 55120 56682
rect 12130 56476 12182 56485
rect 12130 56442 12139 56476
rect 12139 56442 12173 56476
rect 12173 56442 12182 56476
rect 12130 56433 12182 56442
rect 55068 56476 55120 56485
rect 55068 56442 55077 56476
rect 55077 56442 55111 56476
rect 55111 56442 55120 56476
rect 55068 56433 55120 56442
rect 12130 55926 12182 55935
rect 12130 55892 12139 55926
rect 12139 55892 12173 55926
rect 12173 55892 12182 55926
rect 12130 55883 12182 55892
rect 55068 55926 55120 55935
rect 55068 55892 55077 55926
rect 55077 55892 55111 55926
rect 55111 55892 55120 55926
rect 55068 55883 55120 55892
rect 12130 55686 12182 55695
rect 12130 55652 12139 55686
rect 12139 55652 12173 55686
rect 12173 55652 12182 55686
rect 12130 55643 12182 55652
rect 55068 55686 55120 55695
rect 55068 55652 55077 55686
rect 55077 55652 55111 55686
rect 55111 55652 55120 55686
rect 55068 55643 55120 55652
rect 12130 55136 12182 55145
rect 12130 55102 12139 55136
rect 12139 55102 12173 55136
rect 12173 55102 12182 55136
rect 12130 55093 12182 55102
rect 55068 55136 55120 55145
rect 55068 55102 55077 55136
rect 55077 55102 55111 55136
rect 55111 55102 55120 55136
rect 55068 55093 55120 55102
rect 12130 54896 12182 54905
rect 12130 54862 12139 54896
rect 12139 54862 12173 54896
rect 12173 54862 12182 54896
rect 12130 54853 12182 54862
rect 55068 54896 55120 54905
rect 55068 54862 55077 54896
rect 55077 54862 55111 54896
rect 55111 54862 55120 54896
rect 55068 54853 55120 54862
rect 12130 54346 12182 54355
rect 12130 54312 12139 54346
rect 12139 54312 12173 54346
rect 12173 54312 12182 54346
rect 12130 54303 12182 54312
rect 55068 54346 55120 54355
rect 55068 54312 55077 54346
rect 55077 54312 55111 54346
rect 55111 54312 55120 54346
rect 55068 54303 55120 54312
rect 12130 54106 12182 54115
rect 12130 54072 12139 54106
rect 12139 54072 12173 54106
rect 12173 54072 12182 54106
rect 12130 54063 12182 54072
rect 55068 54106 55120 54115
rect 55068 54072 55077 54106
rect 55077 54072 55111 54106
rect 55111 54072 55120 54106
rect 55068 54063 55120 54072
rect 12130 53556 12182 53565
rect 12130 53522 12139 53556
rect 12139 53522 12173 53556
rect 12173 53522 12182 53556
rect 12130 53513 12182 53522
rect 55068 53556 55120 53565
rect 55068 53522 55077 53556
rect 55077 53522 55111 53556
rect 55111 53522 55120 53556
rect 55068 53513 55120 53522
rect 12130 53316 12182 53325
rect 12130 53282 12139 53316
rect 12139 53282 12173 53316
rect 12173 53282 12182 53316
rect 12130 53273 12182 53282
rect 55068 53316 55120 53325
rect 55068 53282 55077 53316
rect 55077 53282 55111 53316
rect 55111 53282 55120 53316
rect 55068 53273 55120 53282
rect 12130 52766 12182 52775
rect 12130 52732 12139 52766
rect 12139 52732 12173 52766
rect 12173 52732 12182 52766
rect 12130 52723 12182 52732
rect 55068 52766 55120 52775
rect 55068 52732 55077 52766
rect 55077 52732 55111 52766
rect 55111 52732 55120 52766
rect 55068 52723 55120 52732
rect 12130 52526 12182 52535
rect 12130 52492 12139 52526
rect 12139 52492 12173 52526
rect 12173 52492 12182 52526
rect 12130 52483 12182 52492
rect 55068 52526 55120 52535
rect 55068 52492 55077 52526
rect 55077 52492 55111 52526
rect 55111 52492 55120 52526
rect 55068 52483 55120 52492
rect 12130 51976 12182 51985
rect 12130 51942 12139 51976
rect 12139 51942 12173 51976
rect 12173 51942 12182 51976
rect 12130 51933 12182 51942
rect 55068 51976 55120 51985
rect 55068 51942 55077 51976
rect 55077 51942 55111 51976
rect 55111 51942 55120 51976
rect 55068 51933 55120 51942
rect 12130 51736 12182 51745
rect 12130 51702 12139 51736
rect 12139 51702 12173 51736
rect 12173 51702 12182 51736
rect 12130 51693 12182 51702
rect 55068 51736 55120 51745
rect 55068 51702 55077 51736
rect 55077 51702 55111 51736
rect 55111 51702 55120 51736
rect 55068 51693 55120 51702
rect 12130 51186 12182 51195
rect 12130 51152 12139 51186
rect 12139 51152 12173 51186
rect 12173 51152 12182 51186
rect 12130 51143 12182 51152
rect 55068 51186 55120 51195
rect 55068 51152 55077 51186
rect 55077 51152 55111 51186
rect 55111 51152 55120 51186
rect 55068 51143 55120 51152
rect 12130 50946 12182 50955
rect 12130 50912 12139 50946
rect 12139 50912 12173 50946
rect 12173 50912 12182 50946
rect 12130 50903 12182 50912
rect 55068 50946 55120 50955
rect 55068 50912 55077 50946
rect 55077 50912 55111 50946
rect 55111 50912 55120 50946
rect 55068 50903 55120 50912
rect 12130 50396 12182 50405
rect 12130 50362 12139 50396
rect 12139 50362 12173 50396
rect 12173 50362 12182 50396
rect 12130 50353 12182 50362
rect 55068 50396 55120 50405
rect 55068 50362 55077 50396
rect 55077 50362 55111 50396
rect 55111 50362 55120 50396
rect 55068 50353 55120 50362
rect 12130 50156 12182 50165
rect 12130 50122 12139 50156
rect 12139 50122 12173 50156
rect 12173 50122 12182 50156
rect 12130 50113 12182 50122
rect 55068 50156 55120 50165
rect 55068 50122 55077 50156
rect 55077 50122 55111 50156
rect 55111 50122 55120 50156
rect 55068 50113 55120 50122
rect 12130 49606 12182 49615
rect 12130 49572 12139 49606
rect 12139 49572 12173 49606
rect 12173 49572 12182 49606
rect 12130 49563 12182 49572
rect 55068 49606 55120 49615
rect 55068 49572 55077 49606
rect 55077 49572 55111 49606
rect 55111 49572 55120 49606
rect 55068 49563 55120 49572
rect 12130 49366 12182 49375
rect 12130 49332 12139 49366
rect 12139 49332 12173 49366
rect 12173 49332 12182 49366
rect 12130 49323 12182 49332
rect 55068 49366 55120 49375
rect 55068 49332 55077 49366
rect 55077 49332 55111 49366
rect 55111 49332 55120 49366
rect 55068 49323 55120 49332
rect 12130 48816 12182 48825
rect 12130 48782 12139 48816
rect 12139 48782 12173 48816
rect 12173 48782 12182 48816
rect 12130 48773 12182 48782
rect 55068 48816 55120 48825
rect 55068 48782 55077 48816
rect 55077 48782 55111 48816
rect 55111 48782 55120 48816
rect 55068 48773 55120 48782
rect 12130 48576 12182 48585
rect 12130 48542 12139 48576
rect 12139 48542 12173 48576
rect 12173 48542 12182 48576
rect 12130 48533 12182 48542
rect 55068 48576 55120 48585
rect 55068 48542 55077 48576
rect 55077 48542 55111 48576
rect 55111 48542 55120 48576
rect 55068 48533 55120 48542
rect 12130 48026 12182 48035
rect 12130 47992 12139 48026
rect 12139 47992 12173 48026
rect 12173 47992 12182 48026
rect 12130 47983 12182 47992
rect 55068 48026 55120 48035
rect 55068 47992 55077 48026
rect 55077 47992 55111 48026
rect 55111 47992 55120 48026
rect 55068 47983 55120 47992
rect 12130 47786 12182 47795
rect 12130 47752 12139 47786
rect 12139 47752 12173 47786
rect 12173 47752 12182 47786
rect 12130 47743 12182 47752
rect 55068 47786 55120 47795
rect 55068 47752 55077 47786
rect 55077 47752 55111 47786
rect 55111 47752 55120 47786
rect 55068 47743 55120 47752
rect 12130 47236 12182 47245
rect 12130 47202 12139 47236
rect 12139 47202 12173 47236
rect 12173 47202 12182 47236
rect 12130 47193 12182 47202
rect 55068 47236 55120 47245
rect 55068 47202 55077 47236
rect 55077 47202 55111 47236
rect 55111 47202 55120 47236
rect 55068 47193 55120 47202
rect 12130 46996 12182 47005
rect 12130 46962 12139 46996
rect 12139 46962 12173 46996
rect 12173 46962 12182 46996
rect 12130 46953 12182 46962
rect 55068 46996 55120 47005
rect 55068 46962 55077 46996
rect 55077 46962 55111 46996
rect 55111 46962 55120 46996
rect 55068 46953 55120 46962
rect 12130 46446 12182 46455
rect 12130 46412 12139 46446
rect 12139 46412 12173 46446
rect 12173 46412 12182 46446
rect 12130 46403 12182 46412
rect 55068 46446 55120 46455
rect 55068 46412 55077 46446
rect 55077 46412 55111 46446
rect 55111 46412 55120 46446
rect 55068 46403 55120 46412
rect 12130 46206 12182 46215
rect 12130 46172 12139 46206
rect 12139 46172 12173 46206
rect 12173 46172 12182 46206
rect 12130 46163 12182 46172
rect 55068 46206 55120 46215
rect 55068 46172 55077 46206
rect 55077 46172 55111 46206
rect 55111 46172 55120 46206
rect 55068 46163 55120 46172
rect 12130 45656 12182 45665
rect 12130 45622 12139 45656
rect 12139 45622 12173 45656
rect 12173 45622 12182 45656
rect 12130 45613 12182 45622
rect 55068 45656 55120 45665
rect 55068 45622 55077 45656
rect 55077 45622 55111 45656
rect 55111 45622 55120 45656
rect 55068 45613 55120 45622
rect 12130 45416 12182 45425
rect 12130 45382 12139 45416
rect 12139 45382 12173 45416
rect 12173 45382 12182 45416
rect 12130 45373 12182 45382
rect 55068 45416 55120 45425
rect 55068 45382 55077 45416
rect 55077 45382 55111 45416
rect 55111 45382 55120 45416
rect 55068 45373 55120 45382
rect 12130 44866 12182 44875
rect 12130 44832 12139 44866
rect 12139 44832 12173 44866
rect 12173 44832 12182 44866
rect 12130 44823 12182 44832
rect 55068 44866 55120 44875
rect 55068 44832 55077 44866
rect 55077 44832 55111 44866
rect 55111 44832 55120 44866
rect 55068 44823 55120 44832
rect 12130 44626 12182 44635
rect 12130 44592 12139 44626
rect 12139 44592 12173 44626
rect 12173 44592 12182 44626
rect 12130 44583 12182 44592
rect 55068 44626 55120 44635
rect 55068 44592 55077 44626
rect 55077 44592 55111 44626
rect 55111 44592 55120 44626
rect 55068 44583 55120 44592
rect 12130 44076 12182 44085
rect 12130 44042 12139 44076
rect 12139 44042 12173 44076
rect 12173 44042 12182 44076
rect 12130 44033 12182 44042
rect 55068 44076 55120 44085
rect 55068 44042 55077 44076
rect 55077 44042 55111 44076
rect 55111 44042 55120 44076
rect 55068 44033 55120 44042
rect 12130 43836 12182 43845
rect 12130 43802 12139 43836
rect 12139 43802 12173 43836
rect 12173 43802 12182 43836
rect 12130 43793 12182 43802
rect 55068 43836 55120 43845
rect 55068 43802 55077 43836
rect 55077 43802 55111 43836
rect 55111 43802 55120 43836
rect 55068 43793 55120 43802
rect 12130 43286 12182 43295
rect 12130 43252 12139 43286
rect 12139 43252 12173 43286
rect 12173 43252 12182 43286
rect 12130 43243 12182 43252
rect 55068 43286 55120 43295
rect 55068 43252 55077 43286
rect 55077 43252 55111 43286
rect 55111 43252 55120 43286
rect 55068 43243 55120 43252
rect 12130 43046 12182 43055
rect 12130 43012 12139 43046
rect 12139 43012 12173 43046
rect 12173 43012 12182 43046
rect 12130 43003 12182 43012
rect 55068 43046 55120 43055
rect 55068 43012 55077 43046
rect 55077 43012 55111 43046
rect 55111 43012 55120 43046
rect 55068 43003 55120 43012
rect 12130 42496 12182 42505
rect 12130 42462 12139 42496
rect 12139 42462 12173 42496
rect 12173 42462 12182 42496
rect 12130 42453 12182 42462
rect 55068 42496 55120 42505
rect 55068 42462 55077 42496
rect 55077 42462 55111 42496
rect 55111 42462 55120 42496
rect 55068 42453 55120 42462
rect 12130 42256 12182 42265
rect 12130 42222 12139 42256
rect 12139 42222 12173 42256
rect 12173 42222 12182 42256
rect 12130 42213 12182 42222
rect 55068 42256 55120 42265
rect 55068 42222 55077 42256
rect 55077 42222 55111 42256
rect 55111 42222 55120 42256
rect 55068 42213 55120 42222
rect 12130 41706 12182 41715
rect 12130 41672 12139 41706
rect 12139 41672 12173 41706
rect 12173 41672 12182 41706
rect 12130 41663 12182 41672
rect 55068 41706 55120 41715
rect 55068 41672 55077 41706
rect 55077 41672 55111 41706
rect 55111 41672 55120 41706
rect 55068 41663 55120 41672
rect 12130 41466 12182 41475
rect 12130 41432 12139 41466
rect 12139 41432 12173 41466
rect 12173 41432 12182 41466
rect 12130 41423 12182 41432
rect 55068 41466 55120 41475
rect 55068 41432 55077 41466
rect 55077 41432 55111 41466
rect 55111 41432 55120 41466
rect 55068 41423 55120 41432
rect 12130 40916 12182 40925
rect 12130 40882 12139 40916
rect 12139 40882 12173 40916
rect 12173 40882 12182 40916
rect 12130 40873 12182 40882
rect 55068 40916 55120 40925
rect 55068 40882 55077 40916
rect 55077 40882 55111 40916
rect 55111 40882 55120 40916
rect 55068 40873 55120 40882
rect 12130 40676 12182 40685
rect 12130 40642 12139 40676
rect 12139 40642 12173 40676
rect 12173 40642 12182 40676
rect 12130 40633 12182 40642
rect 55068 40676 55120 40685
rect 55068 40642 55077 40676
rect 55077 40642 55111 40676
rect 55111 40642 55120 40676
rect 55068 40633 55120 40642
rect 12130 40126 12182 40135
rect 12130 40092 12139 40126
rect 12139 40092 12173 40126
rect 12173 40092 12182 40126
rect 12130 40083 12182 40092
rect 55068 40126 55120 40135
rect 55068 40092 55077 40126
rect 55077 40092 55111 40126
rect 55111 40092 55120 40126
rect 55068 40083 55120 40092
rect 12130 39886 12182 39895
rect 12130 39852 12139 39886
rect 12139 39852 12173 39886
rect 12173 39852 12182 39886
rect 12130 39843 12182 39852
rect 55068 39886 55120 39895
rect 55068 39852 55077 39886
rect 55077 39852 55111 39886
rect 55111 39852 55120 39886
rect 55068 39843 55120 39852
rect 12130 39336 12182 39345
rect 12130 39302 12139 39336
rect 12139 39302 12173 39336
rect 12173 39302 12182 39336
rect 12130 39293 12182 39302
rect 55068 39336 55120 39345
rect 55068 39302 55077 39336
rect 55077 39302 55111 39336
rect 55111 39302 55120 39336
rect 55068 39293 55120 39302
rect 12130 39096 12182 39105
rect 12130 39062 12139 39096
rect 12139 39062 12173 39096
rect 12173 39062 12182 39096
rect 12130 39053 12182 39062
rect 55068 39096 55120 39105
rect 55068 39062 55077 39096
rect 55077 39062 55111 39096
rect 55111 39062 55120 39096
rect 55068 39053 55120 39062
rect 12130 38546 12182 38555
rect 12130 38512 12139 38546
rect 12139 38512 12173 38546
rect 12173 38512 12182 38546
rect 12130 38503 12182 38512
rect 55068 38546 55120 38555
rect 55068 38512 55077 38546
rect 55077 38512 55111 38546
rect 55111 38512 55120 38546
rect 55068 38503 55120 38512
rect 12130 38306 12182 38315
rect 12130 38272 12139 38306
rect 12139 38272 12173 38306
rect 12173 38272 12182 38306
rect 12130 38263 12182 38272
rect 55068 38306 55120 38315
rect 55068 38272 55077 38306
rect 55077 38272 55111 38306
rect 55111 38272 55120 38306
rect 55068 38263 55120 38272
rect 12130 37756 12182 37765
rect 12130 37722 12139 37756
rect 12139 37722 12173 37756
rect 12173 37722 12182 37756
rect 12130 37713 12182 37722
rect 55068 37756 55120 37765
rect 55068 37722 55077 37756
rect 55077 37722 55111 37756
rect 55111 37722 55120 37756
rect 55068 37713 55120 37722
rect 12130 37516 12182 37525
rect 12130 37482 12139 37516
rect 12139 37482 12173 37516
rect 12173 37482 12182 37516
rect 12130 37473 12182 37482
rect 55068 37516 55120 37525
rect 55068 37482 55077 37516
rect 55077 37482 55111 37516
rect 55111 37482 55120 37516
rect 55068 37473 55120 37482
rect 12130 36966 12182 36975
rect 12130 36932 12139 36966
rect 12139 36932 12173 36966
rect 12173 36932 12182 36966
rect 12130 36923 12182 36932
rect 55068 36966 55120 36975
rect 55068 36932 55077 36966
rect 55077 36932 55111 36966
rect 55111 36932 55120 36966
rect 55068 36923 55120 36932
rect 12130 36726 12182 36735
rect 12130 36692 12139 36726
rect 12139 36692 12173 36726
rect 12173 36692 12182 36726
rect 12130 36683 12182 36692
rect 55068 36726 55120 36735
rect 55068 36692 55077 36726
rect 55077 36692 55111 36726
rect 55111 36692 55120 36726
rect 55068 36683 55120 36692
rect 12130 36176 12182 36185
rect 12130 36142 12139 36176
rect 12139 36142 12173 36176
rect 12173 36142 12182 36176
rect 12130 36133 12182 36142
rect 55068 36176 55120 36185
rect 55068 36142 55077 36176
rect 55077 36142 55111 36176
rect 55111 36142 55120 36176
rect 55068 36133 55120 36142
rect 12130 35936 12182 35945
rect 12130 35902 12139 35936
rect 12139 35902 12173 35936
rect 12173 35902 12182 35936
rect 12130 35893 12182 35902
rect 55068 35936 55120 35945
rect 55068 35902 55077 35936
rect 55077 35902 55111 35936
rect 55111 35902 55120 35936
rect 55068 35893 55120 35902
rect 12130 35386 12182 35395
rect 12130 35352 12139 35386
rect 12139 35352 12173 35386
rect 12173 35352 12182 35386
rect 12130 35343 12182 35352
rect 55068 35386 55120 35395
rect 55068 35352 55077 35386
rect 55077 35352 55111 35386
rect 55111 35352 55120 35386
rect 55068 35343 55120 35352
rect 12130 35146 12182 35155
rect 12130 35112 12139 35146
rect 12139 35112 12173 35146
rect 12173 35112 12182 35146
rect 12130 35103 12182 35112
rect 55068 35146 55120 35155
rect 55068 35112 55077 35146
rect 55077 35112 55111 35146
rect 55111 35112 55120 35146
rect 55068 35103 55120 35112
rect 12130 34596 12182 34605
rect 12130 34562 12139 34596
rect 12139 34562 12173 34596
rect 12173 34562 12182 34596
rect 12130 34553 12182 34562
rect 55068 34596 55120 34605
rect 55068 34562 55077 34596
rect 55077 34562 55111 34596
rect 55111 34562 55120 34596
rect 55068 34553 55120 34562
rect 12130 34356 12182 34365
rect 12130 34322 12139 34356
rect 12139 34322 12173 34356
rect 12173 34322 12182 34356
rect 12130 34313 12182 34322
rect 55068 34356 55120 34365
rect 55068 34322 55077 34356
rect 55077 34322 55111 34356
rect 55111 34322 55120 34356
rect 55068 34313 55120 34322
rect 12130 33806 12182 33815
rect 12130 33772 12139 33806
rect 12139 33772 12173 33806
rect 12173 33772 12182 33806
rect 12130 33763 12182 33772
rect 55068 33806 55120 33815
rect 55068 33772 55077 33806
rect 55077 33772 55111 33806
rect 55111 33772 55120 33806
rect 55068 33763 55120 33772
rect 12130 33566 12182 33575
rect 12130 33532 12139 33566
rect 12139 33532 12173 33566
rect 12173 33532 12182 33566
rect 12130 33523 12182 33532
rect 55068 33566 55120 33575
rect 55068 33532 55077 33566
rect 55077 33532 55111 33566
rect 55111 33532 55120 33566
rect 55068 33523 55120 33532
rect 12130 33016 12182 33025
rect 12130 32982 12139 33016
rect 12139 32982 12173 33016
rect 12173 32982 12182 33016
rect 12130 32973 12182 32982
rect 55068 33016 55120 33025
rect 55068 32982 55077 33016
rect 55077 32982 55111 33016
rect 55111 32982 55120 33016
rect 55068 32973 55120 32982
rect 12130 32776 12182 32785
rect 12130 32742 12139 32776
rect 12139 32742 12173 32776
rect 12173 32742 12182 32776
rect 12130 32733 12182 32742
rect 55068 32776 55120 32785
rect 55068 32742 55077 32776
rect 55077 32742 55111 32776
rect 55111 32742 55120 32776
rect 55068 32733 55120 32742
rect 12130 32226 12182 32235
rect 12130 32192 12139 32226
rect 12139 32192 12173 32226
rect 12173 32192 12182 32226
rect 12130 32183 12182 32192
rect 55068 32226 55120 32235
rect 55068 32192 55077 32226
rect 55077 32192 55111 32226
rect 55111 32192 55120 32226
rect 55068 32183 55120 32192
rect 12130 31986 12182 31995
rect 12130 31952 12139 31986
rect 12139 31952 12173 31986
rect 12173 31952 12182 31986
rect 12130 31943 12182 31952
rect 55068 31986 55120 31995
rect 55068 31952 55077 31986
rect 55077 31952 55111 31986
rect 55111 31952 55120 31986
rect 55068 31943 55120 31952
rect 12130 31436 12182 31445
rect 12130 31402 12139 31436
rect 12139 31402 12173 31436
rect 12173 31402 12182 31436
rect 12130 31393 12182 31402
rect 55068 31436 55120 31445
rect 55068 31402 55077 31436
rect 55077 31402 55111 31436
rect 55111 31402 55120 31436
rect 55068 31393 55120 31402
rect 12130 31196 12182 31205
rect 12130 31162 12139 31196
rect 12139 31162 12173 31196
rect 12173 31162 12182 31196
rect 12130 31153 12182 31162
rect 55068 31196 55120 31205
rect 55068 31162 55077 31196
rect 55077 31162 55111 31196
rect 55111 31162 55120 31196
rect 55068 31153 55120 31162
rect 12130 30646 12182 30655
rect 12130 30612 12139 30646
rect 12139 30612 12173 30646
rect 12173 30612 12182 30646
rect 12130 30603 12182 30612
rect 55068 30646 55120 30655
rect 55068 30612 55077 30646
rect 55077 30612 55111 30646
rect 55111 30612 55120 30646
rect 55068 30603 55120 30612
rect 12130 30406 12182 30415
rect 12130 30372 12139 30406
rect 12139 30372 12173 30406
rect 12173 30372 12182 30406
rect 12130 30363 12182 30372
rect 55068 30406 55120 30415
rect 55068 30372 55077 30406
rect 55077 30372 55111 30406
rect 55111 30372 55120 30406
rect 55068 30363 55120 30372
rect 12130 29856 12182 29865
rect 12130 29822 12139 29856
rect 12139 29822 12173 29856
rect 12173 29822 12182 29856
rect 12130 29813 12182 29822
rect 55068 29856 55120 29865
rect 55068 29822 55077 29856
rect 55077 29822 55111 29856
rect 55111 29822 55120 29856
rect 55068 29813 55120 29822
rect 12130 29616 12182 29625
rect 12130 29582 12139 29616
rect 12139 29582 12173 29616
rect 12173 29582 12182 29616
rect 12130 29573 12182 29582
rect 55068 29616 55120 29625
rect 55068 29582 55077 29616
rect 55077 29582 55111 29616
rect 55111 29582 55120 29616
rect 55068 29573 55120 29582
rect 12130 29066 12182 29075
rect 12130 29032 12139 29066
rect 12139 29032 12173 29066
rect 12173 29032 12182 29066
rect 12130 29023 12182 29032
rect 55068 29066 55120 29075
rect 55068 29032 55077 29066
rect 55077 29032 55111 29066
rect 55111 29032 55120 29066
rect 55068 29023 55120 29032
rect 12130 28826 12182 28835
rect 12130 28792 12139 28826
rect 12139 28792 12173 28826
rect 12173 28792 12182 28826
rect 12130 28783 12182 28792
rect 55068 28826 55120 28835
rect 55068 28792 55077 28826
rect 55077 28792 55111 28826
rect 55111 28792 55120 28826
rect 55068 28783 55120 28792
rect 12130 28276 12182 28285
rect 12130 28242 12139 28276
rect 12139 28242 12173 28276
rect 12173 28242 12182 28276
rect 12130 28233 12182 28242
rect 55068 28276 55120 28285
rect 55068 28242 55077 28276
rect 55077 28242 55111 28276
rect 55111 28242 55120 28276
rect 55068 28233 55120 28242
rect 12130 28036 12182 28045
rect 12130 28002 12139 28036
rect 12139 28002 12173 28036
rect 12173 28002 12182 28036
rect 12130 27993 12182 28002
rect 55068 28036 55120 28045
rect 55068 28002 55077 28036
rect 55077 28002 55111 28036
rect 55111 28002 55120 28036
rect 55068 27993 55120 28002
rect 12130 27486 12182 27495
rect 12130 27452 12139 27486
rect 12139 27452 12173 27486
rect 12173 27452 12182 27486
rect 12130 27443 12182 27452
rect 55068 27486 55120 27495
rect 55068 27452 55077 27486
rect 55077 27452 55111 27486
rect 55111 27452 55120 27486
rect 55068 27443 55120 27452
rect 12130 27246 12182 27255
rect 12130 27212 12139 27246
rect 12139 27212 12173 27246
rect 12173 27212 12182 27246
rect 12130 27203 12182 27212
rect 55068 27246 55120 27255
rect 55068 27212 55077 27246
rect 55077 27212 55111 27246
rect 55111 27212 55120 27246
rect 55068 27203 55120 27212
rect 12130 26696 12182 26705
rect 12130 26662 12139 26696
rect 12139 26662 12173 26696
rect 12173 26662 12182 26696
rect 12130 26653 12182 26662
rect 55068 26696 55120 26705
rect 55068 26662 55077 26696
rect 55077 26662 55111 26696
rect 55111 26662 55120 26696
rect 55068 26653 55120 26662
rect 12130 26456 12182 26465
rect 12130 26422 12139 26456
rect 12139 26422 12173 26456
rect 12173 26422 12182 26456
rect 12130 26413 12182 26422
rect 55068 26456 55120 26465
rect 55068 26422 55077 26456
rect 55077 26422 55111 26456
rect 55111 26422 55120 26456
rect 55068 26413 55120 26422
rect 12130 25906 12182 25915
rect 12130 25872 12139 25906
rect 12139 25872 12173 25906
rect 12173 25872 12182 25906
rect 12130 25863 12182 25872
rect 55068 25906 55120 25915
rect 55068 25872 55077 25906
rect 55077 25872 55111 25906
rect 55111 25872 55120 25906
rect 55068 25863 55120 25872
rect 12130 25666 12182 25675
rect 12130 25632 12139 25666
rect 12139 25632 12173 25666
rect 12173 25632 12182 25666
rect 12130 25623 12182 25632
rect 55068 25666 55120 25675
rect 55068 25632 55077 25666
rect 55077 25632 55111 25666
rect 55111 25632 55120 25666
rect 55068 25623 55120 25632
rect 12130 25116 12182 25125
rect 12130 25082 12139 25116
rect 12139 25082 12173 25116
rect 12173 25082 12182 25116
rect 12130 25073 12182 25082
rect 55068 25116 55120 25125
rect 55068 25082 55077 25116
rect 55077 25082 55111 25116
rect 55111 25082 55120 25116
rect 55068 25073 55120 25082
rect 12130 24876 12182 24885
rect 12130 24842 12139 24876
rect 12139 24842 12173 24876
rect 12173 24842 12182 24876
rect 12130 24833 12182 24842
rect 55068 24876 55120 24885
rect 55068 24842 55077 24876
rect 55077 24842 55111 24876
rect 55111 24842 55120 24876
rect 55068 24833 55120 24842
rect 12130 24326 12182 24335
rect 12130 24292 12139 24326
rect 12139 24292 12173 24326
rect 12173 24292 12182 24326
rect 12130 24283 12182 24292
rect 55068 24326 55120 24335
rect 55068 24292 55077 24326
rect 55077 24292 55111 24326
rect 55111 24292 55120 24326
rect 55068 24283 55120 24292
rect 12130 24086 12182 24095
rect 12130 24052 12139 24086
rect 12139 24052 12173 24086
rect 12173 24052 12182 24086
rect 12130 24043 12182 24052
rect 55068 24086 55120 24095
rect 55068 24052 55077 24086
rect 55077 24052 55111 24086
rect 55111 24052 55120 24086
rect 55068 24043 55120 24052
rect 12130 23536 12182 23545
rect 12130 23502 12139 23536
rect 12139 23502 12173 23536
rect 12173 23502 12182 23536
rect 12130 23493 12182 23502
rect 55068 23536 55120 23545
rect 55068 23502 55077 23536
rect 55077 23502 55111 23536
rect 55111 23502 55120 23536
rect 55068 23493 55120 23502
rect 12130 23296 12182 23305
rect 12130 23262 12139 23296
rect 12139 23262 12173 23296
rect 12173 23262 12182 23296
rect 12130 23253 12182 23262
rect 55068 23296 55120 23305
rect 55068 23262 55077 23296
rect 55077 23262 55111 23296
rect 55111 23262 55120 23296
rect 55068 23253 55120 23262
rect 12130 22746 12182 22755
rect 12130 22712 12139 22746
rect 12139 22712 12173 22746
rect 12173 22712 12182 22746
rect 12130 22703 12182 22712
rect 55068 22746 55120 22755
rect 55068 22712 55077 22746
rect 55077 22712 55111 22746
rect 55111 22712 55120 22746
rect 55068 22703 55120 22712
rect 12130 22506 12182 22515
rect 12130 22472 12139 22506
rect 12139 22472 12173 22506
rect 12173 22472 12182 22506
rect 12130 22463 12182 22472
rect 55068 22506 55120 22515
rect 55068 22472 55077 22506
rect 55077 22472 55111 22506
rect 55111 22472 55120 22506
rect 55068 22463 55120 22472
rect 12130 21956 12182 21965
rect 12130 21922 12139 21956
rect 12139 21922 12173 21956
rect 12173 21922 12182 21956
rect 12130 21913 12182 21922
rect 55068 21956 55120 21965
rect 55068 21922 55077 21956
rect 55077 21922 55111 21956
rect 55111 21922 55120 21956
rect 55068 21913 55120 21922
rect 12130 21716 12182 21725
rect 12130 21682 12139 21716
rect 12139 21682 12173 21716
rect 12173 21682 12182 21716
rect 12130 21673 12182 21682
rect 55068 21716 55120 21725
rect 55068 21682 55077 21716
rect 55077 21682 55111 21716
rect 55111 21682 55120 21716
rect 55068 21673 55120 21682
rect 12130 21166 12182 21175
rect 12130 21132 12139 21166
rect 12139 21132 12173 21166
rect 12173 21132 12182 21166
rect 12130 21123 12182 21132
rect 55068 21166 55120 21175
rect 55068 21132 55077 21166
rect 55077 21132 55111 21166
rect 55111 21132 55120 21166
rect 55068 21123 55120 21132
rect 12130 20926 12182 20935
rect 12130 20892 12139 20926
rect 12139 20892 12173 20926
rect 12173 20892 12182 20926
rect 12130 20883 12182 20892
rect 55068 20926 55120 20935
rect 55068 20892 55077 20926
rect 55077 20892 55111 20926
rect 55111 20892 55120 20926
rect 55068 20883 55120 20892
rect 12130 20376 12182 20385
rect 12130 20342 12139 20376
rect 12139 20342 12173 20376
rect 12173 20342 12182 20376
rect 12130 20333 12182 20342
rect 55068 20376 55120 20385
rect 55068 20342 55077 20376
rect 55077 20342 55111 20376
rect 55111 20342 55120 20376
rect 55068 20333 55120 20342
rect 12130 20136 12182 20145
rect 12130 20102 12139 20136
rect 12139 20102 12173 20136
rect 12173 20102 12182 20136
rect 12130 20093 12182 20102
rect 55068 20136 55120 20145
rect 55068 20102 55077 20136
rect 55077 20102 55111 20136
rect 55111 20102 55120 20136
rect 55068 20093 55120 20102
rect 12130 19586 12182 19595
rect 12130 19552 12139 19586
rect 12139 19552 12173 19586
rect 12173 19552 12182 19586
rect 12130 19543 12182 19552
rect 55068 19586 55120 19595
rect 55068 19552 55077 19586
rect 55077 19552 55111 19586
rect 55111 19552 55120 19586
rect 55068 19543 55120 19552
rect 12130 19346 12182 19355
rect 12130 19312 12139 19346
rect 12139 19312 12173 19346
rect 12173 19312 12182 19346
rect 12130 19303 12182 19312
rect 55068 19346 55120 19355
rect 55068 19312 55077 19346
rect 55077 19312 55111 19346
rect 55111 19312 55120 19346
rect 55068 19303 55120 19312
rect 12130 18796 12182 18805
rect 12130 18762 12139 18796
rect 12139 18762 12173 18796
rect 12173 18762 12182 18796
rect 12130 18753 12182 18762
rect 55068 18796 55120 18805
rect 55068 18762 55077 18796
rect 55077 18762 55111 18796
rect 55111 18762 55120 18796
rect 55068 18753 55120 18762
rect 12130 18556 12182 18565
rect 12130 18522 12139 18556
rect 12139 18522 12173 18556
rect 12173 18522 12182 18556
rect 12130 18513 12182 18522
rect 55068 18556 55120 18565
rect 55068 18522 55077 18556
rect 55077 18522 55111 18556
rect 55111 18522 55120 18556
rect 55068 18513 55120 18522
rect 12130 18006 12182 18015
rect 12130 17972 12139 18006
rect 12139 17972 12173 18006
rect 12173 17972 12182 18006
rect 12130 17963 12182 17972
rect 55068 18006 55120 18015
rect 55068 17972 55077 18006
rect 55077 17972 55111 18006
rect 55111 17972 55120 18006
rect 55068 17963 55120 17972
rect 12130 17766 12182 17775
rect 12130 17732 12139 17766
rect 12139 17732 12173 17766
rect 12173 17732 12182 17766
rect 12130 17723 12182 17732
rect 55068 17766 55120 17775
rect 55068 17732 55077 17766
rect 55077 17732 55111 17766
rect 55111 17732 55120 17766
rect 55068 17723 55120 17732
rect 12130 17216 12182 17225
rect 12130 17182 12139 17216
rect 12139 17182 12173 17216
rect 12173 17182 12182 17216
rect 12130 17173 12182 17182
rect 55068 17216 55120 17225
rect 55068 17182 55077 17216
rect 55077 17182 55111 17216
rect 55111 17182 55120 17216
rect 55068 17173 55120 17182
rect 12130 16976 12182 16985
rect 12130 16942 12139 16976
rect 12139 16942 12173 16976
rect 12173 16942 12182 16976
rect 12130 16933 12182 16942
rect 55068 16976 55120 16985
rect 55068 16942 55077 16976
rect 55077 16942 55111 16976
rect 55111 16942 55120 16976
rect 55068 16933 55120 16942
rect 12130 16426 12182 16435
rect 12130 16392 12139 16426
rect 12139 16392 12173 16426
rect 12173 16392 12182 16426
rect 12130 16383 12182 16392
rect 55068 16426 55120 16435
rect 55068 16392 55077 16426
rect 55077 16392 55111 16426
rect 55111 16392 55120 16426
rect 55068 16383 55120 16392
rect 12130 16186 12182 16195
rect 12130 16152 12139 16186
rect 12139 16152 12173 16186
rect 12173 16152 12182 16186
rect 12130 16143 12182 16152
rect 55068 16186 55120 16195
rect 55068 16152 55077 16186
rect 55077 16152 55111 16186
rect 55111 16152 55120 16186
rect 55068 16143 55120 16152
rect 12130 15636 12182 15645
rect 12130 15602 12139 15636
rect 12139 15602 12173 15636
rect 12173 15602 12182 15636
rect 12130 15593 12182 15602
rect 55068 15636 55120 15645
rect 55068 15602 55077 15636
rect 55077 15602 55111 15636
rect 55111 15602 55120 15636
rect 55068 15593 55120 15602
rect 12130 15396 12182 15405
rect 12130 15362 12139 15396
rect 12139 15362 12173 15396
rect 12173 15362 12182 15396
rect 12130 15353 12182 15362
rect 55068 15396 55120 15405
rect 55068 15362 55077 15396
rect 55077 15362 55111 15396
rect 55111 15362 55120 15396
rect 55068 15353 55120 15362
rect 12130 14846 12182 14855
rect 12130 14812 12139 14846
rect 12139 14812 12173 14846
rect 12173 14812 12182 14846
rect 12130 14803 12182 14812
rect 55068 14846 55120 14855
rect 55068 14812 55077 14846
rect 55077 14812 55111 14846
rect 55111 14812 55120 14846
rect 55068 14803 55120 14812
rect 12130 14606 12182 14615
rect 12130 14572 12139 14606
rect 12139 14572 12173 14606
rect 12173 14572 12182 14606
rect 12130 14563 12182 14572
rect 55068 14606 55120 14615
rect 55068 14572 55077 14606
rect 55077 14572 55111 14606
rect 55111 14572 55120 14606
rect 55068 14563 55120 14572
rect 12130 14056 12182 14065
rect 12130 14022 12139 14056
rect 12139 14022 12173 14056
rect 12173 14022 12182 14056
rect 12130 14013 12182 14022
rect 55068 14056 55120 14065
rect 55068 14022 55077 14056
rect 55077 14022 55111 14056
rect 55111 14022 55120 14056
rect 55068 14013 55120 14022
rect 12130 13816 12182 13825
rect 12130 13782 12139 13816
rect 12139 13782 12173 13816
rect 12173 13782 12182 13816
rect 12130 13773 12182 13782
rect 13551 11973 13603 12025
rect 6840 10709 6892 10718
rect 6840 10675 6849 10709
rect 6849 10675 6883 10709
rect 6883 10675 6892 10709
rect 6840 10666 6892 10675
rect 6840 9219 6892 9228
rect 6840 9185 6849 9219
rect 6849 9185 6883 9219
rect 6883 9185 6892 9219
rect 6840 9176 6892 9185
rect 6840 7881 6892 7890
rect 6840 7847 6849 7881
rect 6849 7847 6883 7881
rect 6883 7847 6892 7881
rect 6840 7838 6892 7847
rect 6840 6391 6892 6400
rect 6840 6357 6849 6391
rect 6849 6357 6883 6391
rect 6883 6357 6892 6391
rect 6840 6348 6892 6357
rect 6840 5053 6892 5062
rect 6840 5019 6849 5053
rect 6849 5019 6883 5053
rect 6883 5019 6892 5053
rect 6840 5010 6892 5019
rect 6840 3563 6892 3572
rect 6840 3529 6849 3563
rect 6849 3529 6883 3563
rect 6883 3529 6892 3563
rect 6840 3520 6892 3529
rect 6840 2225 6892 2234
rect 6840 2191 6849 2225
rect 6849 2191 6883 2225
rect 6883 2191 6892 2225
rect 6840 2182 6892 2191
rect 6840 735 6892 744
rect 6840 701 6849 735
rect 6849 701 6883 735
rect 6883 701 6892 735
rect 6840 692 6892 701
<< metal2 >>
rect 55277 69558 55305 78433
rect 55263 69549 55319 69558
rect 55263 69484 55319 69493
rect 53645 66427 53701 66436
rect 53645 66362 53701 66371
rect 55277 65269 55305 69484
rect 55401 66287 55429 78433
rect 59777 77708 59833 77717
rect 59777 77643 59833 77652
rect 60232 77708 60288 77717
rect 60232 77643 60288 77652
rect 59641 76218 59697 76227
rect 59641 76153 59697 76162
rect 59505 74880 59561 74889
rect 59505 74815 59561 74824
rect 59369 73390 59425 73399
rect 59369 73325 59425 73334
rect 59233 72052 59289 72061
rect 59233 71987 59289 71996
rect 58961 70562 59017 70571
rect 58961 70497 59017 70506
rect 58975 68222 59003 70497
rect 59097 69224 59153 69233
rect 59097 69159 59153 69168
rect 58961 68213 59017 68222
rect 58961 68148 59017 68157
rect 59111 68098 59139 69159
rect 59247 68346 59275 71987
rect 59383 68470 59411 73325
rect 59519 68594 59547 74815
rect 59655 68718 59683 76153
rect 59791 68842 59819 77643
rect 60232 76218 60288 76227
rect 60232 76153 60288 76162
rect 60232 74880 60288 74889
rect 60232 74815 60288 74824
rect 60232 73390 60288 73399
rect 60232 73325 60288 73334
rect 60232 72052 60288 72061
rect 60232 71987 60288 71996
rect 60232 70562 60288 70571
rect 60232 70497 60288 70506
rect 60232 69224 60288 69233
rect 60232 69159 60288 69168
rect 59777 68833 59833 68842
rect 59777 68768 59833 68777
rect 59641 68709 59697 68718
rect 59641 68644 59697 68653
rect 59505 68585 59561 68594
rect 59505 68520 59561 68529
rect 59369 68461 59425 68470
rect 59369 68396 59425 68405
rect 59233 68337 59289 68346
rect 59233 68272 59289 68281
rect 59097 68089 59153 68098
rect 59097 68024 59153 68033
rect 58961 67965 59017 67974
rect 58961 67900 59017 67909
rect 58975 67743 59003 67900
rect 58961 67734 59017 67743
rect 58961 67669 59017 67678
rect 60232 67734 60288 67743
rect 60232 67669 60288 67678
rect 55387 66278 55443 66287
rect 55387 66213 55443 66222
rect 55401 65269 55429 66213
rect 59262 64764 59290 64792
rect 55068 64625 55120 64631
rect 54967 64592 55068 64620
rect 55068 64567 55120 64573
rect 12130 64385 12182 64391
rect 55068 64385 55120 64391
rect 54967 64338 55068 64366
rect 12130 64327 12182 64333
rect 55068 64327 55120 64333
rect 12142 64146 12170 64327
rect 12142 64118 12283 64146
rect 12142 64022 12283 64050
rect 12142 63841 12170 64022
rect 12130 63835 12182 63841
rect 55068 63835 55120 63841
rect 54967 63802 55068 63830
rect 12130 63777 12182 63783
rect 55068 63777 55120 63783
rect 12130 63595 12182 63601
rect 55068 63595 55120 63601
rect 54967 63548 55068 63576
rect 12130 63537 12182 63543
rect 55068 63537 55120 63543
rect 12142 63356 12170 63537
rect 12142 63328 12283 63356
rect 12142 63232 12283 63260
rect 12142 63051 12170 63232
rect 12130 63045 12182 63051
rect 55068 63045 55120 63051
rect 54967 63012 55068 63040
rect 12130 62987 12182 62993
rect 55068 62987 55120 62993
rect 12130 62805 12182 62811
rect 55068 62805 55120 62811
rect 54967 62758 55068 62786
rect 12130 62747 12182 62753
rect 55068 62747 55120 62753
rect 12142 62566 12170 62747
rect 12142 62538 12283 62566
rect 12142 62442 12283 62470
rect 12142 62261 12170 62442
rect 12130 62255 12182 62261
rect 55068 62255 55120 62261
rect 54967 62222 55068 62250
rect 12130 62197 12182 62203
rect 55068 62197 55120 62203
rect 12130 62015 12182 62021
rect 55068 62015 55120 62021
rect 54967 61968 55068 61996
rect 12130 61957 12182 61963
rect 55068 61957 55120 61963
rect 12142 61776 12170 61957
rect 12142 61748 12283 61776
rect 12142 61652 12283 61680
rect 12142 61471 12170 61652
rect 12130 61465 12182 61471
rect 55068 61465 55120 61471
rect 54967 61432 55068 61460
rect 12130 61407 12182 61413
rect 55068 61407 55120 61413
rect 12130 61225 12182 61231
rect 55068 61225 55120 61231
rect 54967 61178 55068 61206
rect 12130 61167 12182 61173
rect 55068 61167 55120 61173
rect 12142 60986 12170 61167
rect 12142 60958 12283 60986
rect 12142 60862 12283 60890
rect 12142 60681 12170 60862
rect 12130 60675 12182 60681
rect 55068 60675 55120 60681
rect 54967 60642 55068 60670
rect 12130 60617 12182 60623
rect 55068 60617 55120 60623
rect 12130 60435 12182 60441
rect 55068 60435 55120 60441
rect 54967 60388 55068 60416
rect 12130 60377 12182 60383
rect 55068 60377 55120 60383
rect 12142 60196 12170 60377
rect 12142 60168 12283 60196
rect 12142 60072 12283 60100
rect 12142 59891 12170 60072
rect 12130 59885 12182 59891
rect 55068 59885 55120 59891
rect 54967 59852 55068 59880
rect 12130 59827 12182 59833
rect 55068 59827 55120 59833
rect 12130 59645 12182 59651
rect 55068 59645 55120 59651
rect 54967 59598 55068 59626
rect 12130 59587 12182 59593
rect 55068 59587 55120 59593
rect 12142 59406 12170 59587
rect 12142 59378 12283 59406
rect 12142 59282 12283 59310
rect 12142 59101 12170 59282
rect 12130 59095 12182 59101
rect 55068 59095 55120 59101
rect 54967 59062 55068 59090
rect 12130 59037 12182 59043
rect 55068 59037 55120 59043
rect 12130 58855 12182 58861
rect 55068 58855 55120 58861
rect 54967 58808 55068 58836
rect 12130 58797 12182 58803
rect 55068 58797 55120 58803
rect 12142 58616 12170 58797
rect 12142 58588 12283 58616
rect 12142 58492 12283 58520
rect 12142 58311 12170 58492
rect 12130 58305 12182 58311
rect 55068 58305 55120 58311
rect 54967 58272 55068 58300
rect 12130 58247 12182 58253
rect 55068 58247 55120 58253
rect 12130 58065 12182 58071
rect 55068 58065 55120 58071
rect 54967 58018 55068 58046
rect 12130 58007 12182 58013
rect 55068 58007 55120 58013
rect 12142 57826 12170 58007
rect 12142 57798 12283 57826
rect 12142 57702 12283 57730
rect 12142 57521 12170 57702
rect 12130 57515 12182 57521
rect 55068 57515 55120 57521
rect 54967 57482 55068 57510
rect 12130 57457 12182 57463
rect 55068 57457 55120 57463
rect 12130 57275 12182 57281
rect 55068 57275 55120 57281
rect 54967 57228 55068 57256
rect 12130 57217 12182 57223
rect 55068 57217 55120 57223
rect 12142 57036 12170 57217
rect 12142 57008 12283 57036
rect 12142 56912 12283 56940
rect 12142 56731 12170 56912
rect 12130 56725 12182 56731
rect 55068 56725 55120 56731
rect 54967 56692 55068 56720
rect 12130 56667 12182 56673
rect 55068 56667 55120 56673
rect 12130 56485 12182 56491
rect 55068 56485 55120 56491
rect 54967 56438 55068 56466
rect 12130 56427 12182 56433
rect 55068 56427 55120 56433
rect 12142 56246 12170 56427
rect 12142 56218 12283 56246
rect 12142 56122 12283 56150
rect 12142 55941 12170 56122
rect 12130 55935 12182 55941
rect 55068 55935 55120 55941
rect 54967 55902 55068 55930
rect 12130 55877 12182 55883
rect 55068 55877 55120 55883
rect 12130 55695 12182 55701
rect 55068 55695 55120 55701
rect 54967 55648 55068 55676
rect 12130 55637 12182 55643
rect 55068 55637 55120 55643
rect 12142 55456 12170 55637
rect 12142 55428 12283 55456
rect 12142 55332 12283 55360
rect 12142 55151 12170 55332
rect 12130 55145 12182 55151
rect 55068 55145 55120 55151
rect 54967 55112 55068 55140
rect 12130 55087 12182 55093
rect 55068 55087 55120 55093
rect 12130 54905 12182 54911
rect 55068 54905 55120 54911
rect 54967 54858 55068 54886
rect 12130 54847 12182 54853
rect 55068 54847 55120 54853
rect 12142 54666 12170 54847
rect 12142 54638 12283 54666
rect 12142 54542 12283 54570
rect 12142 54361 12170 54542
rect 12130 54355 12182 54361
rect 55068 54355 55120 54361
rect 54967 54322 55068 54350
rect 12130 54297 12182 54303
rect 55068 54297 55120 54303
rect 12130 54115 12182 54121
rect 55068 54115 55120 54121
rect 54967 54068 55068 54096
rect 12130 54057 12182 54063
rect 55068 54057 55120 54063
rect 12142 53876 12170 54057
rect 12142 53848 12283 53876
rect 12142 53752 12283 53780
rect 12142 53571 12170 53752
rect 12130 53565 12182 53571
rect 55068 53565 55120 53571
rect 54967 53532 55068 53560
rect 12130 53507 12182 53513
rect 55068 53507 55120 53513
rect 12130 53325 12182 53331
rect 55068 53325 55120 53331
rect 54967 53278 55068 53306
rect 12130 53267 12182 53273
rect 55068 53267 55120 53273
rect 12142 53086 12170 53267
rect 12142 53058 12283 53086
rect 12142 52962 12283 52990
rect 12142 52781 12170 52962
rect 12130 52775 12182 52781
rect 55068 52775 55120 52781
rect 54967 52742 55068 52770
rect 12130 52717 12182 52723
rect 55068 52717 55120 52723
rect 12130 52535 12182 52541
rect 55068 52535 55120 52541
rect 54967 52488 55068 52516
rect 12130 52477 12182 52483
rect 55068 52477 55120 52483
rect 12142 52296 12170 52477
rect 12142 52268 12283 52296
rect 12142 52172 12283 52200
rect 12142 51991 12170 52172
rect 12130 51985 12182 51991
rect 55068 51985 55120 51991
rect 54967 51952 55068 51980
rect 12130 51927 12182 51933
rect 55068 51927 55120 51933
rect 12130 51745 12182 51751
rect 55068 51745 55120 51751
rect 54967 51698 55068 51726
rect 12130 51687 12182 51693
rect 55068 51687 55120 51693
rect 12142 51506 12170 51687
rect 12142 51478 12283 51506
rect 12142 51382 12283 51410
rect 12142 51201 12170 51382
rect 12130 51195 12182 51201
rect 55068 51195 55120 51201
rect 54967 51162 55068 51190
rect 12130 51137 12182 51143
rect 55068 51137 55120 51143
rect 12130 50955 12182 50961
rect 55068 50955 55120 50961
rect 54967 50908 55068 50936
rect 12130 50897 12182 50903
rect 55068 50897 55120 50903
rect 12142 50716 12170 50897
rect 12142 50688 12283 50716
rect 12142 50592 12283 50620
rect 12142 50411 12170 50592
rect 12130 50405 12182 50411
rect 55068 50405 55120 50411
rect 54967 50372 55068 50400
rect 12130 50347 12182 50353
rect 55068 50347 55120 50353
rect 12130 50165 12182 50171
rect 55068 50165 55120 50171
rect 54967 50118 55068 50146
rect 12130 50107 12182 50113
rect 55068 50107 55120 50113
rect 12142 49926 12170 50107
rect 12142 49898 12283 49926
rect 12142 49802 12283 49830
rect 12142 49621 12170 49802
rect 12130 49615 12182 49621
rect 55068 49615 55120 49621
rect 54967 49582 55068 49610
rect 12130 49557 12182 49563
rect 55068 49557 55120 49563
rect 12130 49375 12182 49381
rect 55068 49375 55120 49381
rect 54967 49328 55068 49356
rect 12130 49317 12182 49323
rect 55068 49317 55120 49323
rect 12142 49136 12170 49317
rect 12142 49108 12283 49136
rect 12142 49012 12283 49040
rect 12142 48831 12170 49012
rect 12130 48825 12182 48831
rect 55068 48825 55120 48831
rect 54967 48792 55068 48820
rect 12130 48767 12182 48773
rect 55068 48767 55120 48773
rect 12130 48585 12182 48591
rect 55068 48585 55120 48591
rect 54967 48538 55068 48566
rect 12130 48527 12182 48533
rect 55068 48527 55120 48533
rect 12142 48346 12170 48527
rect 12142 48318 12283 48346
rect 12142 48222 12283 48250
rect 12142 48041 12170 48222
rect 12130 48035 12182 48041
rect 55068 48035 55120 48041
rect 54967 48002 55068 48030
rect 12130 47977 12182 47983
rect 55068 47977 55120 47983
rect 12130 47795 12182 47801
rect 55068 47795 55120 47801
rect 54967 47748 55068 47776
rect 12130 47737 12182 47743
rect 55068 47737 55120 47743
rect 12142 47556 12170 47737
rect 12142 47528 12283 47556
rect 12142 47432 12283 47460
rect 12142 47251 12170 47432
rect 12130 47245 12182 47251
rect 55068 47245 55120 47251
rect 54967 47212 55068 47240
rect 12130 47187 12182 47193
rect 55068 47187 55120 47193
rect 12130 47005 12182 47011
rect 55068 47005 55120 47011
rect 54967 46958 55068 46986
rect 12130 46947 12182 46953
rect 55068 46947 55120 46953
rect 12142 46766 12170 46947
rect 12142 46738 12283 46766
rect 12142 46642 12283 46670
rect 12142 46461 12170 46642
rect 12130 46455 12182 46461
rect 55068 46455 55120 46461
rect 54967 46422 55068 46450
rect 12130 46397 12182 46403
rect 55068 46397 55120 46403
rect 12130 46215 12182 46221
rect 55068 46215 55120 46221
rect 54967 46168 55068 46196
rect 12130 46157 12182 46163
rect 55068 46157 55120 46163
rect 12142 45976 12170 46157
rect 12142 45948 12283 45976
rect 12142 45852 12283 45880
rect 12142 45671 12170 45852
rect 12130 45665 12182 45671
rect 55068 45665 55120 45671
rect 54967 45632 55068 45660
rect 12130 45607 12182 45613
rect 55068 45607 55120 45613
rect 12130 45425 12182 45431
rect 55068 45425 55120 45431
rect 54967 45378 55068 45406
rect 12130 45367 12182 45373
rect 55068 45367 55120 45373
rect 12142 45186 12170 45367
rect 12142 45158 12283 45186
rect 12142 45062 12283 45090
rect 12142 44881 12170 45062
rect 12130 44875 12182 44881
rect 55068 44875 55120 44881
rect 54967 44842 55068 44870
rect 12130 44817 12182 44823
rect 55068 44817 55120 44823
rect 12130 44635 12182 44641
rect 55068 44635 55120 44641
rect 54967 44588 55068 44616
rect 12130 44577 12182 44583
rect 55068 44577 55120 44583
rect 12142 44396 12170 44577
rect 12142 44368 12283 44396
rect 12142 44272 12283 44300
rect 12142 44091 12170 44272
rect 12130 44085 12182 44091
rect 55068 44085 55120 44091
rect 54967 44052 55068 44080
rect 12130 44027 12182 44033
rect 55068 44027 55120 44033
rect 12130 43845 12182 43851
rect 55068 43845 55120 43851
rect 54967 43798 55068 43826
rect 12130 43787 12182 43793
rect 55068 43787 55120 43793
rect 12142 43606 12170 43787
rect 12142 43578 12283 43606
rect 12142 43482 12283 43510
rect 12142 43301 12170 43482
rect 12130 43295 12182 43301
rect 55068 43295 55120 43301
rect 54967 43262 55068 43290
rect 12130 43237 12182 43243
rect 55068 43237 55120 43243
rect 12130 43055 12182 43061
rect 55068 43055 55120 43061
rect 54967 43008 55068 43036
rect 12130 42997 12182 43003
rect 55068 42997 55120 43003
rect 12142 42816 12170 42997
rect 12142 42788 12283 42816
rect 12142 42692 12283 42720
rect 12142 42511 12170 42692
rect 12130 42505 12182 42511
rect 55068 42505 55120 42511
rect 54967 42472 55068 42500
rect 12130 42447 12182 42453
rect 55068 42447 55120 42453
rect 12130 42265 12182 42271
rect 55068 42265 55120 42271
rect 54967 42218 55068 42246
rect 12130 42207 12182 42213
rect 55068 42207 55120 42213
rect 12142 42026 12170 42207
rect 12142 41998 12283 42026
rect 12142 41902 12283 41930
rect 12142 41721 12170 41902
rect 12130 41715 12182 41721
rect 55068 41715 55120 41721
rect 54967 41682 55068 41710
rect 12130 41657 12182 41663
rect 55068 41657 55120 41663
rect 12130 41475 12182 41481
rect 55068 41475 55120 41481
rect 54967 41428 55068 41456
rect 12130 41417 12182 41423
rect 55068 41417 55120 41423
rect 12142 41236 12170 41417
rect 12142 41208 12283 41236
rect 12142 41112 12283 41140
rect 12142 40931 12170 41112
rect 12130 40925 12182 40931
rect 55068 40925 55120 40931
rect 54967 40892 55068 40920
rect 12130 40867 12182 40873
rect 55068 40867 55120 40873
rect 12130 40685 12182 40691
rect 55068 40685 55120 40691
rect 54967 40638 55068 40666
rect 12130 40627 12182 40633
rect 55068 40627 55120 40633
rect 12142 40446 12170 40627
rect 12142 40418 12283 40446
rect 12142 40322 12283 40350
rect 12142 40141 12170 40322
rect 12130 40135 12182 40141
rect 55068 40135 55120 40141
rect 54967 40102 55068 40130
rect 12130 40077 12182 40083
rect 55068 40077 55120 40083
rect 12130 39895 12182 39901
rect 55068 39895 55120 39901
rect 54967 39848 55068 39876
rect 12130 39837 12182 39843
rect 55068 39837 55120 39843
rect 12142 39656 12170 39837
rect 12142 39628 12283 39656
rect 12142 39532 12283 39560
rect 12142 39351 12170 39532
rect 12130 39345 12182 39351
rect 55068 39345 55120 39351
rect 54967 39312 55068 39340
rect 12130 39287 12182 39293
rect 55068 39287 55120 39293
rect 12130 39105 12182 39111
rect 55068 39105 55120 39111
rect 54967 39058 55068 39086
rect 12130 39047 12182 39053
rect 55068 39047 55120 39053
rect 12142 38866 12170 39047
rect 12142 38838 12283 38866
rect 12142 38742 12283 38770
rect 12142 38561 12170 38742
rect 12130 38555 12182 38561
rect 55068 38555 55120 38561
rect 54967 38522 55068 38550
rect 12130 38497 12182 38503
rect 55068 38497 55120 38503
rect 12130 38315 12182 38321
rect 55068 38315 55120 38321
rect 54967 38268 55068 38296
rect 12130 38257 12182 38263
rect 55068 38257 55120 38263
rect 12142 38076 12170 38257
rect 12142 38048 12283 38076
rect 12142 37952 12283 37980
rect 12142 37771 12170 37952
rect 12130 37765 12182 37771
rect 55068 37765 55120 37771
rect 54967 37732 55068 37760
rect 12130 37707 12182 37713
rect 55068 37707 55120 37713
rect 12130 37525 12182 37531
rect 55068 37525 55120 37531
rect 54967 37478 55068 37506
rect 12130 37467 12182 37473
rect 55068 37467 55120 37473
rect 12142 37286 12170 37467
rect 12142 37258 12283 37286
rect 12142 37162 12283 37190
rect 12142 36981 12170 37162
rect 12130 36975 12182 36981
rect 55068 36975 55120 36981
rect 54967 36942 55068 36970
rect 12130 36917 12182 36923
rect 55068 36917 55120 36923
rect 12130 36735 12182 36741
rect 55068 36735 55120 36741
rect 54967 36688 55068 36716
rect 12130 36677 12182 36683
rect 55068 36677 55120 36683
rect 12142 36496 12170 36677
rect 12142 36468 12283 36496
rect 12142 36372 12283 36400
rect 12142 36191 12170 36372
rect 12130 36185 12182 36191
rect 55068 36185 55120 36191
rect 54967 36152 55068 36180
rect 12130 36127 12182 36133
rect 55068 36127 55120 36133
rect 12130 35945 12182 35951
rect 55068 35945 55120 35951
rect 54967 35898 55068 35926
rect 12130 35887 12182 35893
rect 55068 35887 55120 35893
rect 12142 35706 12170 35887
rect 12142 35678 12283 35706
rect 12142 35582 12283 35610
rect 12142 35401 12170 35582
rect 12130 35395 12182 35401
rect 55068 35395 55120 35401
rect 54967 35362 55068 35390
rect 12130 35337 12182 35343
rect 55068 35337 55120 35343
rect 12130 35155 12182 35161
rect 55068 35155 55120 35161
rect 54967 35108 55068 35136
rect 12130 35097 12182 35103
rect 55068 35097 55120 35103
rect 12142 34916 12170 35097
rect 12142 34888 12283 34916
rect 12142 34792 12283 34820
rect 12142 34611 12170 34792
rect 12130 34605 12182 34611
rect 55068 34605 55120 34611
rect 54967 34572 55068 34600
rect 12130 34547 12182 34553
rect 55068 34547 55120 34553
rect 12130 34365 12182 34371
rect 55068 34365 55120 34371
rect 54967 34318 55068 34346
rect 12130 34307 12182 34313
rect 55068 34307 55120 34313
rect 12142 34126 12170 34307
rect 12142 34098 12283 34126
rect 12142 34002 12283 34030
rect 12142 33821 12170 34002
rect 12130 33815 12182 33821
rect 55068 33815 55120 33821
rect 54967 33782 55068 33810
rect 12130 33757 12182 33763
rect 55068 33757 55120 33763
rect 12130 33575 12182 33581
rect 55068 33575 55120 33581
rect 54967 33528 55068 33556
rect 12130 33517 12182 33523
rect 55068 33517 55120 33523
rect 12142 33336 12170 33517
rect 12142 33308 12283 33336
rect 12142 33212 12283 33240
rect 12142 33031 12170 33212
rect 12130 33025 12182 33031
rect 55068 33025 55120 33031
rect 54967 32992 55068 33020
rect 12130 32967 12182 32973
rect 55068 32967 55120 32973
rect 12130 32785 12182 32791
rect 55068 32785 55120 32791
rect 54967 32738 55068 32766
rect 12130 32727 12182 32733
rect 55068 32727 55120 32733
rect 12142 32546 12170 32727
rect 12142 32518 12283 32546
rect 12142 32422 12283 32450
rect 12142 32241 12170 32422
rect 12130 32235 12182 32241
rect 55068 32235 55120 32241
rect 54967 32202 55068 32230
rect 12130 32177 12182 32183
rect 55068 32177 55120 32183
rect 12130 31995 12182 32001
rect 55068 31995 55120 32001
rect 54967 31948 55068 31976
rect 12130 31937 12182 31943
rect 55068 31937 55120 31943
rect 12142 31756 12170 31937
rect 12142 31728 12283 31756
rect 12142 31632 12283 31660
rect 12142 31451 12170 31632
rect 12130 31445 12182 31451
rect 55068 31445 55120 31451
rect 54967 31412 55068 31440
rect 12130 31387 12182 31393
rect 55068 31387 55120 31393
rect 12130 31205 12182 31211
rect 55068 31205 55120 31211
rect 54967 31158 55068 31186
rect 12130 31147 12182 31153
rect 55068 31147 55120 31153
rect 12142 30966 12170 31147
rect 12142 30938 12283 30966
rect 12142 30842 12283 30870
rect 12142 30661 12170 30842
rect 12130 30655 12182 30661
rect 55068 30655 55120 30661
rect 54967 30622 55068 30650
rect 12130 30597 12182 30603
rect 55068 30597 55120 30603
rect 12130 30415 12182 30421
rect 55068 30415 55120 30421
rect 54967 30368 55068 30396
rect 12130 30357 12182 30363
rect 55068 30357 55120 30363
rect 12142 30176 12170 30357
rect 12142 30148 12283 30176
rect 12142 30052 12283 30080
rect 12142 29871 12170 30052
rect 12130 29865 12182 29871
rect 55068 29865 55120 29871
rect 54967 29832 55068 29860
rect 12130 29807 12182 29813
rect 55068 29807 55120 29813
rect 12130 29625 12182 29631
rect 55068 29625 55120 29631
rect 54967 29578 55068 29606
rect 12130 29567 12182 29573
rect 55068 29567 55120 29573
rect 12142 29386 12170 29567
rect 12142 29358 12283 29386
rect 12142 29262 12283 29290
rect 12142 29081 12170 29262
rect 12130 29075 12182 29081
rect 55068 29075 55120 29081
rect 54967 29042 55068 29070
rect 12130 29017 12182 29023
rect 55068 29017 55120 29023
rect 12130 28835 12182 28841
rect 55068 28835 55120 28841
rect 54967 28788 55068 28816
rect 12130 28777 12182 28783
rect 55068 28777 55120 28783
rect 12142 28596 12170 28777
rect 12142 28568 12283 28596
rect 12142 28472 12283 28500
rect 12142 28291 12170 28472
rect 12130 28285 12182 28291
rect 55068 28285 55120 28291
rect 54967 28252 55068 28280
rect 12130 28227 12182 28233
rect 55068 28227 55120 28233
rect 12130 28045 12182 28051
rect 55068 28045 55120 28051
rect 54967 27998 55068 28026
rect 12130 27987 12182 27993
rect 55068 27987 55120 27993
rect 12142 27806 12170 27987
rect 12142 27778 12283 27806
rect 12142 27682 12283 27710
rect 12142 27501 12170 27682
rect 12130 27495 12182 27501
rect 55068 27495 55120 27501
rect 54967 27462 55068 27490
rect 12130 27437 12182 27443
rect 55068 27437 55120 27443
rect 12130 27255 12182 27261
rect 55068 27255 55120 27261
rect 54967 27208 55068 27236
rect 12130 27197 12182 27203
rect 55068 27197 55120 27203
rect 12142 27016 12170 27197
rect 12142 26988 12283 27016
rect 12142 26892 12283 26920
rect 12142 26711 12170 26892
rect 12130 26705 12182 26711
rect 55068 26705 55120 26711
rect 54967 26672 55068 26700
rect 12130 26647 12182 26653
rect 55068 26647 55120 26653
rect 12130 26465 12182 26471
rect 55068 26465 55120 26471
rect 54967 26418 55068 26446
rect 12130 26407 12182 26413
rect 55068 26407 55120 26413
rect 12142 26226 12170 26407
rect 12142 26198 12283 26226
rect 12142 26102 12283 26130
rect 12142 25921 12170 26102
rect 12130 25915 12182 25921
rect 55068 25915 55120 25921
rect 54967 25882 55068 25910
rect 12130 25857 12182 25863
rect 55068 25857 55120 25863
rect 12130 25675 12182 25681
rect 55068 25675 55120 25681
rect 54967 25628 55068 25656
rect 12130 25617 12182 25623
rect 55068 25617 55120 25623
rect 12142 25436 12170 25617
rect 12142 25408 12283 25436
rect 12142 25312 12283 25340
rect 12142 25131 12170 25312
rect 12130 25125 12182 25131
rect 55068 25125 55120 25131
rect 54967 25092 55068 25120
rect 12130 25067 12182 25073
rect 55068 25067 55120 25073
rect 12130 24885 12182 24891
rect 55068 24885 55120 24891
rect 54967 24838 55068 24866
rect 12130 24827 12182 24833
rect 55068 24827 55120 24833
rect 12142 24646 12170 24827
rect 12142 24618 12283 24646
rect 12142 24522 12283 24550
rect 12142 24341 12170 24522
rect 12130 24335 12182 24341
rect 55068 24335 55120 24341
rect 54967 24302 55068 24330
rect 12130 24277 12182 24283
rect 55068 24277 55120 24283
rect 12130 24095 12182 24101
rect 55068 24095 55120 24101
rect 54967 24048 55068 24076
rect 12130 24037 12182 24043
rect 55068 24037 55120 24043
rect 12142 23856 12170 24037
rect 12142 23828 12283 23856
rect 12142 23732 12283 23760
rect 12142 23551 12170 23732
rect 12130 23545 12182 23551
rect 55068 23545 55120 23551
rect 54967 23512 55068 23540
rect 12130 23487 12182 23493
rect 55068 23487 55120 23493
rect 12130 23305 12182 23311
rect 55068 23305 55120 23311
rect 54967 23258 55068 23286
rect 12130 23247 12182 23253
rect 55068 23247 55120 23253
rect 12142 23066 12170 23247
rect 12142 23038 12283 23066
rect 12142 22942 12283 22970
rect 12142 22761 12170 22942
rect 12130 22755 12182 22761
rect 55068 22755 55120 22761
rect 54967 22722 55068 22750
rect 12130 22697 12182 22703
rect 55068 22697 55120 22703
rect 12130 22515 12182 22521
rect 55068 22515 55120 22521
rect 54967 22468 55068 22496
rect 12130 22457 12182 22463
rect 55068 22457 55120 22463
rect 12142 22276 12170 22457
rect 12142 22248 12283 22276
rect 12142 22152 12283 22180
rect 12142 21971 12170 22152
rect 12130 21965 12182 21971
rect 55068 21965 55120 21971
rect 54967 21932 55068 21960
rect 12130 21907 12182 21913
rect 55068 21907 55120 21913
rect 12130 21725 12182 21731
rect 55068 21725 55120 21731
rect 54967 21678 55068 21706
rect 12130 21667 12182 21673
rect 55068 21667 55120 21673
rect 12142 21486 12170 21667
rect 12142 21458 12283 21486
rect 12142 21362 12283 21390
rect 12142 21181 12170 21362
rect 12130 21175 12182 21181
rect 55068 21175 55120 21181
rect 54967 21142 55068 21170
rect 12130 21117 12182 21123
rect 55068 21117 55120 21123
rect 12130 20935 12182 20941
rect 55068 20935 55120 20941
rect 54967 20888 55068 20916
rect 12130 20877 12182 20883
rect 55068 20877 55120 20883
rect 12142 20696 12170 20877
rect 12142 20668 12283 20696
rect 12142 20572 12283 20600
rect 12142 20391 12170 20572
rect 12130 20385 12182 20391
rect 55068 20385 55120 20391
rect 54967 20352 55068 20380
rect 12130 20327 12182 20333
rect 55068 20327 55120 20333
rect 12130 20145 12182 20151
rect 55068 20145 55120 20151
rect 54967 20098 55068 20126
rect 12130 20087 12182 20093
rect 55068 20087 55120 20093
rect 12142 19906 12170 20087
rect 12142 19878 12283 19906
rect 12142 19782 12283 19810
rect 12142 19601 12170 19782
rect 12130 19595 12182 19601
rect 55068 19595 55120 19601
rect 54967 19562 55068 19590
rect 12130 19537 12182 19543
rect 55068 19537 55120 19543
rect 12130 19355 12182 19361
rect 55068 19355 55120 19361
rect 54967 19308 55068 19336
rect 12130 19297 12182 19303
rect 55068 19297 55120 19303
rect 12142 19116 12170 19297
rect 12142 19088 12283 19116
rect 12142 18992 12283 19020
rect 12142 18811 12170 18992
rect 12130 18805 12182 18811
rect 55068 18805 55120 18811
rect 54967 18772 55068 18800
rect 12130 18747 12182 18753
rect 55068 18747 55120 18753
rect 12130 18565 12182 18571
rect 55068 18565 55120 18571
rect 54967 18518 55068 18546
rect 12130 18507 12182 18513
rect 55068 18507 55120 18513
rect 12142 18326 12170 18507
rect 12142 18298 12283 18326
rect 12142 18202 12283 18230
rect 12142 18021 12170 18202
rect 12130 18015 12182 18021
rect 55068 18015 55120 18021
rect 54967 17982 55068 18010
rect 12130 17957 12182 17963
rect 55068 17957 55120 17963
rect 12130 17775 12182 17781
rect 55068 17775 55120 17781
rect 54967 17728 55068 17756
rect 12130 17717 12182 17723
rect 55068 17717 55120 17723
rect 12142 17536 12170 17717
rect 12142 17508 12283 17536
rect 12142 17412 12283 17440
rect 12142 17231 12170 17412
rect 12130 17225 12182 17231
rect 55068 17225 55120 17231
rect 54967 17192 55068 17220
rect 12130 17167 12182 17173
rect 55068 17167 55120 17173
rect 12130 16985 12182 16991
rect 55068 16985 55120 16991
rect 54967 16938 55068 16966
rect 12130 16927 12182 16933
rect 55068 16927 55120 16933
rect 12142 16746 12170 16927
rect 12142 16718 12283 16746
rect 12142 16622 12283 16650
rect 12142 16441 12170 16622
rect 12130 16435 12182 16441
rect 55068 16435 55120 16441
rect 54967 16402 55068 16430
rect 12130 16377 12182 16383
rect 55068 16377 55120 16383
rect 12130 16195 12182 16201
rect 55068 16195 55120 16201
rect 54967 16148 55068 16176
rect 12130 16137 12182 16143
rect 55068 16137 55120 16143
rect 12142 15956 12170 16137
rect 12142 15928 12283 15956
rect 12142 15832 12283 15860
rect 12142 15651 12170 15832
rect 12130 15645 12182 15651
rect 55068 15645 55120 15651
rect 54967 15612 55068 15640
rect 12130 15587 12182 15593
rect 55068 15587 55120 15593
rect 12130 15405 12182 15411
rect 55068 15405 55120 15411
rect 54967 15358 55068 15386
rect 12130 15347 12182 15353
rect 55068 15347 55120 15353
rect 12142 15166 12170 15347
rect 12142 15138 12283 15166
rect 12142 15042 12283 15070
rect 12142 14861 12170 15042
rect 12130 14855 12182 14861
rect 55068 14855 55120 14861
rect 54967 14822 55068 14850
rect 12130 14797 12182 14803
rect 55068 14797 55120 14803
rect 12130 14615 12182 14621
rect 55068 14615 55120 14621
rect 54967 14568 55068 14596
rect 12130 14557 12182 14563
rect 55068 14557 55120 14563
rect 12142 14376 12170 14557
rect 12142 14348 12283 14376
rect 12142 14252 12283 14280
rect 12142 14071 12170 14252
rect 12130 14065 12182 14071
rect 55068 14065 55120 14071
rect 54967 14032 55068 14060
rect 12130 14007 12182 14013
rect 55068 14007 55120 14013
rect 12130 13825 12182 13831
rect 12130 13767 12182 13773
rect 7960 13606 7988 13634
rect 12142 13586 12170 13767
rect 12142 13558 12283 13586
rect 11663 12185 11691 13129
rect 11649 12176 11705 12185
rect 11649 12111 11705 12120
rect 6838 10720 6894 10729
rect 6838 10655 6894 10664
rect 7117 10720 7173 10729
rect 7117 10655 7173 10664
rect 7131 10498 7159 10655
rect 7117 10489 7173 10498
rect 7117 10424 7173 10433
rect 7933 10365 7989 10374
rect 7933 10300 7989 10309
rect 7797 10241 7853 10250
rect 7797 10176 7853 10185
rect 7661 10117 7717 10126
rect 7661 10052 7717 10061
rect 7525 9993 7581 10002
rect 7525 9928 7581 9937
rect 7389 9869 7445 9878
rect 7389 9804 7445 9813
rect 7253 9745 7309 9754
rect 7253 9680 7309 9689
rect 7117 9621 7173 9630
rect 7117 9556 7173 9565
rect 6838 9230 6894 9239
rect 6838 9165 6894 9174
rect 6838 7892 6894 7901
rect 6838 7827 6894 7836
rect 6838 6402 6894 6411
rect 6838 6337 6894 6346
rect 6838 5064 6894 5073
rect 6838 4999 6894 5008
rect 6838 3574 6894 3583
rect 6838 3509 6894 3518
rect 6838 2236 6894 2245
rect 6838 2171 6894 2180
rect 7131 755 7159 9556
rect 7267 2245 7295 9680
rect 7403 3583 7431 9804
rect 7539 5073 7567 9928
rect 7675 6411 7703 10052
rect 7811 7901 7839 10176
rect 7947 9239 7975 10300
rect 7933 9230 7989 9239
rect 7933 9165 7989 9174
rect 7797 7892 7853 7901
rect 7797 7827 7853 7836
rect 7661 6402 7717 6411
rect 7661 6337 7717 6346
rect 7525 5064 7581 5073
rect 7525 4999 7581 5008
rect 7389 3574 7445 3583
rect 7389 3509 7445 3518
rect 7253 2236 7309 2245
rect 7253 2171 7309 2180
rect 6838 746 6894 755
rect 6838 681 6894 690
rect 7117 746 7173 755
rect 7117 681 7173 690
rect 11663 49 11691 12111
rect 11787 8914 11815 13129
rect 11773 8905 11829 8914
rect 11773 8840 11829 8849
rect 11787 49 11815 8840
rect 11911 3603 11939 13129
rect 13549 12027 13605 12036
rect 13549 11962 13605 11971
rect 11897 3594 11953 3603
rect 11897 3529 11953 3538
rect 11911 49 11939 3529
rect 13643 3304 13671 3332
<< via2 >>
rect 55263 69493 55319 69549
rect 53645 66425 53701 66427
rect 53645 66373 53647 66425
rect 53647 66373 53699 66425
rect 53699 66373 53701 66425
rect 53645 66371 53701 66373
rect 59777 77652 59833 77708
rect 60232 77706 60288 77708
rect 60232 77654 60234 77706
rect 60234 77654 60286 77706
rect 60286 77654 60288 77706
rect 60232 77652 60288 77654
rect 59641 76162 59697 76218
rect 59505 74824 59561 74880
rect 59369 73334 59425 73390
rect 59233 71996 59289 72052
rect 58961 70506 59017 70562
rect 59097 69168 59153 69224
rect 58961 68157 59017 68213
rect 60232 76216 60288 76218
rect 60232 76164 60234 76216
rect 60234 76164 60286 76216
rect 60286 76164 60288 76216
rect 60232 76162 60288 76164
rect 60232 74878 60288 74880
rect 60232 74826 60234 74878
rect 60234 74826 60286 74878
rect 60286 74826 60288 74878
rect 60232 74824 60288 74826
rect 60232 73388 60288 73390
rect 60232 73336 60234 73388
rect 60234 73336 60286 73388
rect 60286 73336 60288 73388
rect 60232 73334 60288 73336
rect 60232 72050 60288 72052
rect 60232 71998 60234 72050
rect 60234 71998 60286 72050
rect 60286 71998 60288 72050
rect 60232 71996 60288 71998
rect 60232 70560 60288 70562
rect 60232 70508 60234 70560
rect 60234 70508 60286 70560
rect 60286 70508 60288 70560
rect 60232 70506 60288 70508
rect 60232 69222 60288 69224
rect 60232 69170 60234 69222
rect 60234 69170 60286 69222
rect 60286 69170 60288 69222
rect 60232 69168 60288 69170
rect 59777 68777 59833 68833
rect 59641 68653 59697 68709
rect 59505 68529 59561 68585
rect 59369 68405 59425 68461
rect 59233 68281 59289 68337
rect 59097 68033 59153 68089
rect 58961 67909 59017 67965
rect 58961 67678 59017 67734
rect 60232 67732 60288 67734
rect 60232 67680 60234 67732
rect 60234 67680 60286 67732
rect 60286 67680 60288 67732
rect 60232 67678 60288 67680
rect 55387 66222 55443 66278
rect 11649 12120 11705 12176
rect 6838 10718 6894 10720
rect 6838 10666 6840 10718
rect 6840 10666 6892 10718
rect 6892 10666 6894 10718
rect 6838 10664 6894 10666
rect 7117 10664 7173 10720
rect 7117 10433 7173 10489
rect 7933 10309 7989 10365
rect 7797 10185 7853 10241
rect 7661 10061 7717 10117
rect 7525 9937 7581 9993
rect 7389 9813 7445 9869
rect 7253 9689 7309 9745
rect 7117 9565 7173 9621
rect 6838 9228 6894 9230
rect 6838 9176 6840 9228
rect 6840 9176 6892 9228
rect 6892 9176 6894 9228
rect 6838 9174 6894 9176
rect 6838 7890 6894 7892
rect 6838 7838 6840 7890
rect 6840 7838 6892 7890
rect 6892 7838 6894 7890
rect 6838 7836 6894 7838
rect 6838 6400 6894 6402
rect 6838 6348 6840 6400
rect 6840 6348 6892 6400
rect 6892 6348 6894 6400
rect 6838 6346 6894 6348
rect 6838 5062 6894 5064
rect 6838 5010 6840 5062
rect 6840 5010 6892 5062
rect 6892 5010 6894 5062
rect 6838 5008 6894 5010
rect 6838 3572 6894 3574
rect 6838 3520 6840 3572
rect 6840 3520 6892 3572
rect 6892 3520 6894 3572
rect 6838 3518 6894 3520
rect 6838 2234 6894 2236
rect 6838 2182 6840 2234
rect 6840 2182 6892 2234
rect 6892 2182 6894 2234
rect 6838 2180 6894 2182
rect 7933 9174 7989 9230
rect 7797 7836 7853 7892
rect 7661 6346 7717 6402
rect 7525 5008 7581 5064
rect 7389 3518 7445 3574
rect 7253 2180 7309 2236
rect 6838 744 6894 746
rect 6838 692 6840 744
rect 6840 692 6892 744
rect 6892 692 6894 744
rect 6838 690 6894 692
rect 7117 690 7173 746
rect 11773 8849 11829 8905
rect 13549 12025 13605 12027
rect 13549 11973 13551 12025
rect 13551 11973 13603 12025
rect 13603 11973 13605 12025
rect 13549 11971 13605 11973
rect 11897 3538 11953 3594
<< metal3 >>
rect 60992 78300 61090 78398
rect 62352 78300 62450 78398
rect 59772 77710 59838 77713
rect 60227 77710 60293 77713
rect 59772 77708 60293 77710
rect 59772 77652 59777 77708
rect 59833 77652 60232 77708
rect 60288 77652 60293 77708
rect 59772 77650 60293 77652
rect 59772 77647 59838 77650
rect 60227 77647 60293 77650
rect 60992 76886 61090 76984
rect 62352 76886 62450 76984
rect 59636 76220 59702 76223
rect 60227 76220 60293 76223
rect 59636 76218 60293 76220
rect 59636 76162 59641 76218
rect 59697 76162 60232 76218
rect 60288 76162 60293 76218
rect 59636 76160 60293 76162
rect 59636 76157 59702 76160
rect 60227 76157 60293 76160
rect 60992 75472 61090 75570
rect 62352 75472 62450 75570
rect 59500 74882 59566 74885
rect 60227 74882 60293 74885
rect 59500 74880 60293 74882
rect 59500 74824 59505 74880
rect 59561 74824 60232 74880
rect 60288 74824 60293 74880
rect 59500 74822 60293 74824
rect 59500 74819 59566 74822
rect 60227 74819 60293 74822
rect 60992 74058 61090 74156
rect 62352 74058 62450 74156
rect 59364 73392 59430 73395
rect 60227 73392 60293 73395
rect 59364 73390 60293 73392
rect 59364 73334 59369 73390
rect 59425 73334 60232 73390
rect 60288 73334 60293 73390
rect 59364 73332 60293 73334
rect 59364 73329 59430 73332
rect 60227 73329 60293 73332
rect 60992 72644 61090 72742
rect 62352 72644 62450 72742
rect 59228 72054 59294 72057
rect 60227 72054 60293 72057
rect 59228 72052 60293 72054
rect 59228 71996 59233 72052
rect 59289 71996 60232 72052
rect 60288 71996 60293 72052
rect 59228 71994 60293 71996
rect 59228 71991 59294 71994
rect 60227 71991 60293 71994
rect 13989 71558 14087 71656
rect 18981 71558 19079 71656
rect 23973 71558 24071 71656
rect 28965 71558 29063 71656
rect 33957 71558 34055 71656
rect 38949 71558 39047 71656
rect 43941 71558 44039 71656
rect 48933 71558 49031 71656
rect 13989 71236 14087 71334
rect 18981 71236 19079 71334
rect 23973 71236 24071 71334
rect 28965 71236 29063 71334
rect 33957 71236 34055 71334
rect 38949 71236 39047 71334
rect 43941 71236 44039 71334
rect 48933 71236 49031 71334
rect 60992 71230 61090 71328
rect 62352 71230 62450 71328
rect 58956 70564 59022 70567
rect 60227 70564 60293 70567
rect 58956 70562 60293 70564
rect 58956 70506 58961 70562
rect 59017 70506 60232 70562
rect 60288 70506 60293 70562
rect 58956 70504 60293 70506
rect 58956 70501 59022 70504
rect 60227 70501 60293 70504
rect 13977 70398 14075 70496
rect 18969 70398 19067 70496
rect 23961 70398 24059 70496
rect 28953 70398 29051 70496
rect 33945 70398 34043 70496
rect 38937 70398 39035 70496
rect 43929 70398 44027 70496
rect 48921 70398 49019 70496
rect 60992 69816 61090 69914
rect 62352 69816 62450 69914
rect 14059 69624 14157 69722
rect 19051 69624 19149 69722
rect 24043 69624 24141 69722
rect 29035 69624 29133 69722
rect 34027 69624 34125 69722
rect 39019 69624 39117 69722
rect 44011 69624 44109 69722
rect 49003 69624 49101 69722
rect 55258 69551 55324 69554
rect 30692 69549 55324 69551
rect 30692 69493 55263 69549
rect 55319 69493 55324 69549
rect 30692 69491 55324 69493
rect 55258 69488 55324 69491
rect 59092 69226 59158 69229
rect 60227 69226 60293 69229
rect 59092 69224 60293 69226
rect 59092 69168 59097 69224
rect 59153 69168 60232 69224
rect 60288 69168 60293 69224
rect 59092 69166 60293 69168
rect 59092 69163 59158 69166
rect 60227 69163 60293 69166
rect 59772 68835 59838 68838
rect 53563 68833 59838 68835
rect 53563 68777 59777 68833
rect 59833 68777 59838 68833
rect 53563 68775 59838 68777
rect 59772 68772 59838 68775
rect 59636 68711 59702 68714
rect 53563 68709 59702 68711
rect 53563 68653 59641 68709
rect 59697 68653 59702 68709
rect 53563 68651 59702 68653
rect 59636 68648 59702 68651
rect 59500 68587 59566 68590
rect 53563 68585 59566 68587
rect 53563 68529 59505 68585
rect 59561 68529 59566 68585
rect 53563 68527 59566 68529
rect 59500 68524 59566 68527
rect 59364 68463 59430 68466
rect 53563 68461 59430 68463
rect 53563 68405 59369 68461
rect 59425 68405 59430 68461
rect 53563 68403 59430 68405
rect 59364 68400 59430 68403
rect 60992 68402 61090 68500
rect 62352 68402 62450 68500
rect 59228 68339 59294 68342
rect 53563 68337 59294 68339
rect 53563 68281 59233 68337
rect 59289 68281 59294 68337
rect 53563 68279 59294 68281
rect 59228 68276 59294 68279
rect 58956 68215 59022 68218
rect 53563 68213 59022 68215
rect 53563 68157 58961 68213
rect 59017 68157 59022 68213
rect 53563 68155 59022 68157
rect 58956 68152 59022 68155
rect 59092 68091 59158 68094
rect 53563 68089 59158 68091
rect 53563 68033 59097 68089
rect 59153 68033 59158 68089
rect 53563 68031 59158 68033
rect 59092 68028 59158 68031
rect 58956 67967 59022 67970
rect 53563 67965 59022 67967
rect 53563 67909 58961 67965
rect 59017 67909 59022 67965
rect 53563 67907 59022 67909
rect 58956 67904 59022 67907
rect 58956 67736 59022 67739
rect 60227 67736 60293 67739
rect 58956 67734 60293 67736
rect 58956 67678 58961 67734
rect 59017 67678 60232 67734
rect 60288 67678 60293 67734
rect 58956 67676 60293 67678
rect 58956 67673 59022 67676
rect 60227 67673 60293 67676
rect 14232 67131 14330 67229
rect 15480 67131 15578 67229
rect 16728 67131 16826 67229
rect 17976 67131 18074 67229
rect 19224 67131 19322 67229
rect 20472 67131 20570 67229
rect 21720 67131 21818 67229
rect 22968 67131 23066 67229
rect 24216 67131 24314 67229
rect 25464 67131 25562 67229
rect 26712 67131 26810 67229
rect 27960 67131 28058 67229
rect 29208 67131 29306 67229
rect 30456 67131 30554 67229
rect 31704 67131 31802 67229
rect 32952 67131 33050 67229
rect 34200 67131 34298 67229
rect 35448 67131 35546 67229
rect 36696 67131 36794 67229
rect 37944 67131 38042 67229
rect 39192 67131 39290 67229
rect 40440 67131 40538 67229
rect 41688 67131 41786 67229
rect 42936 67131 43034 67229
rect 44184 67131 44282 67229
rect 45432 67131 45530 67229
rect 46680 67131 46778 67229
rect 47928 67131 48026 67229
rect 49176 67131 49274 67229
rect 50424 67131 50522 67229
rect 51672 67131 51770 67229
rect 52920 67131 53018 67229
rect 60992 66988 61090 67086
rect 62352 66988 62450 67086
rect 53640 66429 53706 66432
rect 53640 66427 67334 66429
rect 53640 66371 53645 66427
rect 53701 66371 67334 66427
rect 53640 66369 67334 66371
rect 53640 66366 53706 66369
rect 55382 66280 55448 66283
rect 33250 66278 55448 66280
rect 33250 66222 55387 66278
rect 55443 66222 55448 66278
rect 33250 66220 55448 66222
rect 55382 66217 55448 66220
rect 13801 65582 13899 65680
rect 14663 65582 14761 65680
rect 15049 65582 15147 65680
rect 15911 65582 16009 65680
rect 16297 65582 16395 65680
rect 17159 65582 17257 65680
rect 17545 65582 17643 65680
rect 18407 65582 18505 65680
rect 18793 65582 18891 65680
rect 19655 65582 19753 65680
rect 20041 65582 20139 65680
rect 20903 65582 21001 65680
rect 21289 65582 21387 65680
rect 22151 65582 22249 65680
rect 22537 65582 22635 65680
rect 23399 65582 23497 65680
rect 23785 65582 23883 65680
rect 24647 65582 24745 65680
rect 25033 65582 25131 65680
rect 25895 65582 25993 65680
rect 26281 65582 26379 65680
rect 27143 65582 27241 65680
rect 27529 65582 27627 65680
rect 28391 65582 28489 65680
rect 28777 65582 28875 65680
rect 29639 65582 29737 65680
rect 30025 65582 30123 65680
rect 30887 65582 30985 65680
rect 31273 65582 31371 65680
rect 32135 65582 32233 65680
rect 32521 65582 32619 65680
rect 33383 65582 33481 65680
rect 33769 65582 33867 65680
rect 34631 65582 34729 65680
rect 35017 65582 35115 65680
rect 35879 65582 35977 65680
rect 36265 65582 36363 65680
rect 37127 65582 37225 65680
rect 37513 65582 37611 65680
rect 38375 65582 38473 65680
rect 38761 65582 38859 65680
rect 39623 65582 39721 65680
rect 40009 65582 40107 65680
rect 40871 65582 40969 65680
rect 41257 65582 41355 65680
rect 42119 65582 42217 65680
rect 42505 65582 42603 65680
rect 43367 65582 43465 65680
rect 43753 65582 43851 65680
rect 44615 65582 44713 65680
rect 45001 65582 45099 65680
rect 45863 65582 45961 65680
rect 46249 65582 46347 65680
rect 47111 65582 47209 65680
rect 47497 65582 47595 65680
rect 48359 65582 48457 65680
rect 48745 65582 48843 65680
rect 49607 65582 49705 65680
rect 49993 65582 50091 65680
rect 50855 65582 50953 65680
rect 51241 65582 51339 65680
rect 52103 65582 52201 65680
rect 52489 65582 52587 65680
rect 53351 65582 53449 65680
rect 53737 65582 53835 65680
rect 13296 64991 13394 65089
rect 13920 64991 14018 65089
rect 14544 64991 14642 65089
rect 15168 64991 15266 65089
rect 15792 64991 15890 65089
rect 16416 64991 16514 65089
rect 17040 64991 17138 65089
rect 17664 64991 17762 65089
rect 18288 64991 18386 65089
rect 18912 64991 19010 65089
rect 19536 64991 19634 65089
rect 20160 64991 20258 65089
rect 20784 64991 20882 65089
rect 21408 64991 21506 65089
rect 22032 64991 22130 65089
rect 22656 64991 22754 65089
rect 23280 64991 23378 65089
rect 23904 64991 24002 65089
rect 24528 64991 24626 65089
rect 25152 64991 25250 65089
rect 25776 64991 25874 65089
rect 26400 64991 26498 65089
rect 27024 64991 27122 65089
rect 27648 64991 27746 65089
rect 28272 64991 28370 65089
rect 28896 64991 28994 65089
rect 29520 64991 29618 65089
rect 30144 64991 30242 65089
rect 30768 64991 30866 65089
rect 31392 64991 31490 65089
rect 32016 64991 32114 65089
rect 32640 64991 32738 65089
rect 33264 64991 33362 65089
rect 33888 64991 33986 65089
rect 34512 64991 34610 65089
rect 35136 64991 35234 65089
rect 35760 64991 35858 65089
rect 36384 64991 36482 65089
rect 37008 64991 37106 65089
rect 37632 64991 37730 65089
rect 38256 64991 38354 65089
rect 38880 64991 38978 65089
rect 39504 64991 39602 65089
rect 40128 64991 40226 65089
rect 40752 64991 40850 65089
rect 41376 64991 41474 65089
rect 42000 64991 42098 65089
rect 42624 64991 42722 65089
rect 43248 64991 43346 65089
rect 43872 64991 43970 65089
rect 44496 64991 44594 65089
rect 45120 64991 45218 65089
rect 45744 64991 45842 65089
rect 46368 64991 46466 65089
rect 46992 64991 47090 65089
rect 47616 64991 47714 65089
rect 48240 64991 48338 65089
rect 48864 64991 48962 65089
rect 49488 64991 49586 65089
rect 50112 64991 50210 65089
rect 50736 64991 50834 65089
rect 51360 64991 51458 65089
rect 51984 64991 52082 65089
rect 52608 64991 52706 65089
rect 53232 64991 53330 65089
rect 53856 64991 53954 65089
rect 12234 64777 12332 64875
rect 54918 64777 55016 64875
rect 55944 64627 56042 64725
rect 58635 64615 58733 64713
rect 59467 64621 59565 64719
rect 12600 64430 12698 64528
rect 54552 64430 54650 64528
rect 12600 64193 12698 64291
rect 54552 64193 54650 64291
rect 6025 64058 6123 64156
rect 6450 64058 6548 64156
rect 6882 64058 6980 64156
rect 7264 64035 7362 64133
rect 7660 64035 7758 64133
rect 59492 64035 59590 64133
rect 59888 64035 59986 64133
rect 60270 64058 60368 64156
rect 60702 64058 60800 64156
rect 61127 64058 61225 64156
rect 12600 63877 12698 63975
rect 54552 63877 54650 63975
rect 6025 63684 6123 63782
rect 6450 63626 6548 63724
rect 6882 63626 6980 63724
rect 7264 63640 7362 63738
rect 7660 63640 7758 63738
rect 12600 63640 12698 63738
rect 54552 63640 54650 63738
rect 59492 63640 59590 63738
rect 59888 63640 59986 63738
rect 60270 63626 60368 63724
rect 60702 63626 60800 63724
rect 61127 63684 61225 63782
rect 12600 63403 12698 63501
rect 54552 63403 54650 63501
rect 6025 63268 6123 63366
rect 6450 63268 6548 63366
rect 6882 63268 6980 63366
rect 7264 63245 7362 63343
rect 7660 63245 7758 63343
rect 59492 63245 59590 63343
rect 59888 63245 59986 63343
rect 60270 63268 60368 63366
rect 60702 63268 60800 63366
rect 61127 63268 61225 63366
rect 12600 63087 12698 63185
rect 54552 63087 54650 63185
rect 6025 62894 6123 62992
rect 6450 62836 6548 62934
rect 6882 62836 6980 62934
rect 7264 62850 7362 62948
rect 7660 62850 7758 62948
rect 12600 62850 12698 62948
rect 54552 62850 54650 62948
rect 59492 62850 59590 62948
rect 59888 62850 59986 62948
rect 60270 62836 60368 62934
rect 60702 62836 60800 62934
rect 61127 62894 61225 62992
rect 12600 62613 12698 62711
rect 54552 62613 54650 62711
rect 6025 62478 6123 62576
rect 6450 62478 6548 62576
rect 6882 62478 6980 62576
rect 7264 62455 7362 62553
rect 7660 62455 7758 62553
rect 59492 62455 59590 62553
rect 59888 62455 59986 62553
rect 60270 62478 60368 62576
rect 60702 62478 60800 62576
rect 61127 62478 61225 62576
rect 12600 62297 12698 62395
rect 54552 62297 54650 62395
rect 6025 62104 6123 62202
rect 6450 62046 6548 62144
rect 6882 62046 6980 62144
rect 7264 62060 7362 62158
rect 7660 62060 7758 62158
rect 12600 62060 12698 62158
rect 54552 62060 54650 62158
rect 59492 62060 59590 62158
rect 59888 62060 59986 62158
rect 60270 62046 60368 62144
rect 60702 62046 60800 62144
rect 61127 62104 61225 62202
rect 12600 61823 12698 61921
rect 54552 61823 54650 61921
rect 6025 61688 6123 61786
rect 6450 61688 6548 61786
rect 6882 61688 6980 61786
rect 7264 61665 7362 61763
rect 7660 61665 7758 61763
rect 59492 61665 59590 61763
rect 59888 61665 59986 61763
rect 60270 61688 60368 61786
rect 60702 61688 60800 61786
rect 61127 61688 61225 61786
rect 12600 61507 12698 61605
rect 54552 61507 54650 61605
rect 6025 61314 6123 61412
rect 6450 61256 6548 61354
rect 6882 61256 6980 61354
rect 7264 61270 7362 61368
rect 7660 61270 7758 61368
rect 12600 61270 12698 61368
rect 54552 61270 54650 61368
rect 59492 61270 59590 61368
rect 59888 61270 59986 61368
rect 60270 61256 60368 61354
rect 60702 61256 60800 61354
rect 61127 61314 61225 61412
rect 12600 61033 12698 61131
rect 54552 61033 54650 61131
rect 6025 60898 6123 60996
rect 6450 60898 6548 60996
rect 6882 60898 6980 60996
rect 7264 60875 7362 60973
rect 7660 60875 7758 60973
rect 59492 60875 59590 60973
rect 59888 60875 59986 60973
rect 60270 60898 60368 60996
rect 60702 60898 60800 60996
rect 61127 60898 61225 60996
rect 12600 60717 12698 60815
rect 54552 60717 54650 60815
rect 6025 60524 6123 60622
rect 6450 60466 6548 60564
rect 6882 60466 6980 60564
rect 7264 60480 7362 60578
rect 7660 60480 7758 60578
rect 12600 60480 12698 60578
rect 54552 60480 54650 60578
rect 59492 60480 59590 60578
rect 59888 60480 59986 60578
rect 60270 60466 60368 60564
rect 60702 60466 60800 60564
rect 61127 60524 61225 60622
rect 12600 60243 12698 60341
rect 54552 60243 54650 60341
rect 6025 60108 6123 60206
rect 6450 60108 6548 60206
rect 6882 60108 6980 60206
rect 7264 60085 7362 60183
rect 7660 60085 7758 60183
rect 59492 60085 59590 60183
rect 59888 60085 59986 60183
rect 60270 60108 60368 60206
rect 60702 60108 60800 60206
rect 61127 60108 61225 60206
rect 12600 59927 12698 60025
rect 54552 59927 54650 60025
rect 6025 59734 6123 59832
rect 6450 59676 6548 59774
rect 6882 59676 6980 59774
rect 7264 59690 7362 59788
rect 7660 59690 7758 59788
rect 12600 59690 12698 59788
rect 54552 59690 54650 59788
rect 59492 59690 59590 59788
rect 59888 59690 59986 59788
rect 60270 59676 60368 59774
rect 60702 59676 60800 59774
rect 61127 59734 61225 59832
rect 12600 59453 12698 59551
rect 54552 59453 54650 59551
rect 6025 59318 6123 59416
rect 6450 59318 6548 59416
rect 6882 59318 6980 59416
rect 7264 59295 7362 59393
rect 7660 59295 7758 59393
rect 59492 59295 59590 59393
rect 59888 59295 59986 59393
rect 60270 59318 60368 59416
rect 60702 59318 60800 59416
rect 61127 59318 61225 59416
rect 12600 59137 12698 59235
rect 54552 59137 54650 59235
rect 6025 58944 6123 59042
rect 6450 58886 6548 58984
rect 6882 58886 6980 58984
rect 7264 58900 7362 58998
rect 7660 58900 7758 58998
rect 12600 58900 12698 58998
rect 54552 58900 54650 58998
rect 59492 58900 59590 58998
rect 59888 58900 59986 58998
rect 60270 58886 60368 58984
rect 60702 58886 60800 58984
rect 61127 58944 61225 59042
rect 12600 58663 12698 58761
rect 54552 58663 54650 58761
rect 6025 58528 6123 58626
rect 6450 58528 6548 58626
rect 6882 58528 6980 58626
rect 7264 58505 7362 58603
rect 7660 58505 7758 58603
rect 59492 58505 59590 58603
rect 59888 58505 59986 58603
rect 60270 58528 60368 58626
rect 60702 58528 60800 58626
rect 61127 58528 61225 58626
rect 12600 58347 12698 58445
rect 54552 58347 54650 58445
rect 6025 58154 6123 58252
rect 6450 58096 6548 58194
rect 6882 58096 6980 58194
rect 7264 58110 7362 58208
rect 7660 58110 7758 58208
rect 12600 58110 12698 58208
rect 54552 58110 54650 58208
rect 59492 58110 59590 58208
rect 59888 58110 59986 58208
rect 60270 58096 60368 58194
rect 60702 58096 60800 58194
rect 61127 58154 61225 58252
rect 12600 57873 12698 57971
rect 54552 57873 54650 57971
rect 6025 57738 6123 57836
rect 6450 57738 6548 57836
rect 6882 57738 6980 57836
rect 7264 57715 7362 57813
rect 7660 57715 7758 57813
rect 59492 57715 59590 57813
rect 59888 57715 59986 57813
rect 60270 57738 60368 57836
rect 60702 57738 60800 57836
rect 61127 57738 61225 57836
rect 12600 57557 12698 57655
rect 54552 57557 54650 57655
rect 6025 57364 6123 57462
rect 6450 57306 6548 57404
rect 6882 57306 6980 57404
rect 7264 57320 7362 57418
rect 7660 57320 7758 57418
rect 12600 57320 12698 57418
rect 54552 57320 54650 57418
rect 59492 57320 59590 57418
rect 59888 57320 59986 57418
rect 60270 57306 60368 57404
rect 60702 57306 60800 57404
rect 61127 57364 61225 57462
rect 12600 57083 12698 57181
rect 54552 57083 54650 57181
rect 6025 56948 6123 57046
rect 6450 56948 6548 57046
rect 6882 56948 6980 57046
rect 7264 56925 7362 57023
rect 7660 56925 7758 57023
rect 59492 56925 59590 57023
rect 59888 56925 59986 57023
rect 60270 56948 60368 57046
rect 60702 56948 60800 57046
rect 61127 56948 61225 57046
rect 12600 56767 12698 56865
rect 54552 56767 54650 56865
rect 6025 56574 6123 56672
rect 6450 56516 6548 56614
rect 6882 56516 6980 56614
rect 7264 56530 7362 56628
rect 7660 56530 7758 56628
rect 12600 56530 12698 56628
rect 54552 56530 54650 56628
rect 59492 56530 59590 56628
rect 59888 56530 59986 56628
rect 60270 56516 60368 56614
rect 60702 56516 60800 56614
rect 61127 56574 61225 56672
rect 12600 56293 12698 56391
rect 54552 56293 54650 56391
rect 6025 56158 6123 56256
rect 6450 56158 6548 56256
rect 6882 56158 6980 56256
rect 7264 56135 7362 56233
rect 7660 56135 7758 56233
rect 59492 56135 59590 56233
rect 59888 56135 59986 56233
rect 60270 56158 60368 56256
rect 60702 56158 60800 56256
rect 61127 56158 61225 56256
rect 12600 55977 12698 56075
rect 54552 55977 54650 56075
rect 6025 55784 6123 55882
rect 6450 55726 6548 55824
rect 6882 55726 6980 55824
rect 7264 55740 7362 55838
rect 7660 55740 7758 55838
rect 12600 55740 12698 55838
rect 54552 55740 54650 55838
rect 59492 55740 59590 55838
rect 59888 55740 59986 55838
rect 60270 55726 60368 55824
rect 60702 55726 60800 55824
rect 61127 55784 61225 55882
rect 12600 55503 12698 55601
rect 54552 55503 54650 55601
rect 6025 55368 6123 55466
rect 6450 55368 6548 55466
rect 6882 55368 6980 55466
rect 7264 55345 7362 55443
rect 7660 55345 7758 55443
rect 59492 55345 59590 55443
rect 59888 55345 59986 55443
rect 60270 55368 60368 55466
rect 60702 55368 60800 55466
rect 61127 55368 61225 55466
rect 12600 55187 12698 55285
rect 54552 55187 54650 55285
rect 6025 54994 6123 55092
rect 6450 54936 6548 55034
rect 6882 54936 6980 55034
rect 7264 54950 7362 55048
rect 7660 54950 7758 55048
rect 12600 54950 12698 55048
rect 54552 54950 54650 55048
rect 59492 54950 59590 55048
rect 59888 54950 59986 55048
rect 60270 54936 60368 55034
rect 60702 54936 60800 55034
rect 61127 54994 61225 55092
rect 12600 54713 12698 54811
rect 54552 54713 54650 54811
rect 6025 54578 6123 54676
rect 6450 54578 6548 54676
rect 6882 54578 6980 54676
rect 7264 54555 7362 54653
rect 7660 54555 7758 54653
rect 59492 54555 59590 54653
rect 59888 54555 59986 54653
rect 60270 54578 60368 54676
rect 60702 54578 60800 54676
rect 61127 54578 61225 54676
rect 12600 54397 12698 54495
rect 54552 54397 54650 54495
rect 6025 54204 6123 54302
rect 6450 54146 6548 54244
rect 6882 54146 6980 54244
rect 7264 54160 7362 54258
rect 7660 54160 7758 54258
rect 12600 54160 12698 54258
rect 54552 54160 54650 54258
rect 59492 54160 59590 54258
rect 59888 54160 59986 54258
rect 60270 54146 60368 54244
rect 60702 54146 60800 54244
rect 61127 54204 61225 54302
rect 12600 53923 12698 54021
rect 54552 53923 54650 54021
rect 6025 53788 6123 53886
rect 6450 53788 6548 53886
rect 6882 53788 6980 53886
rect 7264 53765 7362 53863
rect 7660 53765 7758 53863
rect 59492 53765 59590 53863
rect 59888 53765 59986 53863
rect 60270 53788 60368 53886
rect 60702 53788 60800 53886
rect 61127 53788 61225 53886
rect 12600 53607 12698 53705
rect 54552 53607 54650 53705
rect 6025 53414 6123 53512
rect 6450 53356 6548 53454
rect 6882 53356 6980 53454
rect 7264 53370 7362 53468
rect 7660 53370 7758 53468
rect 12600 53370 12698 53468
rect 54552 53370 54650 53468
rect 59492 53370 59590 53468
rect 59888 53370 59986 53468
rect 60270 53356 60368 53454
rect 60702 53356 60800 53454
rect 61127 53414 61225 53512
rect 12600 53133 12698 53231
rect 54552 53133 54650 53231
rect 6025 52998 6123 53096
rect 6450 52998 6548 53096
rect 6882 52998 6980 53096
rect 7264 52975 7362 53073
rect 7660 52975 7758 53073
rect 59492 52975 59590 53073
rect 59888 52975 59986 53073
rect 60270 52998 60368 53096
rect 60702 52998 60800 53096
rect 61127 52998 61225 53096
rect 12600 52817 12698 52915
rect 54552 52817 54650 52915
rect 6025 52624 6123 52722
rect 6450 52566 6548 52664
rect 6882 52566 6980 52664
rect 7264 52580 7362 52678
rect 7660 52580 7758 52678
rect 12600 52580 12698 52678
rect 54552 52580 54650 52678
rect 59492 52580 59590 52678
rect 59888 52580 59986 52678
rect 60270 52566 60368 52664
rect 60702 52566 60800 52664
rect 61127 52624 61225 52722
rect 12600 52343 12698 52441
rect 54552 52343 54650 52441
rect 6025 52208 6123 52306
rect 6450 52208 6548 52306
rect 6882 52208 6980 52306
rect 7264 52185 7362 52283
rect 7660 52185 7758 52283
rect 59492 52185 59590 52283
rect 59888 52185 59986 52283
rect 60270 52208 60368 52306
rect 60702 52208 60800 52306
rect 61127 52208 61225 52306
rect 12600 52027 12698 52125
rect 54552 52027 54650 52125
rect 6025 51834 6123 51932
rect 6450 51776 6548 51874
rect 6882 51776 6980 51874
rect 7264 51790 7362 51888
rect 7660 51790 7758 51888
rect 12600 51790 12698 51888
rect 54552 51790 54650 51888
rect 59492 51790 59590 51888
rect 59888 51790 59986 51888
rect 60270 51776 60368 51874
rect 60702 51776 60800 51874
rect 61127 51834 61225 51932
rect 12600 51553 12698 51651
rect 54552 51553 54650 51651
rect 6025 51418 6123 51516
rect 6450 51418 6548 51516
rect 6882 51418 6980 51516
rect 7264 51395 7362 51493
rect 7660 51395 7758 51493
rect 59492 51395 59590 51493
rect 59888 51395 59986 51493
rect 60270 51418 60368 51516
rect 60702 51418 60800 51516
rect 61127 51418 61225 51516
rect 12600 51237 12698 51335
rect 54552 51237 54650 51335
rect 6025 51044 6123 51142
rect 6450 50986 6548 51084
rect 6882 50986 6980 51084
rect 7264 51000 7362 51098
rect 7660 51000 7758 51098
rect 12600 51000 12698 51098
rect 54552 51000 54650 51098
rect 59492 51000 59590 51098
rect 59888 51000 59986 51098
rect 60270 50986 60368 51084
rect 60702 50986 60800 51084
rect 61127 51044 61225 51142
rect 12600 50763 12698 50861
rect 54552 50763 54650 50861
rect 6025 50628 6123 50726
rect 6450 50628 6548 50726
rect 6882 50628 6980 50726
rect 7264 50605 7362 50703
rect 7660 50605 7758 50703
rect 59492 50605 59590 50703
rect 59888 50605 59986 50703
rect 60270 50628 60368 50726
rect 60702 50628 60800 50726
rect 61127 50628 61225 50726
rect 12600 50447 12698 50545
rect 54552 50447 54650 50545
rect 6025 50254 6123 50352
rect 6450 50196 6548 50294
rect 6882 50196 6980 50294
rect 7264 50210 7362 50308
rect 7660 50210 7758 50308
rect 12600 50210 12698 50308
rect 54552 50210 54650 50308
rect 59492 50210 59590 50308
rect 59888 50210 59986 50308
rect 60270 50196 60368 50294
rect 60702 50196 60800 50294
rect 61127 50254 61225 50352
rect 12600 49973 12698 50071
rect 54552 49973 54650 50071
rect 6025 49838 6123 49936
rect 6450 49838 6548 49936
rect 6882 49838 6980 49936
rect 7264 49815 7362 49913
rect 7660 49815 7758 49913
rect 59492 49815 59590 49913
rect 59888 49815 59986 49913
rect 60270 49838 60368 49936
rect 60702 49838 60800 49936
rect 61127 49838 61225 49936
rect 12600 49657 12698 49755
rect 54552 49657 54650 49755
rect 6025 49464 6123 49562
rect 6450 49406 6548 49504
rect 6882 49406 6980 49504
rect 7264 49420 7362 49518
rect 7660 49420 7758 49518
rect 12600 49420 12698 49518
rect 54552 49420 54650 49518
rect 59492 49420 59590 49518
rect 59888 49420 59986 49518
rect 60270 49406 60368 49504
rect 60702 49406 60800 49504
rect 61127 49464 61225 49562
rect 12600 49183 12698 49281
rect 54552 49183 54650 49281
rect 6025 49048 6123 49146
rect 6450 49048 6548 49146
rect 6882 49048 6980 49146
rect 7264 49025 7362 49123
rect 7660 49025 7758 49123
rect 59492 49025 59590 49123
rect 59888 49025 59986 49123
rect 60270 49048 60368 49146
rect 60702 49048 60800 49146
rect 61127 49048 61225 49146
rect 12600 48867 12698 48965
rect 54552 48867 54650 48965
rect 6025 48674 6123 48772
rect 6450 48616 6548 48714
rect 6882 48616 6980 48714
rect 7264 48630 7362 48728
rect 7660 48630 7758 48728
rect 12600 48630 12698 48728
rect 54552 48630 54650 48728
rect 59492 48630 59590 48728
rect 59888 48630 59986 48728
rect 60270 48616 60368 48714
rect 60702 48616 60800 48714
rect 61127 48674 61225 48772
rect 12600 48393 12698 48491
rect 54552 48393 54650 48491
rect 6025 48258 6123 48356
rect 6450 48258 6548 48356
rect 6882 48258 6980 48356
rect 7264 48235 7362 48333
rect 7660 48235 7758 48333
rect 59492 48235 59590 48333
rect 59888 48235 59986 48333
rect 60270 48258 60368 48356
rect 60702 48258 60800 48356
rect 61127 48258 61225 48356
rect 12600 48077 12698 48175
rect 54552 48077 54650 48175
rect 6025 47884 6123 47982
rect 6450 47826 6548 47924
rect 6882 47826 6980 47924
rect 7264 47840 7362 47938
rect 7660 47840 7758 47938
rect 12600 47840 12698 47938
rect 54552 47840 54650 47938
rect 59492 47840 59590 47938
rect 59888 47840 59986 47938
rect 60270 47826 60368 47924
rect 60702 47826 60800 47924
rect 61127 47884 61225 47982
rect 12600 47603 12698 47701
rect 54552 47603 54650 47701
rect 6025 47468 6123 47566
rect 6450 47468 6548 47566
rect 6882 47468 6980 47566
rect 7264 47445 7362 47543
rect 7660 47445 7758 47543
rect 59492 47445 59590 47543
rect 59888 47445 59986 47543
rect 60270 47468 60368 47566
rect 60702 47468 60800 47566
rect 61127 47468 61225 47566
rect 12600 47287 12698 47385
rect 54552 47287 54650 47385
rect 6025 47094 6123 47192
rect 6450 47036 6548 47134
rect 6882 47036 6980 47134
rect 7264 47050 7362 47148
rect 7660 47050 7758 47148
rect 12600 47050 12698 47148
rect 54552 47050 54650 47148
rect 59492 47050 59590 47148
rect 59888 47050 59986 47148
rect 60270 47036 60368 47134
rect 60702 47036 60800 47134
rect 61127 47094 61225 47192
rect 12600 46813 12698 46911
rect 54552 46813 54650 46911
rect 6025 46678 6123 46776
rect 6450 46678 6548 46776
rect 6882 46678 6980 46776
rect 7264 46655 7362 46753
rect 7660 46655 7758 46753
rect 59492 46655 59590 46753
rect 59888 46655 59986 46753
rect 60270 46678 60368 46776
rect 60702 46678 60800 46776
rect 61127 46678 61225 46776
rect 12600 46497 12698 46595
rect 54552 46497 54650 46595
rect 6025 46304 6123 46402
rect 6450 46246 6548 46344
rect 6882 46246 6980 46344
rect 7264 46260 7362 46358
rect 7660 46260 7758 46358
rect 12600 46260 12698 46358
rect 54552 46260 54650 46358
rect 59492 46260 59590 46358
rect 59888 46260 59986 46358
rect 60270 46246 60368 46344
rect 60702 46246 60800 46344
rect 61127 46304 61225 46402
rect 12600 46023 12698 46121
rect 54552 46023 54650 46121
rect 6025 45888 6123 45986
rect 6450 45888 6548 45986
rect 6882 45888 6980 45986
rect 7264 45865 7362 45963
rect 7660 45865 7758 45963
rect 59492 45865 59590 45963
rect 59888 45865 59986 45963
rect 60270 45888 60368 45986
rect 60702 45888 60800 45986
rect 61127 45888 61225 45986
rect 12600 45707 12698 45805
rect 54552 45707 54650 45805
rect 6025 45514 6123 45612
rect 6450 45456 6548 45554
rect 6882 45456 6980 45554
rect 7264 45470 7362 45568
rect 7660 45470 7758 45568
rect 12600 45470 12698 45568
rect 54552 45470 54650 45568
rect 59492 45470 59590 45568
rect 59888 45470 59986 45568
rect 60270 45456 60368 45554
rect 60702 45456 60800 45554
rect 61127 45514 61225 45612
rect 12600 45233 12698 45331
rect 54552 45233 54650 45331
rect 6025 45098 6123 45196
rect 6450 45098 6548 45196
rect 6882 45098 6980 45196
rect 7264 45075 7362 45173
rect 7660 45075 7758 45173
rect 59492 45075 59590 45173
rect 59888 45075 59986 45173
rect 60270 45098 60368 45196
rect 60702 45098 60800 45196
rect 61127 45098 61225 45196
rect 12600 44917 12698 45015
rect 54552 44917 54650 45015
rect 6025 44724 6123 44822
rect 6450 44666 6548 44764
rect 6882 44666 6980 44764
rect 7264 44680 7362 44778
rect 7660 44680 7758 44778
rect 12600 44680 12698 44778
rect 54552 44680 54650 44778
rect 59492 44680 59590 44778
rect 59888 44680 59986 44778
rect 60270 44666 60368 44764
rect 60702 44666 60800 44764
rect 61127 44724 61225 44822
rect 12600 44443 12698 44541
rect 54552 44443 54650 44541
rect 6025 44308 6123 44406
rect 6450 44308 6548 44406
rect 6882 44308 6980 44406
rect 7264 44285 7362 44383
rect 7660 44285 7758 44383
rect 59492 44285 59590 44383
rect 59888 44285 59986 44383
rect 60270 44308 60368 44406
rect 60702 44308 60800 44406
rect 61127 44308 61225 44406
rect 12600 44127 12698 44225
rect 54552 44127 54650 44225
rect 6025 43934 6123 44032
rect 6450 43876 6548 43974
rect 6882 43876 6980 43974
rect 7264 43890 7362 43988
rect 7660 43890 7758 43988
rect 12600 43890 12698 43988
rect 54552 43890 54650 43988
rect 59492 43890 59590 43988
rect 59888 43890 59986 43988
rect 60270 43876 60368 43974
rect 60702 43876 60800 43974
rect 61127 43934 61225 44032
rect 12600 43653 12698 43751
rect 54552 43653 54650 43751
rect 6025 43518 6123 43616
rect 6450 43518 6548 43616
rect 6882 43518 6980 43616
rect 7264 43495 7362 43593
rect 7660 43495 7758 43593
rect 59492 43495 59590 43593
rect 59888 43495 59986 43593
rect 60270 43518 60368 43616
rect 60702 43518 60800 43616
rect 61127 43518 61225 43616
rect 12600 43337 12698 43435
rect 54552 43337 54650 43435
rect 6025 43144 6123 43242
rect 6450 43086 6548 43184
rect 6882 43086 6980 43184
rect 7264 43100 7362 43198
rect 7660 43100 7758 43198
rect 12600 43100 12698 43198
rect 54552 43100 54650 43198
rect 59492 43100 59590 43198
rect 59888 43100 59986 43198
rect 60270 43086 60368 43184
rect 60702 43086 60800 43184
rect 61127 43144 61225 43242
rect 12600 42863 12698 42961
rect 54552 42863 54650 42961
rect 6025 42728 6123 42826
rect 6450 42728 6548 42826
rect 6882 42728 6980 42826
rect 7264 42705 7362 42803
rect 7660 42705 7758 42803
rect 59492 42705 59590 42803
rect 59888 42705 59986 42803
rect 60270 42728 60368 42826
rect 60702 42728 60800 42826
rect 61127 42728 61225 42826
rect 12600 42547 12698 42645
rect 54552 42547 54650 42645
rect 6025 42354 6123 42452
rect 6450 42296 6548 42394
rect 6882 42296 6980 42394
rect 7264 42310 7362 42408
rect 7660 42310 7758 42408
rect 12600 42310 12698 42408
rect 54552 42310 54650 42408
rect 59492 42310 59590 42408
rect 59888 42310 59986 42408
rect 60270 42296 60368 42394
rect 60702 42296 60800 42394
rect 61127 42354 61225 42452
rect 12600 42073 12698 42171
rect 54552 42073 54650 42171
rect 6025 41938 6123 42036
rect 6450 41938 6548 42036
rect 6882 41938 6980 42036
rect 7264 41915 7362 42013
rect 7660 41915 7758 42013
rect 59492 41915 59590 42013
rect 59888 41915 59986 42013
rect 60270 41938 60368 42036
rect 60702 41938 60800 42036
rect 61127 41938 61225 42036
rect 12600 41757 12698 41855
rect 54552 41757 54650 41855
rect 6025 41564 6123 41662
rect 6450 41506 6548 41604
rect 6882 41506 6980 41604
rect 7264 41520 7362 41618
rect 7660 41520 7758 41618
rect 12600 41520 12698 41618
rect 54552 41520 54650 41618
rect 59492 41520 59590 41618
rect 59888 41520 59986 41618
rect 60270 41506 60368 41604
rect 60702 41506 60800 41604
rect 61127 41564 61225 41662
rect 12600 41283 12698 41381
rect 54552 41283 54650 41381
rect 6025 41148 6123 41246
rect 6450 41148 6548 41246
rect 6882 41148 6980 41246
rect 7264 41125 7362 41223
rect 7660 41125 7758 41223
rect 59492 41125 59590 41223
rect 59888 41125 59986 41223
rect 60270 41148 60368 41246
rect 60702 41148 60800 41246
rect 61127 41148 61225 41246
rect 12600 40967 12698 41065
rect 54552 40967 54650 41065
rect 6025 40774 6123 40872
rect 6450 40716 6548 40814
rect 6882 40716 6980 40814
rect 7264 40730 7362 40828
rect 7660 40730 7758 40828
rect 12600 40730 12698 40828
rect 54552 40730 54650 40828
rect 59492 40730 59590 40828
rect 59888 40730 59986 40828
rect 60270 40716 60368 40814
rect 60702 40716 60800 40814
rect 61127 40774 61225 40872
rect 12600 40493 12698 40591
rect 54552 40493 54650 40591
rect 6025 40358 6123 40456
rect 6450 40358 6548 40456
rect 6882 40358 6980 40456
rect 7264 40335 7362 40433
rect 7660 40335 7758 40433
rect 59492 40335 59590 40433
rect 59888 40335 59986 40433
rect 60270 40358 60368 40456
rect 60702 40358 60800 40456
rect 61127 40358 61225 40456
rect 12600 40177 12698 40275
rect 54552 40177 54650 40275
rect 6025 39984 6123 40082
rect 6450 39926 6548 40024
rect 6882 39926 6980 40024
rect 7264 39940 7362 40038
rect 7660 39940 7758 40038
rect 12600 39940 12698 40038
rect 54552 39940 54650 40038
rect 59492 39940 59590 40038
rect 59888 39940 59986 40038
rect 60270 39926 60368 40024
rect 60702 39926 60800 40024
rect 61127 39984 61225 40082
rect 12600 39703 12698 39801
rect 54552 39703 54650 39801
rect 6025 39568 6123 39666
rect 6450 39568 6548 39666
rect 6882 39568 6980 39666
rect 7264 39545 7362 39643
rect 7660 39545 7758 39643
rect 59492 39545 59590 39643
rect 59888 39545 59986 39643
rect 60270 39568 60368 39666
rect 60702 39568 60800 39666
rect 61127 39568 61225 39666
rect 12600 39387 12698 39485
rect 54552 39387 54650 39485
rect 6025 39194 6123 39292
rect 6450 39136 6548 39234
rect 6882 39136 6980 39234
rect 7264 39150 7362 39248
rect 7660 39150 7758 39248
rect 8092 39135 8190 39233
rect 8517 39134 8615 39232
rect 9560 39150 9658 39248
rect 11208 39150 11306 39248
rect 12600 39150 12698 39248
rect 54552 39150 54650 39248
rect 55944 39150 56042 39248
rect 57592 39150 57690 39248
rect 58635 39134 58733 39232
rect 59060 39135 59158 39233
rect 59492 39150 59590 39248
rect 59888 39150 59986 39248
rect 60270 39136 60368 39234
rect 60702 39136 60800 39234
rect 61127 39194 61225 39292
rect 12600 38913 12698 39011
rect 54552 38913 54650 39011
rect 6025 38778 6123 38876
rect 6450 38778 6548 38876
rect 6882 38778 6980 38876
rect 7264 38755 7362 38853
rect 7660 38755 7758 38853
rect 59492 38755 59590 38853
rect 59888 38755 59986 38853
rect 60270 38778 60368 38876
rect 60702 38778 60800 38876
rect 61127 38778 61225 38876
rect 12600 38597 12698 38695
rect 54552 38597 54650 38695
rect 6025 38404 6123 38502
rect 6450 38346 6548 38444
rect 6882 38346 6980 38444
rect 7264 38360 7362 38458
rect 7660 38360 7758 38458
rect 12600 38360 12698 38458
rect 54552 38360 54650 38458
rect 59492 38360 59590 38458
rect 59888 38360 59986 38458
rect 60270 38346 60368 38444
rect 60702 38346 60800 38444
rect 61127 38404 61225 38502
rect 12600 38123 12698 38221
rect 54552 38123 54650 38221
rect 6025 37988 6123 38086
rect 6450 37988 6548 38086
rect 6882 37988 6980 38086
rect 7264 37965 7362 38063
rect 7660 37965 7758 38063
rect 59492 37965 59590 38063
rect 59888 37965 59986 38063
rect 60270 37988 60368 38086
rect 60702 37988 60800 38086
rect 61127 37988 61225 38086
rect 12600 37807 12698 37905
rect 54552 37807 54650 37905
rect 6025 37614 6123 37712
rect 6450 37556 6548 37654
rect 6882 37556 6980 37654
rect 7264 37570 7362 37668
rect 7660 37570 7758 37668
rect 12600 37570 12698 37668
rect 54552 37570 54650 37668
rect 59492 37570 59590 37668
rect 59888 37570 59986 37668
rect 60270 37556 60368 37654
rect 60702 37556 60800 37654
rect 61127 37614 61225 37712
rect 12600 37333 12698 37431
rect 54552 37333 54650 37431
rect 6025 37198 6123 37296
rect 6450 37198 6548 37296
rect 6882 37198 6980 37296
rect 7264 37175 7362 37273
rect 7660 37175 7758 37273
rect 59492 37175 59590 37273
rect 59888 37175 59986 37273
rect 60270 37198 60368 37296
rect 60702 37198 60800 37296
rect 61127 37198 61225 37296
rect 12600 37017 12698 37115
rect 54552 37017 54650 37115
rect 6025 36824 6123 36922
rect 6450 36766 6548 36864
rect 6882 36766 6980 36864
rect 7264 36780 7362 36878
rect 7660 36780 7758 36878
rect 12600 36780 12698 36878
rect 54552 36780 54650 36878
rect 59492 36780 59590 36878
rect 59888 36780 59986 36878
rect 60270 36766 60368 36864
rect 60702 36766 60800 36864
rect 61127 36824 61225 36922
rect 12600 36543 12698 36641
rect 54552 36543 54650 36641
rect 6025 36408 6123 36506
rect 6450 36408 6548 36506
rect 6882 36408 6980 36506
rect 7264 36385 7362 36483
rect 7660 36385 7758 36483
rect 59492 36385 59590 36483
rect 59888 36385 59986 36483
rect 60270 36408 60368 36506
rect 60702 36408 60800 36506
rect 61127 36408 61225 36506
rect 12600 36227 12698 36325
rect 54552 36227 54650 36325
rect 6025 36034 6123 36132
rect 6450 35976 6548 36074
rect 6882 35976 6980 36074
rect 7264 35990 7362 36088
rect 7660 35990 7758 36088
rect 12600 35990 12698 36088
rect 54552 35990 54650 36088
rect 59492 35990 59590 36088
rect 59888 35990 59986 36088
rect 60270 35976 60368 36074
rect 60702 35976 60800 36074
rect 61127 36034 61225 36132
rect 12600 35753 12698 35851
rect 54552 35753 54650 35851
rect 6025 35618 6123 35716
rect 6450 35618 6548 35716
rect 6882 35618 6980 35716
rect 7264 35595 7362 35693
rect 7660 35595 7758 35693
rect 59492 35595 59590 35693
rect 59888 35595 59986 35693
rect 60270 35618 60368 35716
rect 60702 35618 60800 35716
rect 61127 35618 61225 35716
rect 12600 35437 12698 35535
rect 54552 35437 54650 35535
rect 6025 35244 6123 35342
rect 6450 35186 6548 35284
rect 6882 35186 6980 35284
rect 7264 35200 7362 35298
rect 7660 35200 7758 35298
rect 12600 35200 12698 35298
rect 54552 35200 54650 35298
rect 59492 35200 59590 35298
rect 59888 35200 59986 35298
rect 60270 35186 60368 35284
rect 60702 35186 60800 35284
rect 61127 35244 61225 35342
rect 12600 34963 12698 35061
rect 54552 34963 54650 35061
rect 6025 34828 6123 34926
rect 6450 34828 6548 34926
rect 6882 34828 6980 34926
rect 7264 34805 7362 34903
rect 7660 34805 7758 34903
rect 59492 34805 59590 34903
rect 59888 34805 59986 34903
rect 60270 34828 60368 34926
rect 60702 34828 60800 34926
rect 61127 34828 61225 34926
rect 12600 34647 12698 34745
rect 54552 34647 54650 34745
rect 6025 34454 6123 34552
rect 6450 34396 6548 34494
rect 6882 34396 6980 34494
rect 7264 34410 7362 34508
rect 7660 34410 7758 34508
rect 12600 34410 12698 34508
rect 54552 34410 54650 34508
rect 59492 34410 59590 34508
rect 59888 34410 59986 34508
rect 60270 34396 60368 34494
rect 60702 34396 60800 34494
rect 61127 34454 61225 34552
rect 12600 34173 12698 34271
rect 54552 34173 54650 34271
rect 6025 34038 6123 34136
rect 6450 34038 6548 34136
rect 6882 34038 6980 34136
rect 7264 34015 7362 34113
rect 7660 34015 7758 34113
rect 59492 34015 59590 34113
rect 59888 34015 59986 34113
rect 60270 34038 60368 34136
rect 60702 34038 60800 34136
rect 61127 34038 61225 34136
rect 12600 33857 12698 33955
rect 54552 33857 54650 33955
rect 6025 33664 6123 33762
rect 6450 33606 6548 33704
rect 6882 33606 6980 33704
rect 7264 33620 7362 33718
rect 7660 33620 7758 33718
rect 12600 33620 12698 33718
rect 54552 33620 54650 33718
rect 59492 33620 59590 33718
rect 59888 33620 59986 33718
rect 60270 33606 60368 33704
rect 60702 33606 60800 33704
rect 61127 33664 61225 33762
rect 12600 33383 12698 33481
rect 54552 33383 54650 33481
rect 6025 33248 6123 33346
rect 6450 33248 6548 33346
rect 6882 33248 6980 33346
rect 7264 33225 7362 33323
rect 7660 33225 7758 33323
rect 59492 33225 59590 33323
rect 59888 33225 59986 33323
rect 60270 33248 60368 33346
rect 60702 33248 60800 33346
rect 61127 33248 61225 33346
rect 12600 33067 12698 33165
rect 54552 33067 54650 33165
rect 6025 32874 6123 32972
rect 6450 32816 6548 32914
rect 6882 32816 6980 32914
rect 7264 32830 7362 32928
rect 7660 32830 7758 32928
rect 12600 32830 12698 32928
rect 54552 32830 54650 32928
rect 59492 32830 59590 32928
rect 59888 32830 59986 32928
rect 60270 32816 60368 32914
rect 60702 32816 60800 32914
rect 61127 32874 61225 32972
rect 12600 32593 12698 32691
rect 54552 32593 54650 32691
rect 6025 32458 6123 32556
rect 6450 32458 6548 32556
rect 6882 32458 6980 32556
rect 7264 32435 7362 32533
rect 7660 32435 7758 32533
rect 59492 32435 59590 32533
rect 59888 32435 59986 32533
rect 60270 32458 60368 32556
rect 60702 32458 60800 32556
rect 61127 32458 61225 32556
rect 12600 32277 12698 32375
rect 54552 32277 54650 32375
rect 6025 32084 6123 32182
rect 6450 32026 6548 32124
rect 6882 32026 6980 32124
rect 7264 32040 7362 32138
rect 7660 32040 7758 32138
rect 12600 32040 12698 32138
rect 54552 32040 54650 32138
rect 59492 32040 59590 32138
rect 59888 32040 59986 32138
rect 60270 32026 60368 32124
rect 60702 32026 60800 32124
rect 61127 32084 61225 32182
rect 12600 31803 12698 31901
rect 54552 31803 54650 31901
rect 6025 31668 6123 31766
rect 6450 31668 6548 31766
rect 6882 31668 6980 31766
rect 7264 31645 7362 31743
rect 7660 31645 7758 31743
rect 59492 31645 59590 31743
rect 59888 31645 59986 31743
rect 60270 31668 60368 31766
rect 60702 31668 60800 31766
rect 61127 31668 61225 31766
rect 12600 31487 12698 31585
rect 54552 31487 54650 31585
rect 6025 31294 6123 31392
rect 6450 31236 6548 31334
rect 6882 31236 6980 31334
rect 7264 31250 7362 31348
rect 7660 31250 7758 31348
rect 12600 31250 12698 31348
rect 54552 31250 54650 31348
rect 59492 31250 59590 31348
rect 59888 31250 59986 31348
rect 60270 31236 60368 31334
rect 60702 31236 60800 31334
rect 61127 31294 61225 31392
rect 12600 31013 12698 31111
rect 54552 31013 54650 31111
rect 6025 30878 6123 30976
rect 6450 30878 6548 30976
rect 6882 30878 6980 30976
rect 7264 30855 7362 30953
rect 7660 30855 7758 30953
rect 59492 30855 59590 30953
rect 59888 30855 59986 30953
rect 60270 30878 60368 30976
rect 60702 30878 60800 30976
rect 61127 30878 61225 30976
rect 12600 30697 12698 30795
rect 54552 30697 54650 30795
rect 6025 30504 6123 30602
rect 6450 30446 6548 30544
rect 6882 30446 6980 30544
rect 7264 30460 7362 30558
rect 7660 30460 7758 30558
rect 12600 30460 12698 30558
rect 54552 30460 54650 30558
rect 59492 30460 59590 30558
rect 59888 30460 59986 30558
rect 60270 30446 60368 30544
rect 60702 30446 60800 30544
rect 61127 30504 61225 30602
rect 12600 30223 12698 30321
rect 54552 30223 54650 30321
rect 6025 30088 6123 30186
rect 6450 30088 6548 30186
rect 6882 30088 6980 30186
rect 7264 30065 7362 30163
rect 7660 30065 7758 30163
rect 59492 30065 59590 30163
rect 59888 30065 59986 30163
rect 60270 30088 60368 30186
rect 60702 30088 60800 30186
rect 61127 30088 61225 30186
rect 12600 29907 12698 30005
rect 54552 29907 54650 30005
rect 6025 29714 6123 29812
rect 6450 29656 6548 29754
rect 6882 29656 6980 29754
rect 7264 29670 7362 29768
rect 7660 29670 7758 29768
rect 12600 29670 12698 29768
rect 54552 29670 54650 29768
rect 59492 29670 59590 29768
rect 59888 29670 59986 29768
rect 60270 29656 60368 29754
rect 60702 29656 60800 29754
rect 61127 29714 61225 29812
rect 12600 29433 12698 29531
rect 54552 29433 54650 29531
rect 6025 29298 6123 29396
rect 6450 29298 6548 29396
rect 6882 29298 6980 29396
rect 7264 29275 7362 29373
rect 7660 29275 7758 29373
rect 59492 29275 59590 29373
rect 59888 29275 59986 29373
rect 60270 29298 60368 29396
rect 60702 29298 60800 29396
rect 61127 29298 61225 29396
rect 12600 29117 12698 29215
rect 54552 29117 54650 29215
rect 6025 28924 6123 29022
rect 6450 28866 6548 28964
rect 6882 28866 6980 28964
rect 7264 28880 7362 28978
rect 7660 28880 7758 28978
rect 12600 28880 12698 28978
rect 54552 28880 54650 28978
rect 59492 28880 59590 28978
rect 59888 28880 59986 28978
rect 60270 28866 60368 28964
rect 60702 28866 60800 28964
rect 61127 28924 61225 29022
rect 12600 28643 12698 28741
rect 54552 28643 54650 28741
rect 6025 28508 6123 28606
rect 6450 28508 6548 28606
rect 6882 28508 6980 28606
rect 7264 28485 7362 28583
rect 7660 28485 7758 28583
rect 59492 28485 59590 28583
rect 59888 28485 59986 28583
rect 60270 28508 60368 28606
rect 60702 28508 60800 28606
rect 61127 28508 61225 28606
rect 12600 28327 12698 28425
rect 54552 28327 54650 28425
rect 6025 28134 6123 28232
rect 6450 28076 6548 28174
rect 6882 28076 6980 28174
rect 7264 28090 7362 28188
rect 7660 28090 7758 28188
rect 12600 28090 12698 28188
rect 54552 28090 54650 28188
rect 59492 28090 59590 28188
rect 59888 28090 59986 28188
rect 60270 28076 60368 28174
rect 60702 28076 60800 28174
rect 61127 28134 61225 28232
rect 12600 27853 12698 27951
rect 54552 27853 54650 27951
rect 6025 27718 6123 27816
rect 6450 27718 6548 27816
rect 6882 27718 6980 27816
rect 7264 27695 7362 27793
rect 7660 27695 7758 27793
rect 59492 27695 59590 27793
rect 59888 27695 59986 27793
rect 60270 27718 60368 27816
rect 60702 27718 60800 27816
rect 61127 27718 61225 27816
rect 12600 27537 12698 27635
rect 54552 27537 54650 27635
rect 6025 27344 6123 27442
rect 6450 27286 6548 27384
rect 6882 27286 6980 27384
rect 7264 27300 7362 27398
rect 7660 27300 7758 27398
rect 12600 27300 12698 27398
rect 54552 27300 54650 27398
rect 59492 27300 59590 27398
rect 59888 27300 59986 27398
rect 60270 27286 60368 27384
rect 60702 27286 60800 27384
rect 61127 27344 61225 27442
rect 12600 27063 12698 27161
rect 54552 27063 54650 27161
rect 6025 26928 6123 27026
rect 6450 26928 6548 27026
rect 6882 26928 6980 27026
rect 7264 26905 7362 27003
rect 7660 26905 7758 27003
rect 59492 26905 59590 27003
rect 59888 26905 59986 27003
rect 60270 26928 60368 27026
rect 60702 26928 60800 27026
rect 61127 26928 61225 27026
rect 12600 26747 12698 26845
rect 54552 26747 54650 26845
rect 6025 26554 6123 26652
rect 6450 26496 6548 26594
rect 6882 26496 6980 26594
rect 7264 26510 7362 26608
rect 7660 26510 7758 26608
rect 12600 26510 12698 26608
rect 54552 26510 54650 26608
rect 59492 26510 59590 26608
rect 59888 26510 59986 26608
rect 60270 26496 60368 26594
rect 60702 26496 60800 26594
rect 61127 26554 61225 26652
rect 12600 26273 12698 26371
rect 54552 26273 54650 26371
rect 6025 26138 6123 26236
rect 6450 26138 6548 26236
rect 6882 26138 6980 26236
rect 7264 26115 7362 26213
rect 7660 26115 7758 26213
rect 59492 26115 59590 26213
rect 59888 26115 59986 26213
rect 60270 26138 60368 26236
rect 60702 26138 60800 26236
rect 61127 26138 61225 26236
rect 12600 25957 12698 26055
rect 54552 25957 54650 26055
rect 6025 25764 6123 25862
rect 6450 25706 6548 25804
rect 6882 25706 6980 25804
rect 7264 25720 7362 25818
rect 7660 25720 7758 25818
rect 12600 25720 12698 25818
rect 54552 25720 54650 25818
rect 59492 25720 59590 25818
rect 59888 25720 59986 25818
rect 60270 25706 60368 25804
rect 60702 25706 60800 25804
rect 61127 25764 61225 25862
rect 12600 25483 12698 25581
rect 54552 25483 54650 25581
rect 6025 25348 6123 25446
rect 6450 25348 6548 25446
rect 6882 25348 6980 25446
rect 7264 25325 7362 25423
rect 7660 25325 7758 25423
rect 59492 25325 59590 25423
rect 59888 25325 59986 25423
rect 60270 25348 60368 25446
rect 60702 25348 60800 25446
rect 61127 25348 61225 25446
rect 12600 25167 12698 25265
rect 54552 25167 54650 25265
rect 6025 24974 6123 25072
rect 6450 24916 6548 25014
rect 6882 24916 6980 25014
rect 7264 24930 7362 25028
rect 7660 24930 7758 25028
rect 12600 24930 12698 25028
rect 54552 24930 54650 25028
rect 59492 24930 59590 25028
rect 59888 24930 59986 25028
rect 60270 24916 60368 25014
rect 60702 24916 60800 25014
rect 61127 24974 61225 25072
rect 12600 24693 12698 24791
rect 54552 24693 54650 24791
rect 6025 24558 6123 24656
rect 6450 24558 6548 24656
rect 6882 24558 6980 24656
rect 7264 24535 7362 24633
rect 7660 24535 7758 24633
rect 59492 24535 59590 24633
rect 59888 24535 59986 24633
rect 60270 24558 60368 24656
rect 60702 24558 60800 24656
rect 61127 24558 61225 24656
rect 12600 24377 12698 24475
rect 54552 24377 54650 24475
rect 6025 24184 6123 24282
rect 6450 24126 6548 24224
rect 6882 24126 6980 24224
rect 7264 24140 7362 24238
rect 7660 24140 7758 24238
rect 12600 24140 12698 24238
rect 54552 24140 54650 24238
rect 59492 24140 59590 24238
rect 59888 24140 59986 24238
rect 60270 24126 60368 24224
rect 60702 24126 60800 24224
rect 61127 24184 61225 24282
rect 12600 23903 12698 24001
rect 54552 23903 54650 24001
rect 6025 23768 6123 23866
rect 6450 23768 6548 23866
rect 6882 23768 6980 23866
rect 7264 23745 7362 23843
rect 7660 23745 7758 23843
rect 59492 23745 59590 23843
rect 59888 23745 59986 23843
rect 60270 23768 60368 23866
rect 60702 23768 60800 23866
rect 61127 23768 61225 23866
rect 12600 23587 12698 23685
rect 54552 23587 54650 23685
rect 6025 23394 6123 23492
rect 6450 23336 6548 23434
rect 6882 23336 6980 23434
rect 7264 23350 7362 23448
rect 7660 23350 7758 23448
rect 12600 23350 12698 23448
rect 54552 23350 54650 23448
rect 59492 23350 59590 23448
rect 59888 23350 59986 23448
rect 60270 23336 60368 23434
rect 60702 23336 60800 23434
rect 61127 23394 61225 23492
rect 12600 23113 12698 23211
rect 54552 23113 54650 23211
rect 6025 22978 6123 23076
rect 6450 22978 6548 23076
rect 6882 22978 6980 23076
rect 7264 22955 7362 23053
rect 7660 22955 7758 23053
rect 59492 22955 59590 23053
rect 59888 22955 59986 23053
rect 60270 22978 60368 23076
rect 60702 22978 60800 23076
rect 61127 22978 61225 23076
rect 12600 22797 12698 22895
rect 54552 22797 54650 22895
rect 6025 22604 6123 22702
rect 6450 22546 6548 22644
rect 6882 22546 6980 22644
rect 7264 22560 7362 22658
rect 7660 22560 7758 22658
rect 12600 22560 12698 22658
rect 54552 22560 54650 22658
rect 59492 22560 59590 22658
rect 59888 22560 59986 22658
rect 60270 22546 60368 22644
rect 60702 22546 60800 22644
rect 61127 22604 61225 22702
rect 12600 22323 12698 22421
rect 54552 22323 54650 22421
rect 6025 22188 6123 22286
rect 6450 22188 6548 22286
rect 6882 22188 6980 22286
rect 7264 22165 7362 22263
rect 7660 22165 7758 22263
rect 59492 22165 59590 22263
rect 59888 22165 59986 22263
rect 60270 22188 60368 22286
rect 60702 22188 60800 22286
rect 61127 22188 61225 22286
rect 12600 22007 12698 22105
rect 54552 22007 54650 22105
rect 6025 21814 6123 21912
rect 6450 21756 6548 21854
rect 6882 21756 6980 21854
rect 7264 21770 7362 21868
rect 7660 21770 7758 21868
rect 12600 21770 12698 21868
rect 54552 21770 54650 21868
rect 59492 21770 59590 21868
rect 59888 21770 59986 21868
rect 60270 21756 60368 21854
rect 60702 21756 60800 21854
rect 61127 21814 61225 21912
rect 12600 21533 12698 21631
rect 54552 21533 54650 21631
rect 2611 21398 2709 21496
rect 3036 21398 3134 21496
rect 3468 21398 3566 21496
rect 3850 21375 3948 21473
rect 4246 21375 4344 21473
rect 6025 21398 6123 21496
rect 6450 21398 6548 21496
rect 6882 21398 6980 21496
rect 7264 21375 7362 21473
rect 7660 21375 7758 21473
rect 59492 21375 59590 21473
rect 59888 21375 59986 21473
rect 60270 21398 60368 21496
rect 60702 21398 60800 21496
rect 61127 21398 61225 21496
rect 62906 21375 63004 21473
rect 63302 21375 63400 21473
rect 63684 21398 63782 21496
rect 64116 21398 64214 21496
rect 64541 21398 64639 21496
rect 12600 21217 12698 21315
rect 54552 21217 54650 21315
rect 6025 21024 6123 21122
rect 6450 20966 6548 21064
rect 6882 20966 6980 21064
rect 7264 20980 7362 21078
rect 7660 20980 7758 21078
rect 12600 20980 12698 21078
rect 54552 20980 54650 21078
rect 59492 20980 59590 21078
rect 59888 20980 59986 21078
rect 60270 20966 60368 21064
rect 60702 20966 60800 21064
rect 61127 21024 61225 21122
rect 12600 20743 12698 20841
rect 54552 20743 54650 20841
rect 2611 20608 2709 20706
rect 3036 20608 3134 20706
rect 3468 20608 3566 20706
rect 3850 20585 3948 20683
rect 4246 20585 4344 20683
rect 6025 20608 6123 20706
rect 6450 20608 6548 20706
rect 6882 20608 6980 20706
rect 7264 20585 7362 20683
rect 7660 20585 7758 20683
rect 59492 20585 59590 20683
rect 59888 20585 59986 20683
rect 60270 20608 60368 20706
rect 60702 20608 60800 20706
rect 61127 20608 61225 20706
rect 62906 20585 63004 20683
rect 63302 20585 63400 20683
rect 63684 20608 63782 20706
rect 64116 20608 64214 20706
rect 64541 20608 64639 20706
rect 12600 20427 12698 20525
rect 54552 20427 54650 20525
rect 6025 20234 6123 20332
rect 6450 20176 6548 20274
rect 6882 20176 6980 20274
rect 7264 20190 7362 20288
rect 7660 20190 7758 20288
rect 12600 20190 12698 20288
rect 54552 20190 54650 20288
rect 59492 20190 59590 20288
rect 59888 20190 59986 20288
rect 60270 20176 60368 20274
rect 60702 20176 60800 20274
rect 61127 20234 61225 20332
rect 12600 19953 12698 20051
rect 54552 19953 54650 20051
rect 2611 19818 2709 19916
rect 3036 19818 3134 19916
rect 3468 19818 3566 19916
rect 3850 19795 3948 19893
rect 4246 19795 4344 19893
rect 6025 19818 6123 19916
rect 6450 19818 6548 19916
rect 6882 19818 6980 19916
rect 7264 19795 7362 19893
rect 7660 19795 7758 19893
rect 59492 19795 59590 19893
rect 59888 19795 59986 19893
rect 60270 19818 60368 19916
rect 60702 19818 60800 19916
rect 61127 19818 61225 19916
rect 62906 19795 63004 19893
rect 63302 19795 63400 19893
rect 63684 19818 63782 19916
rect 64116 19818 64214 19916
rect 64541 19818 64639 19916
rect 12600 19637 12698 19735
rect 54552 19637 54650 19735
rect 6025 19444 6123 19542
rect 6450 19386 6548 19484
rect 6882 19386 6980 19484
rect 7264 19400 7362 19498
rect 7660 19400 7758 19498
rect 12600 19400 12698 19498
rect 54552 19400 54650 19498
rect 59492 19400 59590 19498
rect 59888 19400 59986 19498
rect 60270 19386 60368 19484
rect 60702 19386 60800 19484
rect 61127 19444 61225 19542
rect 12600 19163 12698 19261
rect 54552 19163 54650 19261
rect 1156 19005 1254 19103
rect 1552 19005 1650 19103
rect 2611 19028 2709 19126
rect 3036 19028 3134 19126
rect 3468 19028 3566 19126
rect 3850 19005 3948 19103
rect 4246 19005 4344 19103
rect 6025 19028 6123 19126
rect 6450 19028 6548 19126
rect 6882 19028 6980 19126
rect 7264 19005 7362 19103
rect 7660 19005 7758 19103
rect 59492 19005 59590 19103
rect 59888 19005 59986 19103
rect 60270 19028 60368 19126
rect 60702 19028 60800 19126
rect 61127 19028 61225 19126
rect 62906 19005 63004 19103
rect 63302 19005 63400 19103
rect 63684 19028 63782 19126
rect 64116 19028 64214 19126
rect 64541 19028 64639 19126
rect 65600 19005 65698 19103
rect 65996 19005 66094 19103
rect 12600 18847 12698 18945
rect 54552 18847 54650 18945
rect 6025 18654 6123 18752
rect 6450 18596 6548 18694
rect 6882 18596 6980 18694
rect 7264 18610 7362 18708
rect 7660 18610 7758 18708
rect 12600 18610 12698 18708
rect 54552 18610 54650 18708
rect 59492 18610 59590 18708
rect 59888 18610 59986 18708
rect 60270 18596 60368 18694
rect 60702 18596 60800 18694
rect 61127 18654 61225 18752
rect 12600 18373 12698 18471
rect 54552 18373 54650 18471
rect 6025 18238 6123 18336
rect 6450 18238 6548 18336
rect 6882 18238 6980 18336
rect 7264 18215 7362 18313
rect 7660 18215 7758 18313
rect 59492 18215 59590 18313
rect 59888 18215 59986 18313
rect 60270 18238 60368 18336
rect 60702 18238 60800 18336
rect 61127 18238 61225 18336
rect 12600 18057 12698 18155
rect 54552 18057 54650 18155
rect 6025 17864 6123 17962
rect 6450 17806 6548 17904
rect 6882 17806 6980 17904
rect 7264 17820 7362 17918
rect 7660 17820 7758 17918
rect 12600 17820 12698 17918
rect 54552 17820 54650 17918
rect 59492 17820 59590 17918
rect 59888 17820 59986 17918
rect 60270 17806 60368 17904
rect 60702 17806 60800 17904
rect 61127 17864 61225 17962
rect 12600 17583 12698 17681
rect 54552 17583 54650 17681
rect 3046 17432 3144 17530
rect 3471 17432 3569 17530
rect 3850 17425 3948 17523
rect 4246 17425 4344 17523
rect 6025 17448 6123 17546
rect 6450 17448 6548 17546
rect 6882 17448 6980 17546
rect 7264 17425 7362 17523
rect 7660 17425 7758 17523
rect 59492 17425 59590 17523
rect 59888 17425 59986 17523
rect 60270 17448 60368 17546
rect 60702 17448 60800 17546
rect 61127 17448 61225 17546
rect 62906 17425 63004 17523
rect 63302 17425 63400 17523
rect 63681 17432 63779 17530
rect 64106 17432 64204 17530
rect 12600 17267 12698 17365
rect 54552 17267 54650 17365
rect 6025 17074 6123 17172
rect 6450 17016 6548 17114
rect 6882 17016 6980 17114
rect 7264 17030 7362 17128
rect 7660 17030 7758 17128
rect 12600 17030 12698 17128
rect 54552 17030 54650 17128
rect 59492 17030 59590 17128
rect 59888 17030 59986 17128
rect 60270 17016 60368 17114
rect 60702 17016 60800 17114
rect 61127 17074 61225 17172
rect 12600 16793 12698 16891
rect 54552 16793 54650 16891
rect 1752 16635 1850 16733
rect 2148 16635 2246 16733
rect 3046 16642 3144 16740
rect 3471 16642 3569 16740
rect 3850 16635 3948 16733
rect 4246 16635 4344 16733
rect 6025 16658 6123 16756
rect 6450 16658 6548 16756
rect 6882 16658 6980 16756
rect 7264 16635 7362 16733
rect 7660 16635 7758 16733
rect 59492 16635 59590 16733
rect 59888 16635 59986 16733
rect 60270 16658 60368 16756
rect 60702 16658 60800 16756
rect 61127 16658 61225 16756
rect 62906 16635 63004 16733
rect 63302 16635 63400 16733
rect 63681 16642 63779 16740
rect 64106 16642 64204 16740
rect 65004 16635 65102 16733
rect 65400 16635 65498 16733
rect 12600 16477 12698 16575
rect 54552 16477 54650 16575
rect 6025 16284 6123 16382
rect 6450 16226 6548 16324
rect 6882 16226 6980 16324
rect 7264 16240 7362 16338
rect 7660 16240 7758 16338
rect 12600 16240 12698 16338
rect 54552 16240 54650 16338
rect 59492 16240 59590 16338
rect 59888 16240 59986 16338
rect 60270 16226 60368 16324
rect 60702 16226 60800 16324
rect 61127 16284 61225 16382
rect 12600 16003 12698 16101
rect 54552 16003 54650 16101
rect 6025 15868 6123 15966
rect 6450 15868 6548 15966
rect 6882 15868 6980 15966
rect 7264 15845 7362 15943
rect 7660 15845 7758 15943
rect 59492 15845 59590 15943
rect 59888 15845 59986 15943
rect 60270 15868 60368 15966
rect 60702 15868 60800 15966
rect 61127 15868 61225 15966
rect 12600 15687 12698 15785
rect 54552 15687 54650 15785
rect 6025 15494 6123 15592
rect 6450 15436 6548 15534
rect 6882 15436 6980 15534
rect 7264 15450 7362 15548
rect 7660 15450 7758 15548
rect 12600 15450 12698 15548
rect 54552 15450 54650 15548
rect 59492 15450 59590 15548
rect 59888 15450 59986 15548
rect 60270 15436 60368 15534
rect 60702 15436 60800 15534
rect 61127 15494 61225 15592
rect 12600 15213 12698 15311
rect 54552 15213 54650 15311
rect 3046 15062 3144 15160
rect 3471 15062 3569 15160
rect 3850 15055 3948 15153
rect 4246 15055 4344 15153
rect 6025 15078 6123 15176
rect 6450 15078 6548 15176
rect 6882 15078 6980 15176
rect 7264 15055 7362 15153
rect 7660 15055 7758 15153
rect 59492 15055 59590 15153
rect 59888 15055 59986 15153
rect 60270 15078 60368 15176
rect 60702 15078 60800 15176
rect 61127 15078 61225 15176
rect 62906 15055 63004 15153
rect 63302 15055 63400 15153
rect 63681 15062 63779 15160
rect 64106 15062 64204 15160
rect 12600 14897 12698 14995
rect 54552 14897 54650 14995
rect 6025 14704 6123 14802
rect 6450 14646 6548 14744
rect 6882 14646 6980 14744
rect 7264 14660 7362 14758
rect 7660 14660 7758 14758
rect 12600 14660 12698 14758
rect 54552 14660 54650 14758
rect 59492 14660 59590 14758
rect 59888 14660 59986 14758
rect 60270 14646 60368 14744
rect 60702 14646 60800 14744
rect 61127 14704 61225 14802
rect 12600 14423 12698 14521
rect 54552 14423 54650 14521
rect 1752 14265 1850 14363
rect 2148 14265 2246 14363
rect 3046 14272 3144 14370
rect 3471 14272 3569 14370
rect 3850 14265 3948 14363
rect 4246 14265 4344 14363
rect 6025 14288 6123 14386
rect 6450 14288 6548 14386
rect 6882 14288 6980 14386
rect 7264 14265 7362 14363
rect 7660 14265 7758 14363
rect 59492 14265 59590 14363
rect 59888 14265 59986 14363
rect 60270 14288 60368 14386
rect 60702 14288 60800 14386
rect 61127 14288 61225 14386
rect 62906 14265 63004 14363
rect 63302 14265 63400 14363
rect 63681 14272 63779 14370
rect 64106 14272 64204 14370
rect 65004 14265 65102 14363
rect 65400 14265 65498 14363
rect 12600 14107 12698 14205
rect 54552 14107 54650 14205
rect 12600 13870 12698 13968
rect 54552 13870 54650 13968
rect 7685 13679 7783 13777
rect 8517 13685 8615 13783
rect 11208 13673 11306 13771
rect 12234 13743 12332 13841
rect 54918 13743 55016 13841
rect 13296 13309 13394 13407
rect 13920 13309 14018 13407
rect 14544 13309 14642 13407
rect 15168 13309 15266 13407
rect 15792 13309 15890 13407
rect 16416 13309 16514 13407
rect 17040 13309 17138 13407
rect 17664 13309 17762 13407
rect 18288 13309 18386 13407
rect 18912 13309 19010 13407
rect 19536 13309 19634 13407
rect 20160 13309 20258 13407
rect 20784 13309 20882 13407
rect 21408 13309 21506 13407
rect 22032 13309 22130 13407
rect 22656 13309 22754 13407
rect 23280 13309 23378 13407
rect 23904 13309 24002 13407
rect 24528 13309 24626 13407
rect 25152 13309 25250 13407
rect 25776 13309 25874 13407
rect 26400 13309 26498 13407
rect 27024 13309 27122 13407
rect 27648 13309 27746 13407
rect 28272 13309 28370 13407
rect 28896 13309 28994 13407
rect 29520 13309 29618 13407
rect 30144 13309 30242 13407
rect 30768 13309 30866 13407
rect 31392 13309 31490 13407
rect 32016 13309 32114 13407
rect 32640 13309 32738 13407
rect 33264 13309 33362 13407
rect 33888 13309 33986 13407
rect 34512 13309 34610 13407
rect 35136 13309 35234 13407
rect 35760 13309 35858 13407
rect 36384 13309 36482 13407
rect 37008 13309 37106 13407
rect 37632 13309 37730 13407
rect 38256 13309 38354 13407
rect 38880 13309 38978 13407
rect 39504 13309 39602 13407
rect 40128 13309 40226 13407
rect 40752 13309 40850 13407
rect 41376 13309 41474 13407
rect 42000 13309 42098 13407
rect 42624 13309 42722 13407
rect 43248 13309 43346 13407
rect 43872 13309 43970 13407
rect 44496 13309 44594 13407
rect 45120 13309 45218 13407
rect 45744 13309 45842 13407
rect 46368 13309 46466 13407
rect 46992 13309 47090 13407
rect 47616 13309 47714 13407
rect 48240 13309 48338 13407
rect 48864 13309 48962 13407
rect 49488 13309 49586 13407
rect 50112 13309 50210 13407
rect 50736 13309 50834 13407
rect 51360 13309 51458 13407
rect 51984 13309 52082 13407
rect 52608 13309 52706 13407
rect 53232 13309 53330 13407
rect 53856 13309 53954 13407
rect 13415 12718 13513 12816
rect 13801 12718 13899 12816
rect 14663 12718 14761 12816
rect 15049 12718 15147 12816
rect 15911 12718 16009 12816
rect 16297 12718 16395 12816
rect 17159 12718 17257 12816
rect 17545 12718 17643 12816
rect 18407 12718 18505 12816
rect 18793 12718 18891 12816
rect 19655 12718 19753 12816
rect 20041 12718 20139 12816
rect 20903 12718 21001 12816
rect 21289 12718 21387 12816
rect 22151 12718 22249 12816
rect 22537 12718 22635 12816
rect 23399 12718 23497 12816
rect 23785 12718 23883 12816
rect 24647 12718 24745 12816
rect 25033 12718 25131 12816
rect 25895 12718 25993 12816
rect 26281 12718 26379 12816
rect 27143 12718 27241 12816
rect 27529 12718 27627 12816
rect 28391 12718 28489 12816
rect 28777 12718 28875 12816
rect 29639 12718 29737 12816
rect 30025 12718 30123 12816
rect 30887 12718 30985 12816
rect 31273 12718 31371 12816
rect 32135 12718 32233 12816
rect 32521 12718 32619 12816
rect 33383 12718 33481 12816
rect 33769 12718 33867 12816
rect 34631 12718 34729 12816
rect 35017 12718 35115 12816
rect 35879 12718 35977 12816
rect 36265 12718 36363 12816
rect 37127 12718 37225 12816
rect 37513 12718 37611 12816
rect 38375 12718 38473 12816
rect 38761 12718 38859 12816
rect 39623 12718 39721 12816
rect 40009 12718 40107 12816
rect 40871 12718 40969 12816
rect 41257 12718 41355 12816
rect 42119 12718 42217 12816
rect 42505 12718 42603 12816
rect 43367 12718 43465 12816
rect 43753 12718 43851 12816
rect 44615 12718 44713 12816
rect 45001 12718 45099 12816
rect 45863 12718 45961 12816
rect 46249 12718 46347 12816
rect 47111 12718 47209 12816
rect 47497 12718 47595 12816
rect 48359 12718 48457 12816
rect 48745 12718 48843 12816
rect 49607 12718 49705 12816
rect 49993 12718 50091 12816
rect 50855 12718 50953 12816
rect 51241 12718 51339 12816
rect 52103 12718 52201 12816
rect 52489 12718 52587 12816
rect 53351 12718 53449 12816
rect 11644 12178 11710 12181
rect 11644 12176 32938 12178
rect 11644 12120 11649 12176
rect 11705 12120 32938 12176
rect 11644 12118 32938 12120
rect 11644 12115 11710 12118
rect 13544 12029 13610 12032
rect 0 12027 13610 12029
rect 0 11971 13549 12027
rect 13605 11971 13610 12027
rect 0 11969 13610 11971
rect 13544 11966 13610 11969
rect 4676 11312 4774 11410
rect 6036 11312 6134 11410
rect 14232 11169 14330 11267
rect 15480 11169 15578 11267
rect 16728 11169 16826 11267
rect 17976 11169 18074 11267
rect 19224 11169 19322 11267
rect 20472 11169 20570 11267
rect 21720 11169 21818 11267
rect 22968 11169 23066 11267
rect 24216 11169 24314 11267
rect 25464 11169 25562 11267
rect 26712 11169 26810 11267
rect 27960 11169 28058 11267
rect 29208 11169 29306 11267
rect 30456 11169 30554 11267
rect 31704 11169 31802 11267
rect 32952 11169 33050 11267
rect 34200 11169 34298 11267
rect 35448 11169 35546 11267
rect 36696 11169 36794 11267
rect 37944 11169 38042 11267
rect 39192 11169 39290 11267
rect 40440 11169 40538 11267
rect 41688 11169 41786 11267
rect 42936 11169 43034 11267
rect 44184 11169 44282 11267
rect 45432 11169 45530 11267
rect 46680 11169 46778 11267
rect 47928 11169 48026 11267
rect 49176 11169 49274 11267
rect 50424 11169 50522 11267
rect 51672 11169 51770 11267
rect 52920 11169 53018 11267
rect 6833 10722 6899 10725
rect 7112 10722 7178 10725
rect 6833 10720 7178 10722
rect 6833 10664 6838 10720
rect 6894 10664 7117 10720
rect 7173 10664 7178 10720
rect 6833 10662 7178 10664
rect 6833 10659 6899 10662
rect 7112 10659 7178 10662
rect 7112 10491 7178 10494
rect 7112 10489 12313 10491
rect 7112 10433 7117 10489
rect 7173 10433 12313 10489
rect 7112 10431 12313 10433
rect 7112 10428 7178 10431
rect 7928 10367 7994 10370
rect 7928 10365 12313 10367
rect 7928 10309 7933 10365
rect 7989 10309 12313 10365
rect 7928 10307 12313 10309
rect 7928 10304 7994 10307
rect 7792 10243 7858 10246
rect 7792 10241 12313 10243
rect 7792 10185 7797 10241
rect 7853 10185 12313 10241
rect 7792 10183 12313 10185
rect 7792 10180 7858 10183
rect 7656 10119 7722 10122
rect 7656 10117 12313 10119
rect 7656 10061 7661 10117
rect 7717 10061 12313 10117
rect 7656 10059 12313 10061
rect 7656 10056 7722 10059
rect 4676 9898 4774 9996
rect 6036 9898 6134 9996
rect 7520 9995 7586 9998
rect 7520 9993 12313 9995
rect 7520 9937 7525 9993
rect 7581 9937 12313 9993
rect 7520 9935 12313 9937
rect 7520 9932 7586 9935
rect 7384 9871 7450 9874
rect 7384 9869 12313 9871
rect 7384 9813 7389 9869
rect 7445 9813 12313 9869
rect 7384 9811 12313 9813
rect 7384 9808 7450 9811
rect 7248 9747 7314 9750
rect 7248 9745 12313 9747
rect 7248 9689 7253 9745
rect 7309 9689 12313 9745
rect 7248 9687 12313 9689
rect 7248 9684 7314 9687
rect 7112 9623 7178 9626
rect 7112 9621 12313 9623
rect 7112 9565 7117 9621
rect 7173 9565 12313 9621
rect 7112 9563 12313 9565
rect 7112 9560 7178 9563
rect 6833 9232 6899 9235
rect 7928 9232 7994 9235
rect 6833 9230 7994 9232
rect 6833 9174 6838 9230
rect 6894 9174 7933 9230
rect 7989 9174 7994 9230
rect 6833 9172 7994 9174
rect 6833 9169 6899 9172
rect 7928 9169 7994 9172
rect 11768 8907 11834 8910
rect 11768 8905 30692 8907
rect 11768 8849 11773 8905
rect 11829 8849 30692 8905
rect 11768 8847 30692 8849
rect 11768 8844 11834 8847
rect 14059 8676 14157 8774
rect 19051 8676 19149 8774
rect 24043 8676 24141 8774
rect 29035 8676 29133 8774
rect 34027 8676 34125 8774
rect 39019 8676 39117 8774
rect 44011 8676 44109 8774
rect 49003 8676 49101 8774
rect 4676 8484 4774 8582
rect 6036 8484 6134 8582
rect 13977 7902 14075 8000
rect 18969 7902 19067 8000
rect 23961 7902 24059 8000
rect 28953 7902 29051 8000
rect 33945 7902 34043 8000
rect 38937 7902 39035 8000
rect 43929 7902 44027 8000
rect 48921 7902 49019 8000
rect 6833 7894 6899 7897
rect 7792 7894 7858 7897
rect 6833 7892 7858 7894
rect 6833 7836 6838 7892
rect 6894 7836 7797 7892
rect 7853 7836 7858 7892
rect 6833 7834 7858 7836
rect 6833 7831 6899 7834
rect 7792 7831 7858 7834
rect 4676 7070 4774 7168
rect 6036 7070 6134 7168
rect 13989 7064 14087 7162
rect 18981 7064 19079 7162
rect 23973 7064 24071 7162
rect 28965 7064 29063 7162
rect 33957 7064 34055 7162
rect 38949 7064 39047 7162
rect 43941 7064 44039 7162
rect 48933 7064 49031 7162
rect 13989 6742 14087 6840
rect 18981 6742 19079 6840
rect 23973 6742 24071 6840
rect 28965 6742 29063 6840
rect 33957 6742 34055 6840
rect 38949 6742 39047 6840
rect 43941 6742 44039 6840
rect 48933 6742 49031 6840
rect 6833 6404 6899 6407
rect 7656 6404 7722 6407
rect 6833 6402 7722 6404
rect 6833 6346 6838 6402
rect 6894 6346 7661 6402
rect 7717 6346 7722 6402
rect 6833 6344 7722 6346
rect 6833 6341 6899 6344
rect 7656 6341 7722 6344
rect 13875 5949 13973 6047
rect 18867 5949 18965 6047
rect 23859 5949 23957 6047
rect 28851 5949 28949 6047
rect 33843 5949 33941 6047
rect 38835 5949 38933 6047
rect 43827 5949 43925 6047
rect 48819 5949 48917 6047
rect 4676 5656 4774 5754
rect 6036 5656 6134 5754
rect 13864 5512 13962 5610
rect 18856 5512 18954 5610
rect 23848 5512 23946 5610
rect 28840 5512 28938 5610
rect 33832 5512 33930 5610
rect 38824 5512 38922 5610
rect 43816 5512 43914 5610
rect 48808 5512 48906 5610
rect 13985 5180 14083 5278
rect 18977 5180 19075 5278
rect 23969 5180 24067 5278
rect 28961 5180 29059 5278
rect 33953 5180 34051 5278
rect 38945 5180 39043 5278
rect 43937 5180 44035 5278
rect 48929 5180 49027 5278
rect 6833 5066 6899 5069
rect 7520 5066 7586 5069
rect 6833 5064 7586 5066
rect 6833 5008 6838 5064
rect 6894 5008 7525 5064
rect 7581 5008 7586 5064
rect 6833 5006 7586 5008
rect 6833 5003 6899 5006
rect 7520 5003 7586 5006
rect 13870 4978 13968 5076
rect 18862 4978 18960 5076
rect 23854 4978 23952 5076
rect 28846 4978 28944 5076
rect 33838 4978 33936 5076
rect 38830 4978 38928 5076
rect 43822 4978 43920 5076
rect 48814 4978 48912 5076
rect 13884 4562 13982 4660
rect 18876 4562 18974 4660
rect 23868 4562 23966 4660
rect 28860 4562 28958 4660
rect 33852 4562 33950 4660
rect 38844 4562 38942 4660
rect 43836 4562 43934 4660
rect 48828 4562 48926 4660
rect 4676 4242 4774 4340
rect 6036 4242 6134 4340
rect 12234 4119 12332 4217
rect 53544 4119 53642 4217
rect 11892 3596 11958 3599
rect 11892 3594 32938 3596
rect 6833 3576 6899 3579
rect 7384 3576 7450 3579
rect 6833 3574 7450 3576
rect 6833 3518 6838 3574
rect 6894 3518 7389 3574
rect 7445 3518 7450 3574
rect 11892 3538 11897 3594
rect 11953 3538 32938 3594
rect 11892 3536 32938 3538
rect 11892 3533 11958 3536
rect 6833 3516 7450 3518
rect 6833 3513 6899 3516
rect 7384 3513 7450 3516
rect 12234 2999 12332 3097
rect 53544 2999 53642 3097
rect 4676 2828 4774 2926
rect 6036 2828 6134 2926
rect 6833 2238 6899 2241
rect 7248 2238 7314 2241
rect 6833 2236 7314 2238
rect 6833 2180 6838 2236
rect 6894 2180 7253 2236
rect 7309 2180 7314 2236
rect 6833 2178 7314 2180
rect 6833 2175 6899 2178
rect 7248 2175 7314 2178
rect 4676 1414 4774 1512
rect 6036 1414 6134 1512
rect 6833 748 6899 751
rect 7112 748 7178 751
rect 6833 746 7178 748
rect 6833 690 6838 746
rect 6894 690 7117 746
rect 7173 690 7178 746
rect 6833 688 7178 690
rect 6833 685 6899 688
rect 7112 685 7178 688
rect 4676 0 4774 98
rect 6036 0 6134 98
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_0
timestamp 1644511149
transform 1 0 11644 0 1 12111
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_1
timestamp 1644511149
transform 1 0 7928 0 1 10300
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_2
timestamp 1644511149
transform 1 0 6833 0 1 9165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_3
timestamp 1644511149
transform 1 0 7928 0 1 9165
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_4
timestamp 1644511149
transform 1 0 7792 0 1 10176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_5
timestamp 1644511149
transform 1 0 6833 0 1 7827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_6
timestamp 1644511149
transform 1 0 7792 0 1 7827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_7
timestamp 1644511149
transform 1 0 7656 0 1 10052
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_8
timestamp 1644511149
transform 1 0 6833 0 1 6337
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_9
timestamp 1644511149
transform 1 0 7656 0 1 6337
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_10
timestamp 1644511149
transform 1 0 7520 0 1 9928
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_11
timestamp 1644511149
transform 1 0 6833 0 1 4999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_12
timestamp 1644511149
transform 1 0 7520 0 1 4999
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_13
timestamp 1644511149
transform 1 0 7384 0 1 9804
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_14
timestamp 1644511149
transform 1 0 6833 0 1 3509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_15
timestamp 1644511149
transform 1 0 7384 0 1 3509
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_16
timestamp 1644511149
transform 1 0 7248 0 1 9680
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_17
timestamp 1644511149
transform 1 0 6833 0 1 2171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_18
timestamp 1644511149
transform 1 0 7248 0 1 2171
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_19
timestamp 1644511149
transform 1 0 7112 0 1 10424
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_20
timestamp 1644511149
transform 1 0 6833 0 1 10655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_21
timestamp 1644511149
transform 1 0 7112 0 1 10655
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_22
timestamp 1644511149
transform 1 0 7112 0 1 9556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_23
timestamp 1644511149
transform 1 0 6833 0 1 681
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_24
timestamp 1644511149
transform 1 0 7112 0 1 681
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_25
timestamp 1644511149
transform 1 0 13544 0 1 11962
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_26
timestamp 1644511149
transform 1 0 11892 0 1 3529
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_27
timestamp 1644511149
transform 1 0 11768 0 1 8840
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_28
timestamp 1644511149
transform 1 0 55258 0 1 69484
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_29
timestamp 1644511149
transform 1 0 55382 0 1 66213
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_30
timestamp 1644511149
transform 1 0 59772 0 1 68768
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_31
timestamp 1644511149
transform 1 0 60227 0 1 77643
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_32
timestamp 1644511149
transform 1 0 59772 0 1 77643
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_33
timestamp 1644511149
transform 1 0 59636 0 1 68644
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_34
timestamp 1644511149
transform 1 0 60227 0 1 76153
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_35
timestamp 1644511149
transform 1 0 59636 0 1 76153
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_36
timestamp 1644511149
transform 1 0 59500 0 1 68520
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_37
timestamp 1644511149
transform 1 0 60227 0 1 74815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_38
timestamp 1644511149
transform 1 0 59500 0 1 74815
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_39
timestamp 1644511149
transform 1 0 59364 0 1 68396
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_40
timestamp 1644511149
transform 1 0 60227 0 1 73325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_41
timestamp 1644511149
transform 1 0 59364 0 1 73325
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_42
timestamp 1644511149
transform 1 0 59228 0 1 68272
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_43
timestamp 1644511149
transform 1 0 60227 0 1 71987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_44
timestamp 1644511149
transform 1 0 59228 0 1 71987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_45
timestamp 1644511149
transform 1 0 59092 0 1 68024
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_46
timestamp 1644511149
transform 1 0 60227 0 1 69159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_47
timestamp 1644511149
transform 1 0 59092 0 1 69159
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_48
timestamp 1644511149
transform 1 0 58956 0 1 68148
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_49
timestamp 1644511149
transform 1 0 60227 0 1 70497
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_50
timestamp 1644511149
transform 1 0 58956 0 1 70497
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_51
timestamp 1644511149
transform 1 0 58956 0 1 67900
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_52
timestamp 1644511149
transform 1 0 60227 0 1 67669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_53
timestamp 1644511149
transform 1 0 58956 0 1 67669
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_7_54
timestamp 1644511149
transform 1 0 53640 0 1 66362
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_0
timestamp 1644511149
transform 1 0 55065 0 1 16926
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_1
timestamp 1644511149
transform 1 0 55065 0 1 16376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_2
timestamp 1644511149
transform 1 0 55065 0 1 16136
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_3
timestamp 1644511149
transform 1 0 55065 0 1 15586
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_4
timestamp 1644511149
transform 1 0 55065 0 1 15346
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_5
timestamp 1644511149
transform 1 0 55065 0 1 14796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_6
timestamp 1644511149
transform 1 0 55065 0 1 14556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_7
timestamp 1644511149
transform 1 0 55065 0 1 14006
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_8
timestamp 1644511149
transform 1 0 55065 0 1 19296
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_9
timestamp 1644511149
transform 1 0 55065 0 1 18746
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_10
timestamp 1644511149
transform 1 0 55065 0 1 18506
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_11
timestamp 1644511149
transform 1 0 55065 0 1 17956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_12
timestamp 1644511149
transform 1 0 55065 0 1 17716
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_13
timestamp 1644511149
transform 1 0 55065 0 1 17166
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_14
timestamp 1644511149
transform 1 0 55065 0 1 22456
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_15
timestamp 1644511149
transform 1 0 55065 0 1 21906
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_16
timestamp 1644511149
transform 1 0 55065 0 1 21666
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_17
timestamp 1644511149
transform 1 0 55065 0 1 21116
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_18
timestamp 1644511149
transform 1 0 55065 0 1 20876
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_19
timestamp 1644511149
transform 1 0 55065 0 1 20326
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_20
timestamp 1644511149
transform 1 0 55065 0 1 20086
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_21
timestamp 1644511149
transform 1 0 55065 0 1 22696
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_22
timestamp 1644511149
transform 1 0 55065 0 1 39046
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_23
timestamp 1644511149
transform 1 0 55065 0 1 38496
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_24
timestamp 1644511149
transform 1 0 55065 0 1 38256
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_25
timestamp 1644511149
transform 1 0 55065 0 1 37706
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_26
timestamp 1644511149
transform 1 0 55065 0 1 37466
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_27
timestamp 1644511149
transform 1 0 55065 0 1 36916
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_28
timestamp 1644511149
transform 1 0 55065 0 1 36676
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_29
timestamp 1644511149
transform 1 0 55065 0 1 36126
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_30
timestamp 1644511149
transform 1 0 55065 0 1 35886
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_31
timestamp 1644511149
transform 1 0 55065 0 1 35336
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_32
timestamp 1644511149
transform 1 0 55065 0 1 35096
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_33
timestamp 1644511149
transform 1 0 55065 0 1 34546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_34
timestamp 1644511149
transform 1 0 55065 0 1 34306
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_35
timestamp 1644511149
transform 1 0 55065 0 1 33756
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_36
timestamp 1644511149
transform 1 0 55065 0 1 33516
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_37
timestamp 1644511149
transform 1 0 55065 0 1 32966
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_38
timestamp 1644511149
transform 1 0 55065 0 1 32726
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_39
timestamp 1644511149
transform 1 0 55065 0 1 32176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_40
timestamp 1644511149
transform 1 0 55065 0 1 31936
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_41
timestamp 1644511149
transform 1 0 55065 0 1 31386
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_42
timestamp 1644511149
transform 1 0 55065 0 1 31146
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_43
timestamp 1644511149
transform 1 0 55065 0 1 30596
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_44
timestamp 1644511149
transform 1 0 55065 0 1 30356
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_45
timestamp 1644511149
transform 1 0 55065 0 1 29806
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_46
timestamp 1644511149
transform 1 0 55065 0 1 29566
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_47
timestamp 1644511149
transform 1 0 55065 0 1 29016
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_48
timestamp 1644511149
transform 1 0 55065 0 1 28776
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_49
timestamp 1644511149
transform 1 0 55065 0 1 28226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_50
timestamp 1644511149
transform 1 0 55065 0 1 27986
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_51
timestamp 1644511149
transform 1 0 55065 0 1 27436
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_52
timestamp 1644511149
transform 1 0 55065 0 1 27196
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_53
timestamp 1644511149
transform 1 0 55065 0 1 26646
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_54
timestamp 1644511149
transform 1 0 55065 0 1 26406
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_55
timestamp 1644511149
transform 1 0 55065 0 1 25856
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_56
timestamp 1644511149
transform 1 0 55065 0 1 25616
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_57
timestamp 1644511149
transform 1 0 55065 0 1 25066
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_58
timestamp 1644511149
transform 1 0 55065 0 1 24826
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_59
timestamp 1644511149
transform 1 0 55065 0 1 24276
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_60
timestamp 1644511149
transform 1 0 55065 0 1 24036
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_61
timestamp 1644511149
transform 1 0 55065 0 1 23486
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_62
timestamp 1644511149
transform 1 0 55065 0 1 23246
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_63
timestamp 1644511149
transform 1 0 55065 0 1 19536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_64
timestamp 1644511149
transform 1 0 6837 0 1 9169
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_65
timestamp 1644511149
transform 1 0 6837 0 1 7831
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_66
timestamp 1644511149
transform 1 0 6837 0 1 6341
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_67
timestamp 1644511149
transform 1 0 6837 0 1 5003
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_68
timestamp 1644511149
transform 1 0 6837 0 1 3513
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_69
timestamp 1644511149
transform 1 0 6837 0 1 2175
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_70
timestamp 1644511149
transform 1 0 6837 0 1 10659
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_71
timestamp 1644511149
transform 1 0 6837 0 1 685
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_72
timestamp 1644511149
transform 1 0 12127 0 1 13766
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_73
timestamp 1644511149
transform 1 0 12127 0 1 18746
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_74
timestamp 1644511149
transform 1 0 12127 0 1 18506
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_75
timestamp 1644511149
transform 1 0 12127 0 1 17956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_76
timestamp 1644511149
transform 1 0 12127 0 1 17716
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_77
timestamp 1644511149
transform 1 0 12127 0 1 17166
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_78
timestamp 1644511149
transform 1 0 12127 0 1 16926
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_79
timestamp 1644511149
transform 1 0 12127 0 1 16376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_80
timestamp 1644511149
transform 1 0 12127 0 1 16136
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_81
timestamp 1644511149
transform 1 0 12127 0 1 15586
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_82
timestamp 1644511149
transform 1 0 12127 0 1 15346
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_83
timestamp 1644511149
transform 1 0 12127 0 1 14796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_84
timestamp 1644511149
transform 1 0 12127 0 1 14556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_85
timestamp 1644511149
transform 1 0 12127 0 1 14006
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_86
timestamp 1644511149
transform 1 0 12127 0 1 19296
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_87
timestamp 1644511149
transform 1 0 12127 0 1 38496
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_88
timestamp 1644511149
transform 1 0 12127 0 1 38256
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_89
timestamp 1644511149
transform 1 0 12127 0 1 37706
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_90
timestamp 1644511149
transform 1 0 12127 0 1 37466
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_91
timestamp 1644511149
transform 1 0 12127 0 1 36916
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_92
timestamp 1644511149
transform 1 0 12127 0 1 36676
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_93
timestamp 1644511149
transform 1 0 12127 0 1 36126
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_94
timestamp 1644511149
transform 1 0 12127 0 1 35886
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_95
timestamp 1644511149
transform 1 0 12127 0 1 35336
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_96
timestamp 1644511149
transform 1 0 12127 0 1 35096
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_97
timestamp 1644511149
transform 1 0 12127 0 1 34546
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_98
timestamp 1644511149
transform 1 0 12127 0 1 34306
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_99
timestamp 1644511149
transform 1 0 12127 0 1 33756
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_100
timestamp 1644511149
transform 1 0 12127 0 1 33516
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_101
timestamp 1644511149
transform 1 0 12127 0 1 32966
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_102
timestamp 1644511149
transform 1 0 12127 0 1 32726
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_103
timestamp 1644511149
transform 1 0 12127 0 1 32176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_104
timestamp 1644511149
transform 1 0 12127 0 1 31936
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_105
timestamp 1644511149
transform 1 0 12127 0 1 31386
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_106
timestamp 1644511149
transform 1 0 12127 0 1 31146
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_107
timestamp 1644511149
transform 1 0 12127 0 1 30596
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_108
timestamp 1644511149
transform 1 0 12127 0 1 30356
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_109
timestamp 1644511149
transform 1 0 12127 0 1 29806
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_110
timestamp 1644511149
transform 1 0 12127 0 1 29566
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_111
timestamp 1644511149
transform 1 0 12127 0 1 29016
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_112
timestamp 1644511149
transform 1 0 12127 0 1 28776
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_113
timestamp 1644511149
transform 1 0 12127 0 1 28226
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_114
timestamp 1644511149
transform 1 0 12127 0 1 27986
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_115
timestamp 1644511149
transform 1 0 12127 0 1 27436
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_116
timestamp 1644511149
transform 1 0 12127 0 1 27196
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_117
timestamp 1644511149
transform 1 0 12127 0 1 26646
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_118
timestamp 1644511149
transform 1 0 12127 0 1 26406
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_119
timestamp 1644511149
transform 1 0 12127 0 1 25856
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_120
timestamp 1644511149
transform 1 0 12127 0 1 25616
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_121
timestamp 1644511149
transform 1 0 12127 0 1 25066
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_122
timestamp 1644511149
transform 1 0 12127 0 1 24826
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_123
timestamp 1644511149
transform 1 0 12127 0 1 24276
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_124
timestamp 1644511149
transform 1 0 12127 0 1 24036
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_125
timestamp 1644511149
transform 1 0 12127 0 1 23486
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_126
timestamp 1644511149
transform 1 0 12127 0 1 23246
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_127
timestamp 1644511149
transform 1 0 12127 0 1 22696
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_128
timestamp 1644511149
transform 1 0 12127 0 1 22456
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_129
timestamp 1644511149
transform 1 0 12127 0 1 21906
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_130
timestamp 1644511149
transform 1 0 12127 0 1 21666
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_131
timestamp 1644511149
transform 1 0 12127 0 1 21116
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_132
timestamp 1644511149
transform 1 0 12127 0 1 20876
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_133
timestamp 1644511149
transform 1 0 12127 0 1 20326
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_134
timestamp 1644511149
transform 1 0 12127 0 1 20086
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_135
timestamp 1644511149
transform 1 0 12127 0 1 39046
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_136
timestamp 1644511149
transform 1 0 12127 0 1 19536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_137
timestamp 1644511149
transform 1 0 12127 0 1 47976
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_138
timestamp 1644511149
transform 1 0 12127 0 1 47736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_139
timestamp 1644511149
transform 1 0 12127 0 1 47186
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_140
timestamp 1644511149
transform 1 0 12127 0 1 46946
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_141
timestamp 1644511149
transform 1 0 12127 0 1 46396
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_142
timestamp 1644511149
transform 1 0 12127 0 1 46156
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_143
timestamp 1644511149
transform 1 0 12127 0 1 45606
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_144
timestamp 1644511149
transform 1 0 12127 0 1 45366
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_145
timestamp 1644511149
transform 1 0 12127 0 1 44816
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_146
timestamp 1644511149
transform 1 0 12127 0 1 44576
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_147
timestamp 1644511149
transform 1 0 12127 0 1 44026
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_148
timestamp 1644511149
transform 1 0 12127 0 1 43786
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_149
timestamp 1644511149
transform 1 0 12127 0 1 43236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_150
timestamp 1644511149
transform 1 0 12127 0 1 42996
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_151
timestamp 1644511149
transform 1 0 12127 0 1 42446
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_152
timestamp 1644511149
transform 1 0 12127 0 1 42206
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_153
timestamp 1644511149
transform 1 0 12127 0 1 41656
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_154
timestamp 1644511149
transform 1 0 12127 0 1 41416
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_155
timestamp 1644511149
transform 1 0 12127 0 1 40866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_156
timestamp 1644511149
transform 1 0 12127 0 1 40626
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_157
timestamp 1644511149
transform 1 0 12127 0 1 40076
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_158
timestamp 1644511149
transform 1 0 12127 0 1 39836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_159
timestamp 1644511149
transform 1 0 12127 0 1 39286
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_160
timestamp 1644511149
transform 1 0 12127 0 1 54056
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_161
timestamp 1644511149
transform 1 0 12127 0 1 53506
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_162
timestamp 1644511149
transform 1 0 12127 0 1 53266
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_163
timestamp 1644511149
transform 1 0 12127 0 1 52716
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_164
timestamp 1644511149
transform 1 0 12127 0 1 52476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_165
timestamp 1644511149
transform 1 0 12127 0 1 51926
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_166
timestamp 1644511149
transform 1 0 12127 0 1 51686
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_167
timestamp 1644511149
transform 1 0 12127 0 1 51136
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_168
timestamp 1644511149
transform 1 0 12127 0 1 50896
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_169
timestamp 1644511149
transform 1 0 12127 0 1 50346
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_170
timestamp 1644511149
transform 1 0 12127 0 1 50106
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_171
timestamp 1644511149
transform 1 0 12127 0 1 49556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_172
timestamp 1644511149
transform 1 0 12127 0 1 49316
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_173
timestamp 1644511149
transform 1 0 12127 0 1 48766
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_174
timestamp 1644511149
transform 1 0 12127 0 1 48526
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_175
timestamp 1644511149
transform 1 0 12127 0 1 58246
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_176
timestamp 1644511149
transform 1 0 12127 0 1 58006
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_177
timestamp 1644511149
transform 1 0 12127 0 1 57456
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_178
timestamp 1644511149
transform 1 0 12127 0 1 57216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_179
timestamp 1644511149
transform 1 0 12127 0 1 56666
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_180
timestamp 1644511149
transform 1 0 12127 0 1 56426
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_181
timestamp 1644511149
transform 1 0 12127 0 1 55876
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_182
timestamp 1644511149
transform 1 0 12127 0 1 55636
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_183
timestamp 1644511149
transform 1 0 12127 0 1 55086
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_184
timestamp 1644511149
transform 1 0 12127 0 1 54846
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_185
timestamp 1644511149
transform 1 0 12127 0 1 54296
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_186
timestamp 1644511149
transform 1 0 12127 0 1 64326
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_187
timestamp 1644511149
transform 1 0 12127 0 1 63776
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_188
timestamp 1644511149
transform 1 0 12127 0 1 63536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_189
timestamp 1644511149
transform 1 0 12127 0 1 62986
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_190
timestamp 1644511149
transform 1 0 12127 0 1 62746
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_191
timestamp 1644511149
transform 1 0 12127 0 1 62196
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_192
timestamp 1644511149
transform 1 0 12127 0 1 61956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_193
timestamp 1644511149
transform 1 0 12127 0 1 61406
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_194
timestamp 1644511149
transform 1 0 12127 0 1 61166
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_195
timestamp 1644511149
transform 1 0 12127 0 1 60616
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_196
timestamp 1644511149
transform 1 0 12127 0 1 60376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_197
timestamp 1644511149
transform 1 0 12127 0 1 59826
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_198
timestamp 1644511149
transform 1 0 12127 0 1 59586
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_199
timestamp 1644511149
transform 1 0 12127 0 1 59036
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_200
timestamp 1644511149
transform 1 0 12127 0 1 58796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_201
timestamp 1644511149
transform 1 0 55065 0 1 53506
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_202
timestamp 1644511149
transform 1 0 55065 0 1 53266
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_203
timestamp 1644511149
transform 1 0 55065 0 1 52716
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_204
timestamp 1644511149
transform 1 0 55065 0 1 52476
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_205
timestamp 1644511149
transform 1 0 55065 0 1 51926
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_206
timestamp 1644511149
transform 1 0 55065 0 1 51686
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_207
timestamp 1644511149
transform 1 0 55065 0 1 51136
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_208
timestamp 1644511149
transform 1 0 55065 0 1 50896
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_209
timestamp 1644511149
transform 1 0 55065 0 1 50346
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_210
timestamp 1644511149
transform 1 0 55065 0 1 50106
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_211
timestamp 1644511149
transform 1 0 55065 0 1 49556
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_212
timestamp 1644511149
transform 1 0 55065 0 1 49316
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_213
timestamp 1644511149
transform 1 0 55065 0 1 48766
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_214
timestamp 1644511149
transform 1 0 55065 0 1 48526
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_215
timestamp 1644511149
transform 1 0 55065 0 1 47976
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_216
timestamp 1644511149
transform 1 0 55065 0 1 47736
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_217
timestamp 1644511149
transform 1 0 55065 0 1 47186
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_218
timestamp 1644511149
transform 1 0 55065 0 1 46946
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_219
timestamp 1644511149
transform 1 0 55065 0 1 46396
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_220
timestamp 1644511149
transform 1 0 55065 0 1 46156
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_221
timestamp 1644511149
transform 1 0 55065 0 1 45606
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_222
timestamp 1644511149
transform 1 0 55065 0 1 45366
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_223
timestamp 1644511149
transform 1 0 55065 0 1 44816
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_224
timestamp 1644511149
transform 1 0 55065 0 1 44576
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_225
timestamp 1644511149
transform 1 0 55065 0 1 44026
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_226
timestamp 1644511149
transform 1 0 55065 0 1 43786
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_227
timestamp 1644511149
transform 1 0 55065 0 1 43236
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_228
timestamp 1644511149
transform 1 0 55065 0 1 42996
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_229
timestamp 1644511149
transform 1 0 55065 0 1 42446
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_230
timestamp 1644511149
transform 1 0 55065 0 1 42206
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_231
timestamp 1644511149
transform 1 0 55065 0 1 41656
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_232
timestamp 1644511149
transform 1 0 55065 0 1 41416
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_233
timestamp 1644511149
transform 1 0 55065 0 1 40866
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_234
timestamp 1644511149
transform 1 0 55065 0 1 40626
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_235
timestamp 1644511149
transform 1 0 55065 0 1 40076
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_236
timestamp 1644511149
transform 1 0 55065 0 1 39836
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_237
timestamp 1644511149
transform 1 0 55065 0 1 39286
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_238
timestamp 1644511149
transform 1 0 55065 0 1 58246
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_239
timestamp 1644511149
transform 1 0 55065 0 1 58006
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_240
timestamp 1644511149
transform 1 0 55065 0 1 57456
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_241
timestamp 1644511149
transform 1 0 55065 0 1 57216
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_242
timestamp 1644511149
transform 1 0 55065 0 1 56666
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_243
timestamp 1644511149
transform 1 0 55065 0 1 56426
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_244
timestamp 1644511149
transform 1 0 55065 0 1 55876
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_245
timestamp 1644511149
transform 1 0 55065 0 1 55636
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_246
timestamp 1644511149
transform 1 0 55065 0 1 55086
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_247
timestamp 1644511149
transform 1 0 55065 0 1 54846
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_248
timestamp 1644511149
transform 1 0 55065 0 1 54296
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_249
timestamp 1644511149
transform 1 0 55065 0 1 54056
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_250
timestamp 1644511149
transform 1 0 60231 0 1 77647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_251
timestamp 1644511149
transform 1 0 60231 0 1 76157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_252
timestamp 1644511149
transform 1 0 60231 0 1 74819
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_253
timestamp 1644511149
transform 1 0 60231 0 1 73329
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_254
timestamp 1644511149
transform 1 0 60231 0 1 71991
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_255
timestamp 1644511149
transform 1 0 60231 0 1 69163
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_256
timestamp 1644511149
transform 1 0 60231 0 1 70501
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_257
timestamp 1644511149
transform 1 0 60231 0 1 67673
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_258
timestamp 1644511149
transform 1 0 55065 0 1 64566
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_259
timestamp 1644511149
transform 1 0 55065 0 1 64326
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_260
timestamp 1644511149
transform 1 0 55065 0 1 63776
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_261
timestamp 1644511149
transform 1 0 55065 0 1 63536
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_262
timestamp 1644511149
transform 1 0 55065 0 1 62986
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_263
timestamp 1644511149
transform 1 0 55065 0 1 62746
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_264
timestamp 1644511149
transform 1 0 55065 0 1 62196
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_265
timestamp 1644511149
transform 1 0 55065 0 1 61956
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_266
timestamp 1644511149
transform 1 0 55065 0 1 61406
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_267
timestamp 1644511149
transform 1 0 55065 0 1 61166
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_268
timestamp 1644511149
transform 1 0 55065 0 1 60616
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_269
timestamp 1644511149
transform 1 0 55065 0 1 60376
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_270
timestamp 1644511149
transform 1 0 55065 0 1 59826
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_271
timestamp 1644511149
transform 1 0 55065 0 1 59586
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_272
timestamp 1644511149
transform 1 0 55065 0 1 59036
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_14_273
timestamp 1644511149
transform 1 0 55065 0 1 58796
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_0
timestamp 1644511149
transform 1 0 55062 0 1 16927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_1
timestamp 1644511149
transform 1 0 55062 0 1 16377
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_2
timestamp 1644511149
transform 1 0 55062 0 1 16137
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_3
timestamp 1644511149
transform 1 0 55062 0 1 15587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_4
timestamp 1644511149
transform 1 0 55062 0 1 15347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_5
timestamp 1644511149
transform 1 0 55062 0 1 14797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_6
timestamp 1644511149
transform 1 0 55062 0 1 14557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_7
timestamp 1644511149
transform 1 0 55062 0 1 14007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_8
timestamp 1644511149
transform 1 0 55062 0 1 19297
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_9
timestamp 1644511149
transform 1 0 55062 0 1 18747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_10
timestamp 1644511149
transform 1 0 55062 0 1 18507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_11
timestamp 1644511149
transform 1 0 55062 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_12
timestamp 1644511149
transform 1 0 55062 0 1 17717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_13
timestamp 1644511149
transform 1 0 55062 0 1 17167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_14
timestamp 1644511149
transform 1 0 55062 0 1 22457
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_15
timestamp 1644511149
transform 1 0 55062 0 1 21907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_16
timestamp 1644511149
transform 1 0 55062 0 1 21667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_17
timestamp 1644511149
transform 1 0 55062 0 1 21117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_18
timestamp 1644511149
transform 1 0 55062 0 1 20877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_19
timestamp 1644511149
transform 1 0 55062 0 1 20327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_20
timestamp 1644511149
transform 1 0 55062 0 1 20087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_21
timestamp 1644511149
transform 1 0 55062 0 1 22697
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_22
timestamp 1644511149
transform 1 0 55062 0 1 39047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_23
timestamp 1644511149
transform 1 0 55062 0 1 38497
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_24
timestamp 1644511149
transform 1 0 55062 0 1 38257
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_25
timestamp 1644511149
transform 1 0 55062 0 1 37707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_26
timestamp 1644511149
transform 1 0 55062 0 1 37467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_27
timestamp 1644511149
transform 1 0 55062 0 1 36917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_28
timestamp 1644511149
transform 1 0 55062 0 1 36677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_29
timestamp 1644511149
transform 1 0 55062 0 1 36127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_30
timestamp 1644511149
transform 1 0 55062 0 1 35887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_31
timestamp 1644511149
transform 1 0 55062 0 1 35337
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_32
timestamp 1644511149
transform 1 0 55062 0 1 35097
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_33
timestamp 1644511149
transform 1 0 55062 0 1 34547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_34
timestamp 1644511149
transform 1 0 55062 0 1 34307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_35
timestamp 1644511149
transform 1 0 55062 0 1 33757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_36
timestamp 1644511149
transform 1 0 55062 0 1 33517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_37
timestamp 1644511149
transform 1 0 55062 0 1 32967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_38
timestamp 1644511149
transform 1 0 55062 0 1 32727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_39
timestamp 1644511149
transform 1 0 55062 0 1 32177
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_40
timestamp 1644511149
transform 1 0 55062 0 1 31937
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_41
timestamp 1644511149
transform 1 0 55062 0 1 31387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_42
timestamp 1644511149
transform 1 0 55062 0 1 31147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_43
timestamp 1644511149
transform 1 0 55062 0 1 30597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_44
timestamp 1644511149
transform 1 0 55062 0 1 30357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_45
timestamp 1644511149
transform 1 0 55062 0 1 29807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_46
timestamp 1644511149
transform 1 0 55062 0 1 29567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_47
timestamp 1644511149
transform 1 0 55062 0 1 29017
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_48
timestamp 1644511149
transform 1 0 55062 0 1 28777
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_49
timestamp 1644511149
transform 1 0 55062 0 1 28227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_50
timestamp 1644511149
transform 1 0 55062 0 1 27987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_51
timestamp 1644511149
transform 1 0 55062 0 1 27437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_52
timestamp 1644511149
transform 1 0 55062 0 1 27197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_53
timestamp 1644511149
transform 1 0 55062 0 1 26647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_54
timestamp 1644511149
transform 1 0 55062 0 1 26407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_55
timestamp 1644511149
transform 1 0 55062 0 1 25857
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_56
timestamp 1644511149
transform 1 0 55062 0 1 25617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_57
timestamp 1644511149
transform 1 0 55062 0 1 25067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_58
timestamp 1644511149
transform 1 0 55062 0 1 24827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_59
timestamp 1644511149
transform 1 0 55062 0 1 24277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_60
timestamp 1644511149
transform 1 0 55062 0 1 24037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_61
timestamp 1644511149
transform 1 0 55062 0 1 23487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_62
timestamp 1644511149
transform 1 0 55062 0 1 23247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_63
timestamp 1644511149
transform 1 0 55062 0 1 19537
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_64
timestamp 1644511149
transform 1 0 6834 0 1 9170
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_65
timestamp 1644511149
transform 1 0 6834 0 1 7832
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_66
timestamp 1644511149
transform 1 0 6834 0 1 6342
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_67
timestamp 1644511149
transform 1 0 6834 0 1 5004
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_68
timestamp 1644511149
transform 1 0 6834 0 1 3514
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_69
timestamp 1644511149
transform 1 0 6834 0 1 2176
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_70
timestamp 1644511149
transform 1 0 6834 0 1 10660
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_71
timestamp 1644511149
transform 1 0 6834 0 1 686
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_72
timestamp 1644511149
transform 1 0 12124 0 1 13767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_73
timestamp 1644511149
transform 1 0 12124 0 1 18747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_74
timestamp 1644511149
transform 1 0 12124 0 1 18507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_75
timestamp 1644511149
transform 1 0 12124 0 1 17957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_76
timestamp 1644511149
transform 1 0 12124 0 1 17717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_77
timestamp 1644511149
transform 1 0 12124 0 1 17167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_78
timestamp 1644511149
transform 1 0 12124 0 1 16927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_79
timestamp 1644511149
transform 1 0 12124 0 1 16377
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_80
timestamp 1644511149
transform 1 0 12124 0 1 16137
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_81
timestamp 1644511149
transform 1 0 12124 0 1 15587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_82
timestamp 1644511149
transform 1 0 12124 0 1 15347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_83
timestamp 1644511149
transform 1 0 12124 0 1 14797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_84
timestamp 1644511149
transform 1 0 12124 0 1 14557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_85
timestamp 1644511149
transform 1 0 12124 0 1 14007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_86
timestamp 1644511149
transform 1 0 13545 0 1 11967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_87
timestamp 1644511149
transform 1 0 12124 0 1 19297
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_88
timestamp 1644511149
transform 1 0 12124 0 1 38257
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_89
timestamp 1644511149
transform 1 0 12124 0 1 37707
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_90
timestamp 1644511149
transform 1 0 12124 0 1 37467
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_91
timestamp 1644511149
transform 1 0 12124 0 1 36917
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_92
timestamp 1644511149
transform 1 0 12124 0 1 36677
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_93
timestamp 1644511149
transform 1 0 12124 0 1 36127
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_94
timestamp 1644511149
transform 1 0 12124 0 1 35887
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_95
timestamp 1644511149
transform 1 0 12124 0 1 35337
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_96
timestamp 1644511149
transform 1 0 12124 0 1 35097
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_97
timestamp 1644511149
transform 1 0 12124 0 1 34547
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_98
timestamp 1644511149
transform 1 0 12124 0 1 34307
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_99
timestamp 1644511149
transform 1 0 12124 0 1 33757
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_100
timestamp 1644511149
transform 1 0 12124 0 1 33517
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_101
timestamp 1644511149
transform 1 0 12124 0 1 32967
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_102
timestamp 1644511149
transform 1 0 12124 0 1 32727
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_103
timestamp 1644511149
transform 1 0 12124 0 1 32177
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_104
timestamp 1644511149
transform 1 0 12124 0 1 31937
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_105
timestamp 1644511149
transform 1 0 12124 0 1 31387
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_106
timestamp 1644511149
transform 1 0 12124 0 1 31147
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_107
timestamp 1644511149
transform 1 0 12124 0 1 30597
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_108
timestamp 1644511149
transform 1 0 12124 0 1 30357
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_109
timestamp 1644511149
transform 1 0 12124 0 1 29807
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_110
timestamp 1644511149
transform 1 0 12124 0 1 29567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_111
timestamp 1644511149
transform 1 0 12124 0 1 29017
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_112
timestamp 1644511149
transform 1 0 12124 0 1 28777
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_113
timestamp 1644511149
transform 1 0 12124 0 1 28227
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_114
timestamp 1644511149
transform 1 0 12124 0 1 27987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_115
timestamp 1644511149
transform 1 0 12124 0 1 27437
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_116
timestamp 1644511149
transform 1 0 12124 0 1 27197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_117
timestamp 1644511149
transform 1 0 12124 0 1 26647
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_118
timestamp 1644511149
transform 1 0 12124 0 1 26407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_119
timestamp 1644511149
transform 1 0 12124 0 1 25857
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_120
timestamp 1644511149
transform 1 0 12124 0 1 25617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_121
timestamp 1644511149
transform 1 0 12124 0 1 25067
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_122
timestamp 1644511149
transform 1 0 12124 0 1 24827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_123
timestamp 1644511149
transform 1 0 12124 0 1 24277
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_124
timestamp 1644511149
transform 1 0 12124 0 1 24037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_125
timestamp 1644511149
transform 1 0 12124 0 1 23487
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_126
timestamp 1644511149
transform 1 0 12124 0 1 23247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_127
timestamp 1644511149
transform 1 0 12124 0 1 22697
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_128
timestamp 1644511149
transform 1 0 12124 0 1 22457
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_129
timestamp 1644511149
transform 1 0 12124 0 1 21907
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_130
timestamp 1644511149
transform 1 0 12124 0 1 21667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_131
timestamp 1644511149
transform 1 0 12124 0 1 21117
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_132
timestamp 1644511149
transform 1 0 12124 0 1 20877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_133
timestamp 1644511149
transform 1 0 12124 0 1 20327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_134
timestamp 1644511149
transform 1 0 12124 0 1 20087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_135
timestamp 1644511149
transform 1 0 12124 0 1 38497
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_136
timestamp 1644511149
transform 1 0 12124 0 1 39047
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_137
timestamp 1644511149
transform 1 0 12124 0 1 19537
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_138
timestamp 1644511149
transform 1 0 12124 0 1 47977
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_139
timestamp 1644511149
transform 1 0 12124 0 1 47737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_140
timestamp 1644511149
transform 1 0 12124 0 1 47187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_141
timestamp 1644511149
transform 1 0 12124 0 1 46947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_142
timestamp 1644511149
transform 1 0 12124 0 1 46397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_143
timestamp 1644511149
transform 1 0 12124 0 1 46157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_144
timestamp 1644511149
transform 1 0 12124 0 1 45607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_145
timestamp 1644511149
transform 1 0 12124 0 1 45367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_146
timestamp 1644511149
transform 1 0 12124 0 1 44817
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_147
timestamp 1644511149
transform 1 0 12124 0 1 44577
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_148
timestamp 1644511149
transform 1 0 12124 0 1 44027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_149
timestamp 1644511149
transform 1 0 12124 0 1 43787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_150
timestamp 1644511149
transform 1 0 12124 0 1 43237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_151
timestamp 1644511149
transform 1 0 12124 0 1 42997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_152
timestamp 1644511149
transform 1 0 12124 0 1 42447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_153
timestamp 1644511149
transform 1 0 12124 0 1 42207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_154
timestamp 1644511149
transform 1 0 12124 0 1 41657
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_155
timestamp 1644511149
transform 1 0 12124 0 1 41417
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_156
timestamp 1644511149
transform 1 0 12124 0 1 40867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_157
timestamp 1644511149
transform 1 0 12124 0 1 40627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_158
timestamp 1644511149
transform 1 0 12124 0 1 40077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_159
timestamp 1644511149
transform 1 0 12124 0 1 39837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_160
timestamp 1644511149
transform 1 0 12124 0 1 39287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_161
timestamp 1644511149
transform 1 0 12124 0 1 54057
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_162
timestamp 1644511149
transform 1 0 12124 0 1 53507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_163
timestamp 1644511149
transform 1 0 12124 0 1 53267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_164
timestamp 1644511149
transform 1 0 12124 0 1 52717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_165
timestamp 1644511149
transform 1 0 12124 0 1 52477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_166
timestamp 1644511149
transform 1 0 12124 0 1 51927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_167
timestamp 1644511149
transform 1 0 12124 0 1 51687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_168
timestamp 1644511149
transform 1 0 12124 0 1 51137
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_169
timestamp 1644511149
transform 1 0 12124 0 1 50897
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_170
timestamp 1644511149
transform 1 0 12124 0 1 50347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_171
timestamp 1644511149
transform 1 0 12124 0 1 50107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_172
timestamp 1644511149
transform 1 0 12124 0 1 49557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_173
timestamp 1644511149
transform 1 0 12124 0 1 49317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_174
timestamp 1644511149
transform 1 0 12124 0 1 48767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_175
timestamp 1644511149
transform 1 0 12124 0 1 48527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_176
timestamp 1644511149
transform 1 0 12124 0 1 58247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_177
timestamp 1644511149
transform 1 0 12124 0 1 58007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_178
timestamp 1644511149
transform 1 0 12124 0 1 57457
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_179
timestamp 1644511149
transform 1 0 12124 0 1 57217
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_180
timestamp 1644511149
transform 1 0 12124 0 1 56667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_181
timestamp 1644511149
transform 1 0 12124 0 1 56427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_182
timestamp 1644511149
transform 1 0 12124 0 1 55877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_183
timestamp 1644511149
transform 1 0 12124 0 1 55637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_184
timestamp 1644511149
transform 1 0 12124 0 1 55087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_185
timestamp 1644511149
transform 1 0 12124 0 1 54847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_186
timestamp 1644511149
transform 1 0 12124 0 1 54297
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_187
timestamp 1644511149
transform 1 0 12124 0 1 64327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_188
timestamp 1644511149
transform 1 0 12124 0 1 63777
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_189
timestamp 1644511149
transform 1 0 12124 0 1 63537
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_190
timestamp 1644511149
transform 1 0 12124 0 1 62987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_191
timestamp 1644511149
transform 1 0 12124 0 1 62747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_192
timestamp 1644511149
transform 1 0 12124 0 1 62197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_193
timestamp 1644511149
transform 1 0 12124 0 1 61957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_194
timestamp 1644511149
transform 1 0 12124 0 1 61407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_195
timestamp 1644511149
transform 1 0 12124 0 1 61167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_196
timestamp 1644511149
transform 1 0 12124 0 1 60617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_197
timestamp 1644511149
transform 1 0 12124 0 1 60377
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_198
timestamp 1644511149
transform 1 0 12124 0 1 59827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_199
timestamp 1644511149
transform 1 0 12124 0 1 59587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_200
timestamp 1644511149
transform 1 0 12124 0 1 59037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_201
timestamp 1644511149
transform 1 0 12124 0 1 58797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_202
timestamp 1644511149
transform 1 0 55062 0 1 53507
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_203
timestamp 1644511149
transform 1 0 55062 0 1 53267
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_204
timestamp 1644511149
transform 1 0 55062 0 1 52717
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_205
timestamp 1644511149
transform 1 0 55062 0 1 52477
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_206
timestamp 1644511149
transform 1 0 55062 0 1 51927
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_207
timestamp 1644511149
transform 1 0 55062 0 1 51687
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_208
timestamp 1644511149
transform 1 0 55062 0 1 51137
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_209
timestamp 1644511149
transform 1 0 55062 0 1 50897
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_210
timestamp 1644511149
transform 1 0 55062 0 1 50347
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_211
timestamp 1644511149
transform 1 0 55062 0 1 50107
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_212
timestamp 1644511149
transform 1 0 55062 0 1 49557
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_213
timestamp 1644511149
transform 1 0 55062 0 1 49317
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_214
timestamp 1644511149
transform 1 0 55062 0 1 48767
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_215
timestamp 1644511149
transform 1 0 55062 0 1 48527
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_216
timestamp 1644511149
transform 1 0 55062 0 1 47977
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_217
timestamp 1644511149
transform 1 0 55062 0 1 47737
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_218
timestamp 1644511149
transform 1 0 55062 0 1 47187
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_219
timestamp 1644511149
transform 1 0 55062 0 1 46947
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_220
timestamp 1644511149
transform 1 0 55062 0 1 46397
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_221
timestamp 1644511149
transform 1 0 55062 0 1 46157
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_222
timestamp 1644511149
transform 1 0 55062 0 1 45607
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_223
timestamp 1644511149
transform 1 0 55062 0 1 45367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_224
timestamp 1644511149
transform 1 0 55062 0 1 44817
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_225
timestamp 1644511149
transform 1 0 55062 0 1 44577
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_226
timestamp 1644511149
transform 1 0 55062 0 1 44027
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_227
timestamp 1644511149
transform 1 0 55062 0 1 43787
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_228
timestamp 1644511149
transform 1 0 55062 0 1 43237
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_229
timestamp 1644511149
transform 1 0 55062 0 1 42997
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_230
timestamp 1644511149
transform 1 0 55062 0 1 42447
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_231
timestamp 1644511149
transform 1 0 55062 0 1 42207
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_232
timestamp 1644511149
transform 1 0 55062 0 1 41657
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_233
timestamp 1644511149
transform 1 0 55062 0 1 41417
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_234
timestamp 1644511149
transform 1 0 55062 0 1 40867
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_235
timestamp 1644511149
transform 1 0 55062 0 1 40627
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_236
timestamp 1644511149
transform 1 0 55062 0 1 40077
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_237
timestamp 1644511149
transform 1 0 55062 0 1 39837
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_238
timestamp 1644511149
transform 1 0 55062 0 1 39287
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_239
timestamp 1644511149
transform 1 0 55062 0 1 58247
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_240
timestamp 1644511149
transform 1 0 55062 0 1 58007
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_241
timestamp 1644511149
transform 1 0 55062 0 1 57457
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_242
timestamp 1644511149
transform 1 0 55062 0 1 57217
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_243
timestamp 1644511149
transform 1 0 55062 0 1 56667
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_244
timestamp 1644511149
transform 1 0 55062 0 1 56427
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_245
timestamp 1644511149
transform 1 0 55062 0 1 55877
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_246
timestamp 1644511149
transform 1 0 55062 0 1 55637
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_247
timestamp 1644511149
transform 1 0 55062 0 1 55087
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_248
timestamp 1644511149
transform 1 0 55062 0 1 54847
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_249
timestamp 1644511149
transform 1 0 55062 0 1 54297
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_250
timestamp 1644511149
transform 1 0 55062 0 1 54057
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_251
timestamp 1644511149
transform 1 0 60228 0 1 77648
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_252
timestamp 1644511149
transform 1 0 60228 0 1 76158
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_253
timestamp 1644511149
transform 1 0 60228 0 1 74820
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_254
timestamp 1644511149
transform 1 0 60228 0 1 73330
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_255
timestamp 1644511149
transform 1 0 60228 0 1 71992
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_256
timestamp 1644511149
transform 1 0 60228 0 1 69164
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_257
timestamp 1644511149
transform 1 0 60228 0 1 70502
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_258
timestamp 1644511149
transform 1 0 60228 0 1 67674
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_259
timestamp 1644511149
transform 1 0 55062 0 1 64567
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_260
timestamp 1644511149
transform 1 0 55062 0 1 64327
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_261
timestamp 1644511149
transform 1 0 55062 0 1 63777
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_262
timestamp 1644511149
transform 1 0 55062 0 1 63537
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_263
timestamp 1644511149
transform 1 0 55062 0 1 62987
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_264
timestamp 1644511149
transform 1 0 55062 0 1 62747
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_265
timestamp 1644511149
transform 1 0 55062 0 1 62197
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_266
timestamp 1644511149
transform 1 0 55062 0 1 61957
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_267
timestamp 1644511149
transform 1 0 55062 0 1 61407
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_268
timestamp 1644511149
transform 1 0 55062 0 1 61167
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_269
timestamp 1644511149
transform 1 0 55062 0 1 60617
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_270
timestamp 1644511149
transform 1 0 55062 0 1 60377
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_271
timestamp 1644511149
transform 1 0 55062 0 1 59827
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_272
timestamp 1644511149
transform 1 0 55062 0 1 59587
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_273
timestamp 1644511149
transform 1 0 55062 0 1 59037
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_274
timestamp 1644511149
transform 1 0 53641 0 1 66367
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19  sky130_sram_1kbyte_1rw1r_8x1024_8_contact_19_275
timestamp 1644511149
transform 1 0 55062 0 1 58797
box 0 0 1 1
use sky130_sram_1kbyte_1rw1r_8x1024_8_hierarchical_predecode3x8_0  sky130_sram_1kbyte_1rw1r_8x1024_8_hierarchical_predecode3x8_0_0
timestamp 1644511149
transform 1 0 4195 0 1 49
box 0 -49 2862 11361
use sky130_sram_1kbyte_1rw1r_8x1024_8_hierarchical_predecode3x8_0  sky130_sram_1kbyte_1rw1r_8x1024_8_hierarchical_predecode3x8_0_1
timestamp 1644511149
transform -1 0 62931 0 -1 78349
box 0 -49 2862 11361
use sky130_sram_1kbyte_1rw1r_8x1024_8_port_address  sky130_sram_1kbyte_1rw1r_8x1024_8_port_address_0
timestamp 1644511149
transform 1 0 0 0 1 13919
box 0 -490 12011 50620
use sky130_sram_1kbyte_1rw1r_8x1024_8_port_address_0  sky130_sram_1kbyte_1rw1r_8x1024_8_port_address_0_0
timestamp 1644511149
transform -1 0 67250 0 1 13919
box 0 -60 12011 51050
use sky130_sram_1kbyte_1rw1r_8x1024_8_port_data  sky130_sram_1kbyte_1rw1r_8x1024_8_port_data_0
timestamp 1644511149
transform 1 0 12283 0 -1 13129
box -49 238 41359 10130
use sky130_sram_1kbyte_1rw1r_8x1024_8_port_data_0  sky130_sram_1kbyte_1rw1r_8x1024_8_port_data_0_0
timestamp 1644511149
transform 1 0 12283 0 1 65269
box 0 238 41934 6446
use sky130_sram_1kbyte_1rw1r_8x1024_8_replica_bitcell_array  sky130_sram_1kbyte_1rw1r_8x1024_8_replica_bitcell_array_0
timestamp 1644511149
transform 1 0 12283 0 1 13129
box -49 0 42733 52140
<< labels >>
rlabel metal3 s 62352 76886 62450 76984 4 vdd
port 1 nsew
rlabel metal3 s 60992 71230 61090 71328 4 vdd
port 1 nsew
rlabel metal3 s 60992 76886 61090 76984 4 vdd
port 1 nsew
rlabel metal3 s 62352 74058 62450 74156 4 vdd
port 1 nsew
rlabel metal3 s 62352 71230 62450 71328 4 vdd
port 1 nsew
rlabel metal3 s 60992 74058 61090 74156 4 vdd
port 1 nsew
rlabel metal3 s 60992 72644 61090 72742 4 gnd
port 2 nsew
rlabel metal3 s 60992 78300 61090 78398 4 gnd
port 2 nsew
rlabel metal3 s 62352 75472 62450 75570 4 gnd
port 2 nsew
rlabel metal3 s 62352 72644 62450 72742 4 gnd
port 2 nsew
rlabel metal3 s 60992 75472 61090 75570 4 gnd
port 2 nsew
rlabel metal3 s 60992 69816 61090 69914 4 gnd
port 2 nsew
rlabel metal3 s 62352 78300 62450 78398 4 gnd
port 2 nsew
rlabel metal3 s 62352 69816 62450 69914 4 gnd
port 2 nsew
rlabel metal3 s 51360 64991 51458 65089 4 vdd
port 1 nsew
rlabel metal3 s 52489 65582 52587 65680 4 vdd
port 1 nsew
rlabel metal3 s 53351 65582 53449 65680 4 vdd
port 1 nsew
rlabel metal3 s 50855 65582 50953 65680 4 vdd
port 1 nsew
rlabel metal3 s 53232 64991 53330 65089 4 vdd
port 1 nsew
rlabel metal3 s 53856 64991 53954 65089 4 vdd
port 1 nsew
rlabel metal3 s 52608 64991 52706 65089 4 vdd
port 1 nsew
rlabel metal3 s 51984 64991 52082 65089 4 vdd
port 1 nsew
rlabel metal3 s 54552 59690 54650 59788 4 gnd
port 2 nsew
rlabel metal3 s 54552 63877 54650 63975 4 gnd
port 2 nsew
rlabel metal3 s 54918 64777 55016 64875 4 gnd
port 2 nsew
rlabel metal3 s 50736 64991 50834 65089 4 vdd
port 1 nsew
rlabel metal3 s 54552 61033 54650 61131 4 gnd
port 2 nsew
rlabel metal3 s 54552 60480 54650 60578 4 gnd
port 2 nsew
rlabel metal3 s 54552 61507 54650 61605 4 gnd
port 2 nsew
rlabel metal3 s 52920 67131 53018 67229 4 gnd
port 2 nsew
rlabel metal3 s 54552 62613 54650 62711 4 gnd
port 2 nsew
rlabel metal3 s 51672 67131 51770 67229 4 gnd
port 2 nsew
rlabel metal3 s 54552 62060 54650 62158 4 gnd
port 2 nsew
rlabel metal3 s 50424 67131 50522 67229 4 gnd
port 2 nsew
rlabel metal3 s 54552 62850 54650 62948 4 gnd
port 2 nsew
rlabel metal3 s 54552 59137 54650 59235 4 gnd
port 2 nsew
rlabel metal3 s 54552 63640 54650 63738 4 gnd
port 2 nsew
rlabel metal3 s 54552 61823 54650 61921 4 gnd
port 2 nsew
rlabel metal3 s 54552 63087 54650 63185 4 gnd
port 2 nsew
rlabel metal3 s 54552 60717 54650 60815 4 gnd
port 2 nsew
rlabel metal3 s 54552 61270 54650 61368 4 gnd
port 2 nsew
rlabel metal3 s 50112 64991 50210 65089 4 vdd
port 1 nsew
rlabel metal3 s 54552 62297 54650 62395 4 gnd
port 2 nsew
rlabel metal3 s 54552 64430 54650 64528 4 gnd
port 2 nsew
rlabel metal3 s 54552 63403 54650 63501 4 gnd
port 2 nsew
rlabel metal3 s 54552 58900 54650 58998 4 gnd
port 2 nsew
rlabel metal3 s 54552 60243 54650 60341 4 gnd
port 2 nsew
rlabel metal3 s 53737 65582 53835 65680 4 vdd
port 1 nsew
rlabel metal3 s 54552 59927 54650 60025 4 gnd
port 2 nsew
rlabel metal3 s 55944 64627 56042 64725 4 vdd
port 1 nsew
rlabel metal3 s 52103 65582 52201 65680 4 vdd
port 1 nsew
rlabel metal3 s 54552 59453 54650 59551 4 gnd
port 2 nsew
rlabel metal3 s 51241 65582 51339 65680 4 vdd
port 1 nsew
rlabel metal3 s 54552 64193 54650 64291 4 gnd
port 2 nsew
rlabel metal3 s 49993 65582 50091 65680 4 vdd
port 1 nsew
rlabel metal3 s 59492 63640 59590 63738 4 vdd
port 1 nsew
rlabel metal3 s 60702 61688 60800 61786 4 vdd
port 1 nsew
rlabel metal3 s 60702 62836 60800 62934 4 vdd
port 1 nsew
rlabel metal3 s 53673 66369 67334 66429 4 rbl_bl_1_1
port 3 nsew
rlabel metal3 s 58635 64615 58733 64713 4 vdd
port 1 nsew
rlabel metal3 s 60992 68402 61090 68500 4 vdd
port 1 nsew
rlabel metal3 s 60270 59318 60368 59416 4 vdd
port 1 nsew
rlabel metal3 s 60270 60466 60368 60564 4 vdd
port 1 nsew
rlabel metal3 s 59492 62850 59590 62948 4 vdd
port 1 nsew
rlabel metal3 s 59492 60875 59590 60973 4 vdd
port 1 nsew
rlabel metal3 s 60702 62046 60800 62144 4 vdd
port 1 nsew
rlabel metal3 s 59492 60085 59590 60183 4 vdd
port 1 nsew
rlabel metal3 s 60270 64058 60368 64156 4 vdd
port 1 nsew
rlabel metal3 s 59888 64035 59986 64133 4 gnd
port 2 nsew
rlabel metal3 s 60702 59676 60800 59774 4 vdd
port 1 nsew
rlabel metal3 s 60270 59676 60368 59774 4 vdd
port 1 nsew
rlabel metal3 s 61127 63268 61225 63366 4 gnd
port 2 nsew
rlabel metal3 s 61127 64058 61225 64156 4 gnd
port 2 nsew
rlabel metal3 s 60270 61256 60368 61354 4 vdd
port 1 nsew
rlabel metal3 s 59888 60480 59986 60578 4 gnd
port 2 nsew
rlabel metal3 s 61127 58944 61225 59042 4 gnd
port 2 nsew
rlabel metal3 s 60270 60108 60368 60206 4 vdd
port 1 nsew
rlabel metal3 s 61127 63684 61225 63782 4 gnd
port 2 nsew
rlabel metal3 s 59888 60875 59986 60973 4 gnd
port 2 nsew
rlabel metal3 s 60702 63626 60800 63724 4 vdd
port 1 nsew
rlabel metal3 s 59492 61270 59590 61368 4 vdd
port 1 nsew
rlabel metal3 s 59492 63245 59590 63343 4 vdd
port 1 nsew
rlabel metal3 s 59492 61665 59590 61763 4 vdd
port 1 nsew
rlabel metal3 s 62352 68402 62450 68500 4 vdd
port 1 nsew
rlabel metal3 s 60270 62478 60368 62576 4 vdd
port 1 nsew
rlabel metal3 s 59492 64035 59590 64133 4 vdd
port 1 nsew
rlabel metal3 s 59888 62455 59986 62553 4 gnd
port 2 nsew
rlabel metal3 s 59467 64621 59565 64719 4 vdd
port 1 nsew
rlabel metal3 s 60702 58886 60800 58984 4 vdd
port 1 nsew
rlabel metal3 s 59888 63640 59986 63738 4 gnd
port 2 nsew
rlabel metal3 s 59888 59690 59986 59788 4 gnd
port 2 nsew
rlabel metal3 s 59492 62455 59590 62553 4 vdd
port 1 nsew
rlabel metal3 s 59888 59295 59986 59393 4 gnd
port 2 nsew
rlabel metal3 s 61127 62478 61225 62576 4 gnd
port 2 nsew
rlabel metal3 s 59888 61665 59986 61763 4 gnd
port 2 nsew
rlabel metal3 s 60702 60108 60800 60206 4 vdd
port 1 nsew
rlabel metal3 s 61127 59734 61225 59832 4 gnd
port 2 nsew
rlabel metal3 s 60270 63268 60368 63366 4 vdd
port 1 nsew
rlabel metal3 s 59888 61270 59986 61368 4 gnd
port 2 nsew
rlabel metal3 s 59492 59690 59590 59788 4 vdd
port 1 nsew
rlabel metal3 s 61127 60108 61225 60206 4 gnd
port 2 nsew
rlabel metal3 s 60702 62478 60800 62576 4 vdd
port 1 nsew
rlabel metal3 s 60702 64058 60800 64156 4 vdd
port 1 nsew
rlabel metal3 s 59888 62850 59986 62948 4 gnd
port 2 nsew
rlabel metal3 s 59888 62060 59986 62158 4 gnd
port 2 nsew
rlabel metal3 s 61127 62104 61225 62202 4 gnd
port 2 nsew
rlabel metal3 s 60702 63268 60800 63366 4 vdd
port 1 nsew
rlabel metal3 s 60702 60466 60800 60564 4 vdd
port 1 nsew
rlabel metal3 s 59888 63245 59986 63343 4 gnd
port 2 nsew
rlabel metal3 s 60270 60898 60368 60996 4 vdd
port 1 nsew
rlabel metal3 s 59492 60480 59590 60578 4 vdd
port 1 nsew
rlabel metal3 s 59888 60085 59986 60183 4 gnd
port 2 nsew
rlabel metal3 s 62352 66988 62450 67086 4 gnd
port 2 nsew
rlabel metal3 s 59492 59295 59590 59393 4 vdd
port 1 nsew
rlabel metal3 s 60270 61688 60368 61786 4 vdd
port 1 nsew
rlabel metal3 s 59888 58900 59986 58998 4 gnd
port 2 nsew
rlabel metal3 s 61127 60898 61225 60996 4 gnd
port 2 nsew
rlabel metal3 s 61127 61688 61225 61786 4 gnd
port 2 nsew
rlabel metal3 s 60270 62046 60368 62144 4 vdd
port 1 nsew
rlabel metal3 s 59492 62060 59590 62158 4 vdd
port 1 nsew
rlabel metal3 s 60702 60898 60800 60996 4 vdd
port 1 nsew
rlabel metal3 s 59492 58900 59590 58998 4 vdd
port 1 nsew
rlabel metal3 s 60270 62836 60368 62934 4 vdd
port 1 nsew
rlabel metal3 s 61127 60524 61225 60622 4 gnd
port 2 nsew
rlabel metal3 s 60702 61256 60800 61354 4 vdd
port 1 nsew
rlabel metal3 s 60992 66988 61090 67086 4 gnd
port 2 nsew
rlabel metal3 s 61127 61314 61225 61412 4 gnd
port 2 nsew
rlabel metal3 s 60270 58886 60368 58984 4 vdd
port 1 nsew
rlabel metal3 s 61127 62894 61225 62992 4 gnd
port 2 nsew
rlabel metal3 s 60702 59318 60800 59416 4 vdd
port 1 nsew
rlabel metal3 s 61127 59318 61225 59416 4 gnd
port 2 nsew
rlabel metal3 s 60270 63626 60368 63724 4 vdd
port 1 nsew
rlabel metal3 s 35017 65582 35115 65680 4 vdd
port 1 nsew
rlabel metal3 s 47497 65582 47595 65680 4 vdd
port 1 nsew
rlabel metal3 s 36265 65582 36363 65680 4 vdd
port 1 nsew
rlabel metal3 s 42119 65582 42217 65680 4 vdd
port 1 nsew
rlabel metal3 s 38761 65582 38859 65680 4 vdd
port 1 nsew
rlabel metal3 s 39504 64991 39602 65089 4 vdd
port 1 nsew
rlabel metal3 s 47111 65582 47209 65680 4 vdd
port 1 nsew
rlabel metal3 s 43367 65582 43465 65680 4 vdd
port 1 nsew
rlabel metal3 s 48921 70398 49019 70496 4 vdd
port 1 nsew
rlabel metal3 s 33888 64991 33986 65089 4 vdd
port 1 nsew
rlabel metal3 s 41376 64991 41474 65089 4 vdd
port 1 nsew
rlabel metal3 s 39623 65582 39721 65680 4 vdd
port 1 nsew
rlabel metal3 s 43941 71558 44039 71656 4 gnd
port 2 nsew
rlabel metal3 s 48240 64991 48338 65089 4 vdd
port 1 nsew
rlabel metal3 s 41257 65582 41355 65680 4 vdd
port 1 nsew
rlabel metal3 s 34027 69624 34125 69722 4 gnd
port 2 nsew
rlabel metal3 s 38375 65582 38473 65680 4 vdd
port 1 nsew
rlabel metal3 s 37944 67131 38042 67229 4 gnd
port 2 nsew
rlabel metal3 s 36384 64991 36482 65089 4 vdd
port 1 nsew
rlabel metal3 s 43929 70398 44027 70496 4 vdd
port 1 nsew
rlabel metal3 s 49176 67131 49274 67229 4 gnd
port 2 nsew
rlabel metal3 s 33945 70398 34043 70496 4 vdd
port 1 nsew
rlabel metal3 s 35448 67131 35546 67229 4 gnd
port 2 nsew
rlabel metal3 s 41688 67131 41786 67229 4 gnd
port 2 nsew
rlabel metal3 s 37127 65582 37225 65680 4 vdd
port 1 nsew
rlabel metal3 s 39192 67131 39290 67229 4 gnd
port 2 nsew
rlabel metal3 s 36696 67131 36794 67229 4 gnd
port 2 nsew
rlabel metal3 s 46249 65582 46347 65680 4 vdd
port 1 nsew
rlabel metal3 s 34631 65582 34729 65680 4 vdd
port 1 nsew
rlabel metal3 s 45120 64991 45218 65089 4 vdd
port 1 nsew
rlabel metal3 s 43872 64991 43970 65089 4 vdd
port 1 nsew
rlabel metal3 s 38880 64991 38978 65089 4 vdd
port 1 nsew
rlabel metal3 s 48864 64991 48962 65089 4 vdd
port 1 nsew
rlabel metal3 s 35760 64991 35858 65089 4 vdd
port 1 nsew
rlabel metal3 s 44496 64991 44594 65089 4 vdd
port 1 nsew
rlabel metal3 s 37513 65582 37611 65680 4 vdd
port 1 nsew
rlabel metal3 s 47928 67131 48026 67229 4 gnd
port 2 nsew
rlabel metal3 s 35136 64991 35234 65089 4 vdd
port 1 nsew
rlabel metal3 s 43753 65582 43851 65680 4 vdd
port 1 nsew
rlabel metal3 s 48933 71236 49031 71334 4 vdd
port 1 nsew
rlabel metal3 s 38949 71558 39047 71656 4 gnd
port 2 nsew
rlabel metal3 s 49003 69624 49101 69722 4 gnd
port 2 nsew
rlabel metal3 s 48745 65582 48843 65680 4 vdd
port 1 nsew
rlabel metal3 s 44184 67131 44282 67229 4 gnd
port 2 nsew
rlabel metal3 s 42936 67131 43034 67229 4 gnd
port 2 nsew
rlabel metal3 s 39019 69624 39117 69722 4 gnd
port 2 nsew
rlabel metal3 s 40871 65582 40969 65680 4 vdd
port 1 nsew
rlabel metal3 s 46680 67131 46778 67229 4 gnd
port 2 nsew
rlabel metal3 s 35879 65582 35977 65680 4 vdd
port 1 nsew
rlabel metal3 s 49607 65582 49705 65680 4 vdd
port 1 nsew
rlabel metal3 s 38937 70398 39035 70496 4 vdd
port 1 nsew
rlabel metal3 s 33957 71558 34055 71656 4 gnd
port 2 nsew
rlabel metal3 s 44615 65582 44713 65680 4 vdd
port 1 nsew
rlabel metal3 s 48359 65582 48457 65680 4 vdd
port 1 nsew
rlabel metal3 s 38256 64991 38354 65089 4 vdd
port 1 nsew
rlabel metal3 s 42000 64991 42098 65089 4 vdd
port 1 nsew
rlabel metal3 s 42624 64991 42722 65089 4 vdd
port 1 nsew
rlabel metal3 s 34512 64991 34610 65089 4 vdd
port 1 nsew
rlabel metal3 s 45744 64991 45842 65089 4 vdd
port 1 nsew
rlabel metal3 s 45001 65582 45099 65680 4 vdd
port 1 nsew
rlabel metal3 s 49488 64991 49586 65089 4 vdd
port 1 nsew
rlabel metal3 s 40128 64991 40226 65089 4 vdd
port 1 nsew
rlabel metal3 s 38949 71236 39047 71334 4 vdd
port 1 nsew
rlabel metal3 s 40440 67131 40538 67229 4 gnd
port 2 nsew
rlabel metal3 s 46368 64991 46466 65089 4 vdd
port 1 nsew
rlabel metal3 s 44011 69624 44109 69722 4 gnd
port 2 nsew
rlabel metal3 s 33769 65582 33867 65680 4 vdd
port 1 nsew
rlabel metal3 s 40009 65582 40107 65680 4 vdd
port 1 nsew
rlabel metal3 s 34200 67131 34298 67229 4 gnd
port 2 nsew
rlabel metal3 s 48933 71558 49031 71656 4 gnd
port 2 nsew
rlabel metal3 s 46992 64991 47090 65089 4 vdd
port 1 nsew
rlabel metal3 s 37632 64991 37730 65089 4 vdd
port 1 nsew
rlabel metal3 s 42505 65582 42603 65680 4 vdd
port 1 nsew
rlabel metal3 s 37008 64991 37106 65089 4 vdd
port 1 nsew
rlabel metal3 s 45432 67131 45530 67229 4 gnd
port 2 nsew
rlabel metal3 s 45863 65582 45961 65680 4 vdd
port 1 nsew
rlabel metal3 s 43248 64991 43346 65089 4 vdd
port 1 nsew
rlabel metal3 s 40752 64991 40850 65089 4 vdd
port 1 nsew
rlabel metal3 s 43941 71236 44039 71334 4 vdd
port 1 nsew
rlabel metal3 s 47616 64991 47714 65089 4 vdd
port 1 nsew
rlabel metal3 s 33957 71236 34055 71334 4 vdd
port 1 nsew
rlabel metal3 s 60270 58528 60368 58626 4 vdd
port 1 nsew
rlabel metal3 s 59492 54950 59590 55048 4 vdd
port 1 nsew
rlabel metal3 s 60702 58096 60800 58194 4 vdd
port 1 nsew
rlabel metal3 s 60702 57306 60800 57404 4 vdd
port 1 nsew
rlabel metal3 s 60702 55726 60800 55824 4 vdd
port 1 nsew
rlabel metal3 s 60270 56516 60368 56614 4 vdd
port 1 nsew
rlabel metal3 s 59492 58110 59590 58208 4 vdd
port 1 nsew
rlabel metal3 s 60270 54146 60368 54244 4 vdd
port 1 nsew
rlabel metal3 s 60270 57306 60368 57404 4 vdd
port 1 nsew
rlabel metal3 s 60270 56158 60368 56256 4 vdd
port 1 nsew
rlabel metal3 s 60270 58096 60368 58194 4 vdd
port 1 nsew
rlabel metal3 s 60270 55368 60368 55466 4 vdd
port 1 nsew
rlabel metal3 s 61127 56948 61225 57046 4 gnd
port 2 nsew
rlabel metal3 s 61127 54204 61225 54302 4 gnd
port 2 nsew
rlabel metal3 s 59492 56530 59590 56628 4 vdd
port 1 nsew
rlabel metal3 s 60270 57738 60368 57836 4 vdd
port 1 nsew
rlabel metal3 s 60270 55726 60368 55824 4 vdd
port 1 nsew
rlabel metal3 s 59888 54950 59986 55048 4 gnd
port 2 nsew
rlabel metal3 s 59492 54160 59590 54258 4 vdd
port 1 nsew
rlabel metal3 s 60702 57738 60800 57836 4 vdd
port 1 nsew
rlabel metal3 s 60702 56516 60800 56614 4 vdd
port 1 nsew
rlabel metal3 s 61127 56574 61225 56672 4 gnd
port 2 nsew
rlabel metal3 s 59492 57320 59590 57418 4 vdd
port 1 nsew
rlabel metal3 s 60702 58528 60800 58626 4 vdd
port 1 nsew
rlabel metal3 s 59888 54555 59986 54653 4 gnd
port 2 nsew
rlabel metal3 s 61127 55368 61225 55466 4 gnd
port 2 nsew
rlabel metal3 s 59492 55345 59590 55443 4 vdd
port 1 nsew
rlabel metal3 s 60702 56158 60800 56256 4 vdd
port 1 nsew
rlabel metal3 s 60270 56948 60368 57046 4 vdd
port 1 nsew
rlabel metal3 s 59888 55740 59986 55838 4 gnd
port 2 nsew
rlabel metal3 s 59888 55345 59986 55443 4 gnd
port 2 nsew
rlabel metal3 s 61127 58528 61225 58626 4 gnd
port 2 nsew
rlabel metal3 s 61127 55784 61225 55882 4 gnd
port 2 nsew
rlabel metal3 s 59888 58110 59986 58208 4 gnd
port 2 nsew
rlabel metal3 s 59492 56135 59590 56233 4 vdd
port 1 nsew
rlabel metal3 s 59888 57320 59986 57418 4 gnd
port 2 nsew
rlabel metal3 s 59492 55740 59590 55838 4 vdd
port 1 nsew
rlabel metal3 s 60702 54578 60800 54676 4 vdd
port 1 nsew
rlabel metal3 s 59492 56925 59590 57023 4 vdd
port 1 nsew
rlabel metal3 s 61127 57364 61225 57462 4 gnd
port 2 nsew
rlabel metal3 s 59888 56530 59986 56628 4 gnd
port 2 nsew
rlabel metal3 s 59492 57715 59590 57813 4 vdd
port 1 nsew
rlabel metal3 s 59888 57715 59986 57813 4 gnd
port 2 nsew
rlabel metal3 s 60702 54146 60800 54244 4 vdd
port 1 nsew
rlabel metal3 s 60702 56948 60800 57046 4 vdd
port 1 nsew
rlabel metal3 s 60270 54936 60368 55034 4 vdd
port 1 nsew
rlabel metal3 s 61127 57738 61225 57836 4 gnd
port 2 nsew
rlabel metal3 s 60270 54578 60368 54676 4 vdd
port 1 nsew
rlabel metal3 s 61127 58154 61225 58252 4 gnd
port 2 nsew
rlabel metal3 s 59492 54555 59590 54653 4 vdd
port 1 nsew
rlabel metal3 s 61127 54994 61225 55092 4 gnd
port 2 nsew
rlabel metal3 s 61127 54578 61225 54676 4 gnd
port 2 nsew
rlabel metal3 s 59888 56925 59986 57023 4 gnd
port 2 nsew
rlabel metal3 s 60702 54936 60800 55034 4 vdd
port 1 nsew
rlabel metal3 s 59888 54160 59986 54258 4 gnd
port 2 nsew
rlabel metal3 s 59888 56135 59986 56233 4 gnd
port 2 nsew
rlabel metal3 s 60702 55368 60800 55466 4 vdd
port 1 nsew
rlabel metal3 s 61127 56158 61225 56256 4 gnd
port 2 nsew
rlabel metal3 s 59888 58505 59986 58603 4 gnd
port 2 nsew
rlabel metal3 s 59492 58505 59590 58603 4 vdd
port 1 nsew
rlabel metal3 s 60702 51776 60800 51874 4 vdd
port 1 nsew
rlabel metal3 s 59492 51790 59590 51888 4 vdd
port 1 nsew
rlabel metal3 s 59492 51395 59590 51493 4 vdd
port 1 nsew
rlabel metal3 s 59492 50210 59590 50308 4 vdd
port 1 nsew
rlabel metal3 s 59492 52185 59590 52283 4 vdd
port 1 nsew
rlabel metal3 s 59888 49025 59986 49123 4 gnd
port 2 nsew
rlabel metal3 s 59888 52185 59986 52283 4 gnd
port 2 nsew
rlabel metal3 s 60702 53788 60800 53886 4 vdd
port 1 nsew
rlabel metal3 s 59492 52975 59590 53073 4 vdd
port 1 nsew
rlabel metal3 s 60270 49838 60368 49936 4 vdd
port 1 nsew
rlabel metal3 s 60702 52566 60800 52664 4 vdd
port 1 nsew
rlabel metal3 s 60270 50986 60368 51084 4 vdd
port 1 nsew
rlabel metal3 s 60702 49406 60800 49504 4 vdd
port 1 nsew
rlabel metal3 s 61127 50628 61225 50726 4 gnd
port 2 nsew
rlabel metal3 s 59492 53370 59590 53468 4 vdd
port 1 nsew
rlabel metal3 s 61127 53414 61225 53512 4 gnd
port 2 nsew
rlabel metal3 s 60270 53788 60368 53886 4 vdd
port 1 nsew
rlabel metal3 s 59888 51000 59986 51098 4 gnd
port 2 nsew
rlabel metal3 s 59492 50605 59590 50703 4 vdd
port 1 nsew
rlabel metal3 s 60270 52208 60368 52306 4 vdd
port 1 nsew
rlabel metal3 s 59888 52580 59986 52678 4 gnd
port 2 nsew
rlabel metal3 s 59492 53765 59590 53863 4 vdd
port 1 nsew
rlabel metal3 s 60702 49838 60800 49936 4 vdd
port 1 nsew
rlabel metal3 s 61127 52998 61225 53096 4 gnd
port 2 nsew
rlabel metal3 s 60270 52566 60368 52664 4 vdd
port 1 nsew
rlabel metal3 s 61127 49838 61225 49936 4 gnd
port 2 nsew
rlabel metal3 s 59492 49815 59590 49913 4 vdd
port 1 nsew
rlabel metal3 s 59888 53370 59986 53468 4 gnd
port 2 nsew
rlabel metal3 s 60702 52208 60800 52306 4 vdd
port 1 nsew
rlabel metal3 s 59888 49420 59986 49518 4 gnd
port 2 nsew
rlabel metal3 s 59888 50210 59986 50308 4 gnd
port 2 nsew
rlabel metal3 s 60702 53356 60800 53454 4 vdd
port 1 nsew
rlabel metal3 s 61127 52208 61225 52306 4 gnd
port 2 nsew
rlabel metal3 s 60270 53356 60368 53454 4 vdd
port 1 nsew
rlabel metal3 s 59888 53765 59986 53863 4 gnd
port 2 nsew
rlabel metal3 s 59888 50605 59986 50703 4 gnd
port 2 nsew
rlabel metal3 s 61127 50254 61225 50352 4 gnd
port 2 nsew
rlabel metal3 s 59888 49815 59986 49913 4 gnd
port 2 nsew
rlabel metal3 s 61127 49048 61225 49146 4 gnd
port 2 nsew
rlabel metal3 s 60270 51776 60368 51874 4 vdd
port 1 nsew
rlabel metal3 s 61127 52624 61225 52722 4 gnd
port 2 nsew
rlabel metal3 s 60270 50628 60368 50726 4 vdd
port 1 nsew
rlabel metal3 s 59492 49025 59590 49123 4 vdd
port 1 nsew
rlabel metal3 s 60270 49406 60368 49504 4 vdd
port 1 nsew
rlabel metal3 s 60270 49048 60368 49146 4 vdd
port 1 nsew
rlabel metal3 s 59888 52975 59986 53073 4 gnd
port 2 nsew
rlabel metal3 s 60702 51418 60800 51516 4 vdd
port 1 nsew
rlabel metal3 s 59492 49420 59590 49518 4 vdd
port 1 nsew
rlabel metal3 s 60270 50196 60368 50294 4 vdd
port 1 nsew
rlabel metal3 s 60702 50628 60800 50726 4 vdd
port 1 nsew
rlabel metal3 s 60702 52998 60800 53096 4 vdd
port 1 nsew
rlabel metal3 s 59888 51790 59986 51888 4 gnd
port 2 nsew
rlabel metal3 s 60270 52998 60368 53096 4 vdd
port 1 nsew
rlabel metal3 s 59492 51000 59590 51098 4 vdd
port 1 nsew
rlabel metal3 s 61127 53788 61225 53886 4 gnd
port 2 nsew
rlabel metal3 s 60702 50196 60800 50294 4 vdd
port 1 nsew
rlabel metal3 s 60702 50986 60800 51084 4 vdd
port 1 nsew
rlabel metal3 s 61127 49464 61225 49562 4 gnd
port 2 nsew
rlabel metal3 s 61127 51044 61225 51142 4 gnd
port 2 nsew
rlabel metal3 s 61127 51834 61225 51932 4 gnd
port 2 nsew
rlabel metal3 s 61127 51418 61225 51516 4 gnd
port 2 nsew
rlabel metal3 s 59492 52580 59590 52678 4 vdd
port 1 nsew
rlabel metal3 s 59888 51395 59986 51493 4 gnd
port 2 nsew
rlabel metal3 s 60702 49048 60800 49146 4 vdd
port 1 nsew
rlabel metal3 s 60270 51418 60368 51516 4 vdd
port 1 nsew
rlabel metal3 s 54552 57320 54650 57418 4 gnd
port 2 nsew
rlabel metal3 s 54552 54713 54650 54811 4 gnd
port 2 nsew
rlabel metal3 s 54552 50447 54650 50545 4 gnd
port 2 nsew
rlabel metal3 s 54552 49973 54650 50071 4 gnd
port 2 nsew
rlabel metal3 s 54552 56530 54650 56628 4 gnd
port 2 nsew
rlabel metal3 s 54552 50210 54650 50308 4 gnd
port 2 nsew
rlabel metal3 s 54552 53370 54650 53468 4 gnd
port 2 nsew
rlabel metal3 s 54552 55503 54650 55601 4 gnd
port 2 nsew
rlabel metal3 s 54552 56293 54650 56391 4 gnd
port 2 nsew
rlabel metal3 s 54552 58347 54650 58445 4 gnd
port 2 nsew
rlabel metal3 s 54552 54160 54650 54258 4 gnd
port 2 nsew
rlabel metal3 s 54552 51553 54650 51651 4 gnd
port 2 nsew
rlabel metal3 s 54552 51000 54650 51098 4 gnd
port 2 nsew
rlabel metal3 s 54552 57873 54650 57971 4 gnd
port 2 nsew
rlabel metal3 s 54552 58110 54650 58208 4 gnd
port 2 nsew
rlabel metal3 s 54552 53923 54650 54021 4 gnd
port 2 nsew
rlabel metal3 s 54552 52817 54650 52915 4 gnd
port 2 nsew
rlabel metal3 s 54552 51790 54650 51888 4 gnd
port 2 nsew
rlabel metal3 s 54552 49420 54650 49518 4 gnd
port 2 nsew
rlabel metal3 s 54552 51237 54650 51335 4 gnd
port 2 nsew
rlabel metal3 s 54552 57083 54650 57181 4 gnd
port 2 nsew
rlabel metal3 s 54552 49657 54650 49755 4 gnd
port 2 nsew
rlabel metal3 s 54552 55740 54650 55838 4 gnd
port 2 nsew
rlabel metal3 s 54552 56767 54650 56865 4 gnd
port 2 nsew
rlabel metal3 s 54552 50763 54650 50861 4 gnd
port 2 nsew
rlabel metal3 s 54552 55977 54650 56075 4 gnd
port 2 nsew
rlabel metal3 s 54552 49183 54650 49281 4 gnd
port 2 nsew
rlabel metal3 s 54552 54397 54650 54495 4 gnd
port 2 nsew
rlabel metal3 s 54552 58663 54650 58761 4 gnd
port 2 nsew
rlabel metal3 s 54552 52027 54650 52125 4 gnd
port 2 nsew
rlabel metal3 s 54552 53133 54650 53231 4 gnd
port 2 nsew
rlabel metal3 s 54552 57557 54650 57655 4 gnd
port 2 nsew
rlabel metal3 s 54552 52343 54650 52441 4 gnd
port 2 nsew
rlabel metal3 s 54552 55187 54650 55285 4 gnd
port 2 nsew
rlabel metal3 s 54552 52580 54650 52678 4 gnd
port 2 nsew
rlabel metal3 s 54552 54950 54650 55048 4 gnd
port 2 nsew
rlabel metal3 s 54552 53607 54650 53705 4 gnd
port 2 nsew
rlabel metal3 s 54552 48630 54650 48728 4 gnd
port 2 nsew
rlabel metal3 s 54552 46813 54650 46911 4 gnd
port 2 nsew
rlabel metal3 s 54552 48393 54650 48491 4 gnd
port 2 nsew
rlabel metal3 s 54552 43337 54650 43435 4 gnd
port 2 nsew
rlabel metal3 s 54552 46497 54650 46595 4 gnd
port 2 nsew
rlabel metal3 s 54552 39387 54650 39485 4 gnd
port 2 nsew
rlabel metal3 s 54552 48077 54650 48175 4 gnd
port 2 nsew
rlabel metal3 s 54552 42073 54650 42171 4 gnd
port 2 nsew
rlabel metal3 s 54552 43890 54650 43988 4 gnd
port 2 nsew
rlabel metal3 s 54552 44127 54650 44225 4 gnd
port 2 nsew
rlabel metal3 s 54552 40967 54650 41065 4 gnd
port 2 nsew
rlabel metal3 s 54552 45233 54650 45331 4 gnd
port 2 nsew
rlabel metal3 s 54552 42547 54650 42645 4 gnd
port 2 nsew
rlabel metal3 s 54552 41757 54650 41855 4 gnd
port 2 nsew
rlabel metal3 s 54552 39703 54650 39801 4 gnd
port 2 nsew
rlabel metal3 s 54552 47840 54650 47938 4 gnd
port 2 nsew
rlabel metal3 s 54552 48867 54650 48965 4 gnd
port 2 nsew
rlabel metal3 s 54552 47050 54650 47148 4 gnd
port 2 nsew
rlabel metal3 s 54552 43653 54650 43751 4 gnd
port 2 nsew
rlabel metal3 s 54552 46260 54650 46358 4 gnd
port 2 nsew
rlabel metal3 s 54552 40730 54650 40828 4 gnd
port 2 nsew
rlabel metal3 s 54552 39940 54650 40038 4 gnd
port 2 nsew
rlabel metal3 s 54552 47603 54650 47701 4 gnd
port 2 nsew
rlabel metal3 s 54552 46023 54650 46121 4 gnd
port 2 nsew
rlabel metal3 s 54552 45707 54650 45805 4 gnd
port 2 nsew
rlabel metal3 s 54552 40493 54650 40591 4 gnd
port 2 nsew
rlabel metal3 s 54552 42310 54650 42408 4 gnd
port 2 nsew
rlabel metal3 s 54552 42863 54650 42961 4 gnd
port 2 nsew
rlabel metal3 s 54552 44917 54650 45015 4 gnd
port 2 nsew
rlabel metal3 s 54552 43100 54650 43198 4 gnd
port 2 nsew
rlabel metal3 s 54552 41520 54650 41618 4 gnd
port 2 nsew
rlabel metal3 s 54552 44680 54650 44778 4 gnd
port 2 nsew
rlabel metal3 s 54552 45470 54650 45568 4 gnd
port 2 nsew
rlabel metal3 s 54552 47287 54650 47385 4 gnd
port 2 nsew
rlabel metal3 s 54552 41283 54650 41381 4 gnd
port 2 nsew
rlabel metal3 s 54552 44443 54650 44541 4 gnd
port 2 nsew
rlabel metal3 s 54552 40177 54650 40275 4 gnd
port 2 nsew
rlabel metal3 s 59888 46655 59986 46753 4 gnd
port 2 nsew
rlabel metal3 s 59888 44680 59986 44778 4 gnd
port 2 nsew
rlabel metal3 s 60270 45888 60368 45986 4 vdd
port 1 nsew
rlabel metal3 s 59492 48630 59590 48728 4 vdd
port 1 nsew
rlabel metal3 s 60702 47468 60800 47566 4 vdd
port 1 nsew
rlabel metal3 s 59492 45075 59590 45173 4 vdd
port 1 nsew
rlabel metal3 s 60702 45456 60800 45554 4 vdd
port 1 nsew
rlabel metal3 s 60702 47036 60800 47134 4 vdd
port 1 nsew
rlabel metal3 s 61127 47094 61225 47192 4 gnd
port 2 nsew
rlabel metal3 s 61127 48258 61225 48356 4 gnd
port 2 nsew
rlabel metal3 s 60702 46246 60800 46344 4 vdd
port 1 nsew
rlabel metal3 s 59492 47840 59590 47938 4 vdd
port 1 nsew
rlabel metal3 s 60702 48616 60800 48714 4 vdd
port 1 nsew
rlabel metal3 s 59888 47445 59986 47543 4 gnd
port 2 nsew
rlabel metal3 s 60270 45456 60368 45554 4 vdd
port 1 nsew
rlabel metal3 s 60270 48258 60368 48356 4 vdd
port 1 nsew
rlabel metal3 s 61127 44308 61225 44406 4 gnd
port 2 nsew
rlabel metal3 s 59888 44285 59986 44383 4 gnd
port 2 nsew
rlabel metal3 s 61127 45888 61225 45986 4 gnd
port 2 nsew
rlabel metal3 s 60270 45098 60368 45196 4 vdd
port 1 nsew
rlabel metal3 s 60702 48258 60800 48356 4 vdd
port 1 nsew
rlabel metal3 s 59888 48235 59986 48333 4 gnd
port 2 nsew
rlabel metal3 s 59888 45865 59986 45963 4 gnd
port 2 nsew
rlabel metal3 s 60702 47826 60800 47924 4 vdd
port 1 nsew
rlabel metal3 s 59492 44285 59590 44383 4 vdd
port 1 nsew
rlabel metal3 s 60270 44308 60368 44406 4 vdd
port 1 nsew
rlabel metal3 s 60270 46246 60368 46344 4 vdd
port 1 nsew
rlabel metal3 s 61127 47468 61225 47566 4 gnd
port 2 nsew
rlabel metal3 s 59888 45470 59986 45568 4 gnd
port 2 nsew
rlabel metal3 s 61127 47884 61225 47982 4 gnd
port 2 nsew
rlabel metal3 s 59888 47840 59986 47938 4 gnd
port 2 nsew
rlabel metal3 s 59492 44680 59590 44778 4 vdd
port 1 nsew
rlabel metal3 s 60702 44666 60800 44764 4 vdd
port 1 nsew
rlabel metal3 s 60702 45098 60800 45196 4 vdd
port 1 nsew
rlabel metal3 s 60270 48616 60368 48714 4 vdd
port 1 nsew
rlabel metal3 s 61127 45098 61225 45196 4 gnd
port 2 nsew
rlabel metal3 s 60270 44666 60368 44764 4 vdd
port 1 nsew
rlabel metal3 s 61127 45514 61225 45612 4 gnd
port 2 nsew
rlabel metal3 s 61127 48674 61225 48772 4 gnd
port 2 nsew
rlabel metal3 s 60270 47468 60368 47566 4 vdd
port 1 nsew
rlabel metal3 s 60702 45888 60800 45986 4 vdd
port 1 nsew
rlabel metal3 s 60270 46678 60368 46776 4 vdd
port 1 nsew
rlabel metal3 s 59888 48630 59986 48728 4 gnd
port 2 nsew
rlabel metal3 s 59492 46655 59590 46753 4 vdd
port 1 nsew
rlabel metal3 s 59492 46260 59590 46358 4 vdd
port 1 nsew
rlabel metal3 s 61127 46678 61225 46776 4 gnd
port 2 nsew
rlabel metal3 s 59492 47050 59590 47148 4 vdd
port 1 nsew
rlabel metal3 s 60702 44308 60800 44406 4 vdd
port 1 nsew
rlabel metal3 s 60702 46678 60800 46776 4 vdd
port 1 nsew
rlabel metal3 s 59492 48235 59590 48333 4 vdd
port 1 nsew
rlabel metal3 s 59492 47445 59590 47543 4 vdd
port 1 nsew
rlabel metal3 s 59888 46260 59986 46358 4 gnd
port 2 nsew
rlabel metal3 s 60270 47036 60368 47134 4 vdd
port 1 nsew
rlabel metal3 s 59492 45470 59590 45568 4 vdd
port 1 nsew
rlabel metal3 s 59888 47050 59986 47148 4 gnd
port 2 nsew
rlabel metal3 s 61127 44724 61225 44822 4 gnd
port 2 nsew
rlabel metal3 s 61127 46304 61225 46402 4 gnd
port 2 nsew
rlabel metal3 s 59888 45075 59986 45173 4 gnd
port 2 nsew
rlabel metal3 s 59492 45865 59590 45963 4 vdd
port 1 nsew
rlabel metal3 s 60270 47826 60368 47924 4 vdd
port 1 nsew
rlabel metal3 s 59888 39545 59986 39643 4 gnd
port 2 nsew
rlabel metal3 s 59888 41915 59986 42013 4 gnd
port 2 nsew
rlabel metal3 s 59888 40730 59986 40828 4 gnd
port 2 nsew
rlabel metal3 s 61127 43144 61225 43242 4 gnd
port 2 nsew
rlabel metal3 s 61127 41938 61225 42036 4 gnd
port 2 nsew
rlabel metal3 s 59888 42705 59986 42803 4 gnd
port 2 nsew
rlabel metal3 s 59492 40730 59590 40828 4 vdd
port 1 nsew
rlabel metal3 s 59888 43495 59986 43593 4 gnd
port 2 nsew
rlabel metal3 s 61127 40774 61225 40872 4 gnd
port 2 nsew
rlabel metal3 s 59492 42310 59590 42408 4 vdd
port 1 nsew
rlabel metal3 s 60702 40358 60800 40456 4 vdd
port 1 nsew
rlabel metal3 s 60270 43876 60368 43974 4 vdd
port 1 nsew
rlabel metal3 s 60270 41148 60368 41246 4 vdd
port 1 nsew
rlabel metal3 s 60702 41506 60800 41604 4 vdd
port 1 nsew
rlabel metal3 s 59888 43890 59986 43988 4 gnd
port 2 nsew
rlabel metal3 s 60702 43086 60800 43184 4 vdd
port 1 nsew
rlabel metal3 s 60270 39568 60368 39666 4 vdd
port 1 nsew
rlabel metal3 s 59492 39545 59590 39643 4 vdd
port 1 nsew
rlabel metal3 s 59492 43495 59590 43593 4 vdd
port 1 nsew
rlabel metal3 s 61127 40358 61225 40456 4 gnd
port 2 nsew
rlabel metal3 s 59492 41125 59590 41223 4 vdd
port 1 nsew
rlabel metal3 s 59888 43100 59986 43198 4 gnd
port 2 nsew
rlabel metal3 s 61127 42728 61225 42826 4 gnd
port 2 nsew
rlabel metal3 s 60270 42296 60368 42394 4 vdd
port 1 nsew
rlabel metal3 s 60270 39926 60368 40024 4 vdd
port 1 nsew
rlabel metal3 s 60270 41938 60368 42036 4 vdd
port 1 nsew
rlabel metal3 s 61127 41148 61225 41246 4 gnd
port 2 nsew
rlabel metal3 s 61127 43518 61225 43616 4 gnd
port 2 nsew
rlabel metal3 s 60270 40358 60368 40456 4 vdd
port 1 nsew
rlabel metal3 s 61127 43934 61225 44032 4 gnd
port 2 nsew
rlabel metal3 s 60702 41938 60800 42036 4 vdd
port 1 nsew
rlabel metal3 s 59492 42705 59590 42803 4 vdd
port 1 nsew
rlabel metal3 s 59492 40335 59590 40433 4 vdd
port 1 nsew
rlabel metal3 s 60270 43518 60368 43616 4 vdd
port 1 nsew
rlabel metal3 s 59888 40335 59986 40433 4 gnd
port 2 nsew
rlabel metal3 s 60702 39568 60800 39666 4 vdd
port 1 nsew
rlabel metal3 s 60702 43518 60800 43616 4 vdd
port 1 nsew
rlabel metal3 s 61127 41564 61225 41662 4 gnd
port 2 nsew
rlabel metal3 s 59888 41125 59986 41223 4 gnd
port 2 nsew
rlabel metal3 s 60702 42296 60800 42394 4 vdd
port 1 nsew
rlabel metal3 s 59492 39940 59590 40038 4 vdd
port 1 nsew
rlabel metal3 s 60270 40716 60368 40814 4 vdd
port 1 nsew
rlabel metal3 s 61127 42354 61225 42452 4 gnd
port 2 nsew
rlabel metal3 s 61127 39984 61225 40082 4 gnd
port 2 nsew
rlabel metal3 s 60702 43876 60800 43974 4 vdd
port 1 nsew
rlabel metal3 s 60702 39926 60800 40024 4 vdd
port 1 nsew
rlabel metal3 s 59492 41520 59590 41618 4 vdd
port 1 nsew
rlabel metal3 s 60270 41506 60368 41604 4 vdd
port 1 nsew
rlabel metal3 s 59492 43100 59590 43198 4 vdd
port 1 nsew
rlabel metal3 s 60270 42728 60368 42826 4 vdd
port 1 nsew
rlabel metal3 s 61127 39194 61225 39292 4 gnd
port 2 nsew
rlabel metal3 s 60702 40716 60800 40814 4 vdd
port 1 nsew
rlabel metal3 s 60702 41148 60800 41246 4 vdd
port 1 nsew
rlabel metal3 s 59492 43890 59590 43988 4 vdd
port 1 nsew
rlabel metal3 s 61127 39568 61225 39666 4 gnd
port 2 nsew
rlabel metal3 s 59888 41520 59986 41618 4 gnd
port 2 nsew
rlabel metal3 s 60702 42728 60800 42826 4 vdd
port 1 nsew
rlabel metal3 s 59492 41915 59590 42013 4 vdd
port 1 nsew
rlabel metal3 s 60270 43086 60368 43184 4 vdd
port 1 nsew
rlabel metal3 s 59888 39940 59986 40038 4 gnd
port 2 nsew
rlabel metal3 s 59888 42310 59986 42408 4 gnd
port 2 nsew
rlabel metal3 s 17664 64991 17762 65089 4 vdd
port 1 nsew
rlabel metal3 s 21408 64991 21506 65089 4 vdd
port 1 nsew
rlabel metal3 s 30144 64991 30242 65089 4 vdd
port 1 nsew
rlabel metal3 s 33264 64991 33362 65089 4 vdd
port 1 nsew
rlabel metal3 s 20472 67131 20570 67229 4 gnd
port 2 nsew
rlabel metal3 s 30768 64991 30866 65089 4 vdd
port 1 nsew
rlabel metal3 s 28391 65582 28489 65680 4 vdd
port 1 nsew
rlabel metal3 s 24216 67131 24314 67229 4 gnd
port 2 nsew
rlabel metal3 s 23973 71558 24071 71656 4 gnd
port 2 nsew
rlabel metal3 s 25895 65582 25993 65680 4 vdd
port 1 nsew
rlabel metal3 s 22032 64991 22130 65089 4 vdd
port 1 nsew
rlabel metal3 s 27648 64991 27746 65089 4 vdd
port 1 nsew
rlabel metal3 s 19224 67131 19322 67229 4 gnd
port 2 nsew
rlabel metal3 s 26712 67131 26810 67229 4 gnd
port 2 nsew
rlabel metal3 s 30025 65582 30123 65680 4 vdd
port 1 nsew
rlabel metal3 s 18407 65582 18505 65680 4 vdd
port 1 nsew
rlabel metal3 s 32016 64991 32114 65089 4 vdd
port 1 nsew
rlabel metal3 s 22151 65582 22249 65680 4 vdd
port 1 nsew
rlabel metal3 s 25033 65582 25131 65680 4 vdd
port 1 nsew
rlabel metal3 s 18793 65582 18891 65680 4 vdd
port 1 nsew
rlabel metal3 s 22656 64991 22754 65089 4 vdd
port 1 nsew
rlabel metal3 s 27529 65582 27627 65680 4 vdd
port 1 nsew
rlabel metal3 s 26400 64991 26498 65089 4 vdd
port 1 nsew
rlabel metal3 s 27960 67131 28058 67229 4 gnd
port 2 nsew
rlabel metal3 s 30456 67131 30554 67229 4 gnd
port 2 nsew
rlabel metal3 s 20160 64991 20258 65089 4 vdd
port 1 nsew
rlabel metal3 s 18981 71558 19079 71656 4 gnd
port 2 nsew
rlabel metal3 s 24528 64991 24626 65089 4 vdd
port 1 nsew
rlabel metal3 s 25152 64991 25250 65089 4 vdd
port 1 nsew
rlabel metal3 s 23973 71236 24071 71334 4 vdd
port 1 nsew
rlabel metal3 s 18981 71236 19079 71334 4 vdd
port 1 nsew
rlabel metal3 s 26281 65582 26379 65680 4 vdd
port 1 nsew
rlabel metal3 s 28777 65582 28875 65680 4 vdd
port 1 nsew
rlabel metal3 s 23961 70398 24059 70496 4 vdd
port 1 nsew
rlabel metal3 s 29639 65582 29737 65680 4 vdd
port 1 nsew
rlabel metal3 s 24647 65582 24745 65680 4 vdd
port 1 nsew
rlabel metal3 s 22968 67131 23066 67229 4 gnd
port 2 nsew
rlabel metal3 s 20041 65582 20139 65680 4 vdd
port 1 nsew
rlabel metal3 s 32640 64991 32738 65089 4 vdd
port 1 nsew
rlabel metal3 s 30887 65582 30985 65680 4 vdd
port 1 nsew
rlabel metal3 s 23280 64991 23378 65089 4 vdd
port 1 nsew
rlabel metal3 s 32521 65582 32619 65680 4 vdd
port 1 nsew
rlabel metal3 s 20903 65582 21001 65680 4 vdd
port 1 nsew
rlabel metal3 s 28896 64991 28994 65089 4 vdd
port 1 nsew
rlabel metal3 s 18969 70398 19067 70496 4 vdd
port 1 nsew
rlabel metal3 s 20784 64991 20882 65089 4 vdd
port 1 nsew
rlabel metal3 s 33383 65582 33481 65680 4 vdd
port 1 nsew
rlabel metal3 s 31704 67131 31802 67229 4 gnd
port 2 nsew
rlabel metal3 s 28953 70398 29051 70496 4 vdd
port 1 nsew
rlabel metal3 s 32135 65582 32233 65680 4 vdd
port 1 nsew
rlabel metal3 s 18288 64991 18386 65089 4 vdd
port 1 nsew
rlabel metal3 s 28965 71236 29063 71334 4 vdd
port 1 nsew
rlabel metal3 s 22537 65582 22635 65680 4 vdd
port 1 nsew
rlabel metal3 s 31273 65582 31371 65680 4 vdd
port 1 nsew
rlabel metal3 s 28272 64991 28370 65089 4 vdd
port 1 nsew
rlabel metal3 s 31392 64991 31490 65089 4 vdd
port 1 nsew
rlabel metal3 s 29520 64991 29618 65089 4 vdd
port 1 nsew
rlabel metal3 s 24043 69624 24141 69722 4 gnd
port 2 nsew
rlabel metal3 s 23399 65582 23497 65680 4 vdd
port 1 nsew
rlabel metal3 s 21720 67131 21818 67229 4 gnd
port 2 nsew
rlabel metal3 s 23904 64991 24002 65089 4 vdd
port 1 nsew
rlabel metal3 s 18912 64991 19010 65089 4 vdd
port 1 nsew
rlabel metal3 s 23785 65582 23883 65680 4 vdd
port 1 nsew
rlabel metal3 s 19536 64991 19634 65089 4 vdd
port 1 nsew
rlabel metal3 s 19051 69624 19149 69722 4 gnd
port 2 nsew
rlabel metal3 s 29035 69624 29133 69722 4 gnd
port 2 nsew
rlabel metal3 s 25464 67131 25562 67229 4 gnd
port 2 nsew
rlabel metal3 s 32952 67131 33050 67229 4 gnd
port 2 nsew
rlabel metal3 s 29208 67131 29306 67229 4 gnd
port 2 nsew
rlabel metal3 s 21289 65582 21387 65680 4 vdd
port 1 nsew
rlabel metal3 s 27143 65582 27241 65680 4 vdd
port 1 nsew
rlabel metal3 s 27024 64991 27122 65089 4 vdd
port 1 nsew
rlabel metal3 s 19655 65582 19753 65680 4 vdd
port 1 nsew
rlabel metal3 s 17545 65582 17643 65680 4 vdd
port 1 nsew
rlabel metal3 s 25776 64991 25874 65089 4 vdd
port 1 nsew
rlabel metal3 s 28965 71558 29063 71656 4 gnd
port 2 nsew
rlabel metal3 s 17976 67131 18074 67229 4 gnd
port 2 nsew
rlabel metal3 s 13989 71236 14087 71334 4 vdd
port 1 nsew
rlabel metal3 s 14059 69624 14157 69722 4 gnd
port 2 nsew
rlabel metal3 s 13989 71558 14087 71656 4 gnd
port 2 nsew
rlabel metal3 s 13977 70398 14075 70496 4 vdd
port 1 nsew
rlabel metal3 s 6450 58886 6548 58984 4 vdd
port 1 nsew
rlabel metal3 s 7660 64035 7758 64133 4 vdd
port 1 nsew
rlabel metal3 s 7264 63245 7362 63343 4 gnd
port 2 nsew
rlabel metal3 s 6450 63626 6548 63724 4 vdd
port 1 nsew
rlabel metal3 s 7660 63640 7758 63738 4 vdd
port 1 nsew
rlabel metal3 s 7264 61270 7362 61368 4 gnd
port 2 nsew
rlabel metal3 s 7264 58900 7362 58998 4 gnd
port 2 nsew
rlabel metal3 s 6882 60898 6980 60996 4 vdd
port 1 nsew
rlabel metal3 s 6450 60108 6548 60206 4 vdd
port 1 nsew
rlabel metal3 s 7660 62060 7758 62158 4 vdd
port 1 nsew
rlabel metal3 s 7264 59690 7362 59788 4 gnd
port 2 nsew
rlabel metal3 s 6025 62104 6123 62202 4 gnd
port 2 nsew
rlabel metal3 s 6450 63268 6548 63366 4 vdd
port 1 nsew
rlabel metal3 s 6025 63684 6123 63782 4 gnd
port 2 nsew
rlabel metal3 s 6450 62836 6548 62934 4 vdd
port 1 nsew
rlabel metal3 s 6450 61256 6548 61354 4 vdd
port 1 nsew
rlabel metal3 s 7660 62455 7758 62553 4 vdd
port 1 nsew
rlabel metal3 s 7660 59690 7758 59788 4 vdd
port 1 nsew
rlabel metal3 s 7660 61270 7758 61368 4 vdd
port 1 nsew
rlabel metal3 s 6882 59318 6980 59416 4 vdd
port 1 nsew
rlabel metal3 s 6450 62478 6548 62576 4 vdd
port 1 nsew
rlabel metal3 s 6450 61688 6548 61786 4 vdd
port 1 nsew
rlabel metal3 s 6882 62836 6980 62934 4 vdd
port 1 nsew
rlabel metal3 s 6450 59676 6548 59774 4 vdd
port 1 nsew
rlabel metal3 s 6882 60466 6980 60564 4 vdd
port 1 nsew
rlabel metal3 s 6450 60898 6548 60996 4 vdd
port 1 nsew
rlabel metal3 s 6882 62046 6980 62144 4 vdd
port 1 nsew
rlabel metal3 s 6450 62046 6548 62144 4 vdd
port 1 nsew
rlabel metal3 s 7264 59295 7362 59393 4 gnd
port 2 nsew
rlabel metal3 s 6882 61688 6980 61786 4 vdd
port 1 nsew
rlabel metal3 s 6025 58944 6123 59042 4 gnd
port 2 nsew
rlabel metal3 s 7264 62850 7362 62948 4 gnd
port 2 nsew
rlabel metal3 s 6025 60524 6123 60622 4 gnd
port 2 nsew
rlabel metal3 s 7264 63640 7362 63738 4 gnd
port 2 nsew
rlabel metal3 s 6025 60898 6123 60996 4 gnd
port 2 nsew
rlabel metal3 s 6025 62478 6123 62576 4 gnd
port 2 nsew
rlabel metal3 s 7660 62850 7758 62948 4 vdd
port 1 nsew
rlabel metal3 s 7264 60875 7362 60973 4 gnd
port 2 nsew
rlabel metal3 s 7660 59295 7758 59393 4 vdd
port 1 nsew
rlabel metal3 s 6025 59318 6123 59416 4 gnd
port 2 nsew
rlabel metal3 s 7660 60085 7758 60183 4 vdd
port 1 nsew
rlabel metal3 s 7264 60480 7362 60578 4 gnd
port 2 nsew
rlabel metal3 s 6025 61314 6123 61412 4 gnd
port 2 nsew
rlabel metal3 s 6882 59676 6980 59774 4 vdd
port 1 nsew
rlabel metal3 s 7660 60875 7758 60973 4 vdd
port 1 nsew
rlabel metal3 s 7660 58900 7758 58998 4 vdd
port 1 nsew
rlabel metal3 s 6882 58886 6980 58984 4 vdd
port 1 nsew
rlabel metal3 s 7264 62060 7362 62158 4 gnd
port 2 nsew
rlabel metal3 s 7264 61665 7362 61763 4 gnd
port 2 nsew
rlabel metal3 s 6450 59318 6548 59416 4 vdd
port 1 nsew
rlabel metal3 s 7660 60480 7758 60578 4 vdd
port 1 nsew
rlabel metal3 s 6025 60108 6123 60206 4 gnd
port 2 nsew
rlabel metal3 s 6450 60466 6548 60564 4 vdd
port 1 nsew
rlabel metal3 s 6882 61256 6980 61354 4 vdd
port 1 nsew
rlabel metal3 s 6025 59734 6123 59832 4 gnd
port 2 nsew
rlabel metal3 s 6882 63626 6980 63724 4 vdd
port 1 nsew
rlabel metal3 s 7264 64035 7362 64133 4 gnd
port 2 nsew
rlabel metal3 s 7264 60085 7362 60183 4 gnd
port 2 nsew
rlabel metal3 s 6025 64058 6123 64156 4 gnd
port 2 nsew
rlabel metal3 s 7660 63245 7758 63343 4 vdd
port 1 nsew
rlabel metal3 s 6025 62894 6123 62992 4 gnd
port 2 nsew
rlabel metal3 s 7264 62455 7362 62553 4 gnd
port 2 nsew
rlabel metal3 s 6882 60108 6980 60206 4 vdd
port 1 nsew
rlabel metal3 s 6882 63268 6980 63366 4 vdd
port 1 nsew
rlabel metal3 s 6882 62478 6980 62576 4 vdd
port 1 nsew
rlabel metal3 s 6025 61688 6123 61786 4 gnd
port 2 nsew
rlabel metal3 s 6025 63268 6123 63366 4 gnd
port 2 nsew
rlabel metal3 s 6882 64058 6980 64156 4 vdd
port 1 nsew
rlabel metal3 s 7660 61665 7758 61763 4 vdd
port 1 nsew
rlabel metal3 s 6450 64058 6548 64156 4 vdd
port 1 nsew
rlabel metal3 s 12600 63403 12698 63501 4 gnd
port 2 nsew
rlabel metal3 s 15792 64991 15890 65089 4 vdd
port 1 nsew
rlabel metal3 s 12600 61507 12698 61605 4 gnd
port 2 nsew
rlabel metal3 s 17159 65582 17257 65680 4 vdd
port 1 nsew
rlabel metal3 s 15480 67131 15578 67229 4 gnd
port 2 nsew
rlabel metal3 s 14663 65582 14761 65680 4 vdd
port 1 nsew
rlabel metal3 s 12600 64193 12698 64291 4 gnd
port 2 nsew
rlabel metal3 s 12600 61033 12698 61131 4 gnd
port 2 nsew
rlabel metal3 s 14232 67131 14330 67229 4 gnd
port 2 nsew
rlabel metal3 s 12600 61823 12698 61921 4 gnd
port 2 nsew
rlabel metal3 s 12234 64777 12332 64875 4 gnd
port 2 nsew
rlabel metal3 s 12600 64430 12698 64528 4 gnd
port 2 nsew
rlabel metal3 s 12600 59137 12698 59235 4 gnd
port 2 nsew
rlabel metal3 s 17040 64991 17138 65089 4 vdd
port 1 nsew
rlabel metal3 s 12600 63087 12698 63185 4 gnd
port 2 nsew
rlabel metal3 s 12600 62850 12698 62948 4 gnd
port 2 nsew
rlabel metal3 s 12600 62060 12698 62158 4 gnd
port 2 nsew
rlabel metal3 s 12600 60717 12698 60815 4 gnd
port 2 nsew
rlabel metal3 s 12600 59453 12698 59551 4 gnd
port 2 nsew
rlabel metal3 s 12600 61270 12698 61368 4 gnd
port 2 nsew
rlabel metal3 s 13296 64991 13394 65089 4 vdd
port 1 nsew
rlabel metal3 s 15168 64991 15266 65089 4 vdd
port 1 nsew
rlabel metal3 s 16297 65582 16395 65680 4 vdd
port 1 nsew
rlabel metal3 s 12600 62613 12698 62711 4 gnd
port 2 nsew
rlabel metal3 s 16728 67131 16826 67229 4 gnd
port 2 nsew
rlabel metal3 s 12600 60243 12698 60341 4 gnd
port 2 nsew
rlabel metal3 s 13801 65582 13899 65680 4 vdd
port 1 nsew
rlabel metal3 s 12600 58900 12698 58998 4 gnd
port 2 nsew
rlabel metal3 s 13920 64991 14018 65089 4 vdd
port 1 nsew
rlabel metal3 s 16416 64991 16514 65089 4 vdd
port 1 nsew
rlabel metal3 s 12600 62297 12698 62395 4 gnd
port 2 nsew
rlabel metal3 s 15049 65582 15147 65680 4 vdd
port 1 nsew
rlabel metal3 s 12600 63640 12698 63738 4 gnd
port 2 nsew
rlabel metal3 s 15911 65582 16009 65680 4 vdd
port 1 nsew
rlabel metal3 s 12600 63877 12698 63975 4 gnd
port 2 nsew
rlabel metal3 s 12600 59690 12698 59788 4 gnd
port 2 nsew
rlabel metal3 s 12600 59927 12698 60025 4 gnd
port 2 nsew
rlabel metal3 s 12600 60480 12698 60578 4 gnd
port 2 nsew
rlabel metal3 s 14544 64991 14642 65089 4 vdd
port 1 nsew
rlabel metal3 s 12600 57557 12698 57655 4 gnd
port 2 nsew
rlabel metal3 s 12600 56293 12698 56391 4 gnd
port 2 nsew
rlabel metal3 s 12600 49657 12698 49755 4 gnd
port 2 nsew
rlabel metal3 s 12600 58110 12698 58208 4 gnd
port 2 nsew
rlabel metal3 s 12600 55503 12698 55601 4 gnd
port 2 nsew
rlabel metal3 s 12600 50763 12698 50861 4 gnd
port 2 nsew
rlabel metal3 s 12600 55977 12698 56075 4 gnd
port 2 nsew
rlabel metal3 s 12600 51000 12698 51098 4 gnd
port 2 nsew
rlabel metal3 s 12600 57083 12698 57181 4 gnd
port 2 nsew
rlabel metal3 s 12600 52580 12698 52678 4 gnd
port 2 nsew
rlabel metal3 s 12600 52343 12698 52441 4 gnd
port 2 nsew
rlabel metal3 s 12600 53370 12698 53468 4 gnd
port 2 nsew
rlabel metal3 s 12600 51790 12698 51888 4 gnd
port 2 nsew
rlabel metal3 s 12600 56767 12698 56865 4 gnd
port 2 nsew
rlabel metal3 s 12600 54397 12698 54495 4 gnd
port 2 nsew
rlabel metal3 s 12600 58663 12698 58761 4 gnd
port 2 nsew
rlabel metal3 s 12600 50447 12698 50545 4 gnd
port 2 nsew
rlabel metal3 s 12600 53133 12698 53231 4 gnd
port 2 nsew
rlabel metal3 s 12600 52817 12698 52915 4 gnd
port 2 nsew
rlabel metal3 s 12600 55187 12698 55285 4 gnd
port 2 nsew
rlabel metal3 s 12600 54160 12698 54258 4 gnd
port 2 nsew
rlabel metal3 s 12600 56530 12698 56628 4 gnd
port 2 nsew
rlabel metal3 s 12600 52027 12698 52125 4 gnd
port 2 nsew
rlabel metal3 s 12600 49183 12698 49281 4 gnd
port 2 nsew
rlabel metal3 s 12600 50210 12698 50308 4 gnd
port 2 nsew
rlabel metal3 s 12600 49420 12698 49518 4 gnd
port 2 nsew
rlabel metal3 s 12600 58347 12698 58445 4 gnd
port 2 nsew
rlabel metal3 s 12600 49973 12698 50071 4 gnd
port 2 nsew
rlabel metal3 s 12600 53607 12698 53705 4 gnd
port 2 nsew
rlabel metal3 s 12600 54950 12698 55048 4 gnd
port 2 nsew
rlabel metal3 s 12600 57320 12698 57418 4 gnd
port 2 nsew
rlabel metal3 s 12600 54713 12698 54811 4 gnd
port 2 nsew
rlabel metal3 s 12600 55740 12698 55838 4 gnd
port 2 nsew
rlabel metal3 s 12600 53923 12698 54021 4 gnd
port 2 nsew
rlabel metal3 s 12600 57873 12698 57971 4 gnd
port 2 nsew
rlabel metal3 s 12600 51553 12698 51651 4 gnd
port 2 nsew
rlabel metal3 s 12600 51237 12698 51335 4 gnd
port 2 nsew
rlabel metal3 s 6450 55726 6548 55824 4 vdd
port 1 nsew
rlabel metal3 s 6450 56158 6548 56256 4 vdd
port 1 nsew
rlabel metal3 s 6882 57306 6980 57404 4 vdd
port 1 nsew
rlabel metal3 s 6882 58528 6980 58626 4 vdd
port 1 nsew
rlabel metal3 s 7660 56530 7758 56628 4 vdd
port 1 nsew
rlabel metal3 s 6025 54578 6123 54676 4 gnd
port 2 nsew
rlabel metal3 s 6450 58528 6548 58626 4 vdd
port 1 nsew
rlabel metal3 s 6450 57738 6548 57836 4 vdd
port 1 nsew
rlabel metal3 s 7264 55740 7362 55838 4 gnd
port 2 nsew
rlabel metal3 s 6025 56948 6123 57046 4 gnd
port 2 nsew
rlabel metal3 s 7264 57715 7362 57813 4 gnd
port 2 nsew
rlabel metal3 s 7660 56925 7758 57023 4 vdd
port 1 nsew
rlabel metal3 s 6450 54936 6548 55034 4 vdd
port 1 nsew
rlabel metal3 s 7660 58110 7758 58208 4 vdd
port 1 nsew
rlabel metal3 s 7264 57320 7362 57418 4 gnd
port 2 nsew
rlabel metal3 s 6450 58096 6548 58194 4 vdd
port 1 nsew
rlabel metal3 s 7660 57715 7758 57813 4 vdd
port 1 nsew
rlabel metal3 s 6882 56948 6980 57046 4 vdd
port 1 nsew
rlabel metal3 s 7660 57320 7758 57418 4 vdd
port 1 nsew
rlabel metal3 s 6025 55368 6123 55466 4 gnd
port 2 nsew
rlabel metal3 s 7660 55345 7758 55443 4 vdd
port 1 nsew
rlabel metal3 s 6025 56158 6123 56256 4 gnd
port 2 nsew
rlabel metal3 s 6882 54936 6980 55034 4 vdd
port 1 nsew
rlabel metal3 s 6450 56516 6548 56614 4 vdd
port 1 nsew
rlabel metal3 s 7264 58110 7362 58208 4 gnd
port 2 nsew
rlabel metal3 s 6025 56574 6123 56672 4 gnd
port 2 nsew
rlabel metal3 s 7264 58505 7362 58603 4 gnd
port 2 nsew
rlabel metal3 s 6025 54204 6123 54302 4 gnd
port 2 nsew
rlabel metal3 s 6882 55368 6980 55466 4 vdd
port 1 nsew
rlabel metal3 s 7264 54160 7362 54258 4 gnd
port 2 nsew
rlabel metal3 s 6882 56516 6980 56614 4 vdd
port 1 nsew
rlabel metal3 s 7660 56135 7758 56233 4 vdd
port 1 nsew
rlabel metal3 s 7264 56530 7362 56628 4 gnd
port 2 nsew
rlabel metal3 s 7660 54160 7758 54258 4 vdd
port 1 nsew
rlabel metal3 s 6882 57738 6980 57836 4 vdd
port 1 nsew
rlabel metal3 s 6025 58528 6123 58626 4 gnd
port 2 nsew
rlabel metal3 s 6450 54146 6548 54244 4 vdd
port 1 nsew
rlabel metal3 s 6025 55784 6123 55882 4 gnd
port 2 nsew
rlabel metal3 s 6025 58154 6123 58252 4 gnd
port 2 nsew
rlabel metal3 s 7264 54950 7362 55048 4 gnd
port 2 nsew
rlabel metal3 s 7264 54555 7362 54653 4 gnd
port 2 nsew
rlabel metal3 s 6882 54146 6980 54244 4 vdd
port 1 nsew
rlabel metal3 s 6450 56948 6548 57046 4 vdd
port 1 nsew
rlabel metal3 s 7264 56135 7362 56233 4 gnd
port 2 nsew
rlabel metal3 s 6882 55726 6980 55824 4 vdd
port 1 nsew
rlabel metal3 s 6450 54578 6548 54676 4 vdd
port 1 nsew
rlabel metal3 s 7660 58505 7758 58603 4 vdd
port 1 nsew
rlabel metal3 s 6882 54578 6980 54676 4 vdd
port 1 nsew
rlabel metal3 s 7660 54950 7758 55048 4 vdd
port 1 nsew
rlabel metal3 s 6025 57738 6123 57836 4 gnd
port 2 nsew
rlabel metal3 s 6450 57306 6548 57404 4 vdd
port 1 nsew
rlabel metal3 s 7660 54555 7758 54653 4 vdd
port 1 nsew
rlabel metal3 s 6025 54994 6123 55092 4 gnd
port 2 nsew
rlabel metal3 s 7660 55740 7758 55838 4 vdd
port 1 nsew
rlabel metal3 s 6450 55368 6548 55466 4 vdd
port 1 nsew
rlabel metal3 s 7264 55345 7362 55443 4 gnd
port 2 nsew
rlabel metal3 s 6882 56158 6980 56256 4 vdd
port 1 nsew
rlabel metal3 s 6882 58096 6980 58194 4 vdd
port 1 nsew
rlabel metal3 s 6025 57364 6123 57462 4 gnd
port 2 nsew
rlabel metal3 s 7264 56925 7362 57023 4 gnd
port 2 nsew
rlabel metal3 s 7660 52975 7758 53073 4 vdd
port 1 nsew
rlabel metal3 s 7264 52975 7362 53073 4 gnd
port 2 nsew
rlabel metal3 s 6882 53356 6980 53454 4 vdd
port 1 nsew
rlabel metal3 s 6450 52208 6548 52306 4 vdd
port 1 nsew
rlabel metal3 s 7264 50605 7362 50703 4 gnd
port 2 nsew
rlabel metal3 s 7660 53765 7758 53863 4 vdd
port 1 nsew
rlabel metal3 s 6025 51834 6123 51932 4 gnd
port 2 nsew
rlabel metal3 s 7660 52580 7758 52678 4 vdd
port 1 nsew
rlabel metal3 s 6450 49838 6548 49936 4 vdd
port 1 nsew
rlabel metal3 s 6450 49406 6548 49504 4 vdd
port 1 nsew
rlabel metal3 s 7264 53765 7362 53863 4 gnd
port 2 nsew
rlabel metal3 s 6025 49048 6123 49146 4 gnd
port 2 nsew
rlabel metal3 s 7264 52185 7362 52283 4 gnd
port 2 nsew
rlabel metal3 s 6025 52998 6123 53096 4 gnd
port 2 nsew
rlabel metal3 s 7264 50210 7362 50308 4 gnd
port 2 nsew
rlabel metal3 s 6025 49464 6123 49562 4 gnd
port 2 nsew
rlabel metal3 s 6450 52566 6548 52664 4 vdd
port 1 nsew
rlabel metal3 s 6025 51044 6123 51142 4 gnd
port 2 nsew
rlabel metal3 s 6450 49048 6548 49146 4 vdd
port 1 nsew
rlabel metal3 s 7264 51395 7362 51493 4 gnd
port 2 nsew
rlabel metal3 s 6025 53414 6123 53512 4 gnd
port 2 nsew
rlabel metal3 s 7264 49815 7362 49913 4 gnd
port 2 nsew
rlabel metal3 s 7660 51000 7758 51098 4 vdd
port 1 nsew
rlabel metal3 s 7264 51790 7362 51888 4 gnd
port 2 nsew
rlabel metal3 s 6882 52998 6980 53096 4 vdd
port 1 nsew
rlabel metal3 s 6882 49406 6980 49504 4 vdd
port 1 nsew
rlabel metal3 s 6450 50196 6548 50294 4 vdd
port 1 nsew
rlabel metal3 s 6882 52208 6980 52306 4 vdd
port 1 nsew
rlabel metal3 s 6450 50986 6548 51084 4 vdd
port 1 nsew
rlabel metal3 s 6882 52566 6980 52664 4 vdd
port 1 nsew
rlabel metal3 s 6025 50254 6123 50352 4 gnd
port 2 nsew
rlabel metal3 s 7264 51000 7362 51098 4 gnd
port 2 nsew
rlabel metal3 s 7660 53370 7758 53468 4 vdd
port 1 nsew
rlabel metal3 s 6450 50628 6548 50726 4 vdd
port 1 nsew
rlabel metal3 s 6882 50196 6980 50294 4 vdd
port 1 nsew
rlabel metal3 s 6025 51418 6123 51516 4 gnd
port 2 nsew
rlabel metal3 s 7660 51790 7758 51888 4 vdd
port 1 nsew
rlabel metal3 s 6025 50628 6123 50726 4 gnd
port 2 nsew
rlabel metal3 s 7264 49025 7362 49123 4 gnd
port 2 nsew
rlabel metal3 s 7264 52580 7362 52678 4 gnd
port 2 nsew
rlabel metal3 s 6025 53788 6123 53886 4 gnd
port 2 nsew
rlabel metal3 s 6882 51776 6980 51874 4 vdd
port 1 nsew
rlabel metal3 s 6882 50986 6980 51084 4 vdd
port 1 nsew
rlabel metal3 s 6450 52998 6548 53096 4 vdd
port 1 nsew
rlabel metal3 s 6450 51776 6548 51874 4 vdd
port 1 nsew
rlabel metal3 s 7660 49815 7758 49913 4 vdd
port 1 nsew
rlabel metal3 s 7660 51395 7758 51493 4 vdd
port 1 nsew
rlabel metal3 s 6025 49838 6123 49936 4 gnd
port 2 nsew
rlabel metal3 s 7264 49420 7362 49518 4 gnd
port 2 nsew
rlabel metal3 s 6450 53356 6548 53454 4 vdd
port 1 nsew
rlabel metal3 s 7660 52185 7758 52283 4 vdd
port 1 nsew
rlabel metal3 s 7660 49420 7758 49518 4 vdd
port 1 nsew
rlabel metal3 s 6882 49838 6980 49936 4 vdd
port 1 nsew
rlabel metal3 s 7660 49025 7758 49123 4 vdd
port 1 nsew
rlabel metal3 s 6025 52624 6123 52722 4 gnd
port 2 nsew
rlabel metal3 s 7660 50605 7758 50703 4 vdd
port 1 nsew
rlabel metal3 s 7264 53370 7362 53468 4 gnd
port 2 nsew
rlabel metal3 s 6882 51418 6980 51516 4 vdd
port 1 nsew
rlabel metal3 s 7660 50210 7758 50308 4 vdd
port 1 nsew
rlabel metal3 s 6882 50628 6980 50726 4 vdd
port 1 nsew
rlabel metal3 s 6882 53788 6980 53886 4 vdd
port 1 nsew
rlabel metal3 s 6450 53788 6548 53886 4 vdd
port 1 nsew
rlabel metal3 s 6450 51418 6548 51516 4 vdd
port 1 nsew
rlabel metal3 s 6882 49048 6980 49146 4 vdd
port 1 nsew
rlabel metal3 s 6025 52208 6123 52306 4 gnd
port 2 nsew
rlabel metal3 s 6450 47036 6548 47134 4 vdd
port 1 nsew
rlabel metal3 s 6025 45888 6123 45986 4 gnd
port 2 nsew
rlabel metal3 s 6450 47826 6548 47924 4 vdd
port 1 nsew
rlabel metal3 s 6025 46678 6123 46776 4 gnd
port 2 nsew
rlabel metal3 s 6450 48616 6548 48714 4 vdd
port 1 nsew
rlabel metal3 s 6450 44666 6548 44764 4 vdd
port 1 nsew
rlabel metal3 s 7660 45075 7758 45173 4 vdd
port 1 nsew
rlabel metal3 s 7264 45470 7362 45568 4 gnd
port 2 nsew
rlabel metal3 s 6882 47468 6980 47566 4 vdd
port 1 nsew
rlabel metal3 s 6025 44724 6123 44822 4 gnd
port 2 nsew
rlabel metal3 s 6450 46246 6548 46344 4 vdd
port 1 nsew
rlabel metal3 s 6025 47468 6123 47566 4 gnd
port 2 nsew
rlabel metal3 s 7660 44680 7758 44778 4 vdd
port 1 nsew
rlabel metal3 s 7264 46260 7362 46358 4 gnd
port 2 nsew
rlabel metal3 s 7264 47840 7362 47938 4 gnd
port 2 nsew
rlabel metal3 s 7660 45470 7758 45568 4 vdd
port 1 nsew
rlabel metal3 s 6882 45098 6980 45196 4 vdd
port 1 nsew
rlabel metal3 s 6450 45888 6548 45986 4 vdd
port 1 nsew
rlabel metal3 s 7264 47050 7362 47148 4 gnd
port 2 nsew
rlabel metal3 s 7660 45865 7758 45963 4 vdd
port 1 nsew
rlabel metal3 s 6882 46246 6980 46344 4 vdd
port 1 nsew
rlabel metal3 s 7264 45075 7362 45173 4 gnd
port 2 nsew
rlabel metal3 s 6882 47826 6980 47924 4 vdd
port 1 nsew
rlabel metal3 s 6882 47036 6980 47134 4 vdd
port 1 nsew
rlabel metal3 s 6025 48258 6123 48356 4 gnd
port 2 nsew
rlabel metal3 s 6882 44666 6980 44764 4 vdd
port 1 nsew
rlabel metal3 s 7660 44285 7758 44383 4 vdd
port 1 nsew
rlabel metal3 s 6025 46304 6123 46402 4 gnd
port 2 nsew
rlabel metal3 s 6882 48258 6980 48356 4 vdd
port 1 nsew
rlabel metal3 s 7264 44285 7362 44383 4 gnd
port 2 nsew
rlabel metal3 s 7660 48235 7758 48333 4 vdd
port 1 nsew
rlabel metal3 s 7264 44680 7362 44778 4 gnd
port 2 nsew
rlabel metal3 s 6025 45098 6123 45196 4 gnd
port 2 nsew
rlabel metal3 s 6025 47094 6123 47192 4 gnd
port 2 nsew
rlabel metal3 s 7264 45865 7362 45963 4 gnd
port 2 nsew
rlabel metal3 s 7660 46655 7758 46753 4 vdd
port 1 nsew
rlabel metal3 s 7264 46655 7362 46753 4 gnd
port 2 nsew
rlabel metal3 s 6882 44308 6980 44406 4 vdd
port 1 nsew
rlabel metal3 s 7660 46260 7758 46358 4 vdd
port 1 nsew
rlabel metal3 s 6450 45098 6548 45196 4 vdd
port 1 nsew
rlabel metal3 s 7660 47840 7758 47938 4 vdd
port 1 nsew
rlabel metal3 s 6450 48258 6548 48356 4 vdd
port 1 nsew
rlabel metal3 s 6450 46678 6548 46776 4 vdd
port 1 nsew
rlabel metal3 s 7660 47445 7758 47543 4 vdd
port 1 nsew
rlabel metal3 s 7660 48630 7758 48728 4 vdd
port 1 nsew
rlabel metal3 s 6882 46678 6980 46776 4 vdd
port 1 nsew
rlabel metal3 s 6450 47468 6548 47566 4 vdd
port 1 nsew
rlabel metal3 s 6450 44308 6548 44406 4 vdd
port 1 nsew
rlabel metal3 s 6025 48674 6123 48772 4 gnd
port 2 nsew
rlabel metal3 s 6882 48616 6980 48714 4 vdd
port 1 nsew
rlabel metal3 s 6025 47884 6123 47982 4 gnd
port 2 nsew
rlabel metal3 s 7264 48235 7362 48333 4 gnd
port 2 nsew
rlabel metal3 s 6450 45456 6548 45554 4 vdd
port 1 nsew
rlabel metal3 s 6025 44308 6123 44406 4 gnd
port 2 nsew
rlabel metal3 s 6882 45456 6980 45554 4 vdd
port 1 nsew
rlabel metal3 s 6882 45888 6980 45986 4 vdd
port 1 nsew
rlabel metal3 s 6025 45514 6123 45612 4 gnd
port 2 nsew
rlabel metal3 s 7264 48630 7362 48728 4 gnd
port 2 nsew
rlabel metal3 s 7264 47445 7362 47543 4 gnd
port 2 nsew
rlabel metal3 s 7660 47050 7758 47148 4 vdd
port 1 nsew
rlabel metal3 s 6450 42296 6548 42394 4 vdd
port 1 nsew
rlabel metal3 s 6882 42728 6980 42826 4 vdd
port 1 nsew
rlabel metal3 s 7660 39545 7758 39643 4 vdd
port 1 nsew
rlabel metal3 s 7264 39545 7362 39643 4 gnd
port 2 nsew
rlabel metal3 s 6450 40358 6548 40456 4 vdd
port 1 nsew
rlabel metal3 s 7264 41520 7362 41618 4 gnd
port 2 nsew
rlabel metal3 s 6450 43876 6548 43974 4 vdd
port 1 nsew
rlabel metal3 s 6025 43934 6123 44032 4 gnd
port 2 nsew
rlabel metal3 s 6882 41506 6980 41604 4 vdd
port 1 nsew
rlabel metal3 s 7660 41915 7758 42013 4 vdd
port 1 nsew
rlabel metal3 s 6450 42728 6548 42826 4 vdd
port 1 nsew
rlabel metal3 s 7264 41125 7362 41223 4 gnd
port 2 nsew
rlabel metal3 s 6025 43518 6123 43616 4 gnd
port 2 nsew
rlabel metal3 s 7264 43890 7362 43988 4 gnd
port 2 nsew
rlabel metal3 s 6882 41938 6980 42036 4 vdd
port 1 nsew
rlabel metal3 s 6882 41148 6980 41246 4 vdd
port 1 nsew
rlabel metal3 s 7660 41125 7758 41223 4 vdd
port 1 nsew
rlabel metal3 s 6882 43518 6980 43616 4 vdd
port 1 nsew
rlabel metal3 s 6025 43144 6123 43242 4 gnd
port 2 nsew
rlabel metal3 s 6025 42728 6123 42826 4 gnd
port 2 nsew
rlabel metal3 s 6025 41938 6123 42036 4 gnd
port 2 nsew
rlabel metal3 s 7660 40730 7758 40828 4 vdd
port 1 nsew
rlabel metal3 s 6450 39568 6548 39666 4 vdd
port 1 nsew
rlabel metal3 s 6450 41506 6548 41604 4 vdd
port 1 nsew
rlabel metal3 s 6025 41148 6123 41246 4 gnd
port 2 nsew
rlabel metal3 s 7660 43890 7758 43988 4 vdd
port 1 nsew
rlabel metal3 s 6025 42354 6123 42452 4 gnd
port 2 nsew
rlabel metal3 s 7660 43100 7758 43198 4 vdd
port 1 nsew
rlabel metal3 s 6450 39926 6548 40024 4 vdd
port 1 nsew
rlabel metal3 s 7660 42705 7758 42803 4 vdd
port 1 nsew
rlabel metal3 s 7264 39940 7362 40038 4 gnd
port 2 nsew
rlabel metal3 s 7660 41520 7758 41618 4 vdd
port 1 nsew
rlabel metal3 s 6882 43086 6980 43184 4 vdd
port 1 nsew
rlabel metal3 s 7264 42705 7362 42803 4 gnd
port 2 nsew
rlabel metal3 s 6025 39984 6123 40082 4 gnd
port 2 nsew
rlabel metal3 s 6882 42296 6980 42394 4 vdd
port 1 nsew
rlabel metal3 s 6882 40716 6980 40814 4 vdd
port 1 nsew
rlabel metal3 s 7264 40730 7362 40828 4 gnd
port 2 nsew
rlabel metal3 s 6882 43876 6980 43974 4 vdd
port 1 nsew
rlabel metal3 s 6882 40358 6980 40456 4 vdd
port 1 nsew
rlabel metal3 s 7264 43495 7362 43593 4 gnd
port 2 nsew
rlabel metal3 s 6450 41938 6548 42036 4 vdd
port 1 nsew
rlabel metal3 s 6882 39568 6980 39666 4 vdd
port 1 nsew
rlabel metal3 s 7264 42310 7362 42408 4 gnd
port 2 nsew
rlabel metal3 s 6025 39568 6123 39666 4 gnd
port 2 nsew
rlabel metal3 s 6450 41148 6548 41246 4 vdd
port 1 nsew
rlabel metal3 s 6025 40774 6123 40872 4 gnd
port 2 nsew
rlabel metal3 s 6882 39926 6980 40024 4 vdd
port 1 nsew
rlabel metal3 s 7264 41915 7362 42013 4 gnd
port 2 nsew
rlabel metal3 s 7264 43100 7362 43198 4 gnd
port 2 nsew
rlabel metal3 s 6025 39194 6123 39292 4 gnd
port 2 nsew
rlabel metal3 s 6450 43518 6548 43616 4 vdd
port 1 nsew
rlabel metal3 s 6025 41564 6123 41662 4 gnd
port 2 nsew
rlabel metal3 s 7660 42310 7758 42408 4 vdd
port 1 nsew
rlabel metal3 s 6025 40358 6123 40456 4 gnd
port 2 nsew
rlabel metal3 s 7660 40335 7758 40433 4 vdd
port 1 nsew
rlabel metal3 s 6450 43086 6548 43184 4 vdd
port 1 nsew
rlabel metal3 s 7264 40335 7362 40433 4 gnd
port 2 nsew
rlabel metal3 s 7660 39940 7758 40038 4 vdd
port 1 nsew
rlabel metal3 s 7660 43495 7758 43593 4 vdd
port 1 nsew
rlabel metal3 s 6450 40716 6548 40814 4 vdd
port 1 nsew
rlabel metal3 s 12600 46497 12698 46595 4 gnd
port 2 nsew
rlabel metal3 s 12600 39940 12698 40038 4 gnd
port 2 nsew
rlabel metal3 s 12600 43890 12698 43988 4 gnd
port 2 nsew
rlabel metal3 s 12600 42863 12698 42961 4 gnd
port 2 nsew
rlabel metal3 s 12600 42073 12698 42171 4 gnd
port 2 nsew
rlabel metal3 s 12600 48630 12698 48728 4 gnd
port 2 nsew
rlabel metal3 s 12600 46813 12698 46911 4 gnd
port 2 nsew
rlabel metal3 s 12600 47603 12698 47701 4 gnd
port 2 nsew
rlabel metal3 s 12600 45233 12698 45331 4 gnd
port 2 nsew
rlabel metal3 s 12600 47287 12698 47385 4 gnd
port 2 nsew
rlabel metal3 s 12600 48077 12698 48175 4 gnd
port 2 nsew
rlabel metal3 s 12600 41757 12698 41855 4 gnd
port 2 nsew
rlabel metal3 s 12600 46023 12698 46121 4 gnd
port 2 nsew
rlabel metal3 s 12600 45707 12698 45805 4 gnd
port 2 nsew
rlabel metal3 s 12600 39703 12698 39801 4 gnd
port 2 nsew
rlabel metal3 s 12600 44680 12698 44778 4 gnd
port 2 nsew
rlabel metal3 s 12600 43337 12698 43435 4 gnd
port 2 nsew
rlabel metal3 s 12600 46260 12698 46358 4 gnd
port 2 nsew
rlabel metal3 s 12600 42310 12698 42408 4 gnd
port 2 nsew
rlabel metal3 s 12600 48393 12698 48491 4 gnd
port 2 nsew
rlabel metal3 s 12600 48867 12698 48965 4 gnd
port 2 nsew
rlabel metal3 s 12600 45470 12698 45568 4 gnd
port 2 nsew
rlabel metal3 s 12600 40730 12698 40828 4 gnd
port 2 nsew
rlabel metal3 s 12600 43653 12698 43751 4 gnd
port 2 nsew
rlabel metal3 s 12600 47050 12698 47148 4 gnd
port 2 nsew
rlabel metal3 s 12600 43100 12698 43198 4 gnd
port 2 nsew
rlabel metal3 s 12600 42547 12698 42645 4 gnd
port 2 nsew
rlabel metal3 s 12600 40967 12698 41065 4 gnd
port 2 nsew
rlabel metal3 s 12600 44127 12698 44225 4 gnd
port 2 nsew
rlabel metal3 s 12600 41283 12698 41381 4 gnd
port 2 nsew
rlabel metal3 s 12600 41520 12698 41618 4 gnd
port 2 nsew
rlabel metal3 s 12600 44917 12698 45015 4 gnd
port 2 nsew
rlabel metal3 s 12600 47840 12698 47938 4 gnd
port 2 nsew
rlabel metal3 s 12600 40493 12698 40591 4 gnd
port 2 nsew
rlabel metal3 s 12600 39387 12698 39485 4 gnd
port 2 nsew
rlabel metal3 s 12600 40177 12698 40275 4 gnd
port 2 nsew
rlabel metal3 s 12600 44443 12698 44541 4 gnd
port 2 nsew
rlabel metal3 s 12600 35200 12698 35298 4 gnd
port 2 nsew
rlabel metal3 s 12600 29907 12698 30005 4 gnd
port 2 nsew
rlabel metal3 s 12600 38913 12698 39011 4 gnd
port 2 nsew
rlabel metal3 s 12600 30697 12698 30795 4 gnd
port 2 nsew
rlabel metal3 s 12600 35990 12698 36088 4 gnd
port 2 nsew
rlabel metal3 s 12600 36543 12698 36641 4 gnd
port 2 nsew
rlabel metal3 s 12600 39150 12698 39248 4 gnd
port 2 nsew
rlabel metal3 s 12600 31250 12698 31348 4 gnd
port 2 nsew
rlabel metal3 s 12600 35437 12698 35535 4 gnd
port 2 nsew
rlabel metal3 s 12600 35753 12698 35851 4 gnd
port 2 nsew
rlabel metal3 s 12600 33383 12698 33481 4 gnd
port 2 nsew
rlabel metal3 s 12600 29433 12698 29531 4 gnd
port 2 nsew
rlabel metal3 s 12600 38123 12698 38221 4 gnd
port 2 nsew
rlabel metal3 s 12600 34647 12698 34745 4 gnd
port 2 nsew
rlabel metal3 s 12600 29670 12698 29768 4 gnd
port 2 nsew
rlabel metal3 s 12600 33620 12698 33718 4 gnd
port 2 nsew
rlabel metal3 s 11208 39150 11306 39248 4 vdd
port 1 nsew
rlabel metal3 s 12600 33857 12698 33955 4 gnd
port 2 nsew
rlabel metal3 s 12600 32830 12698 32928 4 gnd
port 2 nsew
rlabel metal3 s 12600 32040 12698 32138 4 gnd
port 2 nsew
rlabel metal3 s 12600 38360 12698 38458 4 gnd
port 2 nsew
rlabel metal3 s 12600 37570 12698 37668 4 gnd
port 2 nsew
rlabel metal3 s 12600 36780 12698 36878 4 gnd
port 2 nsew
rlabel metal3 s 12600 31803 12698 31901 4 gnd
port 2 nsew
rlabel metal3 s 12600 36227 12698 36325 4 gnd
port 2 nsew
rlabel metal3 s 12600 34410 12698 34508 4 gnd
port 2 nsew
rlabel metal3 s 9560 39150 9658 39248 4 gnd
port 2 nsew
rlabel metal3 s 12600 30223 12698 30321 4 gnd
port 2 nsew
rlabel metal3 s 12600 31013 12698 31111 4 gnd
port 2 nsew
rlabel metal3 s 12600 31487 12698 31585 4 gnd
port 2 nsew
rlabel metal3 s 12600 37807 12698 37905 4 gnd
port 2 nsew
rlabel metal3 s 12600 37017 12698 37115 4 gnd
port 2 nsew
rlabel metal3 s 12600 30460 12698 30558 4 gnd
port 2 nsew
rlabel metal3 s 12600 37333 12698 37431 4 gnd
port 2 nsew
rlabel metal3 s 12600 32593 12698 32691 4 gnd
port 2 nsew
rlabel metal3 s 12600 34173 12698 34271 4 gnd
port 2 nsew
rlabel metal3 s 12600 38597 12698 38695 4 gnd
port 2 nsew
rlabel metal3 s 12600 33067 12698 33165 4 gnd
port 2 nsew
rlabel metal3 s 12600 34963 12698 35061 4 gnd
port 2 nsew
rlabel metal3 s 12600 32277 12698 32375 4 gnd
port 2 nsew
rlabel metal3 s 7660 39150 7758 39248 4 vdd
port 1 nsew
rlabel metal3 s 6882 35618 6980 35716 4 vdd
port 1 nsew
rlabel metal3 s 6450 37988 6548 38086 4 vdd
port 1 nsew
rlabel metal3 s 6450 38778 6548 38876 4 vdd
port 1 nsew
rlabel metal3 s 7264 38360 7362 38458 4 gnd
port 2 nsew
rlabel metal3 s 6450 38346 6548 38444 4 vdd
port 1 nsew
rlabel metal3 s 6882 37988 6980 38086 4 vdd
port 1 nsew
rlabel metal3 s 7264 35990 7362 36088 4 gnd
port 2 nsew
rlabel metal3 s 6450 35186 6548 35284 4 vdd
port 1 nsew
rlabel metal3 s 6882 34828 6980 34926 4 vdd
port 1 nsew
rlabel metal3 s 6882 38346 6980 38444 4 vdd
port 1 nsew
rlabel metal3 s 6450 37198 6548 37296 4 vdd
port 1 nsew
rlabel metal3 s 6882 39136 6980 39234 4 vdd
port 1 nsew
rlabel metal3 s 6882 35186 6980 35284 4 vdd
port 1 nsew
rlabel metal3 s 7264 34805 7362 34903 4 gnd
port 2 nsew
rlabel metal3 s 7660 34410 7758 34508 4 vdd
port 1 nsew
rlabel metal3 s 7660 35990 7758 36088 4 vdd
port 1 nsew
rlabel metal3 s 6450 39136 6548 39234 4 vdd
port 1 nsew
rlabel metal3 s 7264 37965 7362 38063 4 gnd
port 2 nsew
rlabel metal3 s 6882 36408 6980 36506 4 vdd
port 1 nsew
rlabel metal3 s 6450 37556 6548 37654 4 vdd
port 1 nsew
rlabel metal3 s 7660 34805 7758 34903 4 vdd
port 1 nsew
rlabel metal3 s 6882 35976 6980 36074 4 vdd
port 1 nsew
rlabel metal3 s 7264 37570 7362 37668 4 gnd
port 2 nsew
rlabel metal3 s 7660 36385 7758 36483 4 vdd
port 1 nsew
rlabel metal3 s 7660 38755 7758 38853 4 vdd
port 1 nsew
rlabel metal3 s 7660 35595 7758 35693 4 vdd
port 1 nsew
rlabel metal3 s 6025 37614 6123 37712 4 gnd
port 2 nsew
rlabel metal3 s 7660 37570 7758 37668 4 vdd
port 1 nsew
rlabel metal3 s 7660 37965 7758 38063 4 vdd
port 1 nsew
rlabel metal3 s 6025 34828 6123 34926 4 gnd
port 2 nsew
rlabel metal3 s 6450 36766 6548 36864 4 vdd
port 1 nsew
rlabel metal3 s 7660 37175 7758 37273 4 vdd
port 1 nsew
rlabel metal3 s 6450 34396 6548 34494 4 vdd
port 1 nsew
rlabel metal3 s 6882 36766 6980 36864 4 vdd
port 1 nsew
rlabel metal3 s 7264 39150 7362 39248 4 gnd
port 2 nsew
rlabel metal3 s 6450 34828 6548 34926 4 vdd
port 1 nsew
rlabel metal3 s 6882 37198 6980 37296 4 vdd
port 1 nsew
rlabel metal3 s 6025 38778 6123 38876 4 gnd
port 2 nsew
rlabel metal3 s 7264 38755 7362 38853 4 gnd
port 2 nsew
rlabel metal3 s 6882 37556 6980 37654 4 vdd
port 1 nsew
rlabel metal3 s 6882 34396 6980 34494 4 vdd
port 1 nsew
rlabel metal3 s 6025 34454 6123 34552 4 gnd
port 2 nsew
rlabel metal3 s 6882 38778 6980 38876 4 vdd
port 1 nsew
rlabel metal3 s 7264 37175 7362 37273 4 gnd
port 2 nsew
rlabel metal3 s 7264 36780 7362 36878 4 gnd
port 2 nsew
rlabel metal3 s 6450 36408 6548 36506 4 vdd
port 1 nsew
rlabel metal3 s 7264 34410 7362 34508 4 gnd
port 2 nsew
rlabel metal3 s 6025 35244 6123 35342 4 gnd
port 2 nsew
rlabel metal3 s 7264 35200 7362 35298 4 gnd
port 2 nsew
rlabel metal3 s 6025 37198 6123 37296 4 gnd
port 2 nsew
rlabel metal3 s 6025 36824 6123 36922 4 gnd
port 2 nsew
rlabel metal3 s 6025 36408 6123 36506 4 gnd
port 2 nsew
rlabel metal3 s 7264 35595 7362 35693 4 gnd
port 2 nsew
rlabel metal3 s 6025 35618 6123 35716 4 gnd
port 2 nsew
rlabel metal3 s 7264 36385 7362 36483 4 gnd
port 2 nsew
rlabel metal3 s 8092 39135 8190 39233 4 gnd
port 2 nsew
rlabel metal3 s 6025 36034 6123 36132 4 gnd
port 2 nsew
rlabel metal3 s 7660 36780 7758 36878 4 vdd
port 1 nsew
rlabel metal3 s 8517 39134 8615 39232 4 vdd
port 1 nsew
rlabel metal3 s 6450 35976 6548 36074 4 vdd
port 1 nsew
rlabel metal3 s 7660 35200 7758 35298 4 vdd
port 1 nsew
rlabel metal3 s 6450 35618 6548 35716 4 vdd
port 1 nsew
rlabel metal3 s 7660 38360 7758 38458 4 vdd
port 1 nsew
rlabel metal3 s 6025 37988 6123 38086 4 gnd
port 2 nsew
rlabel metal3 s 6025 38404 6123 38502 4 gnd
port 2 nsew
rlabel metal3 s 6025 31294 6123 31392 4 gnd
port 2 nsew
rlabel metal3 s 7660 33225 7758 33323 4 vdd
port 1 nsew
rlabel metal3 s 7264 31645 7362 31743 4 gnd
port 2 nsew
rlabel metal3 s 6025 31668 6123 31766 4 gnd
port 2 nsew
rlabel metal3 s 7264 32040 7362 32138 4 gnd
port 2 nsew
rlabel metal3 s 6882 31236 6980 31334 4 vdd
port 1 nsew
rlabel metal3 s 7264 29670 7362 29768 4 gnd
port 2 nsew
rlabel metal3 s 6450 32816 6548 32914 4 vdd
port 1 nsew
rlabel metal3 s 6882 32026 6980 32124 4 vdd
port 1 nsew
rlabel metal3 s 6450 31668 6548 31766 4 vdd
port 1 nsew
rlabel metal3 s 6882 33606 6980 33704 4 vdd
port 1 nsew
rlabel metal3 s 6450 29656 6548 29754 4 vdd
port 1 nsew
rlabel metal3 s 6025 34038 6123 34136 4 gnd
port 2 nsew
rlabel metal3 s 6025 30088 6123 30186 4 gnd
port 2 nsew
rlabel metal3 s 7660 33620 7758 33718 4 vdd
port 1 nsew
rlabel metal3 s 6882 32816 6980 32914 4 vdd
port 1 nsew
rlabel metal3 s 7264 30855 7362 30953 4 gnd
port 2 nsew
rlabel metal3 s 6450 32026 6548 32124 4 vdd
port 1 nsew
rlabel metal3 s 7264 30065 7362 30163 4 gnd
port 2 nsew
rlabel metal3 s 6025 30878 6123 30976 4 gnd
port 2 nsew
rlabel metal3 s 7264 33225 7362 33323 4 gnd
port 2 nsew
rlabel metal3 s 7264 32435 7362 32533 4 gnd
port 2 nsew
rlabel metal3 s 7660 30855 7758 30953 4 vdd
port 1 nsew
rlabel metal3 s 7660 30065 7758 30163 4 vdd
port 1 nsew
rlabel metal3 s 7264 34015 7362 34113 4 gnd
port 2 nsew
rlabel metal3 s 6882 30878 6980 30976 4 vdd
port 1 nsew
rlabel metal3 s 6882 29656 6980 29754 4 vdd
port 1 nsew
rlabel metal3 s 6882 31668 6980 31766 4 vdd
port 1 nsew
rlabel metal3 s 6025 32458 6123 32556 4 gnd
port 2 nsew
rlabel metal3 s 6450 30446 6548 30544 4 vdd
port 1 nsew
rlabel metal3 s 6882 30088 6980 30186 4 vdd
port 1 nsew
rlabel metal3 s 7264 31250 7362 31348 4 gnd
port 2 nsew
rlabel metal3 s 6450 34038 6548 34136 4 vdd
port 1 nsew
rlabel metal3 s 7660 30460 7758 30558 4 vdd
port 1 nsew
rlabel metal3 s 6025 32084 6123 32182 4 gnd
port 2 nsew
rlabel metal3 s 7660 31250 7758 31348 4 vdd
port 1 nsew
rlabel metal3 s 6882 32458 6980 32556 4 vdd
port 1 nsew
rlabel metal3 s 6025 29714 6123 29812 4 gnd
port 2 nsew
rlabel metal3 s 7660 29670 7758 29768 4 vdd
port 1 nsew
rlabel metal3 s 7264 32830 7362 32928 4 gnd
port 2 nsew
rlabel metal3 s 7660 32040 7758 32138 4 vdd
port 1 nsew
rlabel metal3 s 6882 30446 6980 30544 4 vdd
port 1 nsew
rlabel metal3 s 6882 33248 6980 33346 4 vdd
port 1 nsew
rlabel metal3 s 6450 33606 6548 33704 4 vdd
port 1 nsew
rlabel metal3 s 6882 34038 6980 34136 4 vdd
port 1 nsew
rlabel metal3 s 6450 31236 6548 31334 4 vdd
port 1 nsew
rlabel metal3 s 6450 32458 6548 32556 4 vdd
port 1 nsew
rlabel metal3 s 6025 30504 6123 30602 4 gnd
port 2 nsew
rlabel metal3 s 6025 32874 6123 32972 4 gnd
port 2 nsew
rlabel metal3 s 6450 30088 6548 30186 4 vdd
port 1 nsew
rlabel metal3 s 6025 33248 6123 33346 4 gnd
port 2 nsew
rlabel metal3 s 7660 32435 7758 32533 4 vdd
port 1 nsew
rlabel metal3 s 6025 33664 6123 33762 4 gnd
port 2 nsew
rlabel metal3 s 6450 33248 6548 33346 4 vdd
port 1 nsew
rlabel metal3 s 7264 33620 7362 33718 4 gnd
port 2 nsew
rlabel metal3 s 7264 30460 7362 30558 4 gnd
port 2 nsew
rlabel metal3 s 7660 32830 7758 32928 4 vdd
port 1 nsew
rlabel metal3 s 6450 30878 6548 30976 4 vdd
port 1 nsew
rlabel metal3 s 7660 34015 7758 34113 4 vdd
port 1 nsew
rlabel metal3 s 7660 31645 7758 31743 4 vdd
port 1 nsew
rlabel metal3 s 7660 26905 7758 27003 4 vdd
port 1 nsew
rlabel metal3 s 6450 26928 6548 27026 4 vdd
port 1 nsew
rlabel metal3 s 7660 29275 7758 29373 4 vdd
port 1 nsew
rlabel metal3 s 6025 28134 6123 28232 4 gnd
port 2 nsew
rlabel metal3 s 7264 27300 7362 27398 4 gnd
port 2 nsew
rlabel metal3 s 7660 27695 7758 27793 4 vdd
port 1 nsew
rlabel metal3 s 7264 28880 7362 28978 4 gnd
port 2 nsew
rlabel metal3 s 7264 24535 7362 24633 4 gnd
port 2 nsew
rlabel metal3 s 6025 27344 6123 27442 4 gnd
port 2 nsew
rlabel metal3 s 6882 25348 6980 25446 4 vdd
port 1 nsew
rlabel metal3 s 7264 26510 7362 26608 4 gnd
port 2 nsew
rlabel metal3 s 6025 26928 6123 27026 4 gnd
port 2 nsew
rlabel metal3 s 6025 26138 6123 26236 4 gnd
port 2 nsew
rlabel metal3 s 7660 28090 7758 28188 4 vdd
port 1 nsew
rlabel metal3 s 6882 26928 6980 27026 4 vdd
port 1 nsew
rlabel metal3 s 6882 27286 6980 27384 4 vdd
port 1 nsew
rlabel metal3 s 6450 29298 6548 29396 4 vdd
port 1 nsew
rlabel metal3 s 6025 28508 6123 28606 4 gnd
port 2 nsew
rlabel metal3 s 7264 27695 7362 27793 4 gnd
port 2 nsew
rlabel metal3 s 6882 26496 6980 26594 4 vdd
port 1 nsew
rlabel metal3 s 6882 28076 6980 28174 4 vdd
port 1 nsew
rlabel metal3 s 6882 25706 6980 25804 4 vdd
port 1 nsew
rlabel metal3 s 6882 24916 6980 25014 4 vdd
port 1 nsew
rlabel metal3 s 6450 28866 6548 28964 4 vdd
port 1 nsew
rlabel metal3 s 6882 28508 6980 28606 4 vdd
port 1 nsew
rlabel metal3 s 7264 24930 7362 25028 4 gnd
port 2 nsew
rlabel metal3 s 7264 25720 7362 25818 4 gnd
port 2 nsew
rlabel metal3 s 6450 28508 6548 28606 4 vdd
port 1 nsew
rlabel metal3 s 6025 28924 6123 29022 4 gnd
port 2 nsew
rlabel metal3 s 7660 28880 7758 28978 4 vdd
port 1 nsew
rlabel metal3 s 7660 27300 7758 27398 4 vdd
port 1 nsew
rlabel metal3 s 6450 26138 6548 26236 4 vdd
port 1 nsew
rlabel metal3 s 6025 25764 6123 25862 4 gnd
port 2 nsew
rlabel metal3 s 6025 29298 6123 29396 4 gnd
port 2 nsew
rlabel metal3 s 7660 26510 7758 26608 4 vdd
port 1 nsew
rlabel metal3 s 7264 29275 7362 29373 4 gnd
port 2 nsew
rlabel metal3 s 6025 25348 6123 25446 4 gnd
port 2 nsew
rlabel metal3 s 7264 26905 7362 27003 4 gnd
port 2 nsew
rlabel metal3 s 6450 28076 6548 28174 4 vdd
port 1 nsew
rlabel metal3 s 6025 26554 6123 26652 4 gnd
port 2 nsew
rlabel metal3 s 7264 25325 7362 25423 4 gnd
port 2 nsew
rlabel metal3 s 6882 27718 6980 27816 4 vdd
port 1 nsew
rlabel metal3 s 7264 28090 7362 28188 4 gnd
port 2 nsew
rlabel metal3 s 6450 24558 6548 24656 4 vdd
port 1 nsew
rlabel metal3 s 6450 25348 6548 25446 4 vdd
port 1 nsew
rlabel metal3 s 6882 29298 6980 29396 4 vdd
port 1 nsew
rlabel metal3 s 6450 26496 6548 26594 4 vdd
port 1 nsew
rlabel metal3 s 7264 26115 7362 26213 4 gnd
port 2 nsew
rlabel metal3 s 6882 26138 6980 26236 4 vdd
port 1 nsew
rlabel metal3 s 6882 28866 6980 28964 4 vdd
port 1 nsew
rlabel metal3 s 6450 27718 6548 27816 4 vdd
port 1 nsew
rlabel metal3 s 7660 26115 7758 26213 4 vdd
port 1 nsew
rlabel metal3 s 7264 28485 7362 28583 4 gnd
port 2 nsew
rlabel metal3 s 7660 24930 7758 25028 4 vdd
port 1 nsew
rlabel metal3 s 6450 25706 6548 25804 4 vdd
port 1 nsew
rlabel metal3 s 6025 24974 6123 25072 4 gnd
port 2 nsew
rlabel metal3 s 7660 24535 7758 24633 4 vdd
port 1 nsew
rlabel metal3 s 6025 24558 6123 24656 4 gnd
port 2 nsew
rlabel metal3 s 6882 24558 6980 24656 4 vdd
port 1 nsew
rlabel metal3 s 7660 25325 7758 25423 4 vdd
port 1 nsew
rlabel metal3 s 6025 27718 6123 27816 4 gnd
port 2 nsew
rlabel metal3 s 7660 25720 7758 25818 4 vdd
port 1 nsew
rlabel metal3 s 6450 27286 6548 27384 4 vdd
port 1 nsew
rlabel metal3 s 6450 24916 6548 25014 4 vdd
port 1 nsew
rlabel metal3 s 7660 28485 7758 28583 4 vdd
port 1 nsew
rlabel metal3 s 3036 21398 3134 21496 4 vdd
port 1 nsew
rlabel metal3 s 2611 21398 2709 21496 4 gnd
port 2 nsew
rlabel metal3 s 3850 21375 3948 21473 4 gnd
port 2 nsew
rlabel metal3 s 2611 20608 2709 20706 4 gnd
port 2 nsew
rlabel metal3 s 4246 20585 4344 20683 4 vdd
port 1 nsew
rlabel metal3 s 3468 21398 3566 21496 4 vdd
port 1 nsew
rlabel metal3 s 3850 19795 3948 19893 4 gnd
port 2 nsew
rlabel metal3 s 3036 19818 3134 19916 4 vdd
port 1 nsew
rlabel metal3 s 4246 19795 4344 19893 4 vdd
port 1 nsew
rlabel metal3 s 4246 21375 4344 21473 4 vdd
port 1 nsew
rlabel metal3 s 3850 20585 3948 20683 4 gnd
port 2 nsew
rlabel metal3 s 3468 20608 3566 20706 4 vdd
port 1 nsew
rlabel metal3 s 3468 19818 3566 19916 4 vdd
port 1 nsew
rlabel metal3 s 2611 19818 2709 19916 4 gnd
port 2 nsew
rlabel metal3 s 3036 20608 3134 20706 4 vdd
port 1 nsew
rlabel metal3 s 6025 20234 6123 20332 4 gnd
port 2 nsew
rlabel metal3 s 6025 23394 6123 23492 4 gnd
port 2 nsew
rlabel metal3 s 6882 20608 6980 20706 4 vdd
port 1 nsew
rlabel metal3 s 7264 21770 7362 21868 4 gnd
port 2 nsew
rlabel metal3 s 7660 22560 7758 22658 4 vdd
port 1 nsew
rlabel metal3 s 6450 21398 6548 21496 4 vdd
port 1 nsew
rlabel metal3 s 7264 22560 7362 22658 4 gnd
port 2 nsew
rlabel metal3 s 6450 21756 6548 21854 4 vdd
port 1 nsew
rlabel metal3 s 6450 19818 6548 19916 4 vdd
port 1 nsew
rlabel metal3 s 6025 19818 6123 19916 4 gnd
port 2 nsew
rlabel metal3 s 6025 21814 6123 21912 4 gnd
port 2 nsew
rlabel metal3 s 6450 20966 6548 21064 4 vdd
port 1 nsew
rlabel metal3 s 6882 20966 6980 21064 4 vdd
port 1 nsew
rlabel metal3 s 6025 22978 6123 23076 4 gnd
port 2 nsew
rlabel metal3 s 7660 22165 7758 22263 4 vdd
port 1 nsew
rlabel metal3 s 7264 20980 7362 21078 4 gnd
port 2 nsew
rlabel metal3 s 7660 21375 7758 21473 4 vdd
port 1 nsew
rlabel metal3 s 6882 23768 6980 23866 4 vdd
port 1 nsew
rlabel metal3 s 6882 21756 6980 21854 4 vdd
port 1 nsew
rlabel metal3 s 7264 20585 7362 20683 4 gnd
port 2 nsew
rlabel metal3 s 6882 24126 6980 24224 4 vdd
port 1 nsew
rlabel metal3 s 6882 22188 6980 22286 4 vdd
port 1 nsew
rlabel metal3 s 6025 23768 6123 23866 4 gnd
port 2 nsew
rlabel metal3 s 6882 22546 6980 22644 4 vdd
port 1 nsew
rlabel metal3 s 7660 20585 7758 20683 4 vdd
port 1 nsew
rlabel metal3 s 6450 22546 6548 22644 4 vdd
port 1 nsew
rlabel metal3 s 6450 22188 6548 22286 4 vdd
port 1 nsew
rlabel metal3 s 7264 19795 7362 19893 4 gnd
port 2 nsew
rlabel metal3 s 7660 22955 7758 23053 4 vdd
port 1 nsew
rlabel metal3 s 6450 20176 6548 20274 4 vdd
port 1 nsew
rlabel metal3 s 6450 20608 6548 20706 4 vdd
port 1 nsew
rlabel metal3 s 7264 23745 7362 23843 4 gnd
port 2 nsew
rlabel metal3 s 7660 21770 7758 21868 4 vdd
port 1 nsew
rlabel metal3 s 7264 20190 7362 20288 4 gnd
port 2 nsew
rlabel metal3 s 6025 21398 6123 21496 4 gnd
port 2 nsew
rlabel metal3 s 6025 21024 6123 21122 4 gnd
port 2 nsew
rlabel metal3 s 7660 23350 7758 23448 4 vdd
port 1 nsew
rlabel metal3 s 7264 24140 7362 24238 4 gnd
port 2 nsew
rlabel metal3 s 6450 23768 6548 23866 4 vdd
port 1 nsew
rlabel metal3 s 6882 21398 6980 21496 4 vdd
port 1 nsew
rlabel metal3 s 7264 23350 7362 23448 4 gnd
port 2 nsew
rlabel metal3 s 6882 23336 6980 23434 4 vdd
port 1 nsew
rlabel metal3 s 7264 21375 7362 21473 4 gnd
port 2 nsew
rlabel metal3 s 7264 22955 7362 23053 4 gnd
port 2 nsew
rlabel metal3 s 6025 22188 6123 22286 4 gnd
port 2 nsew
rlabel metal3 s 6025 22604 6123 22702 4 gnd
port 2 nsew
rlabel metal3 s 6882 20176 6980 20274 4 vdd
port 1 nsew
rlabel metal3 s 7660 20190 7758 20288 4 vdd
port 1 nsew
rlabel metal3 s 6450 23336 6548 23434 4 vdd
port 1 nsew
rlabel metal3 s 6025 24184 6123 24282 4 gnd
port 2 nsew
rlabel metal3 s 6450 24126 6548 24224 4 vdd
port 1 nsew
rlabel metal3 s 7264 22165 7362 22263 4 gnd
port 2 nsew
rlabel metal3 s 6025 20608 6123 20706 4 gnd
port 2 nsew
rlabel metal3 s 7660 23745 7758 23843 4 vdd
port 1 nsew
rlabel metal3 s 6450 22978 6548 23076 4 vdd
port 1 nsew
rlabel metal3 s 7660 20980 7758 21078 4 vdd
port 1 nsew
rlabel metal3 s 7660 24140 7758 24238 4 vdd
port 1 nsew
rlabel metal3 s 7660 19795 7758 19893 4 vdd
port 1 nsew
rlabel metal3 s 6882 19818 6980 19916 4 vdd
port 1 nsew
rlabel metal3 s 6882 22978 6980 23076 4 vdd
port 1 nsew
rlabel metal3 s 12600 20190 12698 20288 4 gnd
port 2 nsew
rlabel metal3 s 12600 27063 12698 27161 4 gnd
port 2 nsew
rlabel metal3 s 12600 25957 12698 26055 4 gnd
port 2 nsew
rlabel metal3 s 12600 20743 12698 20841 4 gnd
port 2 nsew
rlabel metal3 s 12600 22007 12698 22105 4 gnd
port 2 nsew
rlabel metal3 s 12600 26273 12698 26371 4 gnd
port 2 nsew
rlabel metal3 s 12600 22797 12698 22895 4 gnd
port 2 nsew
rlabel metal3 s 12600 29117 12698 29215 4 gnd
port 2 nsew
rlabel metal3 s 12600 27853 12698 27951 4 gnd
port 2 nsew
rlabel metal3 s 12600 28643 12698 28741 4 gnd
port 2 nsew
rlabel metal3 s 12600 24140 12698 24238 4 gnd
port 2 nsew
rlabel metal3 s 12600 25720 12698 25818 4 gnd
port 2 nsew
rlabel metal3 s 12600 25167 12698 25265 4 gnd
port 2 nsew
rlabel metal3 s 12600 22560 12698 22658 4 gnd
port 2 nsew
rlabel metal3 s 12600 23113 12698 23211 4 gnd
port 2 nsew
rlabel metal3 s 12600 28327 12698 28425 4 gnd
port 2 nsew
rlabel metal3 s 12600 21217 12698 21315 4 gnd
port 2 nsew
rlabel metal3 s 12600 24377 12698 24475 4 gnd
port 2 nsew
rlabel metal3 s 12600 26747 12698 26845 4 gnd
port 2 nsew
rlabel metal3 s 12600 19637 12698 19735 4 gnd
port 2 nsew
rlabel metal3 s 12600 21533 12698 21631 4 gnd
port 2 nsew
rlabel metal3 s 12600 23350 12698 23448 4 gnd
port 2 nsew
rlabel metal3 s 12600 21770 12698 21868 4 gnd
port 2 nsew
rlabel metal3 s 12600 27300 12698 27398 4 gnd
port 2 nsew
rlabel metal3 s 12600 20980 12698 21078 4 gnd
port 2 nsew
rlabel metal3 s 12600 23903 12698 24001 4 gnd
port 2 nsew
rlabel metal3 s 12600 28090 12698 28188 4 gnd
port 2 nsew
rlabel metal3 s 12600 27537 12698 27635 4 gnd
port 2 nsew
rlabel metal3 s 12600 24693 12698 24791 4 gnd
port 2 nsew
rlabel metal3 s 12600 23587 12698 23685 4 gnd
port 2 nsew
rlabel metal3 s 12600 19953 12698 20051 4 gnd
port 2 nsew
rlabel metal3 s 12600 22323 12698 22421 4 gnd
port 2 nsew
rlabel metal3 s 12600 26510 12698 26608 4 gnd
port 2 nsew
rlabel metal3 s 12600 20427 12698 20525 4 gnd
port 2 nsew
rlabel metal3 s 12600 25483 12698 25581 4 gnd
port 2 nsew
rlabel metal3 s 12600 28880 12698 28978 4 gnd
port 2 nsew
rlabel metal3 s 12600 24930 12698 25028 4 gnd
port 2 nsew
rlabel metal3 s 17040 13309 17138 13407 4 vdd
port 1 nsew
rlabel metal3 s 13296 13309 13394 13407 4 vdd
port 1 nsew
rlabel metal3 s 12600 15213 12698 15311 4 gnd
port 2 nsew
rlabel metal3 s 11208 13673 11306 13771 4 vdd
port 1 nsew
rlabel metal3 s 12600 18373 12698 18471 4 gnd
port 2 nsew
rlabel metal3 s 14663 12718 14761 12816 4 vdd
port 1 nsew
rlabel metal3 s 12600 16477 12698 16575 4 gnd
port 2 nsew
rlabel metal3 s 12600 14660 12698 14758 4 gnd
port 2 nsew
rlabel metal3 s 15168 13309 15266 13407 4 vdd
port 1 nsew
rlabel metal3 s 12600 18610 12698 18708 4 gnd
port 2 nsew
rlabel metal3 s 15911 12718 16009 12816 4 vdd
port 1 nsew
rlabel metal3 s 12600 17583 12698 17681 4 gnd
port 2 nsew
rlabel metal3 s 12600 14107 12698 14205 4 gnd
port 2 nsew
rlabel metal3 s 12600 19163 12698 19261 4 gnd
port 2 nsew
rlabel metal3 s 12600 18057 12698 18155 4 gnd
port 2 nsew
rlabel metal3 s 15480 11169 15578 11267 4 gnd
port 2 nsew
rlabel metal3 s 16728 11169 16826 11267 4 gnd
port 2 nsew
rlabel metal3 s 12234 13743 12332 13841 4 gnd
port 2 nsew
rlabel metal3 s 12600 15687 12698 15785 4 gnd
port 2 nsew
rlabel metal3 s 12600 17267 12698 17365 4 gnd
port 2 nsew
rlabel metal3 s 16297 12718 16395 12816 4 vdd
port 1 nsew
rlabel metal3 s 13415 12718 13513 12816 4 vdd
port 1 nsew
rlabel metal3 s 13801 12718 13899 12816 4 vdd
port 1 nsew
rlabel metal3 s 12600 14423 12698 14521 4 gnd
port 2 nsew
rlabel metal3 s 14544 13309 14642 13407 4 vdd
port 1 nsew
rlabel metal3 s 15049 12718 15147 12816 4 vdd
port 1 nsew
rlabel metal3 s 15792 13309 15890 13407 4 vdd
port 1 nsew
rlabel metal3 s 17159 12718 17257 12816 4 vdd
port 1 nsew
rlabel metal3 s 12600 13870 12698 13968 4 gnd
port 2 nsew
rlabel metal3 s 12600 16793 12698 16891 4 gnd
port 2 nsew
rlabel metal3 s 12600 14897 12698 14995 4 gnd
port 2 nsew
rlabel metal3 s 12600 18847 12698 18945 4 gnd
port 2 nsew
rlabel metal3 s 14232 11169 14330 11267 4 gnd
port 2 nsew
rlabel metal3 s 12600 17030 12698 17128 4 gnd
port 2 nsew
rlabel metal3 s 12600 16003 12698 16101 4 gnd
port 2 nsew
rlabel metal3 s 12600 15450 12698 15548 4 gnd
port 2 nsew
rlabel metal3 s 12600 16240 12698 16338 4 gnd
port 2 nsew
rlabel metal3 s 13920 13309 14018 13407 4 vdd
port 1 nsew
rlabel metal3 s 12600 19400 12698 19498 4 gnd
port 2 nsew
rlabel metal3 s 16416 13309 16514 13407 4 vdd
port 1 nsew
rlabel metal3 s 12600 17820 12698 17918 4 gnd
port 2 nsew
rlabel metal3 s 6882 16226 6980 16324 4 vdd
port 1 nsew
rlabel metal3 s 7264 18610 7362 18708 4 gnd
port 2 nsew
rlabel metal3 s 6025 14704 6123 14802 4 gnd
port 2 nsew
rlabel metal3 s 7660 18610 7758 18708 4 vdd
port 1 nsew
rlabel metal3 s 6882 18596 6980 18694 4 vdd
port 1 nsew
rlabel metal3 s 6450 17806 6548 17904 4 vdd
port 1 nsew
rlabel metal3 s 6025 18654 6123 18752 4 gnd
port 2 nsew
rlabel metal3 s 7660 17030 7758 17128 4 vdd
port 1 nsew
rlabel metal3 s 7264 19400 7362 19498 4 gnd
port 2 nsew
rlabel metal3 s 7660 16240 7758 16338 4 vdd
port 1 nsew
rlabel metal3 s 7264 16635 7362 16733 4 gnd
port 2 nsew
rlabel metal3 s 7264 16240 7362 16338 4 gnd
port 2 nsew
rlabel metal3 s 6025 17864 6123 17962 4 gnd
port 2 nsew
rlabel metal3 s 6025 17448 6123 17546 4 gnd
port 2 nsew
rlabel metal3 s 6025 16284 6123 16382 4 gnd
port 2 nsew
rlabel metal3 s 6882 15868 6980 15966 4 vdd
port 1 nsew
rlabel metal3 s 6882 15436 6980 15534 4 vdd
port 1 nsew
rlabel metal3 s 6882 16658 6980 16756 4 vdd
port 1 nsew
rlabel metal3 s 6025 15494 6123 15592 4 gnd
port 2 nsew
rlabel metal3 s 6450 15436 6548 15534 4 vdd
port 1 nsew
rlabel metal3 s 7264 18215 7362 18313 4 gnd
port 2 nsew
rlabel metal3 s 7264 19005 7362 19103 4 gnd
port 2 nsew
rlabel metal3 s 7660 15450 7758 15548 4 vdd
port 1 nsew
rlabel metal3 s 6025 16658 6123 16756 4 gnd
port 2 nsew
rlabel metal3 s 6882 17448 6980 17546 4 vdd
port 1 nsew
rlabel metal3 s 6882 19028 6980 19126 4 vdd
port 1 nsew
rlabel metal3 s 6882 17806 6980 17904 4 vdd
port 1 nsew
rlabel metal3 s 7264 15055 7362 15153 4 gnd
port 2 nsew
rlabel metal3 s 6025 19444 6123 19542 4 gnd
port 2 nsew
rlabel metal3 s 6882 19386 6980 19484 4 vdd
port 1 nsew
rlabel metal3 s 7660 19400 7758 19498 4 vdd
port 1 nsew
rlabel metal3 s 6450 17448 6548 17546 4 vdd
port 1 nsew
rlabel metal3 s 6025 15868 6123 15966 4 gnd
port 2 nsew
rlabel metal3 s 6450 19028 6548 19126 4 vdd
port 1 nsew
rlabel metal3 s 6450 15868 6548 15966 4 vdd
port 1 nsew
rlabel metal3 s 7264 17425 7362 17523 4 gnd
port 2 nsew
rlabel metal3 s 6450 18596 6548 18694 4 vdd
port 1 nsew
rlabel metal3 s 6450 19386 6548 19484 4 vdd
port 1 nsew
rlabel metal3 s 6025 17074 6123 17172 4 gnd
port 2 nsew
rlabel metal3 s 7660 16635 7758 16733 4 vdd
port 1 nsew
rlabel metal3 s 7660 17425 7758 17523 4 vdd
port 1 nsew
rlabel metal3 s 6450 18238 6548 18336 4 vdd
port 1 nsew
rlabel metal3 s 6025 19028 6123 19126 4 gnd
port 2 nsew
rlabel metal3 s 6882 17016 6980 17114 4 vdd
port 1 nsew
rlabel metal3 s 7264 17820 7362 17918 4 gnd
port 2 nsew
rlabel metal3 s 7660 18215 7758 18313 4 vdd
port 1 nsew
rlabel metal3 s 6025 18238 6123 18336 4 gnd
port 2 nsew
rlabel metal3 s 6450 17016 6548 17114 4 vdd
port 1 nsew
rlabel metal3 s 7660 15055 7758 15153 4 vdd
port 1 nsew
rlabel metal3 s 7264 17030 7362 17128 4 gnd
port 2 nsew
rlabel metal3 s 6025 15078 6123 15176 4 gnd
port 2 nsew
rlabel metal3 s 7264 15845 7362 15943 4 gnd
port 2 nsew
rlabel metal3 s 7660 19005 7758 19103 4 vdd
port 1 nsew
rlabel metal3 s 7264 15450 7362 15548 4 gnd
port 2 nsew
rlabel metal3 s 6882 15078 6980 15176 4 vdd
port 1 nsew
rlabel metal3 s 7660 17820 7758 17918 4 vdd
port 1 nsew
rlabel metal3 s 6450 16658 6548 16756 4 vdd
port 1 nsew
rlabel metal3 s 7660 15845 7758 15943 4 vdd
port 1 nsew
rlabel metal3 s 6450 16226 6548 16324 4 vdd
port 1 nsew
rlabel metal3 s 6450 15078 6548 15176 4 vdd
port 1 nsew
rlabel metal3 s 6882 18238 6980 18336 4 vdd
port 1 nsew
rlabel metal3 s 3471 16642 3569 16740 4 vdd
port 1 nsew
rlabel metal3 s 4246 17425 4344 17523 4 vdd
port 1 nsew
rlabel metal3 s 3850 16635 3948 16733 4 gnd
port 2 nsew
rlabel metal3 s 3046 16642 3144 16740 4 gnd
port 2 nsew
rlabel metal3 s 1752 16635 1850 16733 4 gnd
port 2 nsew
rlabel metal3 s 4246 15055 4344 15153 4 vdd
port 1 nsew
rlabel metal3 s 3471 15062 3569 15160 4 vdd
port 1 nsew
rlabel metal3 s 3468 19028 3566 19126 4 vdd
port 1 nsew
rlabel metal3 s 2611 19028 2709 19126 4 gnd
port 2 nsew
rlabel metal3 s 4246 19005 4344 19103 4 vdd
port 1 nsew
rlabel metal3 s 2148 16635 2246 16733 4 vdd
port 1 nsew
rlabel metal3 s 1156 19005 1254 19103 4 gnd
port 2 nsew
rlabel metal3 s 1552 19005 1650 19103 4 vdd
port 1 nsew
rlabel metal3 s 3036 19028 3134 19126 4 vdd
port 1 nsew
rlabel metal3 s 3850 19005 3948 19103 4 gnd
port 2 nsew
rlabel metal3 s 3046 17432 3144 17530 4 gnd
port 2 nsew
rlabel metal3 s 3471 17432 3569 17530 4 vdd
port 1 nsew
rlabel metal3 s 3046 15062 3144 15160 4 gnd
port 2 nsew
rlabel metal3 s 3850 17425 3948 17523 4 gnd
port 2 nsew
rlabel metal3 s 3850 15055 3948 15153 4 gnd
port 2 nsew
rlabel metal3 s 4246 16635 4344 16733 4 vdd
port 1 nsew
rlabel metal3 s 4676 9898 4774 9996 4 vdd
port 1 nsew
rlabel metal3 s 4246 14265 4344 14363 4 vdd
port 1 nsew
rlabel metal3 s 2148 14265 2246 14363 4 vdd
port 1 nsew
rlabel metal3 s 1752 14265 1850 14363 4 gnd
port 2 nsew
rlabel metal3 s 3046 14272 3144 14370 4 gnd
port 2 nsew
rlabel metal3 s 3850 14265 3948 14363 4 gnd
port 2 nsew
rlabel metal3 s 3471 14272 3569 14370 4 vdd
port 1 nsew
rlabel metal3 s 4676 11312 4774 11410 4 gnd
port 2 nsew
rlabel metal3 s 6450 14288 6548 14386 4 vdd
port 1 nsew
rlabel metal3 s 7685 13679 7783 13777 4 vdd
port 1 nsew
rlabel metal3 s 6036 11312 6134 11410 4 gnd
port 2 nsew
rlabel metal3 s 6450 14646 6548 14744 4 vdd
port 1 nsew
rlabel metal3 s 6025 14288 6123 14386 4 gnd
port 2 nsew
rlabel metal3 s 6882 14646 6980 14744 4 vdd
port 1 nsew
rlabel metal3 s 6882 14288 6980 14386 4 vdd
port 1 nsew
rlabel metal3 s 7660 14660 7758 14758 4 vdd
port 1 nsew
rlabel metal3 s 0 11969 13577 12029 4 rbl_bl_0_0
port 4 nsew
rlabel metal3 s 7264 14265 7362 14363 4 gnd
port 2 nsew
rlabel metal3 s 6036 9898 6134 9996 4 vdd
port 1 nsew
rlabel metal3 s 7264 14660 7362 14758 4 gnd
port 2 nsew
rlabel metal3 s 7660 14265 7758 14363 4 vdd
port 1 nsew
rlabel metal3 s 8517 13685 8615 13783 4 vdd
port 1 nsew
rlabel metal3 s 6036 0 6134 98 4 gnd
port 2 nsew
rlabel metal3 s 4676 2828 4774 2926 4 gnd
port 2 nsew
rlabel metal3 s 6036 4242 6134 4340 4 vdd
port 1 nsew
rlabel metal3 s 6036 5656 6134 5754 4 gnd
port 2 nsew
rlabel metal3 s 6036 7070 6134 7168 4 vdd
port 1 nsew
rlabel metal3 s 4676 0 4774 98 4 gnd
port 2 nsew
rlabel metal3 s 4676 8484 4774 8582 4 gnd
port 2 nsew
rlabel metal3 s 6036 1414 6134 1512 4 vdd
port 1 nsew
rlabel metal3 s 6036 2828 6134 2926 4 gnd
port 2 nsew
rlabel metal3 s 4676 1414 4774 1512 4 vdd
port 1 nsew
rlabel metal3 s 4676 4242 4774 4340 4 vdd
port 1 nsew
rlabel metal3 s 4676 7070 4774 7168 4 vdd
port 1 nsew
rlabel metal3 s 6036 8484 6134 8582 4 gnd
port 2 nsew
rlabel metal3 s 4676 5656 4774 5754 4 gnd
port 2 nsew
rlabel metal3 s 12234 2999 12332 3097 4 gnd
port 2 nsew
rlabel metal3 s 13977 7902 14075 8000 4 vdd
port 1 nsew
rlabel metal3 s 13870 4978 13968 5076 4 gnd
port 2 nsew
rlabel metal3 s 13864 5512 13962 5610 4 vdd
port 1 nsew
rlabel metal3 s 12234 4119 12332 4217 4 vdd
port 1 nsew
rlabel metal3 s 13989 7064 14087 7162 4 vdd
port 1 nsew
rlabel metal3 s 13985 5180 14083 5278 4 gnd
port 2 nsew
rlabel metal3 s 14059 8676 14157 8774 4 gnd
port 2 nsew
rlabel metal3 s 13884 4562 13982 4660 4 vdd
port 1 nsew
rlabel metal3 s 13875 5949 13973 6047 4 gnd
port 2 nsew
rlabel metal3 s 13989 6742 14087 6840 4 gnd
port 2 nsew
rlabel metal3 s 23961 7902 24059 8000 4 vdd
port 1 nsew
rlabel metal3 s 26281 12718 26379 12816 4 vdd
port 1 nsew
rlabel metal3 s 28846 4978 28944 5076 4 gnd
port 2 nsew
rlabel metal3 s 19051 8676 19149 8774 4 gnd
port 2 nsew
rlabel metal3 s 28777 12718 28875 12816 4 vdd
port 1 nsew
rlabel metal3 s 23859 5949 23957 6047 4 gnd
port 2 nsew
rlabel metal3 s 25895 12718 25993 12816 4 vdd
port 1 nsew
rlabel metal3 s 20784 13309 20882 13407 4 vdd
port 1 nsew
rlabel metal3 s 18793 12718 18891 12816 4 vdd
port 1 nsew
rlabel metal3 s 32952 11169 33050 11267 4 gnd
port 2 nsew
rlabel metal3 s 18969 7902 19067 8000 4 vdd
port 1 nsew
rlabel metal3 s 28391 12718 28489 12816 4 vdd
port 1 nsew
rlabel metal3 s 18407 12718 18505 12816 4 vdd
port 1 nsew
rlabel metal3 s 28965 7064 29063 7162 4 vdd
port 1 nsew
rlabel metal3 s 28953 7902 29051 8000 4 vdd
port 1 nsew
rlabel metal3 s 28272 13309 28370 13407 4 vdd
port 1 nsew
rlabel metal3 s 32135 12718 32233 12816 4 vdd
port 1 nsew
rlabel metal3 s 18876 4562 18974 4660 4 vdd
port 1 nsew
rlabel metal3 s 29520 13309 29618 13407 4 vdd
port 1 nsew
rlabel metal3 s 18288 13309 18386 13407 4 vdd
port 1 nsew
rlabel metal3 s 30144 13309 30242 13407 4 vdd
port 1 nsew
rlabel metal3 s 23868 4562 23966 4660 4 vdd
port 1 nsew
rlabel metal3 s 32521 12718 32619 12816 4 vdd
port 1 nsew
rlabel metal3 s 22537 12718 22635 12816 4 vdd
port 1 nsew
rlabel metal3 s 21720 11169 21818 11267 4 gnd
port 2 nsew
rlabel metal3 s 23399 12718 23497 12816 4 vdd
port 1 nsew
rlabel metal3 s 30768 13309 30866 13407 4 vdd
port 1 nsew
rlabel metal3 s 18867 5949 18965 6047 4 gnd
port 2 nsew
rlabel metal3 s 23785 12718 23883 12816 4 vdd
port 1 nsew
rlabel metal3 s 25776 13309 25874 13407 4 vdd
port 1 nsew
rlabel metal3 s 27648 13309 27746 13407 4 vdd
port 1 nsew
rlabel metal3 s 19536 13309 19634 13407 4 vdd
port 1 nsew
rlabel metal3 s 29208 11169 29306 11267 4 gnd
port 2 nsew
rlabel metal3 s 28961 5180 29059 5278 4 gnd
port 2 nsew
rlabel metal3 s 25464 11169 25562 11267 4 gnd
port 2 nsew
rlabel metal3 s 18977 5180 19075 5278 4 gnd
port 2 nsew
rlabel metal3 s 19655 12718 19753 12816 4 vdd
port 1 nsew
rlabel metal3 s 24216 11169 24314 11267 4 gnd
port 2 nsew
rlabel metal3 s 18981 6742 19079 6840 4 gnd
port 2 nsew
rlabel metal3 s 31704 11169 31802 11267 4 gnd
port 2 nsew
rlabel metal3 s 23973 7064 24071 7162 4 vdd
port 1 nsew
rlabel metal3 s 25152 13309 25250 13407 4 vdd
port 1 nsew
rlabel metal3 s 23848 5512 23946 5610 4 vdd
port 1 nsew
rlabel metal3 s 30025 12718 30123 12816 4 vdd
port 1 nsew
rlabel metal3 s 27024 13309 27122 13407 4 vdd
port 1 nsew
rlabel metal3 s 23280 13309 23378 13407 4 vdd
port 1 nsew
rlabel metal3 s 24528 13309 24626 13407 4 vdd
port 1 nsew
rlabel metal3 s 25033 12718 25131 12816 4 vdd
port 1 nsew
rlabel metal3 s 20472 11169 20570 11267 4 gnd
port 2 nsew
rlabel metal3 s 31273 12718 31371 12816 4 vdd
port 1 nsew
rlabel metal3 s 32640 13309 32738 13407 4 vdd
port 1 nsew
rlabel metal3 s 23904 13309 24002 13407 4 vdd
port 1 nsew
rlabel metal3 s 33383 12718 33481 12816 4 vdd
port 1 nsew
rlabel metal3 s 21408 13309 21506 13407 4 vdd
port 1 nsew
rlabel metal3 s 28965 6742 29063 6840 4 gnd
port 2 nsew
rlabel metal3 s 28840 5512 28938 5610 4 vdd
port 1 nsew
rlabel metal3 s 27143 12718 27241 12816 4 vdd
port 1 nsew
rlabel metal3 s 31392 13309 31490 13407 4 vdd
port 1 nsew
rlabel metal3 s 30887 12718 30985 12816 4 vdd
port 1 nsew
rlabel metal3 s 30456 11169 30554 11267 4 gnd
port 2 nsew
rlabel metal3 s 18856 5512 18954 5610 4 vdd
port 1 nsew
rlabel metal3 s 17545 12718 17643 12816 4 vdd
port 1 nsew
rlabel metal3 s 24647 12718 24745 12816 4 vdd
port 1 nsew
rlabel metal3 s 28896 13309 28994 13407 4 vdd
port 1 nsew
rlabel metal3 s 27960 11169 28058 11267 4 gnd
port 2 nsew
rlabel metal3 s 27529 12718 27627 12816 4 vdd
port 1 nsew
rlabel metal3 s 22656 13309 22754 13407 4 vdd
port 1 nsew
rlabel metal3 s 24043 8676 24141 8774 4 gnd
port 2 nsew
rlabel metal3 s 33264 13309 33362 13407 4 vdd
port 1 nsew
rlabel metal3 s 20041 12718 20139 12816 4 vdd
port 1 nsew
rlabel metal3 s 26400 13309 26498 13407 4 vdd
port 1 nsew
rlabel metal3 s 26712 11169 26810 11267 4 gnd
port 2 nsew
rlabel metal3 s 17976 11169 18074 11267 4 gnd
port 2 nsew
rlabel metal3 s 20903 12718 21001 12816 4 vdd
port 1 nsew
rlabel metal3 s 19224 11169 19322 11267 4 gnd
port 2 nsew
rlabel metal3 s 29639 12718 29737 12816 4 vdd
port 1 nsew
rlabel metal3 s 18862 4978 18960 5076 4 gnd
port 2 nsew
rlabel metal3 s 21289 12718 21387 12816 4 vdd
port 1 nsew
rlabel metal3 s 18981 7064 19079 7162 4 vdd
port 1 nsew
rlabel metal3 s 28851 5949 28949 6047 4 gnd
port 2 nsew
rlabel metal3 s 18912 13309 19010 13407 4 vdd
port 1 nsew
rlabel metal3 s 23973 6742 24071 6840 4 gnd
port 2 nsew
rlabel metal3 s 17664 13309 17762 13407 4 vdd
port 1 nsew
rlabel metal3 s 22151 12718 22249 12816 4 vdd
port 1 nsew
rlabel metal3 s 20160 13309 20258 13407 4 vdd
port 1 nsew
rlabel metal3 s 29035 8676 29133 8774 4 gnd
port 2 nsew
rlabel metal3 s 23969 5180 24067 5278 4 gnd
port 2 nsew
rlabel metal3 s 28860 4562 28958 4660 4 vdd
port 1 nsew
rlabel metal3 s 23854 4978 23952 5076 4 gnd
port 2 nsew
rlabel metal3 s 22032 13309 22130 13407 4 vdd
port 1 nsew
rlabel metal3 s 32016 13309 32114 13407 4 vdd
port 1 nsew
rlabel metal3 s 22968 11169 23066 11267 4 gnd
port 2 nsew
rlabel metal3 s 59888 37175 59986 37273 4 gnd
port 2 nsew
rlabel metal3 s 59492 34410 59590 34508 4 vdd
port 1 nsew
rlabel metal3 s 59888 37965 59986 38063 4 gnd
port 2 nsew
rlabel metal3 s 60270 39136 60368 39234 4 vdd
port 1 nsew
rlabel metal3 s 60702 36408 60800 36506 4 vdd
port 1 nsew
rlabel metal3 s 59492 37965 59590 38063 4 vdd
port 1 nsew
rlabel metal3 s 61127 37988 61225 38086 4 gnd
port 2 nsew
rlabel metal3 s 60702 35186 60800 35284 4 vdd
port 1 nsew
rlabel metal3 s 59888 39150 59986 39248 4 gnd
port 2 nsew
rlabel metal3 s 60270 34828 60368 34926 4 vdd
port 1 nsew
rlabel metal3 s 60702 37988 60800 38086 4 vdd
port 1 nsew
rlabel metal3 s 59888 36780 59986 36878 4 gnd
port 2 nsew
rlabel metal3 s 60270 35186 60368 35284 4 vdd
port 1 nsew
rlabel metal3 s 61127 36034 61225 36132 4 gnd
port 2 nsew
rlabel metal3 s 59492 35200 59590 35298 4 vdd
port 1 nsew
rlabel metal3 s 60702 37198 60800 37296 4 vdd
port 1 nsew
rlabel metal3 s 59888 35595 59986 35693 4 gnd
port 2 nsew
rlabel metal3 s 59888 35200 59986 35298 4 gnd
port 2 nsew
rlabel metal3 s 60270 36408 60368 36506 4 vdd
port 1 nsew
rlabel metal3 s 60270 36766 60368 36864 4 vdd
port 1 nsew
rlabel metal3 s 61127 37614 61225 37712 4 gnd
port 2 nsew
rlabel metal3 s 59492 34805 59590 34903 4 vdd
port 1 nsew
rlabel metal3 s 59492 39150 59590 39248 4 vdd
port 1 nsew
rlabel metal3 s 61127 38778 61225 38876 4 gnd
port 2 nsew
rlabel metal3 s 60702 38346 60800 38444 4 vdd
port 1 nsew
rlabel metal3 s 60702 39136 60800 39234 4 vdd
port 1 nsew
rlabel metal3 s 58635 39134 58733 39232 4 vdd
port 1 nsew
rlabel metal3 s 59888 35990 59986 36088 4 gnd
port 2 nsew
rlabel metal3 s 59888 37570 59986 37668 4 gnd
port 2 nsew
rlabel metal3 s 59492 35595 59590 35693 4 vdd
port 1 nsew
rlabel metal3 s 60702 35976 60800 36074 4 vdd
port 1 nsew
rlabel metal3 s 60702 34828 60800 34926 4 vdd
port 1 nsew
rlabel metal3 s 61127 35244 61225 35342 4 gnd
port 2 nsew
rlabel metal3 s 60270 34396 60368 34494 4 vdd
port 1 nsew
rlabel metal3 s 59492 36385 59590 36483 4 vdd
port 1 nsew
rlabel metal3 s 60270 37988 60368 38086 4 vdd
port 1 nsew
rlabel metal3 s 59888 38360 59986 38458 4 gnd
port 2 nsew
rlabel metal3 s 60270 35618 60368 35716 4 vdd
port 1 nsew
rlabel metal3 s 61127 36408 61225 36506 4 gnd
port 2 nsew
rlabel metal3 s 59492 38360 59590 38458 4 vdd
port 1 nsew
rlabel metal3 s 59492 36780 59590 36878 4 vdd
port 1 nsew
rlabel metal3 s 59888 36385 59986 36483 4 gnd
port 2 nsew
rlabel metal3 s 59888 38755 59986 38853 4 gnd
port 2 nsew
rlabel metal3 s 60270 38346 60368 38444 4 vdd
port 1 nsew
rlabel metal3 s 61127 35618 61225 35716 4 gnd
port 2 nsew
rlabel metal3 s 61127 34454 61225 34552 4 gnd
port 2 nsew
rlabel metal3 s 61127 36824 61225 36922 4 gnd
port 2 nsew
rlabel metal3 s 60270 38778 60368 38876 4 vdd
port 1 nsew
rlabel metal3 s 60702 37556 60800 37654 4 vdd
port 1 nsew
rlabel metal3 s 59060 39135 59158 39233 4 gnd
port 2 nsew
rlabel metal3 s 60270 37198 60368 37296 4 vdd
port 1 nsew
rlabel metal3 s 59492 38755 59590 38853 4 vdd
port 1 nsew
rlabel metal3 s 60702 35618 60800 35716 4 vdd
port 1 nsew
rlabel metal3 s 60702 34396 60800 34494 4 vdd
port 1 nsew
rlabel metal3 s 59888 34805 59986 34903 4 gnd
port 2 nsew
rlabel metal3 s 60270 35976 60368 36074 4 vdd
port 1 nsew
rlabel metal3 s 59492 37175 59590 37273 4 vdd
port 1 nsew
rlabel metal3 s 59492 37570 59590 37668 4 vdd
port 1 nsew
rlabel metal3 s 59888 34410 59986 34508 4 gnd
port 2 nsew
rlabel metal3 s 61127 38404 61225 38502 4 gnd
port 2 nsew
rlabel metal3 s 59492 35990 59590 36088 4 vdd
port 1 nsew
rlabel metal3 s 60270 37556 60368 37654 4 vdd
port 1 nsew
rlabel metal3 s 60702 38778 60800 38876 4 vdd
port 1 nsew
rlabel metal3 s 61127 34828 61225 34926 4 gnd
port 2 nsew
rlabel metal3 s 61127 37198 61225 37296 4 gnd
port 2 nsew
rlabel metal3 s 60702 36766 60800 36864 4 vdd
port 1 nsew
rlabel metal3 s 61127 30878 61225 30976 4 gnd
port 2 nsew
rlabel metal3 s 59492 30065 59590 30163 4 vdd
port 1 nsew
rlabel metal3 s 60270 33606 60368 33704 4 vdd
port 1 nsew
rlabel metal3 s 60702 32816 60800 32914 4 vdd
port 1 nsew
rlabel metal3 s 60270 32816 60368 32914 4 vdd
port 1 nsew
rlabel metal3 s 60270 30446 60368 30544 4 vdd
port 1 nsew
rlabel metal3 s 60702 32458 60800 32556 4 vdd
port 1 nsew
rlabel metal3 s 60270 32458 60368 32556 4 vdd
port 1 nsew
rlabel metal3 s 59888 32830 59986 32928 4 gnd
port 2 nsew
rlabel metal3 s 60270 30088 60368 30186 4 vdd
port 1 nsew
rlabel metal3 s 61127 30088 61225 30186 4 gnd
port 2 nsew
rlabel metal3 s 60702 34038 60800 34136 4 vdd
port 1 nsew
rlabel metal3 s 60270 31236 60368 31334 4 vdd
port 1 nsew
rlabel metal3 s 59888 33620 59986 33718 4 gnd
port 2 nsew
rlabel metal3 s 60702 33248 60800 33346 4 vdd
port 1 nsew
rlabel metal3 s 60270 31668 60368 31766 4 vdd
port 1 nsew
rlabel metal3 s 61127 34038 61225 34136 4 gnd
port 2 nsew
rlabel metal3 s 59888 29670 59986 29768 4 gnd
port 2 nsew
rlabel metal3 s 60702 30878 60800 30976 4 vdd
port 1 nsew
rlabel metal3 s 61127 32084 61225 32182 4 gnd
port 2 nsew
rlabel metal3 s 60702 31668 60800 31766 4 vdd
port 1 nsew
rlabel metal3 s 59888 33225 59986 33323 4 gnd
port 2 nsew
rlabel metal3 s 59492 32830 59590 32928 4 vdd
port 1 nsew
rlabel metal3 s 59888 32040 59986 32138 4 gnd
port 2 nsew
rlabel metal3 s 59492 32040 59590 32138 4 vdd
port 1 nsew
rlabel metal3 s 60702 30446 60800 30544 4 vdd
port 1 nsew
rlabel metal3 s 60702 33606 60800 33704 4 vdd
port 1 nsew
rlabel metal3 s 59492 33620 59590 33718 4 vdd
port 1 nsew
rlabel metal3 s 59888 30855 59986 30953 4 gnd
port 2 nsew
rlabel metal3 s 59888 30065 59986 30163 4 gnd
port 2 nsew
rlabel metal3 s 59492 29670 59590 29768 4 vdd
port 1 nsew
rlabel metal3 s 60270 34038 60368 34136 4 vdd
port 1 nsew
rlabel metal3 s 59492 31645 59590 31743 4 vdd
port 1 nsew
rlabel metal3 s 60702 30088 60800 30186 4 vdd
port 1 nsew
rlabel metal3 s 60270 29656 60368 29754 4 vdd
port 1 nsew
rlabel metal3 s 59888 31645 59986 31743 4 gnd
port 2 nsew
rlabel metal3 s 59888 31250 59986 31348 4 gnd
port 2 nsew
rlabel metal3 s 59492 31250 59590 31348 4 vdd
port 1 nsew
rlabel metal3 s 60270 30878 60368 30976 4 vdd
port 1 nsew
rlabel metal3 s 60702 29656 60800 29754 4 vdd
port 1 nsew
rlabel metal3 s 61127 31294 61225 31392 4 gnd
port 2 nsew
rlabel metal3 s 59492 30460 59590 30558 4 vdd
port 1 nsew
rlabel metal3 s 61127 33664 61225 33762 4 gnd
port 2 nsew
rlabel metal3 s 59888 30460 59986 30558 4 gnd
port 2 nsew
rlabel metal3 s 60270 32026 60368 32124 4 vdd
port 1 nsew
rlabel metal3 s 59492 32435 59590 32533 4 vdd
port 1 nsew
rlabel metal3 s 61127 32874 61225 32972 4 gnd
port 2 nsew
rlabel metal3 s 61127 30504 61225 30602 4 gnd
port 2 nsew
rlabel metal3 s 59492 33225 59590 33323 4 vdd
port 1 nsew
rlabel metal3 s 61127 33248 61225 33346 4 gnd
port 2 nsew
rlabel metal3 s 59888 34015 59986 34113 4 gnd
port 2 nsew
rlabel metal3 s 61127 32458 61225 32556 4 gnd
port 2 nsew
rlabel metal3 s 60702 31236 60800 31334 4 vdd
port 1 nsew
rlabel metal3 s 59492 30855 59590 30953 4 vdd
port 1 nsew
rlabel metal3 s 59492 34015 59590 34113 4 vdd
port 1 nsew
rlabel metal3 s 61127 31668 61225 31766 4 gnd
port 2 nsew
rlabel metal3 s 60270 33248 60368 33346 4 vdd
port 1 nsew
rlabel metal3 s 60702 32026 60800 32124 4 vdd
port 1 nsew
rlabel metal3 s 61127 29714 61225 29812 4 gnd
port 2 nsew
rlabel metal3 s 59888 32435 59986 32533 4 gnd
port 2 nsew
rlabel metal3 s 54552 33857 54650 33955 4 gnd
port 2 nsew
rlabel metal3 s 54552 30460 54650 30558 4 gnd
port 2 nsew
rlabel metal3 s 54552 34173 54650 34271 4 gnd
port 2 nsew
rlabel metal3 s 54552 34963 54650 35061 4 gnd
port 2 nsew
rlabel metal3 s 54552 36227 54650 36325 4 gnd
port 2 nsew
rlabel metal3 s 54552 38597 54650 38695 4 gnd
port 2 nsew
rlabel metal3 s 54552 33383 54650 33481 4 gnd
port 2 nsew
rlabel metal3 s 54552 32040 54650 32138 4 gnd
port 2 nsew
rlabel metal3 s 54552 38913 54650 39011 4 gnd
port 2 nsew
rlabel metal3 s 54552 38123 54650 38221 4 gnd
port 2 nsew
rlabel metal3 s 54552 39150 54650 39248 4 gnd
port 2 nsew
rlabel metal3 s 57592 39150 57690 39248 4 gnd
port 2 nsew
rlabel metal3 s 54552 37570 54650 37668 4 gnd
port 2 nsew
rlabel metal3 s 54552 30223 54650 30321 4 gnd
port 2 nsew
rlabel metal3 s 54552 34647 54650 34745 4 gnd
port 2 nsew
rlabel metal3 s 54552 37017 54650 37115 4 gnd
port 2 nsew
rlabel metal3 s 54552 34410 54650 34508 4 gnd
port 2 nsew
rlabel metal3 s 54552 32593 54650 32691 4 gnd
port 2 nsew
rlabel metal3 s 54552 29433 54650 29531 4 gnd
port 2 nsew
rlabel metal3 s 55944 39150 56042 39248 4 vdd
port 1 nsew
rlabel metal3 s 54552 30697 54650 30795 4 gnd
port 2 nsew
rlabel metal3 s 54552 35753 54650 35851 4 gnd
port 2 nsew
rlabel metal3 s 54552 29907 54650 30005 4 gnd
port 2 nsew
rlabel metal3 s 54552 33067 54650 33165 4 gnd
port 2 nsew
rlabel metal3 s 54552 31250 54650 31348 4 gnd
port 2 nsew
rlabel metal3 s 54552 36780 54650 36878 4 gnd
port 2 nsew
rlabel metal3 s 54552 35990 54650 36088 4 gnd
port 2 nsew
rlabel metal3 s 54552 38360 54650 38458 4 gnd
port 2 nsew
rlabel metal3 s 54552 32830 54650 32928 4 gnd
port 2 nsew
rlabel metal3 s 54552 36543 54650 36641 4 gnd
port 2 nsew
rlabel metal3 s 54552 35200 54650 35298 4 gnd
port 2 nsew
rlabel metal3 s 54552 31487 54650 31585 4 gnd
port 2 nsew
rlabel metal3 s 54552 32277 54650 32375 4 gnd
port 2 nsew
rlabel metal3 s 54552 37333 54650 37431 4 gnd
port 2 nsew
rlabel metal3 s 54552 31803 54650 31901 4 gnd
port 2 nsew
rlabel metal3 s 54552 31013 54650 31111 4 gnd
port 2 nsew
rlabel metal3 s 54552 29670 54650 29768 4 gnd
port 2 nsew
rlabel metal3 s 54552 37807 54650 37905 4 gnd
port 2 nsew
rlabel metal3 s 54552 33620 54650 33718 4 gnd
port 2 nsew
rlabel metal3 s 54552 35437 54650 35535 4 gnd
port 2 nsew
rlabel metal3 s 54552 24140 54650 24238 4 gnd
port 2 nsew
rlabel metal3 s 54552 24930 54650 25028 4 gnd
port 2 nsew
rlabel metal3 s 54552 28880 54650 28978 4 gnd
port 2 nsew
rlabel metal3 s 54552 22797 54650 22895 4 gnd
port 2 nsew
rlabel metal3 s 54552 29117 54650 29215 4 gnd
port 2 nsew
rlabel metal3 s 54552 23350 54650 23448 4 gnd
port 2 nsew
rlabel metal3 s 54552 23113 54650 23211 4 gnd
port 2 nsew
rlabel metal3 s 54552 25167 54650 25265 4 gnd
port 2 nsew
rlabel metal3 s 54552 22007 54650 22105 4 gnd
port 2 nsew
rlabel metal3 s 54552 22560 54650 22658 4 gnd
port 2 nsew
rlabel metal3 s 54552 22323 54650 22421 4 gnd
port 2 nsew
rlabel metal3 s 54552 26510 54650 26608 4 gnd
port 2 nsew
rlabel metal3 s 54552 25483 54650 25581 4 gnd
port 2 nsew
rlabel metal3 s 54552 27063 54650 27161 4 gnd
port 2 nsew
rlabel metal3 s 54552 19953 54650 20051 4 gnd
port 2 nsew
rlabel metal3 s 54552 27300 54650 27398 4 gnd
port 2 nsew
rlabel metal3 s 54552 21533 54650 21631 4 gnd
port 2 nsew
rlabel metal3 s 54552 25957 54650 26055 4 gnd
port 2 nsew
rlabel metal3 s 54552 21217 54650 21315 4 gnd
port 2 nsew
rlabel metal3 s 54552 20743 54650 20841 4 gnd
port 2 nsew
rlabel metal3 s 54552 27537 54650 27635 4 gnd
port 2 nsew
rlabel metal3 s 54552 26273 54650 26371 4 gnd
port 2 nsew
rlabel metal3 s 54552 28643 54650 28741 4 gnd
port 2 nsew
rlabel metal3 s 54552 26747 54650 26845 4 gnd
port 2 nsew
rlabel metal3 s 54552 28327 54650 28425 4 gnd
port 2 nsew
rlabel metal3 s 54552 28090 54650 28188 4 gnd
port 2 nsew
rlabel metal3 s 54552 23903 54650 24001 4 gnd
port 2 nsew
rlabel metal3 s 54552 23587 54650 23685 4 gnd
port 2 nsew
rlabel metal3 s 54552 20980 54650 21078 4 gnd
port 2 nsew
rlabel metal3 s 54552 24377 54650 24475 4 gnd
port 2 nsew
rlabel metal3 s 54552 20427 54650 20525 4 gnd
port 2 nsew
rlabel metal3 s 54552 19637 54650 19735 4 gnd
port 2 nsew
rlabel metal3 s 54552 20190 54650 20288 4 gnd
port 2 nsew
rlabel metal3 s 54552 21770 54650 21868 4 gnd
port 2 nsew
rlabel metal3 s 54552 25720 54650 25818 4 gnd
port 2 nsew
rlabel metal3 s 54552 24693 54650 24791 4 gnd
port 2 nsew
rlabel metal3 s 54552 27853 54650 27951 4 gnd
port 2 nsew
rlabel metal3 s 59888 27300 59986 27398 4 gnd
port 2 nsew
rlabel metal3 s 59888 29275 59986 29373 4 gnd
port 2 nsew
rlabel metal3 s 59492 28485 59590 28583 4 vdd
port 1 nsew
rlabel metal3 s 59492 25325 59590 25423 4 vdd
port 1 nsew
rlabel metal3 s 61127 26554 61225 26652 4 gnd
port 2 nsew
rlabel metal3 s 60702 26928 60800 27026 4 vdd
port 1 nsew
rlabel metal3 s 60702 26138 60800 26236 4 vdd
port 1 nsew
rlabel metal3 s 60702 28508 60800 28606 4 vdd
port 1 nsew
rlabel metal3 s 59492 29275 59590 29373 4 vdd
port 1 nsew
rlabel metal3 s 60702 24558 60800 24656 4 vdd
port 1 nsew
rlabel metal3 s 59888 25325 59986 25423 4 gnd
port 2 nsew
rlabel metal3 s 60270 26928 60368 27026 4 vdd
port 1 nsew
rlabel metal3 s 59888 24930 59986 25028 4 gnd
port 2 nsew
rlabel metal3 s 59888 24535 59986 24633 4 gnd
port 2 nsew
rlabel metal3 s 59888 26905 59986 27003 4 gnd
port 2 nsew
rlabel metal3 s 59492 27695 59590 27793 4 vdd
port 1 nsew
rlabel metal3 s 60270 24916 60368 25014 4 vdd
port 1 nsew
rlabel metal3 s 60270 25348 60368 25446 4 vdd
port 1 nsew
rlabel metal3 s 59492 27300 59590 27398 4 vdd
port 1 nsew
rlabel metal3 s 60702 29298 60800 29396 4 vdd
port 1 nsew
rlabel metal3 s 59492 26510 59590 26608 4 vdd
port 1 nsew
rlabel metal3 s 61127 24974 61225 25072 4 gnd
port 2 nsew
rlabel metal3 s 60270 25706 60368 25804 4 vdd
port 1 nsew
rlabel metal3 s 59888 26510 59986 26608 4 gnd
port 2 nsew
rlabel metal3 s 59492 26115 59590 26213 4 vdd
port 1 nsew
rlabel metal3 s 59492 24930 59590 25028 4 vdd
port 1 nsew
rlabel metal3 s 60270 28076 60368 28174 4 vdd
port 1 nsew
rlabel metal3 s 61127 28508 61225 28606 4 gnd
port 2 nsew
rlabel metal3 s 59492 28880 59590 28978 4 vdd
port 1 nsew
rlabel metal3 s 61127 29298 61225 29396 4 gnd
port 2 nsew
rlabel metal3 s 60702 28866 60800 28964 4 vdd
port 1 nsew
rlabel metal3 s 61127 25764 61225 25862 4 gnd
port 2 nsew
rlabel metal3 s 60270 26496 60368 26594 4 vdd
port 1 nsew
rlabel metal3 s 60702 28076 60800 28174 4 vdd
port 1 nsew
rlabel metal3 s 59888 26115 59986 26213 4 gnd
port 2 nsew
rlabel metal3 s 59888 25720 59986 25818 4 gnd
port 2 nsew
rlabel metal3 s 60270 26138 60368 26236 4 vdd
port 1 nsew
rlabel metal3 s 60702 27286 60800 27384 4 vdd
port 1 nsew
rlabel metal3 s 60270 28508 60368 28606 4 vdd
port 1 nsew
rlabel metal3 s 61127 27344 61225 27442 4 gnd
port 2 nsew
rlabel metal3 s 61127 24558 61225 24656 4 gnd
port 2 nsew
rlabel metal3 s 60702 26496 60800 26594 4 vdd
port 1 nsew
rlabel metal3 s 60702 24916 60800 25014 4 vdd
port 1 nsew
rlabel metal3 s 59492 28090 59590 28188 4 vdd
port 1 nsew
rlabel metal3 s 61127 28134 61225 28232 4 gnd
port 2 nsew
rlabel metal3 s 59888 28485 59986 28583 4 gnd
port 2 nsew
rlabel metal3 s 60270 27286 60368 27384 4 vdd
port 1 nsew
rlabel metal3 s 59888 28090 59986 28188 4 gnd
port 2 nsew
rlabel metal3 s 60702 25348 60800 25446 4 vdd
port 1 nsew
rlabel metal3 s 61127 27718 61225 27816 4 gnd
port 2 nsew
rlabel metal3 s 61127 28924 61225 29022 4 gnd
port 2 nsew
rlabel metal3 s 60702 27718 60800 27816 4 vdd
port 1 nsew
rlabel metal3 s 59492 25720 59590 25818 4 vdd
port 1 nsew
rlabel metal3 s 59492 24535 59590 24633 4 vdd
port 1 nsew
rlabel metal3 s 60270 28866 60368 28964 4 vdd
port 1 nsew
rlabel metal3 s 60270 29298 60368 29396 4 vdd
port 1 nsew
rlabel metal3 s 60702 25706 60800 25804 4 vdd
port 1 nsew
rlabel metal3 s 60270 24558 60368 24656 4 vdd
port 1 nsew
rlabel metal3 s 61127 25348 61225 25446 4 gnd
port 2 nsew
rlabel metal3 s 61127 26928 61225 27026 4 gnd
port 2 nsew
rlabel metal3 s 59888 28880 59986 28978 4 gnd
port 2 nsew
rlabel metal3 s 60270 27718 60368 27816 4 vdd
port 1 nsew
rlabel metal3 s 59888 27695 59986 27793 4 gnd
port 2 nsew
rlabel metal3 s 59492 26905 59590 27003 4 vdd
port 1 nsew
rlabel metal3 s 61127 26138 61225 26236 4 gnd
port 2 nsew
rlabel metal3 s 60270 23336 60368 23434 4 vdd
port 1 nsew
rlabel metal3 s 60270 22546 60368 22644 4 vdd
port 1 nsew
rlabel metal3 s 59888 21375 59986 21473 4 gnd
port 2 nsew
rlabel metal3 s 59492 19795 59590 19893 4 vdd
port 1 nsew
rlabel metal3 s 61127 22188 61225 22286 4 gnd
port 2 nsew
rlabel metal3 s 60270 20608 60368 20706 4 vdd
port 1 nsew
rlabel metal3 s 59492 22165 59590 22263 4 vdd
port 1 nsew
rlabel metal3 s 60702 24126 60800 24224 4 vdd
port 1 nsew
rlabel metal3 s 61127 23768 61225 23866 4 gnd
port 2 nsew
rlabel metal3 s 60702 21398 60800 21496 4 vdd
port 1 nsew
rlabel metal3 s 59492 22560 59590 22658 4 vdd
port 1 nsew
rlabel metal3 s 59492 23350 59590 23448 4 vdd
port 1 nsew
rlabel metal3 s 61127 22978 61225 23076 4 gnd
port 2 nsew
rlabel metal3 s 61127 22604 61225 22702 4 gnd
port 2 nsew
rlabel metal3 s 59888 21770 59986 21868 4 gnd
port 2 nsew
rlabel metal3 s 60270 19818 60368 19916 4 vdd
port 1 nsew
rlabel metal3 s 60270 21398 60368 21496 4 vdd
port 1 nsew
rlabel metal3 s 59492 20190 59590 20288 4 vdd
port 1 nsew
rlabel metal3 s 61127 20234 61225 20332 4 gnd
port 2 nsew
rlabel metal3 s 60702 20176 60800 20274 4 vdd
port 1 nsew
rlabel metal3 s 59888 20980 59986 21078 4 gnd
port 2 nsew
rlabel metal3 s 59492 20980 59590 21078 4 vdd
port 1 nsew
rlabel metal3 s 60702 21756 60800 21854 4 vdd
port 1 nsew
rlabel metal3 s 59888 19795 59986 19893 4 gnd
port 2 nsew
rlabel metal3 s 59492 24140 59590 24238 4 vdd
port 1 nsew
rlabel metal3 s 60270 22188 60368 22286 4 vdd
port 1 nsew
rlabel metal3 s 61127 21398 61225 21496 4 gnd
port 2 nsew
rlabel metal3 s 61127 21024 61225 21122 4 gnd
port 2 nsew
rlabel metal3 s 60702 23336 60800 23434 4 vdd
port 1 nsew
rlabel metal3 s 61127 20608 61225 20706 4 gnd
port 2 nsew
rlabel metal3 s 60270 24126 60368 24224 4 vdd
port 1 nsew
rlabel metal3 s 59492 21770 59590 21868 4 vdd
port 1 nsew
rlabel metal3 s 60702 22978 60800 23076 4 vdd
port 1 nsew
rlabel metal3 s 59492 21375 59590 21473 4 vdd
port 1 nsew
rlabel metal3 s 59888 24140 59986 24238 4 gnd
port 2 nsew
rlabel metal3 s 60270 20176 60368 20274 4 vdd
port 1 nsew
rlabel metal3 s 60270 20966 60368 21064 4 vdd
port 1 nsew
rlabel metal3 s 60702 22546 60800 22644 4 vdd
port 1 nsew
rlabel metal3 s 59888 22165 59986 22263 4 gnd
port 2 nsew
rlabel metal3 s 59888 20190 59986 20288 4 gnd
port 2 nsew
rlabel metal3 s 60270 23768 60368 23866 4 vdd
port 1 nsew
rlabel metal3 s 59888 23350 59986 23448 4 gnd
port 2 nsew
rlabel metal3 s 60702 22188 60800 22286 4 vdd
port 1 nsew
rlabel metal3 s 60702 19818 60800 19916 4 vdd
port 1 nsew
rlabel metal3 s 61127 19818 61225 19916 4 gnd
port 2 nsew
rlabel metal3 s 61127 23394 61225 23492 4 gnd
port 2 nsew
rlabel metal3 s 59888 20585 59986 20683 4 gnd
port 2 nsew
rlabel metal3 s 59492 22955 59590 23053 4 vdd
port 1 nsew
rlabel metal3 s 59888 22955 59986 23053 4 gnd
port 2 nsew
rlabel metal3 s 60702 23768 60800 23866 4 vdd
port 1 nsew
rlabel metal3 s 60702 20608 60800 20706 4 vdd
port 1 nsew
rlabel metal3 s 59888 23745 59986 23843 4 gnd
port 2 nsew
rlabel metal3 s 60702 20966 60800 21064 4 vdd
port 1 nsew
rlabel metal3 s 59492 20585 59590 20683 4 vdd
port 1 nsew
rlabel metal3 s 59492 23745 59590 23843 4 vdd
port 1 nsew
rlabel metal3 s 60270 22978 60368 23076 4 vdd
port 1 nsew
rlabel metal3 s 61127 21814 61225 21912 4 gnd
port 2 nsew
rlabel metal3 s 60270 21756 60368 21854 4 vdd
port 1 nsew
rlabel metal3 s 59888 22560 59986 22658 4 gnd
port 2 nsew
rlabel metal3 s 61127 24184 61225 24282 4 gnd
port 2 nsew
rlabel metal3 s 64541 20608 64639 20706 4 gnd
port 2 nsew
rlabel metal3 s 62906 20585 63004 20683 4 vdd
port 1 nsew
rlabel metal3 s 64116 21398 64214 21496 4 vdd
port 1 nsew
rlabel metal3 s 63302 21375 63400 21473 4 gnd
port 2 nsew
rlabel metal3 s 63302 19795 63400 19893 4 gnd
port 2 nsew
rlabel metal3 s 63684 19818 63782 19916 4 vdd
port 1 nsew
rlabel metal3 s 63302 20585 63400 20683 4 gnd
port 2 nsew
rlabel metal3 s 64541 19818 64639 19916 4 gnd
port 2 nsew
rlabel metal3 s 63684 21398 63782 21496 4 vdd
port 1 nsew
rlabel metal3 s 63684 20608 63782 20706 4 vdd
port 1 nsew
rlabel metal3 s 64541 21398 64639 21496 4 gnd
port 2 nsew
rlabel metal3 s 62906 21375 63004 21473 4 vdd
port 1 nsew
rlabel metal3 s 64116 20608 64214 20706 4 vdd
port 1 nsew
rlabel metal3 s 64116 19818 64214 19916 4 vdd
port 1 nsew
rlabel metal3 s 62906 19795 63004 19893 4 vdd
port 1 nsew
rlabel metal3 s 42505 12718 42603 12816 4 vdd
port 1 nsew
rlabel metal3 s 45432 11169 45530 11267 4 gnd
port 2 nsew
rlabel metal3 s 48240 13309 48338 13407 4 vdd
port 1 nsew
rlabel metal3 s 48864 13309 48962 13407 4 vdd
port 1 nsew
rlabel metal3 s 49488 13309 49586 13407 4 vdd
port 1 nsew
rlabel metal3 s 46680 11169 46778 11267 4 gnd
port 2 nsew
rlabel metal3 s 49607 12718 49705 12816 4 vdd
port 1 nsew
rlabel metal3 s 46992 13309 47090 13407 4 vdd
port 1 nsew
rlabel metal3 s 44496 13309 44594 13407 4 vdd
port 1 nsew
rlabel metal3 s 47616 13309 47714 13407 4 vdd
port 1 nsew
rlabel metal3 s 42936 11169 43034 11267 4 gnd
port 2 nsew
rlabel metal3 s 45863 12718 45961 12816 4 vdd
port 1 nsew
rlabel metal3 s 43872 13309 43970 13407 4 vdd
port 1 nsew
rlabel metal3 s 44184 11169 44282 11267 4 gnd
port 2 nsew
rlabel metal3 s 43367 12718 43465 12816 4 vdd
port 1 nsew
rlabel metal3 s 47497 12718 47595 12816 4 vdd
port 1 nsew
rlabel metal3 s 42624 13309 42722 13407 4 vdd
port 1 nsew
rlabel metal3 s 43753 12718 43851 12816 4 vdd
port 1 nsew
rlabel metal3 s 48745 12718 48843 12816 4 vdd
port 1 nsew
rlabel metal3 s 47928 11169 48026 11267 4 gnd
port 2 nsew
rlabel metal3 s 44615 12718 44713 12816 4 vdd
port 1 nsew
rlabel metal3 s 42000 13309 42098 13407 4 vdd
port 1 nsew
rlabel metal3 s 48359 12718 48457 12816 4 vdd
port 1 nsew
rlabel metal3 s 41688 11169 41786 11267 4 gnd
port 2 nsew
rlabel metal3 s 45744 13309 45842 13407 4 vdd
port 1 nsew
rlabel metal3 s 43248 13309 43346 13407 4 vdd
port 1 nsew
rlabel metal3 s 42119 12718 42217 12816 4 vdd
port 1 nsew
rlabel metal3 s 46368 13309 46466 13407 4 vdd
port 1 nsew
rlabel metal3 s 47111 12718 47209 12816 4 vdd
port 1 nsew
rlabel metal3 s 46249 12718 46347 12816 4 vdd
port 1 nsew
rlabel metal3 s 45001 12718 45099 12816 4 vdd
port 1 nsew
rlabel metal3 s 45120 13309 45218 13407 4 vdd
port 1 nsew
rlabel metal3 s 49176 11169 49274 11267 4 gnd
port 2 nsew
rlabel metal3 s 37632 13309 37730 13407 4 vdd
port 1 nsew
rlabel metal3 s 38256 13309 38354 13407 4 vdd
port 1 nsew
rlabel metal3 s 40128 13309 40226 13407 4 vdd
port 1 nsew
rlabel metal3 s 37008 13309 37106 13407 4 vdd
port 1 nsew
rlabel metal3 s 36696 11169 36794 11267 4 gnd
port 2 nsew
rlabel metal3 s 40440 11169 40538 11267 4 gnd
port 2 nsew
rlabel metal3 s 35760 13309 35858 13407 4 vdd
port 1 nsew
rlabel metal3 s 35448 11169 35546 11267 4 gnd
port 2 nsew
rlabel metal3 s 37127 12718 37225 12816 4 vdd
port 1 nsew
rlabel metal3 s 41257 12718 41355 12816 4 vdd
port 1 nsew
rlabel metal3 s 39504 13309 39602 13407 4 vdd
port 1 nsew
rlabel metal3 s 36265 12718 36363 12816 4 vdd
port 1 nsew
rlabel metal3 s 38880 13309 38978 13407 4 vdd
port 1 nsew
rlabel metal3 s 33769 12718 33867 12816 4 vdd
port 1 nsew
rlabel metal3 s 41376 13309 41474 13407 4 vdd
port 1 nsew
rlabel metal3 s 34200 11169 34298 11267 4 gnd
port 2 nsew
rlabel metal3 s 33888 13309 33986 13407 4 vdd
port 1 nsew
rlabel metal3 s 38375 12718 38473 12816 4 vdd
port 1 nsew
rlabel metal3 s 37944 11169 38042 11267 4 gnd
port 2 nsew
rlabel metal3 s 40871 12718 40969 12816 4 vdd
port 1 nsew
rlabel metal3 s 36384 13309 36482 13407 4 vdd
port 1 nsew
rlabel metal3 s 34631 12718 34729 12816 4 vdd
port 1 nsew
rlabel metal3 s 38761 12718 38859 12816 4 vdd
port 1 nsew
rlabel metal3 s 35017 12718 35115 12816 4 vdd
port 1 nsew
rlabel metal3 s 39192 11169 39290 11267 4 gnd
port 2 nsew
rlabel metal3 s 37513 12718 37611 12816 4 vdd
port 1 nsew
rlabel metal3 s 35136 13309 35234 13407 4 vdd
port 1 nsew
rlabel metal3 s 40009 12718 40107 12816 4 vdd
port 1 nsew
rlabel metal3 s 34512 13309 34610 13407 4 vdd
port 1 nsew
rlabel metal3 s 40752 13309 40850 13407 4 vdd
port 1 nsew
rlabel metal3 s 39623 12718 39721 12816 4 vdd
port 1 nsew
rlabel metal3 s 35879 12718 35977 12816 4 vdd
port 1 nsew
rlabel metal3 s 34027 8676 34125 8774 4 gnd
port 2 nsew
rlabel metal3 s 33953 5180 34051 5278 4 gnd
port 2 nsew
rlabel metal3 s 33838 4978 33936 5076 4 gnd
port 2 nsew
rlabel metal3 s 38830 4978 38928 5076 4 gnd
port 2 nsew
rlabel metal3 s 38945 5180 39043 5278 4 gnd
port 2 nsew
rlabel metal3 s 38937 7902 39035 8000 4 vdd
port 1 nsew
rlabel metal3 s 33832 5512 33930 5610 4 vdd
port 1 nsew
rlabel metal3 s 38949 6742 39047 6840 4 gnd
port 2 nsew
rlabel metal3 s 38824 5512 38922 5610 4 vdd
port 1 nsew
rlabel metal3 s 38835 5949 38933 6047 4 gnd
port 2 nsew
rlabel metal3 s 33957 7064 34055 7162 4 vdd
port 1 nsew
rlabel metal3 s 33843 5949 33941 6047 4 gnd
port 2 nsew
rlabel metal3 s 33945 7902 34043 8000 4 vdd
port 1 nsew
rlabel metal3 s 33852 4562 33950 4660 4 vdd
port 1 nsew
rlabel metal3 s 38949 7064 39047 7162 4 vdd
port 1 nsew
rlabel metal3 s 38844 4562 38942 4660 4 vdd
port 1 nsew
rlabel metal3 s 39019 8676 39117 8774 4 gnd
port 2 nsew
rlabel metal3 s 33957 6742 34055 6840 4 gnd
port 2 nsew
rlabel metal3 s 43822 4978 43920 5076 4 gnd
port 2 nsew
rlabel metal3 s 44011 8676 44109 8774 4 gnd
port 2 nsew
rlabel metal3 s 48933 6742 49031 6840 4 gnd
port 2 nsew
rlabel metal3 s 43941 6742 44039 6840 4 gnd
port 2 nsew
rlabel metal3 s 48828 4562 48926 4660 4 vdd
port 1 nsew
rlabel metal3 s 48819 5949 48917 6047 4 gnd
port 2 nsew
rlabel metal3 s 43836 4562 43934 4660 4 vdd
port 1 nsew
rlabel metal3 s 49003 8676 49101 8774 4 gnd
port 2 nsew
rlabel metal3 s 43816 5512 43914 5610 4 vdd
port 1 nsew
rlabel metal3 s 43937 5180 44035 5278 4 gnd
port 2 nsew
rlabel metal3 s 43929 7902 44027 8000 4 vdd
port 1 nsew
rlabel metal3 s 43941 7064 44039 7162 4 vdd
port 1 nsew
rlabel metal3 s 48929 5180 49027 5278 4 gnd
port 2 nsew
rlabel metal3 s 48808 5512 48906 5610 4 vdd
port 1 nsew
rlabel metal3 s 48921 7902 49019 8000 4 vdd
port 1 nsew
rlabel metal3 s 48933 7064 49031 7162 4 vdd
port 1 nsew
rlabel metal3 s 48814 4978 48912 5076 4 gnd
port 2 nsew
rlabel metal3 s 43827 5949 43925 6047 4 gnd
port 2 nsew
rlabel metal3 s 62906 16635 63004 16733 4 vdd
port 1 nsew
rlabel metal3 s 62906 17425 63004 17523 4 vdd
port 1 nsew
rlabel metal3 s 60702 14288 60800 14386 4 vdd
port 1 nsew
rlabel metal3 s 60270 16658 60368 16756 4 vdd
port 1 nsew
rlabel metal3 s 65400 14265 65498 14363 4 gnd
port 2 nsew
rlabel metal3 s 59888 15055 59986 15153 4 gnd
port 2 nsew
rlabel metal3 s 59492 18610 59590 18708 4 vdd
port 1 nsew
rlabel metal3 s 60702 14646 60800 14744 4 vdd
port 1 nsew
rlabel metal3 s 63302 17425 63400 17523 4 gnd
port 2 nsew
rlabel metal3 s 61127 16658 61225 16756 4 gnd
port 2 nsew
rlabel metal3 s 60270 17448 60368 17546 4 vdd
port 1 nsew
rlabel metal3 s 60702 18238 60800 18336 4 vdd
port 1 nsew
rlabel metal3 s 59492 16635 59590 16733 4 vdd
port 1 nsew
rlabel metal3 s 61127 14288 61225 14386 4 gnd
port 2 nsew
rlabel metal3 s 61127 17074 61225 17172 4 gnd
port 2 nsew
rlabel metal3 s 59492 18215 59590 18313 4 vdd
port 1 nsew
rlabel metal3 s 60702 17448 60800 17546 4 vdd
port 1 nsew
rlabel metal3 s 60702 15868 60800 15966 4 vdd
port 1 nsew
rlabel metal3 s 59492 15450 59590 15548 4 vdd
port 1 nsew
rlabel metal3 s 63681 17432 63779 17530 4 vdd
port 1 nsew
rlabel metal3 s 60702 17806 60800 17904 4 vdd
port 1 nsew
rlabel metal3 s 60270 17016 60368 17114 4 vdd
port 1 nsew
rlabel metal3 s 61127 17448 61225 17546 4 gnd
port 2 nsew
rlabel metal3 s 59492 15845 59590 15943 4 vdd
port 1 nsew
rlabel metal3 s 63681 14272 63779 14370 4 vdd
port 1 nsew
rlabel metal3 s 59888 16635 59986 16733 4 gnd
port 2 nsew
rlabel metal3 s 60270 19386 60368 19484 4 vdd
port 1 nsew
rlabel metal3 s 59888 15845 59986 15943 4 gnd
port 2 nsew
rlabel metal3 s 61127 18238 61225 18336 4 gnd
port 2 nsew
rlabel metal3 s 59492 16240 59590 16338 4 vdd
port 1 nsew
rlabel metal3 s 59492 17030 59590 17128 4 vdd
port 1 nsew
rlabel metal3 s 60702 16658 60800 16756 4 vdd
port 1 nsew
rlabel metal3 s 60270 14646 60368 14744 4 vdd
port 1 nsew
rlabel metal3 s 62906 19005 63004 19103 4 vdd
port 1 nsew
rlabel metal3 s 59888 17820 59986 17918 4 gnd
port 2 nsew
rlabel metal3 s 61127 17864 61225 17962 4 gnd
port 2 nsew
rlabel metal3 s 63302 19005 63400 19103 4 gnd
port 2 nsew
rlabel metal3 s 61127 15078 61225 15176 4 gnd
port 2 nsew
rlabel metal3 s 64106 15062 64204 15160 4 gnd
port 2 nsew
rlabel metal3 s 61127 15494 61225 15592 4 gnd
port 2 nsew
rlabel metal3 s 60702 19386 60800 19484 4 vdd
port 1 nsew
rlabel metal3 s 65400 16635 65498 16733 4 gnd
port 2 nsew
rlabel metal3 s 61127 19444 61225 19542 4 gnd
port 2 nsew
rlabel metal3 s 62906 14265 63004 14363 4 vdd
port 1 nsew
rlabel metal3 s 59492 14265 59590 14363 4 vdd
port 1 nsew
rlabel metal3 s 59888 18610 59986 18708 4 gnd
port 2 nsew
rlabel metal3 s 63302 14265 63400 14363 4 gnd
port 2 nsew
rlabel metal3 s 60702 16226 60800 16324 4 vdd
port 1 nsew
rlabel metal3 s 60270 15868 60368 15966 4 vdd
port 1 nsew
rlabel metal3 s 60702 17016 60800 17114 4 vdd
port 1 nsew
rlabel metal3 s 63681 15062 63779 15160 4 vdd
port 1 nsew
rlabel metal3 s 63684 19028 63782 19126 4 vdd
port 1 nsew
rlabel metal3 s 61127 14704 61225 14802 4 gnd
port 2 nsew
rlabel metal3 s 64116 19028 64214 19126 4 vdd
port 1 nsew
rlabel metal3 s 59888 17030 59986 17128 4 gnd
port 2 nsew
rlabel metal3 s 60270 17806 60368 17904 4 vdd
port 1 nsew
rlabel metal3 s 65996 19005 66094 19103 4 gnd
port 2 nsew
rlabel metal3 s 60702 15436 60800 15534 4 vdd
port 1 nsew
rlabel metal3 s 63302 16635 63400 16733 4 gnd
port 2 nsew
rlabel metal3 s 60270 15436 60368 15534 4 vdd
port 1 nsew
rlabel metal3 s 59492 19005 59590 19103 4 vdd
port 1 nsew
rlabel metal3 s 64106 16642 64204 16740 4 gnd
port 2 nsew
rlabel metal3 s 59888 14265 59986 14363 4 gnd
port 2 nsew
rlabel metal3 s 63302 15055 63400 15153 4 gnd
port 2 nsew
rlabel metal3 s 61127 19028 61225 19126 4 gnd
port 2 nsew
rlabel metal3 s 59888 15450 59986 15548 4 gnd
port 2 nsew
rlabel metal3 s 63681 16642 63779 16740 4 vdd
port 1 nsew
rlabel metal3 s 59888 19005 59986 19103 4 gnd
port 2 nsew
rlabel metal3 s 61127 16284 61225 16382 4 gnd
port 2 nsew
rlabel metal3 s 60702 19028 60800 19126 4 vdd
port 1 nsew
rlabel metal3 s 64541 19028 64639 19126 4 gnd
port 2 nsew
rlabel metal3 s 60702 15078 60800 15176 4 vdd
port 1 nsew
rlabel metal3 s 59888 17425 59986 17523 4 gnd
port 2 nsew
rlabel metal3 s 59888 18215 59986 18313 4 gnd
port 2 nsew
rlabel metal3 s 62906 15055 63004 15153 4 vdd
port 1 nsew
rlabel metal3 s 59492 14660 59590 14758 4 vdd
port 1 nsew
rlabel metal3 s 60270 14288 60368 14386 4 vdd
port 1 nsew
rlabel metal3 s 60270 18238 60368 18336 4 vdd
port 1 nsew
rlabel metal3 s 64106 17432 64204 17530 4 gnd
port 2 nsew
rlabel metal3 s 60270 15078 60368 15176 4 vdd
port 1 nsew
rlabel metal3 s 61127 18654 61225 18752 4 gnd
port 2 nsew
rlabel metal3 s 59492 19400 59590 19498 4 vdd
port 1 nsew
rlabel metal3 s 60270 18596 60368 18694 4 vdd
port 1 nsew
rlabel metal3 s 59888 14660 59986 14758 4 gnd
port 2 nsew
rlabel metal3 s 65004 14265 65102 14363 4 vdd
port 1 nsew
rlabel metal3 s 64106 14272 64204 14370 4 gnd
port 2 nsew
rlabel metal3 s 60702 18596 60800 18694 4 vdd
port 1 nsew
rlabel metal3 s 59492 17820 59590 17918 4 vdd
port 1 nsew
rlabel metal3 s 59492 15055 59590 15153 4 vdd
port 1 nsew
rlabel metal3 s 59888 19400 59986 19498 4 gnd
port 2 nsew
rlabel metal3 s 65600 19005 65698 19103 4 vdd
port 1 nsew
rlabel metal3 s 59492 17425 59590 17523 4 vdd
port 1 nsew
rlabel metal3 s 61127 15868 61225 15966 4 gnd
port 2 nsew
rlabel metal3 s 60270 19028 60368 19126 4 vdd
port 1 nsew
rlabel metal3 s 59888 16240 59986 16338 4 gnd
port 2 nsew
rlabel metal3 s 65004 16635 65102 16733 4 vdd
port 1 nsew
rlabel metal3 s 60270 16226 60368 16324 4 vdd
port 1 nsew
rlabel metal3 s 50855 12718 50953 12816 4 vdd
port 1 nsew
rlabel metal3 s 54552 16240 54650 16338 4 gnd
port 2 nsew
rlabel metal3 s 54552 14107 54650 14205 4 gnd
port 2 nsew
rlabel metal3 s 52608 13309 52706 13407 4 vdd
port 1 nsew
rlabel metal3 s 52920 11169 53018 11267 4 gnd
port 2 nsew
rlabel metal3 s 54552 19163 54650 19261 4 gnd
port 2 nsew
rlabel metal3 s 51984 13309 52082 13407 4 vdd
port 1 nsew
rlabel metal3 s 54552 18057 54650 18155 4 gnd
port 2 nsew
rlabel metal3 s 53232 13309 53330 13407 4 vdd
port 1 nsew
rlabel metal3 s 51241 12718 51339 12816 4 vdd
port 1 nsew
rlabel metal3 s 54552 13870 54650 13968 4 gnd
port 2 nsew
rlabel metal3 s 53856 13309 53954 13407 4 vdd
port 1 nsew
rlabel metal3 s 54552 19400 54650 19498 4 gnd
port 2 nsew
rlabel metal3 s 54552 16793 54650 16891 4 gnd
port 2 nsew
rlabel metal3 s 51672 11169 51770 11267 4 gnd
port 2 nsew
rlabel metal3 s 54552 15687 54650 15785 4 gnd
port 2 nsew
rlabel metal3 s 52103 12718 52201 12816 4 vdd
port 1 nsew
rlabel metal3 s 54552 17267 54650 17365 4 gnd
port 2 nsew
rlabel metal3 s 54552 18847 54650 18945 4 gnd
port 2 nsew
rlabel metal3 s 54552 17583 54650 17681 4 gnd
port 2 nsew
rlabel metal3 s 54552 17820 54650 17918 4 gnd
port 2 nsew
rlabel metal3 s 54552 14897 54650 14995 4 gnd
port 2 nsew
rlabel metal3 s 54552 18610 54650 18708 4 gnd
port 2 nsew
rlabel metal3 s 54552 16003 54650 16101 4 gnd
port 2 nsew
rlabel metal3 s 54552 17030 54650 17128 4 gnd
port 2 nsew
rlabel metal3 s 54552 15450 54650 15548 4 gnd
port 2 nsew
rlabel metal3 s 54552 15213 54650 15311 4 gnd
port 2 nsew
rlabel metal3 s 49993 12718 50091 12816 4 vdd
port 1 nsew
rlabel metal3 s 54918 13743 55016 13841 4 gnd
port 2 nsew
rlabel metal3 s 53351 12718 53449 12816 4 vdd
port 1 nsew
rlabel metal3 s 54552 14423 54650 14521 4 gnd
port 2 nsew
rlabel metal3 s 50736 13309 50834 13407 4 vdd
port 1 nsew
rlabel metal3 s 51360 13309 51458 13407 4 vdd
port 1 nsew
rlabel metal3 s 54552 14660 54650 14758 4 gnd
port 2 nsew
rlabel metal3 s 54552 18373 54650 18471 4 gnd
port 2 nsew
rlabel metal3 s 54552 16477 54650 16575 4 gnd
port 2 nsew
rlabel metal3 s 50112 13309 50210 13407 4 vdd
port 1 nsew
rlabel metal3 s 50424 11169 50522 11267 4 gnd
port 2 nsew
rlabel metal3 s 52489 12718 52587 12816 4 vdd
port 1 nsew
rlabel metal3 s 53544 2999 53642 3097 4 gnd
port 2 nsew
rlabel metal3 s 53544 4119 53642 4217 4 vdd
port 1 nsew
rlabel metal2 s 11663 49 11691 13129 4 p_en_bar0
port 5 nsew
rlabel metal2 s 11787 49 11815 13129 4 s_en0
port 6 nsew
rlabel metal2 s 11911 49 11939 13129 4 w_en0
port 7 nsew
rlabel metal2 s 7960 13606 7988 13634 4 wl_en0
port 8 nsew
rlabel metal2 s 55277 65269 55305 78433 4 s_en1
port 9 nsew
rlabel metal2 s 55401 65269 55429 78433 4 p_en_bar1
port 10 nsew
rlabel metal2 s 59262 64764 59290 64792 4 wl_en1
port 11 nsew
rlabel metal2 s 13643 3304 13671 3332 4 bank_wmask0_0
port 12 nsew
rlabel metal1 s 13912 4424 13972 4480 4 din0_0
port 13 nsew
rlabel metal1 s 18904 4424 18964 4480 4 din0_1
port 14 nsew
rlabel metal1 s 23896 4424 23956 4480 4 din0_2
port 15 nsew
rlabel metal1 s 28888 4424 28948 4480 4 din0_3
port 16 nsew
rlabel metal1 s 33880 4424 33940 4480 4 din0_4
port 17 nsew
rlabel metal1 s 38872 4424 38932 4480 4 din0_5
port 18 nsew
rlabel metal1 s 43864 4424 43924 4480 4 din0_6
port 19 nsew
rlabel metal1 s 48856 4424 48916 4480 4 din0_7
port 20 nsew
rlabel metal1 s 13761 6683 13807 6937 4 dout0_0
port 21 nsew
rlabel metal1 s 18753 6683 18799 6937 4 dout0_1
port 22 nsew
rlabel metal1 s 23745 6683 23791 6937 4 dout0_2
port 23 nsew
rlabel metal1 s 28737 6683 28783 6937 4 dout0_3
port 24 nsew
rlabel metal1 s 33729 6683 33775 6937 4 dout0_4
port 25 nsew
rlabel metal1 s 38721 6683 38767 6937 4 dout0_5
port 26 nsew
rlabel metal1 s 43713 6683 43759 6937 4 dout0_6
port 27 nsew
rlabel metal1 s 48705 6683 48751 6937 4 dout0_7
port 28 nsew
rlabel metal1 s 19 13919 47 21819 4 addr0_3
port 29 nsew
rlabel metal1 s 99 13919 127 21819 4 addr0_4
port 30 nsew
rlabel metal1 s 179 13919 207 21819 4 addr0_5
port 31 nsew
rlabel metal1 s 259 13919 287 21819 4 addr0_6
port 32 nsew
rlabel metal1 s 339 13919 367 21819 4 addr0_7
port 33 nsew
rlabel metal1 s 419 13919 447 21819 4 addr0_8
port 34 nsew
rlabel metal1 s 499 13919 527 21819 4 addr0_9
port 35 nsew
rlabel metal1 s 4310 689 4356 747 4 addr0_0
port 36 nsew
rlabel metal1 s 4434 2179 4480 2237 4 addr0_1
port 37 nsew
rlabel metal1 s 4558 3517 4604 3575 4 addr0_2
port 38 nsew
rlabel metal1 s 13761 71461 13807 71715 4 dout1_0
port 39 nsew
rlabel metal1 s 18753 71461 18799 71715 4 dout1_1
port 40 nsew
rlabel metal1 s 23745 71461 23791 71715 4 dout1_2
port 41 nsew
rlabel metal1 s 28737 71461 28783 71715 4 dout1_3
port 42 nsew
rlabel metal1 s 33729 71461 33775 71715 4 dout1_4
port 43 nsew
rlabel metal1 s 38721 71461 38767 71715 4 dout1_5
port 44 nsew
rlabel metal1 s 43713 71461 43759 71715 4 dout1_6
port 45 nsew
rlabel metal1 s 48705 71461 48751 71715 4 dout1_7
port 46 nsew
rlabel metal1 s 67203 13919 67231 21819 4 addr1_3
port 47 nsew
rlabel metal1 s 67123 13919 67151 21819 4 addr1_4
port 48 nsew
rlabel metal1 s 67043 13919 67071 21819 4 addr1_5
port 49 nsew
rlabel metal1 s 66963 13919 66991 21819 4 addr1_6
port 50 nsew
rlabel metal1 s 66883 13919 66911 21819 4 addr1_7
port 51 nsew
rlabel metal1 s 66803 13919 66831 21819 4 addr1_8
port 52 nsew
rlabel metal1 s 66723 13919 66751 21819 4 addr1_9
port 53 nsew
rlabel metal1 s 62770 77651 62816 77709 4 addr1_0
port 54 nsew
rlabel metal1 s 62646 76161 62692 76219 4 addr1_1
port 55 nsew
rlabel metal1 s 62522 74823 62568 74881 4 addr1_2
port 56 nsew
<< properties >>
string FIXED_BBOX 0 0 67334 78384
string GDS_END 7724530
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 7109278
<< end >>
