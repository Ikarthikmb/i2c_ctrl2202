magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -36 679 404 1471
<< locali >>
rect 0 1397 368 1431
rect 64 636 98 702
rect 179 652 213 686
rect 0 -17 368 17
use sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_0  sky130_sram_1kbyte_1rw1r_8x1024_8_pinv_0_0
timestamp 1644511149
transform 1 0 0 0 1 0
box -36 -17 404 1471
<< labels >>
rlabel locali s 196 669 196 669 4 Z
port 1 nsew
rlabel locali s 81 669 81 669 4 A
port 2 nsew
rlabel locali s 184 0 184 0 4 gnd
port 3 nsew
rlabel locali s 184 1414 184 1414 4 vdd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 368 1414
string GDS_END 146574
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 145744
<< end >>
