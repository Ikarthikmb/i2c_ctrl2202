/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/rf_nfet_20v0_withptap_iso/sky130_fd_pr__rf_nfet_20v0_withptap_iso.spice