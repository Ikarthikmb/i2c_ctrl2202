/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/cap_var_hvt/sky130_fd_pr__cap_var_hvt.model.spice