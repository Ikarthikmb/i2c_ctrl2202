magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect 5751 816 6885 1140
rect 5751 600 6245 816
<< pwell >>
rect 3531 1277 4802 1415
rect 3486 625 4804 1277
rect 4990 698 5684 950
<< mvnmos >>
rect 3565 651 3665 1251
rect 3721 651 3821 1251
rect 3877 651 3977 1251
rect 4033 651 4133 1251
rect 4189 651 4289 1251
rect 4345 651 4445 1251
rect 4625 651 4725 1251
rect 5069 724 5169 924
rect 5225 724 5325 924
rect 5505 724 5605 924
<< mvpmos >>
rect 5870 666 5970 966
rect 6026 666 6126 966
rect 6310 882 6510 966
rect 6566 882 6766 966
<< mvndiff >>
rect 3512 1239 3565 1251
rect 3512 1205 3520 1239
rect 3554 1205 3565 1239
rect 3512 1171 3565 1205
rect 3512 1137 3520 1171
rect 3554 1137 3565 1171
rect 3512 1103 3565 1137
rect 3512 1069 3520 1103
rect 3554 1069 3565 1103
rect 3512 1035 3565 1069
rect 3512 1001 3520 1035
rect 3554 1001 3565 1035
rect 3512 967 3565 1001
rect 3512 933 3520 967
rect 3554 933 3565 967
rect 3512 899 3565 933
rect 3512 865 3520 899
rect 3554 865 3565 899
rect 3512 831 3565 865
rect 3512 797 3520 831
rect 3554 797 3565 831
rect 3512 763 3565 797
rect 3512 729 3520 763
rect 3554 729 3565 763
rect 3512 651 3565 729
rect 3665 1239 3721 1251
rect 3665 1205 3676 1239
rect 3710 1205 3721 1239
rect 3665 1171 3721 1205
rect 3665 1137 3676 1171
rect 3710 1137 3721 1171
rect 3665 1103 3721 1137
rect 3665 1069 3676 1103
rect 3710 1069 3721 1103
rect 3665 1035 3721 1069
rect 3665 1001 3676 1035
rect 3710 1001 3721 1035
rect 3665 967 3721 1001
rect 3665 933 3676 967
rect 3710 933 3721 967
rect 3665 899 3721 933
rect 3665 865 3676 899
rect 3710 865 3721 899
rect 3665 831 3721 865
rect 3665 797 3676 831
rect 3710 797 3721 831
rect 3665 763 3721 797
rect 3665 729 3676 763
rect 3710 729 3721 763
rect 3665 651 3721 729
rect 3821 1239 3877 1251
rect 3821 1205 3832 1239
rect 3866 1205 3877 1239
rect 3821 1171 3877 1205
rect 3821 1137 3832 1171
rect 3866 1137 3877 1171
rect 3821 1103 3877 1137
rect 3821 1069 3832 1103
rect 3866 1069 3877 1103
rect 3821 1035 3877 1069
rect 3821 1001 3832 1035
rect 3866 1001 3877 1035
rect 3821 967 3877 1001
rect 3821 933 3832 967
rect 3866 933 3877 967
rect 3821 899 3877 933
rect 3821 865 3832 899
rect 3866 865 3877 899
rect 3821 831 3877 865
rect 3821 797 3832 831
rect 3866 797 3877 831
rect 3821 763 3877 797
rect 3821 729 3832 763
rect 3866 729 3877 763
rect 3821 651 3877 729
rect 3977 1239 4033 1251
rect 3977 1205 3988 1239
rect 4022 1205 4033 1239
rect 3977 1171 4033 1205
rect 3977 1137 3988 1171
rect 4022 1137 4033 1171
rect 3977 1103 4033 1137
rect 3977 1069 3988 1103
rect 4022 1069 4033 1103
rect 3977 1035 4033 1069
rect 3977 1001 3988 1035
rect 4022 1001 4033 1035
rect 3977 967 4033 1001
rect 3977 933 3988 967
rect 4022 933 4033 967
rect 3977 899 4033 933
rect 3977 865 3988 899
rect 4022 865 4033 899
rect 3977 831 4033 865
rect 3977 797 3988 831
rect 4022 797 4033 831
rect 3977 763 4033 797
rect 3977 729 3988 763
rect 4022 729 4033 763
rect 3977 651 4033 729
rect 4133 1239 4189 1251
rect 4133 1205 4144 1239
rect 4178 1205 4189 1239
rect 4133 1171 4189 1205
rect 4133 1137 4144 1171
rect 4178 1137 4189 1171
rect 4133 1103 4189 1137
rect 4133 1069 4144 1103
rect 4178 1069 4189 1103
rect 4133 1035 4189 1069
rect 4133 1001 4144 1035
rect 4178 1001 4189 1035
rect 4133 967 4189 1001
rect 4133 933 4144 967
rect 4178 933 4189 967
rect 4133 899 4189 933
rect 4133 865 4144 899
rect 4178 865 4189 899
rect 4133 831 4189 865
rect 4133 797 4144 831
rect 4178 797 4189 831
rect 4133 763 4189 797
rect 4133 729 4144 763
rect 4178 729 4189 763
rect 4133 651 4189 729
rect 4289 1239 4345 1251
rect 4289 1205 4300 1239
rect 4334 1205 4345 1239
rect 4289 1171 4345 1205
rect 4289 1137 4300 1171
rect 4334 1137 4345 1171
rect 4289 1103 4345 1137
rect 4289 1069 4300 1103
rect 4334 1069 4345 1103
rect 4289 1035 4345 1069
rect 4289 1001 4300 1035
rect 4334 1001 4345 1035
rect 4289 967 4345 1001
rect 4289 933 4300 967
rect 4334 933 4345 967
rect 4289 899 4345 933
rect 4289 865 4300 899
rect 4334 865 4345 899
rect 4289 831 4345 865
rect 4289 797 4300 831
rect 4334 797 4345 831
rect 4289 763 4345 797
rect 4289 729 4300 763
rect 4334 729 4345 763
rect 4289 651 4345 729
rect 4445 1239 4498 1251
rect 4445 1205 4456 1239
rect 4490 1205 4498 1239
rect 4445 1171 4498 1205
rect 4445 1137 4456 1171
rect 4490 1137 4498 1171
rect 4445 1103 4498 1137
rect 4445 1069 4456 1103
rect 4490 1069 4498 1103
rect 4445 1035 4498 1069
rect 4445 1001 4456 1035
rect 4490 1001 4498 1035
rect 4445 967 4498 1001
rect 4445 933 4456 967
rect 4490 933 4498 967
rect 4445 899 4498 933
rect 4445 865 4456 899
rect 4490 865 4498 899
rect 4445 831 4498 865
rect 4445 797 4456 831
rect 4490 797 4498 831
rect 4445 763 4498 797
rect 4445 729 4456 763
rect 4490 729 4498 763
rect 4445 651 4498 729
rect 4572 1239 4625 1251
rect 4572 1205 4580 1239
rect 4614 1205 4625 1239
rect 4572 1171 4625 1205
rect 4572 1137 4580 1171
rect 4614 1137 4625 1171
rect 4572 1103 4625 1137
rect 4572 1069 4580 1103
rect 4614 1069 4625 1103
rect 4572 1035 4625 1069
rect 4572 1001 4580 1035
rect 4614 1001 4625 1035
rect 4572 967 4625 1001
rect 4572 933 4580 967
rect 4614 933 4625 967
rect 4572 899 4625 933
rect 4572 865 4580 899
rect 4614 865 4625 899
rect 4572 831 4625 865
rect 4572 797 4580 831
rect 4614 797 4625 831
rect 4572 763 4625 797
rect 4572 729 4580 763
rect 4614 729 4625 763
rect 4572 651 4625 729
rect 4725 1239 4778 1251
rect 4725 1205 4736 1239
rect 4770 1205 4778 1239
rect 4725 1171 4778 1205
rect 4725 1137 4736 1171
rect 4770 1137 4778 1171
rect 4725 1103 4778 1137
rect 4725 1069 4736 1103
rect 4770 1069 4778 1103
rect 4725 1035 4778 1069
rect 4725 1001 4736 1035
rect 4770 1001 4778 1035
rect 4725 967 4778 1001
rect 4725 933 4736 967
rect 4770 933 4778 967
rect 4725 899 4778 933
rect 4725 865 4736 899
rect 4770 865 4778 899
rect 4725 831 4778 865
rect 4725 797 4736 831
rect 4770 797 4778 831
rect 4725 763 4778 797
rect 4725 729 4736 763
rect 4770 729 4778 763
rect 4725 651 4778 729
rect 5016 912 5069 924
rect 5016 878 5024 912
rect 5058 878 5069 912
rect 5016 844 5069 878
rect 5016 810 5024 844
rect 5058 810 5069 844
rect 5016 776 5069 810
rect 5016 742 5024 776
rect 5058 742 5069 776
rect 5016 724 5069 742
rect 5169 912 5225 924
rect 5169 878 5180 912
rect 5214 878 5225 912
rect 5169 844 5225 878
rect 5169 810 5180 844
rect 5214 810 5225 844
rect 5169 776 5225 810
rect 5169 742 5180 776
rect 5214 742 5225 776
rect 5169 724 5225 742
rect 5325 912 5378 924
rect 5325 878 5336 912
rect 5370 878 5378 912
rect 5325 844 5378 878
rect 5325 810 5336 844
rect 5370 810 5378 844
rect 5325 776 5378 810
rect 5325 742 5336 776
rect 5370 742 5378 776
rect 5325 724 5378 742
rect 5452 912 5505 924
rect 5452 878 5460 912
rect 5494 878 5505 912
rect 5452 844 5505 878
rect 5452 810 5460 844
rect 5494 810 5505 844
rect 5452 776 5505 810
rect 5452 742 5460 776
rect 5494 742 5505 776
rect 5452 724 5505 742
rect 5605 912 5658 924
rect 5605 878 5616 912
rect 5650 878 5658 912
rect 5605 844 5658 878
rect 5605 810 5616 844
rect 5650 810 5658 844
rect 5605 776 5658 810
rect 5605 742 5616 776
rect 5650 742 5658 776
rect 5605 724 5658 742
<< mvpdiff >>
rect 5817 954 5870 966
rect 5817 920 5825 954
rect 5859 920 5870 954
rect 5817 886 5870 920
rect 5817 852 5825 886
rect 5859 852 5870 886
rect 5817 818 5870 852
rect 5817 784 5825 818
rect 5859 784 5870 818
rect 5817 750 5870 784
rect 5817 716 5825 750
rect 5859 716 5870 750
rect 5817 666 5870 716
rect 5970 954 6026 966
rect 5970 920 5981 954
rect 6015 920 6026 954
rect 5970 886 6026 920
rect 5970 852 5981 886
rect 6015 852 6026 886
rect 5970 818 6026 852
rect 5970 784 5981 818
rect 6015 784 6026 818
rect 5970 750 6026 784
rect 5970 716 5981 750
rect 6015 716 6026 750
rect 5970 666 6026 716
rect 6126 954 6179 966
rect 6126 920 6137 954
rect 6171 920 6179 954
rect 6126 886 6179 920
rect 6126 852 6137 886
rect 6171 852 6179 886
rect 6257 928 6310 966
rect 6257 894 6265 928
rect 6299 894 6310 928
rect 6257 882 6310 894
rect 6510 928 6566 966
rect 6510 894 6521 928
rect 6555 894 6566 928
rect 6510 882 6566 894
rect 6766 928 6819 966
rect 6766 894 6777 928
rect 6811 894 6819 928
rect 6766 882 6819 894
rect 6126 818 6179 852
rect 6126 784 6137 818
rect 6171 784 6179 818
rect 6126 750 6179 784
rect 6126 716 6137 750
rect 6171 716 6179 750
rect 6126 666 6179 716
<< mvndiffc >>
rect 3520 1205 3554 1239
rect 3520 1137 3554 1171
rect 3520 1069 3554 1103
rect 3520 1001 3554 1035
rect 3520 933 3554 967
rect 3520 865 3554 899
rect 3520 797 3554 831
rect 3520 729 3554 763
rect 3676 1205 3710 1239
rect 3676 1137 3710 1171
rect 3676 1069 3710 1103
rect 3676 1001 3710 1035
rect 3676 933 3710 967
rect 3676 865 3710 899
rect 3676 797 3710 831
rect 3676 729 3710 763
rect 3832 1205 3866 1239
rect 3832 1137 3866 1171
rect 3832 1069 3866 1103
rect 3832 1001 3866 1035
rect 3832 933 3866 967
rect 3832 865 3866 899
rect 3832 797 3866 831
rect 3832 729 3866 763
rect 3988 1205 4022 1239
rect 3988 1137 4022 1171
rect 3988 1069 4022 1103
rect 3988 1001 4022 1035
rect 3988 933 4022 967
rect 3988 865 4022 899
rect 3988 797 4022 831
rect 3988 729 4022 763
rect 4144 1205 4178 1239
rect 4144 1137 4178 1171
rect 4144 1069 4178 1103
rect 4144 1001 4178 1035
rect 4144 933 4178 967
rect 4144 865 4178 899
rect 4144 797 4178 831
rect 4144 729 4178 763
rect 4300 1205 4334 1239
rect 4300 1137 4334 1171
rect 4300 1069 4334 1103
rect 4300 1001 4334 1035
rect 4300 933 4334 967
rect 4300 865 4334 899
rect 4300 797 4334 831
rect 4300 729 4334 763
rect 4456 1205 4490 1239
rect 4456 1137 4490 1171
rect 4456 1069 4490 1103
rect 4456 1001 4490 1035
rect 4456 933 4490 967
rect 4456 865 4490 899
rect 4456 797 4490 831
rect 4456 729 4490 763
rect 4580 1205 4614 1239
rect 4580 1137 4614 1171
rect 4580 1069 4614 1103
rect 4580 1001 4614 1035
rect 4580 933 4614 967
rect 4580 865 4614 899
rect 4580 797 4614 831
rect 4580 729 4614 763
rect 4736 1205 4770 1239
rect 4736 1137 4770 1171
rect 4736 1069 4770 1103
rect 4736 1001 4770 1035
rect 4736 933 4770 967
rect 4736 865 4770 899
rect 4736 797 4770 831
rect 4736 729 4770 763
rect 5024 878 5058 912
rect 5024 810 5058 844
rect 5024 742 5058 776
rect 5180 878 5214 912
rect 5180 810 5214 844
rect 5180 742 5214 776
rect 5336 878 5370 912
rect 5336 810 5370 844
rect 5336 742 5370 776
rect 5460 878 5494 912
rect 5460 810 5494 844
rect 5460 742 5494 776
rect 5616 878 5650 912
rect 5616 810 5650 844
rect 5616 742 5650 776
<< mvpdiffc >>
rect 5825 920 5859 954
rect 5825 852 5859 886
rect 5825 784 5859 818
rect 5825 716 5859 750
rect 5981 920 6015 954
rect 5981 852 6015 886
rect 5981 784 6015 818
rect 5981 716 6015 750
rect 6137 920 6171 954
rect 6137 852 6171 886
rect 6265 894 6299 928
rect 6521 894 6555 928
rect 6777 894 6811 928
rect 6137 784 6171 818
rect 6137 716 6171 750
<< psubdiff >>
rect 3557 1355 3581 1389
rect 3615 1355 3653 1389
rect 3687 1355 3724 1389
rect 3758 1355 3795 1389
rect 3829 1355 3866 1389
rect 3900 1355 3937 1389
rect 3971 1355 4008 1389
rect 4042 1355 4079 1389
rect 4113 1355 4150 1389
rect 4184 1355 4221 1389
rect 4255 1355 4292 1389
rect 4326 1355 4363 1389
rect 4397 1355 4434 1389
rect 4468 1355 4505 1389
rect 4539 1355 4576 1389
rect 4610 1355 4647 1389
rect 4681 1355 4718 1389
rect 4752 1355 4776 1389
<< mvnsubdiff >>
rect 5817 1040 5841 1074
rect 5875 1040 5912 1074
rect 5946 1040 5983 1074
rect 6017 1040 6054 1074
rect 6088 1040 6125 1074
rect 6159 1040 6196 1074
rect 6230 1040 6267 1074
rect 6301 1040 6338 1074
rect 6372 1040 6409 1074
rect 6443 1040 6480 1074
rect 6514 1040 6551 1074
rect 6585 1040 6621 1074
rect 6655 1040 6691 1074
rect 6725 1040 6761 1074
rect 6795 1040 6819 1074
<< psubdiffcont >>
rect 3581 1355 3615 1389
rect 3653 1355 3687 1389
rect 3724 1355 3758 1389
rect 3795 1355 3829 1389
rect 3866 1355 3900 1389
rect 3937 1355 3971 1389
rect 4008 1355 4042 1389
rect 4079 1355 4113 1389
rect 4150 1355 4184 1389
rect 4221 1355 4255 1389
rect 4292 1355 4326 1389
rect 4363 1355 4397 1389
rect 4434 1355 4468 1389
rect 4505 1355 4539 1389
rect 4576 1355 4610 1389
rect 4647 1355 4681 1389
rect 4718 1355 4752 1389
<< mvnsubdiffcont >>
rect 5841 1040 5875 1074
rect 5912 1040 5946 1074
rect 5983 1040 6017 1074
rect 6054 1040 6088 1074
rect 6125 1040 6159 1074
rect 6196 1040 6230 1074
rect 6267 1040 6301 1074
rect 6338 1040 6372 1074
rect 6409 1040 6443 1074
rect 6480 1040 6514 1074
rect 6551 1040 6585 1074
rect 6621 1040 6655 1074
rect 6691 1040 6725 1074
rect 6761 1040 6795 1074
<< poly >>
rect 3565 1251 3665 1277
rect 3721 1251 3821 1277
rect 3877 1251 3977 1277
rect 4033 1251 4133 1277
rect 4189 1251 4289 1277
rect 4345 1251 4445 1277
rect 4625 1251 4725 1277
rect 5870 966 5970 998
rect 6026 966 6126 998
rect 6310 966 6510 998
rect 6566 966 6766 998
rect 5069 924 5169 950
rect 5225 924 5325 950
rect 5505 924 5605 950
rect 5069 692 5169 724
rect 5035 676 5169 692
rect 3565 625 3665 651
rect 3721 625 3821 651
rect 3877 625 3977 651
rect 3565 609 3977 625
rect 3565 575 3581 609
rect 3615 575 3651 609
rect 3685 575 3720 609
rect 3754 575 3789 609
rect 3823 575 3858 609
rect 3892 575 3927 609
rect 3961 575 3977 609
rect 3565 559 3977 575
rect 4033 625 4133 651
rect 4189 625 4289 651
rect 4345 625 4445 651
rect 4625 625 4725 651
rect 5035 642 5051 676
rect 5085 642 5119 676
rect 5153 642 5169 676
rect 5035 626 5169 642
rect 5225 692 5325 724
rect 5505 698 5605 724
rect 5225 676 5359 692
rect 5225 642 5241 676
rect 5275 642 5309 676
rect 5343 642 5359 676
rect 5225 626 5359 642
rect 5493 682 5627 698
rect 5493 648 5509 682
rect 5543 648 5577 682
rect 5611 648 5627 682
rect 6310 834 6510 882
rect 6310 800 6326 834
rect 6360 800 6460 834
rect 6494 800 6510 834
rect 6310 784 6510 800
rect 6566 834 6766 882
rect 6566 800 6582 834
rect 6616 800 6716 834
rect 6750 800 6766 834
rect 6566 784 6766 800
rect 5493 632 5627 648
rect 5870 634 5970 666
rect 6026 634 6126 666
rect 4033 609 4445 625
rect 4033 575 4049 609
rect 4083 575 4118 609
rect 4152 575 4187 609
rect 4221 575 4256 609
rect 4290 575 4325 609
rect 4359 575 4395 609
rect 4429 575 4445 609
rect 4033 559 4445 575
rect 4607 609 4749 625
rect 4607 575 4623 609
rect 4657 575 4699 609
rect 4733 575 4749 609
rect 4607 559 4749 575
rect 5837 618 5971 634
rect 5837 584 5853 618
rect 5887 584 5921 618
rect 5955 584 5971 618
rect 5837 568 5971 584
rect 6026 618 6160 634
rect 6026 584 6042 618
rect 6076 584 6110 618
rect 6144 584 6160 618
rect 6026 568 6160 584
<< polycont >>
rect 3581 575 3615 609
rect 3651 575 3685 609
rect 3720 575 3754 609
rect 3789 575 3823 609
rect 3858 575 3892 609
rect 3927 575 3961 609
rect 5051 642 5085 676
rect 5119 642 5153 676
rect 5241 642 5275 676
rect 5309 642 5343 676
rect 5509 648 5543 682
rect 5577 648 5611 682
rect 6326 800 6360 834
rect 6460 800 6494 834
rect 6582 800 6616 834
rect 6716 800 6750 834
rect 4049 575 4083 609
rect 4118 575 4152 609
rect 4187 575 4221 609
rect 4256 575 4290 609
rect 4325 575 4359 609
rect 4395 575 4429 609
rect 4623 575 4657 609
rect 4699 575 4733 609
rect 5853 584 5887 618
rect 5921 584 5955 618
rect 6042 584 6076 618
rect 6110 584 6144 618
<< locali >>
rect 3591 1389 3631 1420
rect 3665 1389 3705 1420
rect 3739 1389 3779 1420
rect 3813 1389 3853 1420
rect 3887 1389 3927 1420
rect 3961 1389 4001 1420
rect 4035 1389 4075 1420
rect 4109 1389 4149 1420
rect 4183 1389 4223 1420
rect 4257 1389 4297 1420
rect 4331 1389 4371 1420
rect 4405 1389 4445 1420
rect 4479 1389 4519 1420
rect 4553 1389 4593 1420
rect 4627 1389 4667 1420
rect 4701 1389 4742 1420
rect 3615 1386 3631 1389
rect 3687 1386 3705 1389
rect 3758 1386 3779 1389
rect 3829 1386 3853 1389
rect 3900 1386 3927 1389
rect 3971 1386 4001 1389
rect 4042 1386 4075 1389
rect 4113 1386 4149 1389
rect 3557 1355 3581 1386
rect 3615 1355 3653 1386
rect 3687 1355 3724 1386
rect 3758 1355 3795 1386
rect 3829 1355 3866 1386
rect 3900 1355 3937 1386
rect 3971 1355 4008 1386
rect 4042 1355 4079 1386
rect 4113 1355 4150 1386
rect 4184 1355 4221 1389
rect 4257 1386 4292 1389
rect 4331 1386 4363 1389
rect 4405 1386 4434 1389
rect 4479 1386 4505 1389
rect 4553 1386 4576 1389
rect 4627 1386 4647 1389
rect 4701 1386 4718 1389
rect 4255 1355 4292 1386
rect 4326 1355 4363 1386
rect 4397 1355 4434 1386
rect 4468 1355 4505 1386
rect 4539 1355 4576 1386
rect 4610 1355 4647 1386
rect 4681 1355 4718 1386
rect 4752 1355 4776 1386
rect 3520 1239 3554 1255
rect 3520 1171 3554 1205
rect 3520 1103 3554 1137
rect 3520 1035 3554 1069
rect 3520 967 3554 1001
rect 3520 899 3554 933
rect 3676 1239 3710 1255
rect 3676 1171 3710 1205
rect 3676 1103 3710 1137
rect 3676 1035 3710 1069
rect 3676 967 3710 1001
rect 3676 928 3710 933
rect 3832 1239 3866 1255
rect 3832 1171 3866 1205
rect 3832 1103 3866 1137
rect 3832 1035 3866 1069
rect 3832 967 3866 1001
rect 3675 899 3713 928
rect 3675 894 3676 899
rect 3520 831 3554 865
rect 3520 763 3554 797
rect 3710 894 3713 899
rect 3832 899 3866 933
rect 3988 1239 4022 1255
rect 3988 1171 4022 1205
rect 3988 1103 4022 1137
rect 3988 1035 4022 1069
rect 3988 967 4022 1001
rect 3988 928 4022 933
rect 4144 1239 4178 1255
rect 4144 1171 4178 1205
rect 4144 1103 4178 1137
rect 4144 1035 4178 1069
rect 4144 967 4178 1001
rect 3676 831 3710 865
rect 3676 763 3710 797
rect 3554 729 3576 745
rect 3538 711 3576 729
rect 3986 899 4024 928
rect 3986 894 3988 899
rect 3832 831 3866 865
rect 3832 763 3866 797
rect 4022 894 4024 899
rect 4144 899 4178 933
rect 4300 1239 4334 1255
rect 4300 1171 4334 1205
rect 4300 1103 4334 1137
rect 4300 1035 4334 1069
rect 4300 967 4334 1001
rect 4300 928 4334 933
rect 4456 1239 4490 1255
rect 4456 1171 4490 1205
rect 4456 1103 4490 1137
rect 4456 1035 4490 1069
rect 4456 967 4490 1001
rect 3988 831 4022 865
rect 4298 899 4336 928
rect 4298 894 4300 899
rect 4144 831 4178 865
rect 3988 763 4022 797
rect 4142 797 4144 821
rect 4334 894 4336 899
rect 4456 899 4490 933
rect 4300 831 4334 865
rect 4178 797 4180 821
rect 4142 787 4180 797
rect 4456 831 4490 865
rect 3676 713 3710 729
rect 3819 729 3832 745
rect 3819 711 3857 729
rect 3988 713 4022 729
rect 4144 763 4178 787
rect 4144 713 4178 729
rect 4300 763 4334 797
rect 4454 797 4456 821
rect 4580 1239 4614 1255
rect 4725 1251 4775 1355
rect 4580 1171 4614 1205
rect 4580 1103 4614 1137
rect 4580 1035 4614 1069
rect 4580 967 4614 1001
rect 4580 928 4614 933
rect 4736 1239 4770 1251
rect 4736 1171 4770 1205
rect 4736 1103 4770 1137
rect 4736 1035 4770 1069
rect 5817 1040 5829 1074
rect 5875 1040 5902 1074
rect 5946 1040 5975 1074
rect 6017 1040 6048 1074
rect 6088 1040 6121 1074
rect 6159 1040 6194 1074
rect 6230 1040 6267 1074
rect 6301 1040 6338 1074
rect 6374 1040 6409 1074
rect 6446 1040 6480 1074
rect 6518 1040 6551 1074
rect 6590 1040 6621 1074
rect 6662 1040 6691 1074
rect 6734 1040 6761 1074
rect 6806 1040 6819 1074
rect 4736 967 4770 980
rect 4614 894 4652 928
rect 5180 942 5214 980
rect 4736 899 4770 908
rect 4580 831 4614 865
rect 4490 797 4492 821
rect 4454 787 4492 797
rect 4300 713 4334 729
rect 4456 763 4490 787
rect 4456 713 4490 729
rect 4580 763 4614 797
rect 4580 713 4614 729
rect 4736 831 4770 865
rect 4736 763 4770 797
rect 5024 912 5058 928
rect 5024 844 5058 878
rect 5024 776 5058 810
rect 5460 942 5494 980
rect 5180 844 5214 878
rect 5180 776 5214 810
rect 4736 713 4770 729
rect 5006 742 5024 745
rect 5006 711 5044 742
rect 5336 912 5370 928
rect 5336 844 5370 878
rect 5336 776 5370 810
rect 5825 954 5859 970
rect 5616 920 5825 928
rect 5616 912 5859 920
rect 5650 910 5859 912
rect 5460 844 5494 878
rect 5460 776 5494 810
rect 5180 726 5214 742
rect 5370 742 5392 745
rect 5354 711 5392 742
rect 5460 726 5494 742
rect 5528 865 5540 899
rect 5574 865 5582 899
rect 5528 827 5582 865
rect 5528 793 5540 827
rect 5574 793 5582 827
rect 5528 682 5582 793
rect 5616 876 5648 878
rect 5682 876 5720 910
rect 5754 886 5859 910
rect 6014 962 6015 970
rect 5980 954 6015 962
rect 5980 924 5981 954
rect 6014 890 6015 920
rect 5754 876 5825 886
rect 5616 852 5825 876
rect 5616 844 5859 852
rect 5650 818 5859 844
rect 5650 810 5825 818
rect 5616 784 5825 810
rect 5616 776 5859 784
rect 5650 750 5859 776
rect 5650 742 5825 750
rect 5616 726 5825 742
rect 5825 700 5859 716
rect 5981 886 6015 890
rect 5981 818 6015 852
rect 5981 750 6015 784
rect 6137 954 6171 970
rect 6520 944 6554 960
rect 6137 886 6171 920
rect 6137 818 6171 852
rect 6137 750 6171 784
rect 5981 700 6015 716
rect 6098 711 6136 745
rect 6170 711 6171 716
rect 6137 700 6171 711
rect 6215 928 6299 944
rect 6215 894 6265 928
rect 6215 878 6299 894
rect 6520 928 6555 944
rect 6520 922 6521 928
rect 6554 888 6555 894
rect 6521 878 6555 888
rect 6777 928 6906 944
rect 6811 894 6906 928
rect 6777 878 6906 894
rect 6215 749 6272 878
rect 6310 800 6326 834
rect 6360 831 6460 834
rect 6494 831 6510 834
rect 6360 800 6391 831
rect 6425 800 6460 831
rect 6497 800 6510 831
rect 6566 800 6582 834
rect 6616 800 6716 834
rect 6750 800 6766 834
rect 6425 797 6463 800
rect 6566 749 6766 800
rect 6800 831 6906 878
rect 6834 797 6872 831
rect 5035 671 5051 676
rect 5085 671 5119 676
rect 5035 642 5046 671
rect 5085 642 5118 671
rect 5153 642 5169 676
rect 5225 651 5241 676
rect 5275 651 5309 676
rect 5080 637 5118 642
rect 5225 617 5232 651
rect 5275 642 5304 651
rect 5343 642 5359 676
rect 5266 617 5304 642
rect 5338 617 5359 642
rect 5493 648 5509 682
rect 5543 648 5577 682
rect 5611 648 5677 682
rect 6215 676 6766 749
rect 6215 666 6312 676
rect 5493 634 5677 648
rect 6026 651 6312 666
rect 5493 618 5972 634
rect 3565 575 3581 609
rect 3615 575 3651 609
rect 3685 575 3720 609
rect 3754 575 3789 609
rect 3823 575 3858 609
rect 3897 575 3927 609
rect 3969 575 3977 609
rect 4033 575 4049 609
rect 4083 575 4118 609
rect 4152 575 4187 609
rect 4221 575 4256 609
rect 4290 575 4325 609
rect 4364 575 4395 609
rect 4436 575 4445 609
rect 4607 575 4623 609
rect 4661 575 4699 609
rect 4733 575 4749 609
rect 5493 584 5853 618
rect 5887 584 5921 618
rect 5955 584 5972 618
rect 6026 617 6035 651
rect 6069 618 6107 651
rect 6141 618 6312 651
rect 6076 617 6107 618
rect 6026 584 6042 617
rect 6076 584 6110 617
rect 6144 584 6312 618
rect 5493 568 5972 584
<< viali >>
rect 3557 1389 3591 1420
rect 3631 1389 3665 1420
rect 3705 1389 3739 1420
rect 3779 1389 3813 1420
rect 3853 1389 3887 1420
rect 3927 1389 3961 1420
rect 4001 1389 4035 1420
rect 4075 1389 4109 1420
rect 4149 1389 4183 1420
rect 4223 1389 4257 1420
rect 4297 1389 4331 1420
rect 4371 1389 4405 1420
rect 4445 1389 4479 1420
rect 4519 1389 4553 1420
rect 4593 1389 4627 1420
rect 4667 1389 4701 1420
rect 4742 1389 4776 1420
rect 3557 1386 3581 1389
rect 3581 1386 3591 1389
rect 3631 1386 3653 1389
rect 3653 1386 3665 1389
rect 3705 1386 3724 1389
rect 3724 1386 3739 1389
rect 3779 1386 3795 1389
rect 3795 1386 3813 1389
rect 3853 1386 3866 1389
rect 3866 1386 3887 1389
rect 3927 1386 3937 1389
rect 3937 1386 3961 1389
rect 4001 1386 4008 1389
rect 4008 1386 4035 1389
rect 4075 1386 4079 1389
rect 4079 1386 4109 1389
rect 4149 1386 4150 1389
rect 4150 1386 4183 1389
rect 4223 1386 4255 1389
rect 4255 1386 4257 1389
rect 4297 1386 4326 1389
rect 4326 1386 4331 1389
rect 4371 1386 4397 1389
rect 4397 1386 4405 1389
rect 4445 1386 4468 1389
rect 4468 1386 4479 1389
rect 4519 1386 4539 1389
rect 4539 1386 4553 1389
rect 4593 1386 4610 1389
rect 4610 1386 4627 1389
rect 4667 1386 4681 1389
rect 4681 1386 4701 1389
rect 4742 1386 4752 1389
rect 4752 1386 4776 1389
rect 3641 894 3675 928
rect 3713 894 3747 928
rect 3504 729 3520 745
rect 3520 729 3538 745
rect 3504 711 3538 729
rect 3576 711 3610 745
rect 3952 894 3986 928
rect 4024 894 4058 928
rect 4264 894 4298 928
rect 4108 787 4142 821
rect 4336 894 4370 928
rect 4180 787 4214 821
rect 3785 711 3819 745
rect 3857 729 3866 745
rect 3866 729 3891 745
rect 3857 711 3891 729
rect 4420 787 4454 821
rect 5829 1040 5841 1074
rect 5841 1040 5863 1074
rect 5902 1040 5912 1074
rect 5912 1040 5936 1074
rect 5975 1040 5983 1074
rect 5983 1040 6009 1074
rect 6048 1040 6054 1074
rect 6054 1040 6082 1074
rect 6121 1040 6125 1074
rect 6125 1040 6155 1074
rect 6194 1040 6196 1074
rect 6196 1040 6228 1074
rect 6267 1040 6301 1074
rect 6340 1040 6372 1074
rect 6372 1040 6374 1074
rect 6412 1040 6443 1074
rect 6443 1040 6446 1074
rect 6484 1040 6514 1074
rect 6514 1040 6518 1074
rect 6556 1040 6585 1074
rect 6585 1040 6590 1074
rect 6628 1040 6655 1074
rect 6655 1040 6662 1074
rect 6700 1040 6725 1074
rect 6725 1040 6734 1074
rect 6772 1040 6795 1074
rect 6795 1040 6806 1074
rect 4736 1001 4770 1014
rect 4736 980 4770 1001
rect 4736 933 4770 942
rect 4580 899 4614 928
rect 4580 894 4614 899
rect 4652 894 4686 928
rect 4736 908 4770 933
rect 5180 980 5214 1014
rect 4492 787 4526 821
rect 5180 912 5214 942
rect 5460 980 5494 1014
rect 5180 908 5214 912
rect 4972 711 5006 745
rect 5044 742 5058 745
rect 5058 742 5078 745
rect 5044 711 5078 742
rect 5460 912 5494 942
rect 5460 908 5494 912
rect 5320 742 5336 745
rect 5336 742 5354 745
rect 5320 711 5354 742
rect 5392 711 5426 745
rect 5540 865 5574 899
rect 5540 793 5574 827
rect 5648 878 5650 910
rect 5650 878 5682 910
rect 5648 876 5682 878
rect 5720 876 5754 910
rect 5980 962 6014 996
rect 5980 920 5981 924
rect 5981 920 6014 924
rect 5980 890 6014 920
rect 6520 960 6554 994
rect 6064 711 6098 745
rect 6136 716 6137 745
rect 6137 716 6170 745
rect 6136 711 6170 716
rect 6520 894 6521 922
rect 6521 894 6554 922
rect 6520 888 6554 894
rect 6391 797 6425 831
rect 6463 800 6494 831
rect 6494 800 6497 831
rect 6463 797 6497 800
rect 6800 797 6834 831
rect 6872 797 6906 831
rect 5046 642 5051 671
rect 5051 642 5080 671
rect 5118 642 5119 671
rect 5119 642 5152 671
rect 5046 637 5080 642
rect 5118 637 5152 642
rect 5232 642 5241 651
rect 5241 642 5266 651
rect 5304 642 5309 651
rect 5309 642 5338 651
rect 5232 617 5266 642
rect 5304 617 5338 642
rect 3863 575 3892 609
rect 3892 575 3897 609
rect 3935 575 3961 609
rect 3961 575 3969 609
rect 4330 575 4359 609
rect 4359 575 4364 609
rect 4402 575 4429 609
rect 4429 575 4436 609
rect 4627 575 4657 609
rect 4657 575 4661 609
rect 4699 575 4733 609
rect 6035 618 6069 651
rect 6107 618 6141 651
rect 6035 617 6042 618
rect 6042 617 6069 618
rect 6107 617 6110 618
rect 6110 617 6141 618
<< metal1 >>
tri 4292 1426 4295 1429 se
rect 4295 1426 4301 1429
rect 3545 1420 4301 1426
rect 3545 1386 3557 1420
rect 3591 1386 3631 1420
rect 3665 1386 3705 1420
rect 3739 1386 3779 1420
rect 3813 1386 3853 1420
rect 3887 1386 3927 1420
rect 3961 1386 4001 1420
rect 4035 1386 4075 1420
rect 4109 1386 4149 1420
rect 4183 1386 4223 1420
rect 4257 1386 4297 1420
rect 3545 1380 4301 1386
tri 4292 1377 4295 1380 ne
rect 4295 1377 4301 1380
rect 4353 1377 4365 1429
rect 4417 1426 4423 1429
tri 4423 1426 4426 1429 sw
rect 4417 1420 4788 1426
rect 4417 1386 4445 1420
rect 4479 1386 4519 1420
rect 4553 1386 4593 1420
rect 4627 1386 4667 1420
rect 4701 1386 4742 1420
rect 4776 1386 4788 1420
rect 4417 1380 4788 1386
rect 4417 1377 4423 1380
tri 4423 1377 4426 1380 nw
rect 5817 1074 6818 1080
rect 5817 1040 5829 1074
rect 5863 1040 5902 1074
rect 5936 1040 5975 1074
rect 6009 1040 6048 1074
rect 6082 1040 6121 1074
rect 6155 1040 6194 1074
rect 6228 1040 6267 1074
rect 6301 1040 6340 1074
rect 6374 1040 6412 1074
rect 6446 1040 6484 1074
rect 6518 1040 6556 1074
rect 6590 1040 6628 1074
rect 6662 1040 6700 1074
rect 6734 1040 6772 1074
rect 6806 1040 6818 1074
rect 4730 1014 5500 1026
rect 4730 980 4736 1014
rect 4770 980 5180 1014
rect 5214 980 5460 1014
rect 5494 980 5500 1014
rect 4730 942 5500 980
rect 5817 996 6818 1040
rect 5817 970 5980 996
rect 3629 928 4698 934
rect 3629 894 3641 928
rect 3675 894 3713 928
rect 3747 894 3952 928
rect 3986 894 4024 928
rect 4058 894 4264 928
rect 4298 894 4336 928
rect 4370 894 4580 928
rect 4614 894 4652 928
rect 4686 894 4698 928
rect 4730 908 4736 942
rect 4770 908 5180 942
rect 5214 908 5460 942
rect 5494 908 5500 942
rect 5974 962 5980 970
rect 6014 994 6818 996
rect 6014 970 6520 994
rect 6014 962 6020 970
rect 5974 924 6020 962
rect 4730 896 5500 908
rect 5534 899 5580 911
rect 3629 888 4698 894
rect 5534 865 5540 899
rect 5574 865 5580 899
rect 5636 910 5766 916
rect 5636 876 5648 910
rect 5682 876 5720 910
rect 5754 876 5766 910
rect 5974 890 5980 924
rect 6014 890 6020 924
rect 5974 878 6020 890
rect 6514 960 6520 970
rect 6554 970 6818 994
rect 6554 960 6560 970
rect 6514 922 6560 960
rect 6514 888 6520 922
rect 6554 888 6560 922
rect 6514 876 6560 888
rect 5636 870 5766 876
rect 5534 837 5580 865
rect 5534 831 6918 837
rect 5534 827 6391 831
rect 4096 821 5540 827
rect 4096 787 4108 821
rect 4142 787 4180 821
rect 4214 787 4420 821
rect 4454 787 4492 821
rect 4526 793 5540 821
rect 5574 797 6391 827
rect 6425 797 6463 831
rect 6497 797 6800 831
rect 6834 797 6872 831
rect 6906 797 6918 831
rect 5574 793 6918 797
rect 4526 791 6918 793
rect 4526 787 5580 791
rect 4096 781 5580 787
rect 3492 745 5266 751
rect 3492 711 3504 745
rect 3538 711 3576 745
rect 3610 711 3785 745
rect 3819 711 3857 745
rect 3891 711 4972 745
rect 5006 711 5044 745
rect 5078 711 5266 745
rect 3492 705 5266 711
rect 5308 745 6182 751
rect 5308 711 5320 745
rect 5354 711 5392 745
rect 5426 711 6064 745
rect 6098 711 6136 745
rect 6170 711 6182 745
rect 5308 705 6182 711
rect 5034 671 5164 677
rect 5034 637 5046 671
rect 5080 637 5118 671
rect 5152 637 5164 671
rect 5034 631 5164 637
rect 5220 657 5266 705
rect 5220 651 6153 657
rect 5220 617 5232 651
rect 5266 617 5304 651
rect 5338 617 6035 651
rect 6069 617 6107 651
rect 6141 617 6153 651
rect 3851 609 3981 615
rect 3851 575 3863 609
rect 3897 575 3935 609
rect 3969 575 3981 609
rect 3851 569 3981 575
rect 4318 609 4448 615
rect 4318 575 4330 609
rect 4364 575 4402 609
rect 4436 575 4448 609
rect 4318 569 4448 575
rect 4615 609 4745 615
rect 5220 611 6153 617
rect 4615 575 4627 609
rect 4661 575 4699 609
rect 4733 575 4745 609
rect 4615 569 4745 575
<< via1 >>
rect 4301 1420 4353 1429
rect 4301 1386 4331 1420
rect 4331 1386 4353 1420
rect 4301 1377 4353 1386
rect 4365 1420 4417 1429
rect 4365 1386 4371 1420
rect 4371 1386 4405 1420
rect 4405 1386 4417 1420
rect 4365 1377 4417 1386
<< metal2 >>
rect 4295 1377 4301 1429
rect 4353 1377 4365 1429
rect 4417 1377 4423 1429
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_0
timestamp 1644511149
transform -1 0 3977 0 -1 1251
box -28 0 440 267
use sky130_fd_pr__nfet_01v8__example_55959141808569  sky130_fd_pr__nfet_01v8__example_55959141808569_1
timestamp 1644511149
transform 1 0 4033 0 -1 1251
box -28 0 440 267
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_0
timestamp 1644511149
transform -1 0 5169 0 -1 924
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_1
timestamp 1644511149
transform 1 0 5505 0 -1 924
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808570  sky130_fd_pr__nfet_01v8__example_55959141808570_2
timestamp 1644511149
transform 1 0 5225 0 -1 924
box -28 0 128 97
use sky130_fd_pr__nfet_01v8__example_55959141808589  sky130_fd_pr__nfet_01v8__example_55959141808589_0
timestamp 1644511149
transform -1 0 4725 0 -1 1251
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808475  sky130_fd_pr__pfet_01v8__example_55959141808475_0
timestamp 1644511149
transform -1 0 5970 0 -1 966
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808475  sky130_fd_pr__pfet_01v8__example_55959141808475_1
timestamp 1644511149
transform 1 0 6026 0 -1 966
box -28 0 128 131
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_0
timestamp 1644511149
transform 1 0 6566 0 1 882
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808477  sky130_fd_pr__pfet_01v8__example_55959141808477_1
timestamp 1644511149
transform -1 0 6510 0 1 882
box -28 0 228 29
<< labels >>
flabel metal1 s 3928 577 3956 605 3 FreeSans 520 180 0 0 IN_B
port 1 nsew
flabel metal1 s 4355 578 4383 606 3 FreeSans 520 0 0 0 IN
port 2 nsew
flabel metal1 s 5105 642 5133 670 3 FreeSans 520 0 0 0 RST_H
port 3 nsew
flabel metal1 s 5339 716 5367 744 3 FreeSans 520 0 0 0 OUT_H_N
port 4 nsew
flabel metal1 s 5687 880 5715 908 3 FreeSans 520 90 0 0 OUT_H
port 5 nsew
flabel metal1 s 5979 1001 6007 1029 3 FreeSans 520 0 0 0 VPWR_HV
port 6 nsew
flabel metal1 s 4661 576 4689 604 3 FreeSans 520 0 0 0 HLD_H
port 7 nsew
flabel metal1 s 5261 949 5289 977 3 FreeSans 520 0 0 0 VGND
port 8 nsew
<< properties >>
string GDS_END 8409684
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8390554
<< end >>
