magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 8 157 283 203
rect 637 157 827 203
rect 8 67 827 157
rect 29 -17 63 67
rect 285 21 827 67
<< locali >>
rect 85 199 155 339
rect 189 199 247 265
rect 496 425 624 491
rect 756 299 811 493
rect 523 199 654 265
rect 777 152 811 299
rect 756 83 811 152
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 17 407 69 491
rect 103 441 169 527
rect 302 441 451 475
rect 17 373 383 407
rect 17 165 51 373
rect 198 305 315 339
rect 281 249 315 305
rect 349 317 383 373
rect 417 391 451 441
rect 417 357 624 391
rect 658 367 714 527
rect 590 333 624 357
rect 349 283 479 317
rect 590 299 722 333
rect 281 215 366 249
rect 281 165 315 215
rect 445 199 479 283
rect 688 265 722 299
rect 688 199 743 265
rect 688 165 722 199
rect 17 90 80 165
rect 131 17 165 165
rect 215 131 315 165
rect 403 131 722 165
rect 215 90 249 131
rect 294 17 369 97
rect 403 61 437 131
rect 474 17 540 97
rect 574 61 608 131
rect 642 17 718 97
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
rlabel locali s 523 199 654 265 6 A
port 1 nsew signal input
rlabel locali s 496 425 624 491 6 B
port 2 nsew signal input
rlabel locali s 85 199 155 339 6 C_N
port 3 nsew signal input
rlabel locali s 189 199 247 265 6 D_N
port 4 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 285 21 827 67 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 29 -17 63 67 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 8 67 827 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 637 157 827 203 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 8 157 283 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 756 83 811 152 6 X
port 9 nsew signal output
rlabel locali s 777 152 811 299 6 X
port 9 nsew signal output
rlabel locali s 756 299 811 493 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1106760
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1099712
<< end >>
