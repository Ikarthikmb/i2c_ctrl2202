magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< dnwell >>
rect 26 30 11991 1672
<< nwell >>
rect -54 1466 12071 1753
rect -54 236 232 1466
rect 1839 236 2075 1466
rect 6817 236 7053 1466
rect 11835 236 12071 1466
rect -54 -50 12071 236
rect 6350 -2111 8843 -1087
<< pwell >>
rect 331 296 1735 1380
rect 2166 296 6746 1406
rect 7170 296 11744 1406
<< mvnmos >>
rect 558 1087 1558 1187
rect 558 931 1558 1031
rect 558 645 1558 745
rect 558 489 1558 589
rect 2393 1113 4393 1213
rect 4499 1113 6499 1213
rect 2393 957 4393 1057
rect 4499 957 6499 1057
rect 2393 801 4393 901
rect 4499 801 6499 901
rect 2393 645 4393 745
rect 4499 645 6499 745
rect 2393 489 4393 589
rect 4499 489 6499 589
rect 7412 1113 9412 1213
rect 9518 1113 11518 1213
rect 7412 957 9412 1057
rect 9518 957 11518 1057
rect 7412 801 9412 901
rect 9518 801 11518 901
rect 7412 645 9412 745
rect 9518 645 11518 745
rect 7412 489 9412 589
rect 9518 489 11518 589
<< mvpmos >>
rect 6616 -1415 8616 -1315
rect 6616 -1571 8616 -1471
rect 6616 -1727 8616 -1627
rect 6616 -1883 8616 -1783
<< mvndiff >>
rect 558 1232 1558 1240
rect 558 1198 570 1232
rect 604 1198 638 1232
rect 672 1198 706 1232
rect 740 1198 774 1232
rect 808 1198 842 1232
rect 876 1198 910 1232
rect 944 1198 978 1232
rect 1012 1198 1046 1232
rect 1080 1198 1114 1232
rect 1148 1198 1182 1232
rect 1216 1198 1250 1232
rect 1284 1198 1318 1232
rect 1352 1198 1386 1232
rect 1420 1198 1454 1232
rect 1488 1198 1558 1232
rect 558 1187 1558 1198
rect 558 1076 1558 1087
rect 558 1042 570 1076
rect 604 1042 638 1076
rect 672 1042 706 1076
rect 740 1042 774 1076
rect 808 1042 842 1076
rect 876 1042 910 1076
rect 944 1042 978 1076
rect 1012 1042 1046 1076
rect 1080 1042 1114 1076
rect 1148 1042 1182 1076
rect 1216 1042 1250 1076
rect 1284 1042 1318 1076
rect 1352 1042 1386 1076
rect 1420 1042 1454 1076
rect 1488 1042 1558 1076
rect 558 1031 1558 1042
rect 558 920 1558 931
rect 558 886 570 920
rect 604 886 638 920
rect 672 886 706 920
rect 740 886 774 920
rect 808 886 842 920
rect 876 886 910 920
rect 944 886 978 920
rect 1012 886 1046 920
rect 1080 886 1114 920
rect 1148 886 1182 920
rect 1216 886 1250 920
rect 1284 886 1318 920
rect 1352 886 1386 920
rect 1420 886 1454 920
rect 1488 886 1558 920
rect 558 878 1558 886
rect 558 790 1558 798
rect 558 756 570 790
rect 604 756 638 790
rect 672 756 706 790
rect 740 756 774 790
rect 808 756 842 790
rect 876 756 910 790
rect 944 756 978 790
rect 1012 756 1046 790
rect 1080 756 1114 790
rect 1148 756 1182 790
rect 1216 756 1250 790
rect 1284 756 1318 790
rect 1352 756 1386 790
rect 1420 756 1454 790
rect 1488 756 1558 790
rect 558 745 1558 756
rect 558 634 1558 645
rect 558 600 570 634
rect 604 600 638 634
rect 672 600 706 634
rect 740 600 774 634
rect 808 600 842 634
rect 876 600 910 634
rect 944 600 978 634
rect 1012 600 1046 634
rect 1080 600 1114 634
rect 1148 600 1182 634
rect 1216 600 1250 634
rect 1284 600 1318 634
rect 1352 600 1386 634
rect 1420 600 1454 634
rect 1488 600 1558 634
rect 558 589 1558 600
rect 558 478 1558 489
rect 558 444 570 478
rect 604 444 638 478
rect 672 444 706 478
rect 740 444 774 478
rect 808 444 842 478
rect 876 444 910 478
rect 944 444 978 478
rect 1012 444 1046 478
rect 1080 444 1114 478
rect 1148 444 1182 478
rect 1216 444 1250 478
rect 1284 444 1318 478
rect 1352 444 1386 478
rect 1420 444 1454 478
rect 1488 444 1558 478
rect 558 436 1558 444
rect 2393 1258 4393 1266
rect 2393 1224 2405 1258
rect 2439 1224 2473 1258
rect 2507 1224 2541 1258
rect 2575 1224 2609 1258
rect 2643 1224 2677 1258
rect 2711 1224 2745 1258
rect 2779 1224 2813 1258
rect 2847 1224 2881 1258
rect 2915 1224 2949 1258
rect 2983 1224 3017 1258
rect 3051 1224 3085 1258
rect 3119 1224 3153 1258
rect 3187 1224 3221 1258
rect 3255 1224 3289 1258
rect 3323 1224 3357 1258
rect 3391 1224 3425 1258
rect 3459 1224 3493 1258
rect 3527 1224 3561 1258
rect 3595 1224 3629 1258
rect 3663 1224 3697 1258
rect 3731 1224 3765 1258
rect 3799 1224 3833 1258
rect 3867 1224 3901 1258
rect 3935 1224 3969 1258
rect 4003 1224 4037 1258
rect 4071 1224 4105 1258
rect 4139 1224 4173 1258
rect 4207 1224 4241 1258
rect 4275 1224 4309 1258
rect 4343 1224 4393 1258
rect 2393 1213 4393 1224
rect 4499 1258 6499 1266
rect 4499 1224 4549 1258
rect 4583 1224 4617 1258
rect 4651 1224 4685 1258
rect 4719 1224 4753 1258
rect 4787 1224 4821 1258
rect 4855 1224 4889 1258
rect 4923 1224 4957 1258
rect 4991 1224 5025 1258
rect 5059 1224 5093 1258
rect 5127 1224 5161 1258
rect 5195 1224 5229 1258
rect 5263 1224 5297 1258
rect 5331 1224 5365 1258
rect 5399 1224 5433 1258
rect 5467 1224 5501 1258
rect 5535 1224 5569 1258
rect 5603 1224 5637 1258
rect 5671 1224 5705 1258
rect 5739 1224 5773 1258
rect 5807 1224 5841 1258
rect 5875 1224 5909 1258
rect 5943 1224 5977 1258
rect 6011 1224 6045 1258
rect 6079 1224 6113 1258
rect 6147 1224 6181 1258
rect 6215 1224 6249 1258
rect 6283 1224 6317 1258
rect 6351 1224 6385 1258
rect 6419 1224 6453 1258
rect 6487 1224 6499 1258
rect 4499 1213 6499 1224
rect 2393 1102 4393 1113
rect 2393 1068 2405 1102
rect 2439 1068 2473 1102
rect 2507 1068 2541 1102
rect 2575 1068 2609 1102
rect 2643 1068 2677 1102
rect 2711 1068 2745 1102
rect 2779 1068 2813 1102
rect 2847 1068 2881 1102
rect 2915 1068 2949 1102
rect 2983 1068 3017 1102
rect 3051 1068 3085 1102
rect 3119 1068 3153 1102
rect 3187 1068 3221 1102
rect 3255 1068 3289 1102
rect 3323 1068 3357 1102
rect 3391 1068 3425 1102
rect 3459 1068 3493 1102
rect 3527 1068 3561 1102
rect 3595 1068 3629 1102
rect 3663 1068 3697 1102
rect 3731 1068 3765 1102
rect 3799 1068 3833 1102
rect 3867 1068 3901 1102
rect 3935 1068 3969 1102
rect 4003 1068 4037 1102
rect 4071 1068 4105 1102
rect 4139 1068 4173 1102
rect 4207 1068 4241 1102
rect 4275 1068 4309 1102
rect 4343 1068 4393 1102
rect 2393 1057 4393 1068
rect 4499 1102 6499 1113
rect 4499 1068 4549 1102
rect 4583 1068 4617 1102
rect 4651 1068 4685 1102
rect 4719 1068 4753 1102
rect 4787 1068 4821 1102
rect 4855 1068 4889 1102
rect 4923 1068 4957 1102
rect 4991 1068 5025 1102
rect 5059 1068 5093 1102
rect 5127 1068 5161 1102
rect 5195 1068 5229 1102
rect 5263 1068 5297 1102
rect 5331 1068 5365 1102
rect 5399 1068 5433 1102
rect 5467 1068 5501 1102
rect 5535 1068 5569 1102
rect 5603 1068 5637 1102
rect 5671 1068 5705 1102
rect 5739 1068 5773 1102
rect 5807 1068 5841 1102
rect 5875 1068 5909 1102
rect 5943 1068 5977 1102
rect 6011 1068 6045 1102
rect 6079 1068 6113 1102
rect 6147 1068 6181 1102
rect 6215 1068 6249 1102
rect 6283 1068 6317 1102
rect 6351 1068 6385 1102
rect 6419 1068 6453 1102
rect 6487 1068 6499 1102
rect 4499 1057 6499 1068
rect 2393 946 4393 957
rect 2393 912 2405 946
rect 2439 912 2473 946
rect 2507 912 2541 946
rect 2575 912 2609 946
rect 2643 912 2677 946
rect 2711 912 2745 946
rect 2779 912 2813 946
rect 2847 912 2881 946
rect 2915 912 2949 946
rect 2983 912 3017 946
rect 3051 912 3085 946
rect 3119 912 3153 946
rect 3187 912 3221 946
rect 3255 912 3289 946
rect 3323 912 3357 946
rect 3391 912 3425 946
rect 3459 912 3493 946
rect 3527 912 3561 946
rect 3595 912 3629 946
rect 3663 912 3697 946
rect 3731 912 3765 946
rect 3799 912 3833 946
rect 3867 912 3901 946
rect 3935 912 3969 946
rect 4003 912 4037 946
rect 4071 912 4105 946
rect 4139 912 4173 946
rect 4207 912 4241 946
rect 4275 912 4309 946
rect 4343 912 4393 946
rect 2393 901 4393 912
rect 4499 946 6499 957
rect 4499 912 4549 946
rect 4583 912 4617 946
rect 4651 912 4685 946
rect 4719 912 4753 946
rect 4787 912 4821 946
rect 4855 912 4889 946
rect 4923 912 4957 946
rect 4991 912 5025 946
rect 5059 912 5093 946
rect 5127 912 5161 946
rect 5195 912 5229 946
rect 5263 912 5297 946
rect 5331 912 5365 946
rect 5399 912 5433 946
rect 5467 912 5501 946
rect 5535 912 5569 946
rect 5603 912 5637 946
rect 5671 912 5705 946
rect 5739 912 5773 946
rect 5807 912 5841 946
rect 5875 912 5909 946
rect 5943 912 5977 946
rect 6011 912 6045 946
rect 6079 912 6113 946
rect 6147 912 6181 946
rect 6215 912 6249 946
rect 6283 912 6317 946
rect 6351 912 6385 946
rect 6419 912 6453 946
rect 6487 912 6499 946
rect 4499 901 6499 912
rect 2393 790 4393 801
rect 2393 756 2405 790
rect 2439 756 2473 790
rect 2507 756 2541 790
rect 2575 756 2609 790
rect 2643 756 2677 790
rect 2711 756 2745 790
rect 2779 756 2813 790
rect 2847 756 2881 790
rect 2915 756 2949 790
rect 2983 756 3017 790
rect 3051 756 3085 790
rect 3119 756 3153 790
rect 3187 756 3221 790
rect 3255 756 3289 790
rect 3323 756 3357 790
rect 3391 756 3425 790
rect 3459 756 3493 790
rect 3527 756 3561 790
rect 3595 756 3629 790
rect 3663 756 3697 790
rect 3731 756 3765 790
rect 3799 756 3833 790
rect 3867 756 3901 790
rect 3935 756 3969 790
rect 4003 756 4037 790
rect 4071 756 4105 790
rect 4139 756 4173 790
rect 4207 756 4241 790
rect 4275 756 4309 790
rect 4343 756 4393 790
rect 2393 745 4393 756
rect 4499 790 6499 801
rect 4499 756 4549 790
rect 4583 756 4617 790
rect 4651 756 4685 790
rect 4719 756 4753 790
rect 4787 756 4821 790
rect 4855 756 4889 790
rect 4923 756 4957 790
rect 4991 756 5025 790
rect 5059 756 5093 790
rect 5127 756 5161 790
rect 5195 756 5229 790
rect 5263 756 5297 790
rect 5331 756 5365 790
rect 5399 756 5433 790
rect 5467 756 5501 790
rect 5535 756 5569 790
rect 5603 756 5637 790
rect 5671 756 5705 790
rect 5739 756 5773 790
rect 5807 756 5841 790
rect 5875 756 5909 790
rect 5943 756 5977 790
rect 6011 756 6045 790
rect 6079 756 6113 790
rect 6147 756 6181 790
rect 6215 756 6249 790
rect 6283 756 6317 790
rect 6351 756 6385 790
rect 6419 756 6453 790
rect 6487 756 6499 790
rect 4499 745 6499 756
rect 2393 634 4393 645
rect 2393 600 2405 634
rect 2439 600 2473 634
rect 2507 600 2541 634
rect 2575 600 2609 634
rect 2643 600 2677 634
rect 2711 600 2745 634
rect 2779 600 2813 634
rect 2847 600 2881 634
rect 2915 600 2949 634
rect 2983 600 3017 634
rect 3051 600 3085 634
rect 3119 600 3153 634
rect 3187 600 3221 634
rect 3255 600 3289 634
rect 3323 600 3357 634
rect 3391 600 3425 634
rect 3459 600 3493 634
rect 3527 600 3561 634
rect 3595 600 3629 634
rect 3663 600 3697 634
rect 3731 600 3765 634
rect 3799 600 3833 634
rect 3867 600 3901 634
rect 3935 600 3969 634
rect 4003 600 4037 634
rect 4071 600 4105 634
rect 4139 600 4173 634
rect 4207 600 4241 634
rect 4275 600 4309 634
rect 4343 600 4393 634
rect 2393 589 4393 600
rect 4499 634 6499 645
rect 4499 600 4549 634
rect 4583 600 4617 634
rect 4651 600 4685 634
rect 4719 600 4753 634
rect 4787 600 4821 634
rect 4855 600 4889 634
rect 4923 600 4957 634
rect 4991 600 5025 634
rect 5059 600 5093 634
rect 5127 600 5161 634
rect 5195 600 5229 634
rect 5263 600 5297 634
rect 5331 600 5365 634
rect 5399 600 5433 634
rect 5467 600 5501 634
rect 5535 600 5569 634
rect 5603 600 5637 634
rect 5671 600 5705 634
rect 5739 600 5773 634
rect 5807 600 5841 634
rect 5875 600 5909 634
rect 5943 600 5977 634
rect 6011 600 6045 634
rect 6079 600 6113 634
rect 6147 600 6181 634
rect 6215 600 6249 634
rect 6283 600 6317 634
rect 6351 600 6385 634
rect 6419 600 6453 634
rect 6487 600 6499 634
rect 4499 589 6499 600
rect 2393 478 4393 489
rect 2393 444 2405 478
rect 2439 444 2473 478
rect 2507 444 2541 478
rect 2575 444 2609 478
rect 2643 444 2677 478
rect 2711 444 2745 478
rect 2779 444 2813 478
rect 2847 444 2881 478
rect 2915 444 2949 478
rect 2983 444 3017 478
rect 3051 444 3085 478
rect 3119 444 3153 478
rect 3187 444 3221 478
rect 3255 444 3289 478
rect 3323 444 3357 478
rect 3391 444 3425 478
rect 3459 444 3493 478
rect 3527 444 3561 478
rect 3595 444 3629 478
rect 3663 444 3697 478
rect 3731 444 3765 478
rect 3799 444 3833 478
rect 3867 444 3901 478
rect 3935 444 3969 478
rect 4003 444 4037 478
rect 4071 444 4105 478
rect 4139 444 4173 478
rect 4207 444 4241 478
rect 4275 444 4309 478
rect 4343 444 4393 478
rect 2393 436 4393 444
rect 4499 478 6499 489
rect 4499 444 4549 478
rect 4583 444 4617 478
rect 4651 444 4685 478
rect 4719 444 4753 478
rect 4787 444 4821 478
rect 4855 444 4889 478
rect 4923 444 4957 478
rect 4991 444 5025 478
rect 5059 444 5093 478
rect 5127 444 5161 478
rect 5195 444 5229 478
rect 5263 444 5297 478
rect 5331 444 5365 478
rect 5399 444 5433 478
rect 5467 444 5501 478
rect 5535 444 5569 478
rect 5603 444 5637 478
rect 5671 444 5705 478
rect 5739 444 5773 478
rect 5807 444 5841 478
rect 5875 444 5909 478
rect 5943 444 5977 478
rect 6011 444 6045 478
rect 6079 444 6113 478
rect 6147 444 6181 478
rect 6215 444 6249 478
rect 6283 444 6317 478
rect 6351 444 6385 478
rect 6419 444 6453 478
rect 6487 444 6499 478
rect 4499 436 6499 444
rect 7412 1258 9412 1266
rect 7412 1224 7462 1258
rect 7496 1224 7530 1258
rect 7564 1224 7598 1258
rect 7632 1224 7666 1258
rect 7700 1224 7734 1258
rect 7768 1224 7802 1258
rect 7836 1224 7870 1258
rect 7904 1224 7938 1258
rect 7972 1224 8006 1258
rect 8040 1224 8074 1258
rect 8108 1224 8142 1258
rect 8176 1224 8210 1258
rect 8244 1224 8278 1258
rect 8312 1224 8346 1258
rect 8380 1224 8414 1258
rect 8448 1224 8482 1258
rect 8516 1224 8550 1258
rect 8584 1224 8618 1258
rect 8652 1224 8686 1258
rect 8720 1224 8754 1258
rect 8788 1224 8822 1258
rect 8856 1224 8890 1258
rect 8924 1224 8958 1258
rect 8992 1224 9026 1258
rect 9060 1224 9094 1258
rect 9128 1224 9162 1258
rect 9196 1224 9230 1258
rect 9264 1224 9298 1258
rect 9332 1224 9366 1258
rect 9400 1224 9412 1258
rect 7412 1213 9412 1224
rect 9518 1258 11518 1266
rect 9518 1224 9568 1258
rect 9602 1224 9636 1258
rect 9670 1224 9704 1258
rect 9738 1224 9772 1258
rect 9806 1224 9840 1258
rect 9874 1224 9908 1258
rect 9942 1224 9976 1258
rect 10010 1224 10044 1258
rect 10078 1224 10112 1258
rect 10146 1224 10180 1258
rect 10214 1224 10248 1258
rect 10282 1224 10316 1258
rect 10350 1224 10384 1258
rect 10418 1224 10452 1258
rect 10486 1224 10520 1258
rect 10554 1224 10588 1258
rect 10622 1224 10656 1258
rect 10690 1224 10724 1258
rect 10758 1224 10792 1258
rect 10826 1224 10860 1258
rect 10894 1224 10928 1258
rect 10962 1224 10996 1258
rect 11030 1224 11064 1258
rect 11098 1224 11132 1258
rect 11166 1224 11200 1258
rect 11234 1224 11268 1258
rect 11302 1224 11336 1258
rect 11370 1224 11404 1258
rect 11438 1224 11472 1258
rect 11506 1224 11518 1258
rect 9518 1213 11518 1224
rect 7412 1102 9412 1113
rect 7412 1068 7462 1102
rect 7496 1068 7530 1102
rect 7564 1068 7598 1102
rect 7632 1068 7666 1102
rect 7700 1068 7734 1102
rect 7768 1068 7802 1102
rect 7836 1068 7870 1102
rect 7904 1068 7938 1102
rect 7972 1068 8006 1102
rect 8040 1068 8074 1102
rect 8108 1068 8142 1102
rect 8176 1068 8210 1102
rect 8244 1068 8278 1102
rect 8312 1068 8346 1102
rect 8380 1068 8414 1102
rect 8448 1068 8482 1102
rect 8516 1068 8550 1102
rect 8584 1068 8618 1102
rect 8652 1068 8686 1102
rect 8720 1068 8754 1102
rect 8788 1068 8822 1102
rect 8856 1068 8890 1102
rect 8924 1068 8958 1102
rect 8992 1068 9026 1102
rect 9060 1068 9094 1102
rect 9128 1068 9162 1102
rect 9196 1068 9230 1102
rect 9264 1068 9298 1102
rect 9332 1068 9366 1102
rect 9400 1068 9412 1102
rect 7412 1057 9412 1068
rect 9518 1102 11518 1113
rect 9518 1068 9568 1102
rect 9602 1068 9636 1102
rect 9670 1068 9704 1102
rect 9738 1068 9772 1102
rect 9806 1068 9840 1102
rect 9874 1068 9908 1102
rect 9942 1068 9976 1102
rect 10010 1068 10044 1102
rect 10078 1068 10112 1102
rect 10146 1068 10180 1102
rect 10214 1068 10248 1102
rect 10282 1068 10316 1102
rect 10350 1068 10384 1102
rect 10418 1068 10452 1102
rect 10486 1068 10520 1102
rect 10554 1068 10588 1102
rect 10622 1068 10656 1102
rect 10690 1068 10724 1102
rect 10758 1068 10792 1102
rect 10826 1068 10860 1102
rect 10894 1068 10928 1102
rect 10962 1068 10996 1102
rect 11030 1068 11064 1102
rect 11098 1068 11132 1102
rect 11166 1068 11200 1102
rect 11234 1068 11268 1102
rect 11302 1068 11336 1102
rect 11370 1068 11404 1102
rect 11438 1068 11472 1102
rect 11506 1068 11518 1102
rect 9518 1057 11518 1068
rect 7412 946 9412 957
rect 7412 912 7462 946
rect 7496 912 7530 946
rect 7564 912 7598 946
rect 7632 912 7666 946
rect 7700 912 7734 946
rect 7768 912 7802 946
rect 7836 912 7870 946
rect 7904 912 7938 946
rect 7972 912 8006 946
rect 8040 912 8074 946
rect 8108 912 8142 946
rect 8176 912 8210 946
rect 8244 912 8278 946
rect 8312 912 8346 946
rect 8380 912 8414 946
rect 8448 912 8482 946
rect 8516 912 8550 946
rect 8584 912 8618 946
rect 8652 912 8686 946
rect 8720 912 8754 946
rect 8788 912 8822 946
rect 8856 912 8890 946
rect 8924 912 8958 946
rect 8992 912 9026 946
rect 9060 912 9094 946
rect 9128 912 9162 946
rect 9196 912 9230 946
rect 9264 912 9298 946
rect 9332 912 9366 946
rect 9400 912 9412 946
rect 7412 901 9412 912
rect 9518 946 11518 957
rect 9518 912 9568 946
rect 9602 912 9636 946
rect 9670 912 9704 946
rect 9738 912 9772 946
rect 9806 912 9840 946
rect 9874 912 9908 946
rect 9942 912 9976 946
rect 10010 912 10044 946
rect 10078 912 10112 946
rect 10146 912 10180 946
rect 10214 912 10248 946
rect 10282 912 10316 946
rect 10350 912 10384 946
rect 10418 912 10452 946
rect 10486 912 10520 946
rect 10554 912 10588 946
rect 10622 912 10656 946
rect 10690 912 10724 946
rect 10758 912 10792 946
rect 10826 912 10860 946
rect 10894 912 10928 946
rect 10962 912 10996 946
rect 11030 912 11064 946
rect 11098 912 11132 946
rect 11166 912 11200 946
rect 11234 912 11268 946
rect 11302 912 11336 946
rect 11370 912 11404 946
rect 11438 912 11472 946
rect 11506 912 11518 946
rect 9518 901 11518 912
rect 7412 790 9412 801
rect 7412 756 7462 790
rect 7496 756 7530 790
rect 7564 756 7598 790
rect 7632 756 7666 790
rect 7700 756 7734 790
rect 7768 756 7802 790
rect 7836 756 7870 790
rect 7904 756 7938 790
rect 7972 756 8006 790
rect 8040 756 8074 790
rect 8108 756 8142 790
rect 8176 756 8210 790
rect 8244 756 8278 790
rect 8312 756 8346 790
rect 8380 756 8414 790
rect 8448 756 8482 790
rect 8516 756 8550 790
rect 8584 756 8618 790
rect 8652 756 8686 790
rect 8720 756 8754 790
rect 8788 756 8822 790
rect 8856 756 8890 790
rect 8924 756 8958 790
rect 8992 756 9026 790
rect 9060 756 9094 790
rect 9128 756 9162 790
rect 9196 756 9230 790
rect 9264 756 9298 790
rect 9332 756 9366 790
rect 9400 756 9412 790
rect 7412 745 9412 756
rect 9518 790 11518 801
rect 9518 756 9568 790
rect 9602 756 9636 790
rect 9670 756 9704 790
rect 9738 756 9772 790
rect 9806 756 9840 790
rect 9874 756 9908 790
rect 9942 756 9976 790
rect 10010 756 10044 790
rect 10078 756 10112 790
rect 10146 756 10180 790
rect 10214 756 10248 790
rect 10282 756 10316 790
rect 10350 756 10384 790
rect 10418 756 10452 790
rect 10486 756 10520 790
rect 10554 756 10588 790
rect 10622 756 10656 790
rect 10690 756 10724 790
rect 10758 756 10792 790
rect 10826 756 10860 790
rect 10894 756 10928 790
rect 10962 756 10996 790
rect 11030 756 11064 790
rect 11098 756 11132 790
rect 11166 756 11200 790
rect 11234 756 11268 790
rect 11302 756 11336 790
rect 11370 756 11404 790
rect 11438 756 11472 790
rect 11506 756 11518 790
rect 9518 745 11518 756
rect 7412 634 9412 645
rect 7412 600 7462 634
rect 7496 600 7530 634
rect 7564 600 7598 634
rect 7632 600 7666 634
rect 7700 600 7734 634
rect 7768 600 7802 634
rect 7836 600 7870 634
rect 7904 600 7938 634
rect 7972 600 8006 634
rect 8040 600 8074 634
rect 8108 600 8142 634
rect 8176 600 8210 634
rect 8244 600 8278 634
rect 8312 600 8346 634
rect 8380 600 8414 634
rect 8448 600 8482 634
rect 8516 600 8550 634
rect 8584 600 8618 634
rect 8652 600 8686 634
rect 8720 600 8754 634
rect 8788 600 8822 634
rect 8856 600 8890 634
rect 8924 600 8958 634
rect 8992 600 9026 634
rect 9060 600 9094 634
rect 9128 600 9162 634
rect 9196 600 9230 634
rect 9264 600 9298 634
rect 9332 600 9366 634
rect 9400 600 9412 634
rect 7412 589 9412 600
rect 9518 634 11518 645
rect 9518 600 9568 634
rect 9602 600 9636 634
rect 9670 600 9704 634
rect 9738 600 9772 634
rect 9806 600 9840 634
rect 9874 600 9908 634
rect 9942 600 9976 634
rect 10010 600 10044 634
rect 10078 600 10112 634
rect 10146 600 10180 634
rect 10214 600 10248 634
rect 10282 600 10316 634
rect 10350 600 10384 634
rect 10418 600 10452 634
rect 10486 600 10520 634
rect 10554 600 10588 634
rect 10622 600 10656 634
rect 10690 600 10724 634
rect 10758 600 10792 634
rect 10826 600 10860 634
rect 10894 600 10928 634
rect 10962 600 10996 634
rect 11030 600 11064 634
rect 11098 600 11132 634
rect 11166 600 11200 634
rect 11234 600 11268 634
rect 11302 600 11336 634
rect 11370 600 11404 634
rect 11438 600 11472 634
rect 11506 600 11518 634
rect 9518 589 11518 600
rect 7412 478 9412 489
rect 7412 444 7462 478
rect 7496 444 7530 478
rect 7564 444 7598 478
rect 7632 444 7666 478
rect 7700 444 7734 478
rect 7768 444 7802 478
rect 7836 444 7870 478
rect 7904 444 7938 478
rect 7972 444 8006 478
rect 8040 444 8074 478
rect 8108 444 8142 478
rect 8176 444 8210 478
rect 8244 444 8278 478
rect 8312 444 8346 478
rect 8380 444 8414 478
rect 8448 444 8482 478
rect 8516 444 8550 478
rect 8584 444 8618 478
rect 8652 444 8686 478
rect 8720 444 8754 478
rect 8788 444 8822 478
rect 8856 444 8890 478
rect 8924 444 8958 478
rect 8992 444 9026 478
rect 9060 444 9094 478
rect 9128 444 9162 478
rect 9196 444 9230 478
rect 9264 444 9298 478
rect 9332 444 9366 478
rect 9400 444 9412 478
rect 7412 436 9412 444
rect 9518 478 11518 489
rect 9518 444 9568 478
rect 9602 444 9636 478
rect 9670 444 9704 478
rect 9738 444 9772 478
rect 9806 444 9840 478
rect 9874 444 9908 478
rect 9942 444 9976 478
rect 10010 444 10044 478
rect 10078 444 10112 478
rect 10146 444 10180 478
rect 10214 444 10248 478
rect 10282 444 10316 478
rect 10350 444 10384 478
rect 10418 444 10452 478
rect 10486 444 10520 478
rect 10554 444 10588 478
rect 10622 444 10656 478
rect 10690 444 10724 478
rect 10758 444 10792 478
rect 10826 444 10860 478
rect 10894 444 10928 478
rect 10962 444 10996 478
rect 11030 444 11064 478
rect 11098 444 11132 478
rect 11166 444 11200 478
rect 11234 444 11268 478
rect 11302 444 11336 478
rect 11370 444 11404 478
rect 11438 444 11472 478
rect 11506 444 11518 478
rect 9518 436 11518 444
<< mvpdiff >>
rect 6616 -1270 8616 -1262
rect 6616 -1304 6666 -1270
rect 6700 -1304 6734 -1270
rect 6768 -1304 6802 -1270
rect 6836 -1304 6870 -1270
rect 6904 -1304 6938 -1270
rect 6972 -1304 7006 -1270
rect 7040 -1304 7074 -1270
rect 7108 -1304 7142 -1270
rect 7176 -1304 7210 -1270
rect 7244 -1304 7278 -1270
rect 7312 -1304 7346 -1270
rect 7380 -1304 7414 -1270
rect 7448 -1304 7482 -1270
rect 7516 -1304 7550 -1270
rect 7584 -1304 7618 -1270
rect 7652 -1304 7686 -1270
rect 7720 -1304 7754 -1270
rect 7788 -1304 7822 -1270
rect 7856 -1304 7890 -1270
rect 7924 -1304 7958 -1270
rect 7992 -1304 8026 -1270
rect 8060 -1304 8094 -1270
rect 8128 -1304 8162 -1270
rect 8196 -1304 8230 -1270
rect 8264 -1304 8298 -1270
rect 8332 -1304 8366 -1270
rect 8400 -1304 8434 -1270
rect 8468 -1304 8502 -1270
rect 8536 -1304 8570 -1270
rect 8604 -1304 8616 -1270
rect 6616 -1315 8616 -1304
rect 6616 -1426 8616 -1415
rect 6616 -1460 6666 -1426
rect 6700 -1460 6734 -1426
rect 6768 -1460 6802 -1426
rect 6836 -1460 6870 -1426
rect 6904 -1460 6938 -1426
rect 6972 -1460 7006 -1426
rect 7040 -1460 7074 -1426
rect 7108 -1460 7142 -1426
rect 7176 -1460 7210 -1426
rect 7244 -1460 7278 -1426
rect 7312 -1460 7346 -1426
rect 7380 -1460 7414 -1426
rect 7448 -1460 7482 -1426
rect 7516 -1460 7550 -1426
rect 7584 -1460 7618 -1426
rect 7652 -1460 7686 -1426
rect 7720 -1460 7754 -1426
rect 7788 -1460 7822 -1426
rect 7856 -1460 7890 -1426
rect 7924 -1460 7958 -1426
rect 7992 -1460 8026 -1426
rect 8060 -1460 8094 -1426
rect 8128 -1460 8162 -1426
rect 8196 -1460 8230 -1426
rect 8264 -1460 8298 -1426
rect 8332 -1460 8366 -1426
rect 8400 -1460 8434 -1426
rect 8468 -1460 8502 -1426
rect 8536 -1460 8570 -1426
rect 8604 -1460 8616 -1426
rect 6616 -1471 8616 -1460
rect 6616 -1582 8616 -1571
rect 6616 -1616 6666 -1582
rect 6700 -1616 6734 -1582
rect 6768 -1616 6802 -1582
rect 6836 -1616 6870 -1582
rect 6904 -1616 6938 -1582
rect 6972 -1616 7006 -1582
rect 7040 -1616 7074 -1582
rect 7108 -1616 7142 -1582
rect 7176 -1616 7210 -1582
rect 7244 -1616 7278 -1582
rect 7312 -1616 7346 -1582
rect 7380 -1616 7414 -1582
rect 7448 -1616 7482 -1582
rect 7516 -1616 7550 -1582
rect 7584 -1616 7618 -1582
rect 7652 -1616 7686 -1582
rect 7720 -1616 7754 -1582
rect 7788 -1616 7822 -1582
rect 7856 -1616 7890 -1582
rect 7924 -1616 7958 -1582
rect 7992 -1616 8026 -1582
rect 8060 -1616 8094 -1582
rect 8128 -1616 8162 -1582
rect 8196 -1616 8230 -1582
rect 8264 -1616 8298 -1582
rect 8332 -1616 8366 -1582
rect 8400 -1616 8434 -1582
rect 8468 -1616 8502 -1582
rect 8536 -1616 8570 -1582
rect 8604 -1616 8616 -1582
rect 6616 -1627 8616 -1616
rect 6616 -1738 8616 -1727
rect 6616 -1772 6666 -1738
rect 6700 -1772 6734 -1738
rect 6768 -1772 6802 -1738
rect 6836 -1772 6870 -1738
rect 6904 -1772 6938 -1738
rect 6972 -1772 7006 -1738
rect 7040 -1772 7074 -1738
rect 7108 -1772 7142 -1738
rect 7176 -1772 7210 -1738
rect 7244 -1772 7278 -1738
rect 7312 -1772 7346 -1738
rect 7380 -1772 7414 -1738
rect 7448 -1772 7482 -1738
rect 7516 -1772 7550 -1738
rect 7584 -1772 7618 -1738
rect 7652 -1772 7686 -1738
rect 7720 -1772 7754 -1738
rect 7788 -1772 7822 -1738
rect 7856 -1772 7890 -1738
rect 7924 -1772 7958 -1738
rect 7992 -1772 8026 -1738
rect 8060 -1772 8094 -1738
rect 8128 -1772 8162 -1738
rect 8196 -1772 8230 -1738
rect 8264 -1772 8298 -1738
rect 8332 -1772 8366 -1738
rect 8400 -1772 8434 -1738
rect 8468 -1772 8502 -1738
rect 8536 -1772 8570 -1738
rect 8604 -1772 8616 -1738
rect 6616 -1783 8616 -1772
rect 6616 -1894 8616 -1883
rect 6616 -1928 6666 -1894
rect 6700 -1928 6734 -1894
rect 6768 -1928 6802 -1894
rect 6836 -1928 6870 -1894
rect 6904 -1928 6938 -1894
rect 6972 -1928 7006 -1894
rect 7040 -1928 7074 -1894
rect 7108 -1928 7142 -1894
rect 7176 -1928 7210 -1894
rect 7244 -1928 7278 -1894
rect 7312 -1928 7346 -1894
rect 7380 -1928 7414 -1894
rect 7448 -1928 7482 -1894
rect 7516 -1928 7550 -1894
rect 7584 -1928 7618 -1894
rect 7652 -1928 7686 -1894
rect 7720 -1928 7754 -1894
rect 7788 -1928 7822 -1894
rect 7856 -1928 7890 -1894
rect 7924 -1928 7958 -1894
rect 7992 -1928 8026 -1894
rect 8060 -1928 8094 -1894
rect 8128 -1928 8162 -1894
rect 8196 -1928 8230 -1894
rect 8264 -1928 8298 -1894
rect 8332 -1928 8366 -1894
rect 8400 -1928 8434 -1894
rect 8468 -1928 8502 -1894
rect 8536 -1928 8570 -1894
rect 8604 -1928 8616 -1894
rect 6616 -1936 8616 -1928
<< mvndiffc >>
rect 570 1198 604 1232
rect 638 1198 672 1232
rect 706 1198 740 1232
rect 774 1198 808 1232
rect 842 1198 876 1232
rect 910 1198 944 1232
rect 978 1198 1012 1232
rect 1046 1198 1080 1232
rect 1114 1198 1148 1232
rect 1182 1198 1216 1232
rect 1250 1198 1284 1232
rect 1318 1198 1352 1232
rect 1386 1198 1420 1232
rect 1454 1198 1488 1232
rect 570 1042 604 1076
rect 638 1042 672 1076
rect 706 1042 740 1076
rect 774 1042 808 1076
rect 842 1042 876 1076
rect 910 1042 944 1076
rect 978 1042 1012 1076
rect 1046 1042 1080 1076
rect 1114 1042 1148 1076
rect 1182 1042 1216 1076
rect 1250 1042 1284 1076
rect 1318 1042 1352 1076
rect 1386 1042 1420 1076
rect 1454 1042 1488 1076
rect 570 886 604 920
rect 638 886 672 920
rect 706 886 740 920
rect 774 886 808 920
rect 842 886 876 920
rect 910 886 944 920
rect 978 886 1012 920
rect 1046 886 1080 920
rect 1114 886 1148 920
rect 1182 886 1216 920
rect 1250 886 1284 920
rect 1318 886 1352 920
rect 1386 886 1420 920
rect 1454 886 1488 920
rect 570 756 604 790
rect 638 756 672 790
rect 706 756 740 790
rect 774 756 808 790
rect 842 756 876 790
rect 910 756 944 790
rect 978 756 1012 790
rect 1046 756 1080 790
rect 1114 756 1148 790
rect 1182 756 1216 790
rect 1250 756 1284 790
rect 1318 756 1352 790
rect 1386 756 1420 790
rect 1454 756 1488 790
rect 570 600 604 634
rect 638 600 672 634
rect 706 600 740 634
rect 774 600 808 634
rect 842 600 876 634
rect 910 600 944 634
rect 978 600 1012 634
rect 1046 600 1080 634
rect 1114 600 1148 634
rect 1182 600 1216 634
rect 1250 600 1284 634
rect 1318 600 1352 634
rect 1386 600 1420 634
rect 1454 600 1488 634
rect 570 444 604 478
rect 638 444 672 478
rect 706 444 740 478
rect 774 444 808 478
rect 842 444 876 478
rect 910 444 944 478
rect 978 444 1012 478
rect 1046 444 1080 478
rect 1114 444 1148 478
rect 1182 444 1216 478
rect 1250 444 1284 478
rect 1318 444 1352 478
rect 1386 444 1420 478
rect 1454 444 1488 478
rect 2405 1224 2439 1258
rect 2473 1224 2507 1258
rect 2541 1224 2575 1258
rect 2609 1224 2643 1258
rect 2677 1224 2711 1258
rect 2745 1224 2779 1258
rect 2813 1224 2847 1258
rect 2881 1224 2915 1258
rect 2949 1224 2983 1258
rect 3017 1224 3051 1258
rect 3085 1224 3119 1258
rect 3153 1224 3187 1258
rect 3221 1224 3255 1258
rect 3289 1224 3323 1258
rect 3357 1224 3391 1258
rect 3425 1224 3459 1258
rect 3493 1224 3527 1258
rect 3561 1224 3595 1258
rect 3629 1224 3663 1258
rect 3697 1224 3731 1258
rect 3765 1224 3799 1258
rect 3833 1224 3867 1258
rect 3901 1224 3935 1258
rect 3969 1224 4003 1258
rect 4037 1224 4071 1258
rect 4105 1224 4139 1258
rect 4173 1224 4207 1258
rect 4241 1224 4275 1258
rect 4309 1224 4343 1258
rect 4549 1224 4583 1258
rect 4617 1224 4651 1258
rect 4685 1224 4719 1258
rect 4753 1224 4787 1258
rect 4821 1224 4855 1258
rect 4889 1224 4923 1258
rect 4957 1224 4991 1258
rect 5025 1224 5059 1258
rect 5093 1224 5127 1258
rect 5161 1224 5195 1258
rect 5229 1224 5263 1258
rect 5297 1224 5331 1258
rect 5365 1224 5399 1258
rect 5433 1224 5467 1258
rect 5501 1224 5535 1258
rect 5569 1224 5603 1258
rect 5637 1224 5671 1258
rect 5705 1224 5739 1258
rect 5773 1224 5807 1258
rect 5841 1224 5875 1258
rect 5909 1224 5943 1258
rect 5977 1224 6011 1258
rect 6045 1224 6079 1258
rect 6113 1224 6147 1258
rect 6181 1224 6215 1258
rect 6249 1224 6283 1258
rect 6317 1224 6351 1258
rect 6385 1224 6419 1258
rect 6453 1224 6487 1258
rect 2405 1068 2439 1102
rect 2473 1068 2507 1102
rect 2541 1068 2575 1102
rect 2609 1068 2643 1102
rect 2677 1068 2711 1102
rect 2745 1068 2779 1102
rect 2813 1068 2847 1102
rect 2881 1068 2915 1102
rect 2949 1068 2983 1102
rect 3017 1068 3051 1102
rect 3085 1068 3119 1102
rect 3153 1068 3187 1102
rect 3221 1068 3255 1102
rect 3289 1068 3323 1102
rect 3357 1068 3391 1102
rect 3425 1068 3459 1102
rect 3493 1068 3527 1102
rect 3561 1068 3595 1102
rect 3629 1068 3663 1102
rect 3697 1068 3731 1102
rect 3765 1068 3799 1102
rect 3833 1068 3867 1102
rect 3901 1068 3935 1102
rect 3969 1068 4003 1102
rect 4037 1068 4071 1102
rect 4105 1068 4139 1102
rect 4173 1068 4207 1102
rect 4241 1068 4275 1102
rect 4309 1068 4343 1102
rect 4549 1068 4583 1102
rect 4617 1068 4651 1102
rect 4685 1068 4719 1102
rect 4753 1068 4787 1102
rect 4821 1068 4855 1102
rect 4889 1068 4923 1102
rect 4957 1068 4991 1102
rect 5025 1068 5059 1102
rect 5093 1068 5127 1102
rect 5161 1068 5195 1102
rect 5229 1068 5263 1102
rect 5297 1068 5331 1102
rect 5365 1068 5399 1102
rect 5433 1068 5467 1102
rect 5501 1068 5535 1102
rect 5569 1068 5603 1102
rect 5637 1068 5671 1102
rect 5705 1068 5739 1102
rect 5773 1068 5807 1102
rect 5841 1068 5875 1102
rect 5909 1068 5943 1102
rect 5977 1068 6011 1102
rect 6045 1068 6079 1102
rect 6113 1068 6147 1102
rect 6181 1068 6215 1102
rect 6249 1068 6283 1102
rect 6317 1068 6351 1102
rect 6385 1068 6419 1102
rect 6453 1068 6487 1102
rect 2405 912 2439 946
rect 2473 912 2507 946
rect 2541 912 2575 946
rect 2609 912 2643 946
rect 2677 912 2711 946
rect 2745 912 2779 946
rect 2813 912 2847 946
rect 2881 912 2915 946
rect 2949 912 2983 946
rect 3017 912 3051 946
rect 3085 912 3119 946
rect 3153 912 3187 946
rect 3221 912 3255 946
rect 3289 912 3323 946
rect 3357 912 3391 946
rect 3425 912 3459 946
rect 3493 912 3527 946
rect 3561 912 3595 946
rect 3629 912 3663 946
rect 3697 912 3731 946
rect 3765 912 3799 946
rect 3833 912 3867 946
rect 3901 912 3935 946
rect 3969 912 4003 946
rect 4037 912 4071 946
rect 4105 912 4139 946
rect 4173 912 4207 946
rect 4241 912 4275 946
rect 4309 912 4343 946
rect 4549 912 4583 946
rect 4617 912 4651 946
rect 4685 912 4719 946
rect 4753 912 4787 946
rect 4821 912 4855 946
rect 4889 912 4923 946
rect 4957 912 4991 946
rect 5025 912 5059 946
rect 5093 912 5127 946
rect 5161 912 5195 946
rect 5229 912 5263 946
rect 5297 912 5331 946
rect 5365 912 5399 946
rect 5433 912 5467 946
rect 5501 912 5535 946
rect 5569 912 5603 946
rect 5637 912 5671 946
rect 5705 912 5739 946
rect 5773 912 5807 946
rect 5841 912 5875 946
rect 5909 912 5943 946
rect 5977 912 6011 946
rect 6045 912 6079 946
rect 6113 912 6147 946
rect 6181 912 6215 946
rect 6249 912 6283 946
rect 6317 912 6351 946
rect 6385 912 6419 946
rect 6453 912 6487 946
rect 2405 756 2439 790
rect 2473 756 2507 790
rect 2541 756 2575 790
rect 2609 756 2643 790
rect 2677 756 2711 790
rect 2745 756 2779 790
rect 2813 756 2847 790
rect 2881 756 2915 790
rect 2949 756 2983 790
rect 3017 756 3051 790
rect 3085 756 3119 790
rect 3153 756 3187 790
rect 3221 756 3255 790
rect 3289 756 3323 790
rect 3357 756 3391 790
rect 3425 756 3459 790
rect 3493 756 3527 790
rect 3561 756 3595 790
rect 3629 756 3663 790
rect 3697 756 3731 790
rect 3765 756 3799 790
rect 3833 756 3867 790
rect 3901 756 3935 790
rect 3969 756 4003 790
rect 4037 756 4071 790
rect 4105 756 4139 790
rect 4173 756 4207 790
rect 4241 756 4275 790
rect 4309 756 4343 790
rect 4549 756 4583 790
rect 4617 756 4651 790
rect 4685 756 4719 790
rect 4753 756 4787 790
rect 4821 756 4855 790
rect 4889 756 4923 790
rect 4957 756 4991 790
rect 5025 756 5059 790
rect 5093 756 5127 790
rect 5161 756 5195 790
rect 5229 756 5263 790
rect 5297 756 5331 790
rect 5365 756 5399 790
rect 5433 756 5467 790
rect 5501 756 5535 790
rect 5569 756 5603 790
rect 5637 756 5671 790
rect 5705 756 5739 790
rect 5773 756 5807 790
rect 5841 756 5875 790
rect 5909 756 5943 790
rect 5977 756 6011 790
rect 6045 756 6079 790
rect 6113 756 6147 790
rect 6181 756 6215 790
rect 6249 756 6283 790
rect 6317 756 6351 790
rect 6385 756 6419 790
rect 6453 756 6487 790
rect 2405 600 2439 634
rect 2473 600 2507 634
rect 2541 600 2575 634
rect 2609 600 2643 634
rect 2677 600 2711 634
rect 2745 600 2779 634
rect 2813 600 2847 634
rect 2881 600 2915 634
rect 2949 600 2983 634
rect 3017 600 3051 634
rect 3085 600 3119 634
rect 3153 600 3187 634
rect 3221 600 3255 634
rect 3289 600 3323 634
rect 3357 600 3391 634
rect 3425 600 3459 634
rect 3493 600 3527 634
rect 3561 600 3595 634
rect 3629 600 3663 634
rect 3697 600 3731 634
rect 3765 600 3799 634
rect 3833 600 3867 634
rect 3901 600 3935 634
rect 3969 600 4003 634
rect 4037 600 4071 634
rect 4105 600 4139 634
rect 4173 600 4207 634
rect 4241 600 4275 634
rect 4309 600 4343 634
rect 4549 600 4583 634
rect 4617 600 4651 634
rect 4685 600 4719 634
rect 4753 600 4787 634
rect 4821 600 4855 634
rect 4889 600 4923 634
rect 4957 600 4991 634
rect 5025 600 5059 634
rect 5093 600 5127 634
rect 5161 600 5195 634
rect 5229 600 5263 634
rect 5297 600 5331 634
rect 5365 600 5399 634
rect 5433 600 5467 634
rect 5501 600 5535 634
rect 5569 600 5603 634
rect 5637 600 5671 634
rect 5705 600 5739 634
rect 5773 600 5807 634
rect 5841 600 5875 634
rect 5909 600 5943 634
rect 5977 600 6011 634
rect 6045 600 6079 634
rect 6113 600 6147 634
rect 6181 600 6215 634
rect 6249 600 6283 634
rect 6317 600 6351 634
rect 6385 600 6419 634
rect 6453 600 6487 634
rect 2405 444 2439 478
rect 2473 444 2507 478
rect 2541 444 2575 478
rect 2609 444 2643 478
rect 2677 444 2711 478
rect 2745 444 2779 478
rect 2813 444 2847 478
rect 2881 444 2915 478
rect 2949 444 2983 478
rect 3017 444 3051 478
rect 3085 444 3119 478
rect 3153 444 3187 478
rect 3221 444 3255 478
rect 3289 444 3323 478
rect 3357 444 3391 478
rect 3425 444 3459 478
rect 3493 444 3527 478
rect 3561 444 3595 478
rect 3629 444 3663 478
rect 3697 444 3731 478
rect 3765 444 3799 478
rect 3833 444 3867 478
rect 3901 444 3935 478
rect 3969 444 4003 478
rect 4037 444 4071 478
rect 4105 444 4139 478
rect 4173 444 4207 478
rect 4241 444 4275 478
rect 4309 444 4343 478
rect 4549 444 4583 478
rect 4617 444 4651 478
rect 4685 444 4719 478
rect 4753 444 4787 478
rect 4821 444 4855 478
rect 4889 444 4923 478
rect 4957 444 4991 478
rect 5025 444 5059 478
rect 5093 444 5127 478
rect 5161 444 5195 478
rect 5229 444 5263 478
rect 5297 444 5331 478
rect 5365 444 5399 478
rect 5433 444 5467 478
rect 5501 444 5535 478
rect 5569 444 5603 478
rect 5637 444 5671 478
rect 5705 444 5739 478
rect 5773 444 5807 478
rect 5841 444 5875 478
rect 5909 444 5943 478
rect 5977 444 6011 478
rect 6045 444 6079 478
rect 6113 444 6147 478
rect 6181 444 6215 478
rect 6249 444 6283 478
rect 6317 444 6351 478
rect 6385 444 6419 478
rect 6453 444 6487 478
rect 7462 1224 7496 1258
rect 7530 1224 7564 1258
rect 7598 1224 7632 1258
rect 7666 1224 7700 1258
rect 7734 1224 7768 1258
rect 7802 1224 7836 1258
rect 7870 1224 7904 1258
rect 7938 1224 7972 1258
rect 8006 1224 8040 1258
rect 8074 1224 8108 1258
rect 8142 1224 8176 1258
rect 8210 1224 8244 1258
rect 8278 1224 8312 1258
rect 8346 1224 8380 1258
rect 8414 1224 8448 1258
rect 8482 1224 8516 1258
rect 8550 1224 8584 1258
rect 8618 1224 8652 1258
rect 8686 1224 8720 1258
rect 8754 1224 8788 1258
rect 8822 1224 8856 1258
rect 8890 1224 8924 1258
rect 8958 1224 8992 1258
rect 9026 1224 9060 1258
rect 9094 1224 9128 1258
rect 9162 1224 9196 1258
rect 9230 1224 9264 1258
rect 9298 1224 9332 1258
rect 9366 1224 9400 1258
rect 9568 1224 9602 1258
rect 9636 1224 9670 1258
rect 9704 1224 9738 1258
rect 9772 1224 9806 1258
rect 9840 1224 9874 1258
rect 9908 1224 9942 1258
rect 9976 1224 10010 1258
rect 10044 1224 10078 1258
rect 10112 1224 10146 1258
rect 10180 1224 10214 1258
rect 10248 1224 10282 1258
rect 10316 1224 10350 1258
rect 10384 1224 10418 1258
rect 10452 1224 10486 1258
rect 10520 1224 10554 1258
rect 10588 1224 10622 1258
rect 10656 1224 10690 1258
rect 10724 1224 10758 1258
rect 10792 1224 10826 1258
rect 10860 1224 10894 1258
rect 10928 1224 10962 1258
rect 10996 1224 11030 1258
rect 11064 1224 11098 1258
rect 11132 1224 11166 1258
rect 11200 1224 11234 1258
rect 11268 1224 11302 1258
rect 11336 1224 11370 1258
rect 11404 1224 11438 1258
rect 11472 1224 11506 1258
rect 7462 1068 7496 1102
rect 7530 1068 7564 1102
rect 7598 1068 7632 1102
rect 7666 1068 7700 1102
rect 7734 1068 7768 1102
rect 7802 1068 7836 1102
rect 7870 1068 7904 1102
rect 7938 1068 7972 1102
rect 8006 1068 8040 1102
rect 8074 1068 8108 1102
rect 8142 1068 8176 1102
rect 8210 1068 8244 1102
rect 8278 1068 8312 1102
rect 8346 1068 8380 1102
rect 8414 1068 8448 1102
rect 8482 1068 8516 1102
rect 8550 1068 8584 1102
rect 8618 1068 8652 1102
rect 8686 1068 8720 1102
rect 8754 1068 8788 1102
rect 8822 1068 8856 1102
rect 8890 1068 8924 1102
rect 8958 1068 8992 1102
rect 9026 1068 9060 1102
rect 9094 1068 9128 1102
rect 9162 1068 9196 1102
rect 9230 1068 9264 1102
rect 9298 1068 9332 1102
rect 9366 1068 9400 1102
rect 9568 1068 9602 1102
rect 9636 1068 9670 1102
rect 9704 1068 9738 1102
rect 9772 1068 9806 1102
rect 9840 1068 9874 1102
rect 9908 1068 9942 1102
rect 9976 1068 10010 1102
rect 10044 1068 10078 1102
rect 10112 1068 10146 1102
rect 10180 1068 10214 1102
rect 10248 1068 10282 1102
rect 10316 1068 10350 1102
rect 10384 1068 10418 1102
rect 10452 1068 10486 1102
rect 10520 1068 10554 1102
rect 10588 1068 10622 1102
rect 10656 1068 10690 1102
rect 10724 1068 10758 1102
rect 10792 1068 10826 1102
rect 10860 1068 10894 1102
rect 10928 1068 10962 1102
rect 10996 1068 11030 1102
rect 11064 1068 11098 1102
rect 11132 1068 11166 1102
rect 11200 1068 11234 1102
rect 11268 1068 11302 1102
rect 11336 1068 11370 1102
rect 11404 1068 11438 1102
rect 11472 1068 11506 1102
rect 7462 912 7496 946
rect 7530 912 7564 946
rect 7598 912 7632 946
rect 7666 912 7700 946
rect 7734 912 7768 946
rect 7802 912 7836 946
rect 7870 912 7904 946
rect 7938 912 7972 946
rect 8006 912 8040 946
rect 8074 912 8108 946
rect 8142 912 8176 946
rect 8210 912 8244 946
rect 8278 912 8312 946
rect 8346 912 8380 946
rect 8414 912 8448 946
rect 8482 912 8516 946
rect 8550 912 8584 946
rect 8618 912 8652 946
rect 8686 912 8720 946
rect 8754 912 8788 946
rect 8822 912 8856 946
rect 8890 912 8924 946
rect 8958 912 8992 946
rect 9026 912 9060 946
rect 9094 912 9128 946
rect 9162 912 9196 946
rect 9230 912 9264 946
rect 9298 912 9332 946
rect 9366 912 9400 946
rect 9568 912 9602 946
rect 9636 912 9670 946
rect 9704 912 9738 946
rect 9772 912 9806 946
rect 9840 912 9874 946
rect 9908 912 9942 946
rect 9976 912 10010 946
rect 10044 912 10078 946
rect 10112 912 10146 946
rect 10180 912 10214 946
rect 10248 912 10282 946
rect 10316 912 10350 946
rect 10384 912 10418 946
rect 10452 912 10486 946
rect 10520 912 10554 946
rect 10588 912 10622 946
rect 10656 912 10690 946
rect 10724 912 10758 946
rect 10792 912 10826 946
rect 10860 912 10894 946
rect 10928 912 10962 946
rect 10996 912 11030 946
rect 11064 912 11098 946
rect 11132 912 11166 946
rect 11200 912 11234 946
rect 11268 912 11302 946
rect 11336 912 11370 946
rect 11404 912 11438 946
rect 11472 912 11506 946
rect 7462 756 7496 790
rect 7530 756 7564 790
rect 7598 756 7632 790
rect 7666 756 7700 790
rect 7734 756 7768 790
rect 7802 756 7836 790
rect 7870 756 7904 790
rect 7938 756 7972 790
rect 8006 756 8040 790
rect 8074 756 8108 790
rect 8142 756 8176 790
rect 8210 756 8244 790
rect 8278 756 8312 790
rect 8346 756 8380 790
rect 8414 756 8448 790
rect 8482 756 8516 790
rect 8550 756 8584 790
rect 8618 756 8652 790
rect 8686 756 8720 790
rect 8754 756 8788 790
rect 8822 756 8856 790
rect 8890 756 8924 790
rect 8958 756 8992 790
rect 9026 756 9060 790
rect 9094 756 9128 790
rect 9162 756 9196 790
rect 9230 756 9264 790
rect 9298 756 9332 790
rect 9366 756 9400 790
rect 9568 756 9602 790
rect 9636 756 9670 790
rect 9704 756 9738 790
rect 9772 756 9806 790
rect 9840 756 9874 790
rect 9908 756 9942 790
rect 9976 756 10010 790
rect 10044 756 10078 790
rect 10112 756 10146 790
rect 10180 756 10214 790
rect 10248 756 10282 790
rect 10316 756 10350 790
rect 10384 756 10418 790
rect 10452 756 10486 790
rect 10520 756 10554 790
rect 10588 756 10622 790
rect 10656 756 10690 790
rect 10724 756 10758 790
rect 10792 756 10826 790
rect 10860 756 10894 790
rect 10928 756 10962 790
rect 10996 756 11030 790
rect 11064 756 11098 790
rect 11132 756 11166 790
rect 11200 756 11234 790
rect 11268 756 11302 790
rect 11336 756 11370 790
rect 11404 756 11438 790
rect 11472 756 11506 790
rect 7462 600 7496 634
rect 7530 600 7564 634
rect 7598 600 7632 634
rect 7666 600 7700 634
rect 7734 600 7768 634
rect 7802 600 7836 634
rect 7870 600 7904 634
rect 7938 600 7972 634
rect 8006 600 8040 634
rect 8074 600 8108 634
rect 8142 600 8176 634
rect 8210 600 8244 634
rect 8278 600 8312 634
rect 8346 600 8380 634
rect 8414 600 8448 634
rect 8482 600 8516 634
rect 8550 600 8584 634
rect 8618 600 8652 634
rect 8686 600 8720 634
rect 8754 600 8788 634
rect 8822 600 8856 634
rect 8890 600 8924 634
rect 8958 600 8992 634
rect 9026 600 9060 634
rect 9094 600 9128 634
rect 9162 600 9196 634
rect 9230 600 9264 634
rect 9298 600 9332 634
rect 9366 600 9400 634
rect 9568 600 9602 634
rect 9636 600 9670 634
rect 9704 600 9738 634
rect 9772 600 9806 634
rect 9840 600 9874 634
rect 9908 600 9942 634
rect 9976 600 10010 634
rect 10044 600 10078 634
rect 10112 600 10146 634
rect 10180 600 10214 634
rect 10248 600 10282 634
rect 10316 600 10350 634
rect 10384 600 10418 634
rect 10452 600 10486 634
rect 10520 600 10554 634
rect 10588 600 10622 634
rect 10656 600 10690 634
rect 10724 600 10758 634
rect 10792 600 10826 634
rect 10860 600 10894 634
rect 10928 600 10962 634
rect 10996 600 11030 634
rect 11064 600 11098 634
rect 11132 600 11166 634
rect 11200 600 11234 634
rect 11268 600 11302 634
rect 11336 600 11370 634
rect 11404 600 11438 634
rect 11472 600 11506 634
rect 7462 444 7496 478
rect 7530 444 7564 478
rect 7598 444 7632 478
rect 7666 444 7700 478
rect 7734 444 7768 478
rect 7802 444 7836 478
rect 7870 444 7904 478
rect 7938 444 7972 478
rect 8006 444 8040 478
rect 8074 444 8108 478
rect 8142 444 8176 478
rect 8210 444 8244 478
rect 8278 444 8312 478
rect 8346 444 8380 478
rect 8414 444 8448 478
rect 8482 444 8516 478
rect 8550 444 8584 478
rect 8618 444 8652 478
rect 8686 444 8720 478
rect 8754 444 8788 478
rect 8822 444 8856 478
rect 8890 444 8924 478
rect 8958 444 8992 478
rect 9026 444 9060 478
rect 9094 444 9128 478
rect 9162 444 9196 478
rect 9230 444 9264 478
rect 9298 444 9332 478
rect 9366 444 9400 478
rect 9568 444 9602 478
rect 9636 444 9670 478
rect 9704 444 9738 478
rect 9772 444 9806 478
rect 9840 444 9874 478
rect 9908 444 9942 478
rect 9976 444 10010 478
rect 10044 444 10078 478
rect 10112 444 10146 478
rect 10180 444 10214 478
rect 10248 444 10282 478
rect 10316 444 10350 478
rect 10384 444 10418 478
rect 10452 444 10486 478
rect 10520 444 10554 478
rect 10588 444 10622 478
rect 10656 444 10690 478
rect 10724 444 10758 478
rect 10792 444 10826 478
rect 10860 444 10894 478
rect 10928 444 10962 478
rect 10996 444 11030 478
rect 11064 444 11098 478
rect 11132 444 11166 478
rect 11200 444 11234 478
rect 11268 444 11302 478
rect 11336 444 11370 478
rect 11404 444 11438 478
rect 11472 444 11506 478
<< mvpdiffc >>
rect 6666 -1304 6700 -1270
rect 6734 -1304 6768 -1270
rect 6802 -1304 6836 -1270
rect 6870 -1304 6904 -1270
rect 6938 -1304 6972 -1270
rect 7006 -1304 7040 -1270
rect 7074 -1304 7108 -1270
rect 7142 -1304 7176 -1270
rect 7210 -1304 7244 -1270
rect 7278 -1304 7312 -1270
rect 7346 -1304 7380 -1270
rect 7414 -1304 7448 -1270
rect 7482 -1304 7516 -1270
rect 7550 -1304 7584 -1270
rect 7618 -1304 7652 -1270
rect 7686 -1304 7720 -1270
rect 7754 -1304 7788 -1270
rect 7822 -1304 7856 -1270
rect 7890 -1304 7924 -1270
rect 7958 -1304 7992 -1270
rect 8026 -1304 8060 -1270
rect 8094 -1304 8128 -1270
rect 8162 -1304 8196 -1270
rect 8230 -1304 8264 -1270
rect 8298 -1304 8332 -1270
rect 8366 -1304 8400 -1270
rect 8434 -1304 8468 -1270
rect 8502 -1304 8536 -1270
rect 8570 -1304 8604 -1270
rect 6666 -1460 6700 -1426
rect 6734 -1460 6768 -1426
rect 6802 -1460 6836 -1426
rect 6870 -1460 6904 -1426
rect 6938 -1460 6972 -1426
rect 7006 -1460 7040 -1426
rect 7074 -1460 7108 -1426
rect 7142 -1460 7176 -1426
rect 7210 -1460 7244 -1426
rect 7278 -1460 7312 -1426
rect 7346 -1460 7380 -1426
rect 7414 -1460 7448 -1426
rect 7482 -1460 7516 -1426
rect 7550 -1460 7584 -1426
rect 7618 -1460 7652 -1426
rect 7686 -1460 7720 -1426
rect 7754 -1460 7788 -1426
rect 7822 -1460 7856 -1426
rect 7890 -1460 7924 -1426
rect 7958 -1460 7992 -1426
rect 8026 -1460 8060 -1426
rect 8094 -1460 8128 -1426
rect 8162 -1460 8196 -1426
rect 8230 -1460 8264 -1426
rect 8298 -1460 8332 -1426
rect 8366 -1460 8400 -1426
rect 8434 -1460 8468 -1426
rect 8502 -1460 8536 -1426
rect 8570 -1460 8604 -1426
rect 6666 -1616 6700 -1582
rect 6734 -1616 6768 -1582
rect 6802 -1616 6836 -1582
rect 6870 -1616 6904 -1582
rect 6938 -1616 6972 -1582
rect 7006 -1616 7040 -1582
rect 7074 -1616 7108 -1582
rect 7142 -1616 7176 -1582
rect 7210 -1616 7244 -1582
rect 7278 -1616 7312 -1582
rect 7346 -1616 7380 -1582
rect 7414 -1616 7448 -1582
rect 7482 -1616 7516 -1582
rect 7550 -1616 7584 -1582
rect 7618 -1616 7652 -1582
rect 7686 -1616 7720 -1582
rect 7754 -1616 7788 -1582
rect 7822 -1616 7856 -1582
rect 7890 -1616 7924 -1582
rect 7958 -1616 7992 -1582
rect 8026 -1616 8060 -1582
rect 8094 -1616 8128 -1582
rect 8162 -1616 8196 -1582
rect 8230 -1616 8264 -1582
rect 8298 -1616 8332 -1582
rect 8366 -1616 8400 -1582
rect 8434 -1616 8468 -1582
rect 8502 -1616 8536 -1582
rect 8570 -1616 8604 -1582
rect 6666 -1772 6700 -1738
rect 6734 -1772 6768 -1738
rect 6802 -1772 6836 -1738
rect 6870 -1772 6904 -1738
rect 6938 -1772 6972 -1738
rect 7006 -1772 7040 -1738
rect 7074 -1772 7108 -1738
rect 7142 -1772 7176 -1738
rect 7210 -1772 7244 -1738
rect 7278 -1772 7312 -1738
rect 7346 -1772 7380 -1738
rect 7414 -1772 7448 -1738
rect 7482 -1772 7516 -1738
rect 7550 -1772 7584 -1738
rect 7618 -1772 7652 -1738
rect 7686 -1772 7720 -1738
rect 7754 -1772 7788 -1738
rect 7822 -1772 7856 -1738
rect 7890 -1772 7924 -1738
rect 7958 -1772 7992 -1738
rect 8026 -1772 8060 -1738
rect 8094 -1772 8128 -1738
rect 8162 -1772 8196 -1738
rect 8230 -1772 8264 -1738
rect 8298 -1772 8332 -1738
rect 8366 -1772 8400 -1738
rect 8434 -1772 8468 -1738
rect 8502 -1772 8536 -1738
rect 8570 -1772 8604 -1738
rect 6666 -1928 6700 -1894
rect 6734 -1928 6768 -1894
rect 6802 -1928 6836 -1894
rect 6870 -1928 6904 -1894
rect 6938 -1928 6972 -1894
rect 7006 -1928 7040 -1894
rect 7074 -1928 7108 -1894
rect 7142 -1928 7176 -1894
rect 7210 -1928 7244 -1894
rect 7278 -1928 7312 -1894
rect 7346 -1928 7380 -1894
rect 7414 -1928 7448 -1894
rect 7482 -1928 7516 -1894
rect 7550 -1928 7584 -1894
rect 7618 -1928 7652 -1894
rect 7686 -1928 7720 -1894
rect 7754 -1928 7788 -1894
rect 7822 -1928 7856 -1894
rect 7890 -1928 7924 -1894
rect 7958 -1928 7992 -1894
rect 8026 -1928 8060 -1894
rect 8094 -1928 8128 -1894
rect 8162 -1928 8196 -1894
rect 8230 -1928 8264 -1894
rect 8298 -1928 8332 -1894
rect 8366 -1928 8400 -1894
rect 8434 -1928 8468 -1894
rect 8502 -1928 8536 -1894
rect 8570 -1928 8604 -1894
<< mvpsubdiff >>
rect 357 1351 1709 1354
rect 357 1317 458 1351
rect 492 1317 526 1351
rect 560 1317 594 1351
rect 628 1317 662 1351
rect 696 1317 730 1351
rect 764 1317 798 1351
rect 832 1317 866 1351
rect 900 1317 934 1351
rect 968 1317 1002 1351
rect 1036 1317 1131 1351
rect 1165 1317 1199 1351
rect 1233 1317 1267 1351
rect 1301 1317 1335 1351
rect 1369 1317 1403 1351
rect 1437 1317 1471 1351
rect 1505 1317 1539 1351
rect 1573 1317 1607 1351
rect 1641 1317 1709 1351
rect 357 1314 1709 1317
rect 357 1286 397 1314
rect 357 1252 360 1286
rect 394 1252 397 1286
rect 357 1218 397 1252
rect 1669 1240 1709 1314
rect 357 1184 360 1218
rect 394 1184 397 1218
rect 1669 1206 1672 1240
rect 1706 1206 1709 1240
rect 357 1150 397 1184
rect 357 1116 360 1150
rect 394 1116 397 1150
rect 357 1082 397 1116
rect 357 1048 360 1082
rect 394 1048 397 1082
rect 357 1014 397 1048
rect 357 980 360 1014
rect 394 980 397 1014
rect 357 946 397 980
rect 357 912 360 946
rect 394 912 397 946
rect 357 878 397 912
rect 357 844 360 878
rect 394 844 397 878
rect 357 810 397 844
rect 357 776 360 810
rect 394 776 397 810
rect 357 742 397 776
rect 357 708 360 742
rect 394 708 397 742
rect 357 674 397 708
rect 357 640 360 674
rect 394 640 397 674
rect 357 606 397 640
rect 357 572 360 606
rect 394 572 397 606
rect 357 538 397 572
rect 357 504 360 538
rect 394 504 397 538
rect 357 470 397 504
rect 1669 1172 1709 1206
rect 1669 1138 1672 1172
rect 1706 1138 1709 1172
rect 1669 1104 1709 1138
rect 1669 1070 1672 1104
rect 1706 1070 1709 1104
rect 1669 1036 1709 1070
rect 1669 1002 1672 1036
rect 1706 1002 1709 1036
rect 1669 968 1709 1002
rect 1669 934 1672 968
rect 1706 934 1709 968
rect 1669 900 1709 934
rect 1669 866 1672 900
rect 1706 866 1709 900
rect 1669 832 1709 866
rect 1669 798 1672 832
rect 1706 798 1709 832
rect 1669 764 1709 798
rect 1669 730 1672 764
rect 1706 730 1709 764
rect 1669 696 1709 730
rect 1669 662 1672 696
rect 1706 662 1709 696
rect 1669 628 1709 662
rect 1669 594 1672 628
rect 1706 594 1709 628
rect 1669 560 1709 594
rect 1669 526 1672 560
rect 1706 526 1709 560
rect 1669 492 1709 526
rect 357 436 360 470
rect 394 436 397 470
rect 1669 458 1672 492
rect 1706 458 1709 492
rect 357 362 397 436
rect 1669 424 1709 458
rect 1669 390 1672 424
rect 1706 390 1709 424
rect 1669 362 1709 390
rect 357 359 1709 362
rect 357 325 425 359
rect 459 325 493 359
rect 527 325 561 359
rect 595 325 629 359
rect 663 325 697 359
rect 731 325 765 359
rect 799 325 833 359
rect 867 325 901 359
rect 935 325 969 359
rect 1003 325 1037 359
rect 1071 325 1105 359
rect 1139 325 1173 359
rect 1207 325 1241 359
rect 1275 325 1309 359
rect 1343 325 1377 359
rect 1411 325 1445 359
rect 1479 325 1513 359
rect 1547 325 1581 359
rect 1615 325 1709 359
rect 357 322 1709 325
rect 2192 1377 6720 1380
rect 2192 1343 2287 1377
rect 2321 1343 2355 1377
rect 2389 1343 2423 1377
rect 2457 1343 2491 1377
rect 2525 1343 2559 1377
rect 2593 1343 2627 1377
rect 2661 1343 2695 1377
rect 2729 1343 2763 1377
rect 2797 1343 2831 1377
rect 2865 1343 2899 1377
rect 2933 1343 2967 1377
rect 3001 1343 3035 1377
rect 3069 1343 3103 1377
rect 3137 1343 3171 1377
rect 3205 1343 3239 1377
rect 3273 1343 3307 1377
rect 3341 1343 3375 1377
rect 3409 1343 3443 1377
rect 3477 1343 3511 1377
rect 3545 1343 3579 1377
rect 3613 1343 3647 1377
rect 3681 1343 3715 1377
rect 3749 1343 3783 1377
rect 3817 1343 3851 1377
rect 3885 1343 3919 1377
rect 3953 1343 3987 1377
rect 4021 1343 4055 1377
rect 4089 1343 4123 1377
rect 4157 1343 4191 1377
rect 4225 1343 4259 1377
rect 4293 1343 4327 1377
rect 4361 1343 4395 1377
rect 4429 1343 4510 1377
rect 4544 1343 4578 1377
rect 4612 1343 4646 1377
rect 4680 1343 4714 1377
rect 4748 1343 4782 1377
rect 4816 1343 4850 1377
rect 4884 1343 4918 1377
rect 4952 1343 4986 1377
rect 5020 1343 5054 1377
rect 5088 1343 5122 1377
rect 5156 1343 5190 1377
rect 5224 1343 5258 1377
rect 5292 1343 5326 1377
rect 5360 1343 5394 1377
rect 5428 1343 5462 1377
rect 5496 1343 5530 1377
rect 5564 1343 5598 1377
rect 5632 1343 5666 1377
rect 5700 1343 5734 1377
rect 5768 1343 5802 1377
rect 5836 1343 5870 1377
rect 5904 1343 5938 1377
rect 5972 1343 6006 1377
rect 6040 1343 6074 1377
rect 6108 1343 6142 1377
rect 6176 1343 6210 1377
rect 6244 1343 6278 1377
rect 6312 1343 6346 1377
rect 6380 1343 6414 1377
rect 6448 1343 6482 1377
rect 6516 1343 6550 1377
rect 6584 1343 6618 1377
rect 6652 1343 6720 1377
rect 2192 1340 6720 1343
rect 2192 1312 2232 1340
rect 2192 1278 2195 1312
rect 2229 1278 2232 1312
rect 2192 1244 2232 1278
rect 6680 1308 6720 1340
rect 6680 1274 6683 1308
rect 6717 1274 6720 1308
rect 2192 1210 2195 1244
rect 2229 1210 2232 1244
rect 6680 1240 6720 1274
rect 2192 1176 2232 1210
rect 2192 1142 2195 1176
rect 2229 1142 2232 1176
rect 2192 1108 2232 1142
rect 2192 1074 2195 1108
rect 2229 1074 2232 1108
rect 2192 1040 2232 1074
rect 2192 1006 2195 1040
rect 2229 1006 2232 1040
rect 2192 972 2232 1006
rect 2192 938 2195 972
rect 2229 938 2232 972
rect 2192 904 2232 938
rect 2192 870 2195 904
rect 2229 870 2232 904
rect 2192 836 2232 870
rect 2192 802 2195 836
rect 2229 802 2232 836
rect 2192 768 2232 802
rect 2192 734 2195 768
rect 2229 734 2232 768
rect 2192 700 2232 734
rect 2192 666 2195 700
rect 2229 666 2232 700
rect 2192 632 2232 666
rect 2192 598 2195 632
rect 2229 598 2232 632
rect 2192 564 2232 598
rect 2192 530 2195 564
rect 2229 530 2232 564
rect 2192 496 2232 530
rect 2192 462 2195 496
rect 2229 462 2232 496
rect 6680 1206 6683 1240
rect 6717 1206 6720 1240
rect 6680 1172 6720 1206
rect 6680 1138 6683 1172
rect 6717 1138 6720 1172
rect 6680 1104 6720 1138
rect 6680 1070 6683 1104
rect 6717 1070 6720 1104
rect 6680 1036 6720 1070
rect 6680 1002 6683 1036
rect 6717 1002 6720 1036
rect 6680 968 6720 1002
rect 6680 934 6683 968
rect 6717 934 6720 968
rect 6680 900 6720 934
rect 6680 866 6683 900
rect 6717 866 6720 900
rect 6680 832 6720 866
rect 6680 798 6683 832
rect 6717 798 6720 832
rect 6680 764 6720 798
rect 6680 730 6683 764
rect 6717 730 6720 764
rect 6680 696 6720 730
rect 6680 662 6683 696
rect 6717 662 6720 696
rect 6680 628 6720 662
rect 6680 594 6683 628
rect 6717 594 6720 628
rect 6680 560 6720 594
rect 6680 526 6683 560
rect 6717 526 6720 560
rect 6680 492 6720 526
rect 2192 428 2232 462
rect 6680 458 6683 492
rect 6717 458 6720 492
rect 2192 394 2195 428
rect 2229 394 2232 428
rect 2192 362 2232 394
rect 6680 424 6720 458
rect 6680 390 6683 424
rect 6717 390 6720 424
rect 6680 362 6720 390
rect 2192 359 6720 362
rect 2192 325 2260 359
rect 2294 325 2328 359
rect 2362 325 2396 359
rect 2430 325 2464 359
rect 2498 325 2532 359
rect 2566 325 2600 359
rect 2634 325 2668 359
rect 2702 325 2736 359
rect 2770 325 2804 359
rect 2838 325 2872 359
rect 2906 325 2940 359
rect 2974 325 3008 359
rect 3042 325 3076 359
rect 3110 325 3144 359
rect 3178 325 3212 359
rect 3246 325 3280 359
rect 3314 325 3348 359
rect 3382 325 3416 359
rect 3450 325 3484 359
rect 3518 325 3552 359
rect 3586 325 3620 359
rect 3654 325 3688 359
rect 3722 325 3756 359
rect 3790 325 3824 359
rect 3858 325 3892 359
rect 3926 325 3960 359
rect 3994 325 4028 359
rect 4062 325 4096 359
rect 4130 325 4164 359
rect 4198 325 4232 359
rect 4266 325 4300 359
rect 4334 325 4368 359
rect 4402 325 4436 359
rect 4470 325 4504 359
rect 4538 325 4572 359
rect 4606 325 4640 359
rect 4674 325 4708 359
rect 4742 325 4776 359
rect 4810 325 4844 359
rect 4878 325 4912 359
rect 4946 325 4980 359
rect 5014 325 5048 359
rect 5082 325 5116 359
rect 5150 325 5184 359
rect 5218 325 5252 359
rect 5286 325 5320 359
rect 5354 325 5388 359
rect 5422 325 5456 359
rect 5490 325 5524 359
rect 5558 325 5592 359
rect 5626 325 5660 359
rect 5694 325 5728 359
rect 5762 325 5796 359
rect 5830 325 5864 359
rect 5898 325 5932 359
rect 5966 325 6000 359
rect 6034 325 6068 359
rect 6102 325 6136 359
rect 6170 325 6204 359
rect 6238 325 6272 359
rect 6306 325 6340 359
rect 6374 325 6408 359
rect 6442 325 6476 359
rect 6510 325 6544 359
rect 6578 325 6612 359
rect 6646 325 6720 359
rect 2192 322 6720 325
rect 7196 1377 11718 1380
rect 7196 1343 7264 1377
rect 7298 1343 7332 1377
rect 7366 1343 7400 1377
rect 7434 1343 7468 1377
rect 7502 1343 7536 1377
rect 7570 1343 7604 1377
rect 7638 1343 7672 1377
rect 7706 1343 7740 1377
rect 7774 1343 7808 1377
rect 7842 1343 7876 1377
rect 7910 1343 7944 1377
rect 7978 1343 8012 1377
rect 8046 1343 8080 1377
rect 8114 1343 8148 1377
rect 8182 1343 8216 1377
rect 8250 1343 8284 1377
rect 8318 1343 8352 1377
rect 8386 1343 8420 1377
rect 8454 1343 8488 1377
rect 8522 1343 8556 1377
rect 8590 1343 8624 1377
rect 8658 1343 8692 1377
rect 8726 1343 8760 1377
rect 8794 1343 8828 1377
rect 8862 1343 8896 1377
rect 8930 1343 8964 1377
rect 8998 1343 9032 1377
rect 9066 1343 9100 1377
rect 9134 1343 9168 1377
rect 9202 1343 9236 1377
rect 9270 1343 9304 1377
rect 9338 1343 9372 1377
rect 9406 1343 9500 1377
rect 9534 1343 9568 1377
rect 9602 1343 9636 1377
rect 9670 1343 9704 1377
rect 9738 1343 9772 1377
rect 9806 1343 9840 1377
rect 9874 1343 9908 1377
rect 9942 1343 9976 1377
rect 10010 1343 10044 1377
rect 10078 1343 10112 1377
rect 10146 1343 10180 1377
rect 10214 1343 10248 1377
rect 10282 1343 10316 1377
rect 10350 1343 10384 1377
rect 10418 1343 10452 1377
rect 10486 1343 10520 1377
rect 10554 1343 10588 1377
rect 10622 1343 10656 1377
rect 10690 1343 10724 1377
rect 10758 1343 10792 1377
rect 10826 1343 10860 1377
rect 10894 1343 10928 1377
rect 10962 1343 10996 1377
rect 11030 1343 11064 1377
rect 11098 1343 11132 1377
rect 11166 1343 11200 1377
rect 11234 1343 11268 1377
rect 11302 1343 11336 1377
rect 11370 1343 11404 1377
rect 11438 1343 11472 1377
rect 11506 1343 11540 1377
rect 11574 1343 11608 1377
rect 11642 1343 11718 1377
rect 7196 1340 11718 1343
rect 7196 1308 7236 1340
rect 7196 1274 7199 1308
rect 7233 1274 7236 1308
rect 7196 1240 7236 1274
rect 11678 1312 11718 1340
rect 11678 1278 11681 1312
rect 11715 1278 11718 1312
rect 7196 1206 7199 1240
rect 7233 1206 7236 1240
rect 11678 1244 11718 1278
rect 7196 1172 7236 1206
rect 7196 1138 7199 1172
rect 7233 1138 7236 1172
rect 7196 1104 7236 1138
rect 7196 1070 7199 1104
rect 7233 1070 7236 1104
rect 7196 1036 7236 1070
rect 7196 1002 7199 1036
rect 7233 1002 7236 1036
rect 7196 968 7236 1002
rect 7196 934 7199 968
rect 7233 934 7236 968
rect 7196 900 7236 934
rect 7196 866 7199 900
rect 7233 866 7236 900
rect 7196 832 7236 866
rect 7196 798 7199 832
rect 7233 798 7236 832
rect 7196 764 7236 798
rect 7196 730 7199 764
rect 7233 730 7236 764
rect 7196 696 7236 730
rect 7196 662 7199 696
rect 7233 662 7236 696
rect 7196 628 7236 662
rect 7196 594 7199 628
rect 7233 594 7236 628
rect 7196 560 7236 594
rect 7196 526 7199 560
rect 7233 526 7236 560
rect 7196 492 7236 526
rect 7196 458 7199 492
rect 7233 458 7236 492
rect 11678 1210 11681 1244
rect 11715 1210 11718 1244
rect 11678 1176 11718 1210
rect 11678 1142 11681 1176
rect 11715 1142 11718 1176
rect 11678 1108 11718 1142
rect 11678 1074 11681 1108
rect 11715 1074 11718 1108
rect 11678 1040 11718 1074
rect 11678 1006 11681 1040
rect 11715 1006 11718 1040
rect 11678 972 11718 1006
rect 11678 938 11681 972
rect 11715 938 11718 972
rect 11678 904 11718 938
rect 11678 870 11681 904
rect 11715 870 11718 904
rect 11678 836 11718 870
rect 11678 802 11681 836
rect 11715 802 11718 836
rect 11678 768 11718 802
rect 11678 734 11681 768
rect 11715 734 11718 768
rect 11678 700 11718 734
rect 11678 666 11681 700
rect 11715 666 11718 700
rect 11678 632 11718 666
rect 11678 598 11681 632
rect 11715 598 11718 632
rect 11678 564 11718 598
rect 11678 530 11681 564
rect 11715 530 11718 564
rect 11678 496 11718 530
rect 7196 424 7236 458
rect 11678 462 11681 496
rect 11715 462 11718 496
rect 7196 390 7199 424
rect 7233 390 7236 424
rect 7196 362 7236 390
rect 11678 428 11718 462
rect 11678 394 11681 428
rect 11715 394 11718 428
rect 11678 362 11718 394
rect 7196 359 11718 362
rect 7196 325 7264 359
rect 7298 325 7332 359
rect 7366 325 7400 359
rect 7434 325 7468 359
rect 7502 325 7536 359
rect 7570 325 7604 359
rect 7638 325 7672 359
rect 7706 325 7740 359
rect 7774 325 7808 359
rect 7842 325 7876 359
rect 7910 325 7944 359
rect 7978 325 8012 359
rect 8046 325 8080 359
rect 8114 325 8148 359
rect 8182 325 8216 359
rect 8250 325 8284 359
rect 8318 325 8352 359
rect 8386 325 8420 359
rect 8454 325 8488 359
rect 8522 325 8556 359
rect 8590 325 8624 359
rect 8658 325 8692 359
rect 8726 325 8760 359
rect 8794 325 8828 359
rect 8862 325 8896 359
rect 8930 325 8964 359
rect 8998 325 9032 359
rect 9066 325 9100 359
rect 9134 325 9168 359
rect 9202 325 9236 359
rect 9270 325 9304 359
rect 9338 325 9372 359
rect 9406 325 9440 359
rect 9474 325 9508 359
rect 9542 325 9576 359
rect 9610 325 9644 359
rect 9678 325 9712 359
rect 9746 325 9780 359
rect 9814 325 9848 359
rect 9882 325 9916 359
rect 9950 325 9984 359
rect 10018 325 10052 359
rect 10086 325 10120 359
rect 10154 325 10188 359
rect 10222 325 10256 359
rect 10290 325 10324 359
rect 10358 325 10392 359
rect 10426 325 10460 359
rect 10494 325 10528 359
rect 10562 325 10596 359
rect 10630 325 10664 359
rect 10698 325 10732 359
rect 10766 325 10800 359
rect 10834 325 10868 359
rect 10902 325 10936 359
rect 10970 325 11004 359
rect 11038 325 11072 359
rect 11106 325 11140 359
rect 11174 325 11208 359
rect 11242 325 11276 359
rect 11310 325 11344 359
rect 11378 325 11412 359
rect 11446 325 11480 359
rect 11514 325 11548 359
rect 11582 325 11616 359
rect 11650 325 11718 359
rect 7196 322 11718 325
<< mvnsubdiff >>
rect 63 1535 12004 1637
rect 63 1461 165 1535
rect 1906 1461 2008 1535
rect 165 135 206 169
rect 63 101 206 135
rect 63 67 138 101
rect 172 67 206 101
rect 1872 135 1906 169
rect 6884 1434 6986 1535
rect 11902 1393 12004 1535
rect 6884 169 6986 312
rect 2008 135 2103 169
rect 1872 101 2103 135
rect 1872 67 2035 101
rect 2069 67 2103 101
rect 6897 67 7020 169
rect 11814 135 11902 169
rect 11814 101 12004 135
rect 11814 67 11848 101
rect 11882 67 12004 101
rect 6417 -1188 6498 -1154
rect 6532 -1188 6566 -1154
rect 6600 -1188 6634 -1154
rect 6668 -1188 6702 -1154
rect 6736 -1188 6770 -1154
rect 6804 -1188 6838 -1154
rect 6872 -1188 6906 -1154
rect 6940 -1188 6974 -1154
rect 7008 -1188 7042 -1154
rect 7076 -1188 7110 -1154
rect 7144 -1188 7178 -1154
rect 7212 -1188 7246 -1154
rect 7280 -1188 7314 -1154
rect 7348 -1188 7382 -1154
rect 7416 -1188 7450 -1154
rect 7484 -1188 7518 -1154
rect 7552 -1188 7586 -1154
rect 7620 -1188 7654 -1154
rect 7688 -1188 7722 -1154
rect 7756 -1188 7790 -1154
rect 7824 -1188 7858 -1154
rect 7892 -1188 7926 -1154
rect 7960 -1188 7994 -1154
rect 8028 -1188 8062 -1154
rect 8096 -1188 8130 -1154
rect 8164 -1188 8198 -1154
rect 8232 -1188 8266 -1154
rect 8300 -1188 8334 -1154
rect 8368 -1188 8402 -1154
rect 8436 -1188 8470 -1154
rect 8504 -1188 8538 -1154
rect 8572 -1188 8606 -1154
rect 8640 -1188 8674 -1154
rect 8708 -1188 8776 -1154
rect 6417 -1222 6451 -1188
rect 6417 -1290 6451 -1256
rect 8742 -1262 8776 -1188
rect 6417 -1358 6451 -1324
rect 6417 -1426 6451 -1392
rect 6417 -1494 6451 -1460
rect 6417 -1562 6451 -1528
rect 6417 -1724 6451 -1596
rect 6417 -1792 6451 -1758
rect 6417 -1860 6451 -1826
rect 8742 -1330 8776 -1296
rect 8742 -1398 8776 -1364
rect 8742 -1466 8776 -1432
rect 8742 -1534 8776 -1500
rect 8742 -1602 8776 -1568
rect 8742 -1670 8776 -1636
rect 8742 -1738 8776 -1704
rect 8742 -1806 8776 -1772
rect 8742 -1874 8776 -1840
rect 6417 -1928 6451 -1894
rect 6417 -2010 6451 -1962
rect 8742 -1942 8776 -1908
rect 8742 -2010 8776 -1976
rect 6417 -2044 6485 -2010
rect 6519 -2044 6553 -2010
rect 6587 -2044 6621 -2010
rect 6655 -2044 6689 -2010
rect 6723 -2044 6757 -2010
rect 6791 -2044 6825 -2010
rect 6859 -2044 6893 -2010
rect 6927 -2044 6961 -2010
rect 6995 -2044 7029 -2010
rect 7063 -2044 7097 -2010
rect 7131 -2044 7165 -2010
rect 7199 -2044 7233 -2010
rect 7267 -2044 7301 -2010
rect 7335 -2044 7369 -2010
rect 7403 -2044 7437 -2010
rect 7471 -2044 7505 -2010
rect 7539 -2044 7573 -2010
rect 7607 -2044 7641 -2010
rect 7675 -2044 7709 -2010
rect 7743 -2044 7777 -2010
rect 7811 -2044 7845 -2010
rect 7879 -2044 7913 -2010
rect 7947 -2044 7981 -2010
rect 8015 -2044 8049 -2010
rect 8083 -2044 8117 -2010
rect 8151 -2044 8185 -2010
rect 8219 -2044 8253 -2010
rect 8287 -2044 8321 -2010
rect 8355 -2044 8389 -2010
rect 8423 -2044 8457 -2010
rect 8491 -2044 8525 -2010
rect 8559 -2044 8593 -2010
rect 8627 -2044 8661 -2010
rect 8695 -2044 8776 -2010
<< mvpsubdiffcont >>
rect 458 1317 492 1351
rect 526 1317 560 1351
rect 594 1317 628 1351
rect 662 1317 696 1351
rect 730 1317 764 1351
rect 798 1317 832 1351
rect 866 1317 900 1351
rect 934 1317 968 1351
rect 1002 1317 1036 1351
rect 1131 1317 1165 1351
rect 1199 1317 1233 1351
rect 1267 1317 1301 1351
rect 1335 1317 1369 1351
rect 1403 1317 1437 1351
rect 1471 1317 1505 1351
rect 1539 1317 1573 1351
rect 1607 1317 1641 1351
rect 360 1252 394 1286
rect 360 1184 394 1218
rect 1672 1206 1706 1240
rect 360 1116 394 1150
rect 360 1048 394 1082
rect 360 980 394 1014
rect 360 912 394 946
rect 360 844 394 878
rect 360 776 394 810
rect 360 708 394 742
rect 360 640 394 674
rect 360 572 394 606
rect 360 504 394 538
rect 1672 1138 1706 1172
rect 1672 1070 1706 1104
rect 1672 1002 1706 1036
rect 1672 934 1706 968
rect 1672 866 1706 900
rect 1672 798 1706 832
rect 1672 730 1706 764
rect 1672 662 1706 696
rect 1672 594 1706 628
rect 1672 526 1706 560
rect 360 436 394 470
rect 1672 458 1706 492
rect 1672 390 1706 424
rect 425 325 459 359
rect 493 325 527 359
rect 561 325 595 359
rect 629 325 663 359
rect 697 325 731 359
rect 765 325 799 359
rect 833 325 867 359
rect 901 325 935 359
rect 969 325 1003 359
rect 1037 325 1071 359
rect 1105 325 1139 359
rect 1173 325 1207 359
rect 1241 325 1275 359
rect 1309 325 1343 359
rect 1377 325 1411 359
rect 1445 325 1479 359
rect 1513 325 1547 359
rect 1581 325 1615 359
rect 2287 1343 2321 1377
rect 2355 1343 2389 1377
rect 2423 1343 2457 1377
rect 2491 1343 2525 1377
rect 2559 1343 2593 1377
rect 2627 1343 2661 1377
rect 2695 1343 2729 1377
rect 2763 1343 2797 1377
rect 2831 1343 2865 1377
rect 2899 1343 2933 1377
rect 2967 1343 3001 1377
rect 3035 1343 3069 1377
rect 3103 1343 3137 1377
rect 3171 1343 3205 1377
rect 3239 1343 3273 1377
rect 3307 1343 3341 1377
rect 3375 1343 3409 1377
rect 3443 1343 3477 1377
rect 3511 1343 3545 1377
rect 3579 1343 3613 1377
rect 3647 1343 3681 1377
rect 3715 1343 3749 1377
rect 3783 1343 3817 1377
rect 3851 1343 3885 1377
rect 3919 1343 3953 1377
rect 3987 1343 4021 1377
rect 4055 1343 4089 1377
rect 4123 1343 4157 1377
rect 4191 1343 4225 1377
rect 4259 1343 4293 1377
rect 4327 1343 4361 1377
rect 4395 1343 4429 1377
rect 4510 1343 4544 1377
rect 4578 1343 4612 1377
rect 4646 1343 4680 1377
rect 4714 1343 4748 1377
rect 4782 1343 4816 1377
rect 4850 1343 4884 1377
rect 4918 1343 4952 1377
rect 4986 1343 5020 1377
rect 5054 1343 5088 1377
rect 5122 1343 5156 1377
rect 5190 1343 5224 1377
rect 5258 1343 5292 1377
rect 5326 1343 5360 1377
rect 5394 1343 5428 1377
rect 5462 1343 5496 1377
rect 5530 1343 5564 1377
rect 5598 1343 5632 1377
rect 5666 1343 5700 1377
rect 5734 1343 5768 1377
rect 5802 1343 5836 1377
rect 5870 1343 5904 1377
rect 5938 1343 5972 1377
rect 6006 1343 6040 1377
rect 6074 1343 6108 1377
rect 6142 1343 6176 1377
rect 6210 1343 6244 1377
rect 6278 1343 6312 1377
rect 6346 1343 6380 1377
rect 6414 1343 6448 1377
rect 6482 1343 6516 1377
rect 6550 1343 6584 1377
rect 6618 1343 6652 1377
rect 2195 1278 2229 1312
rect 6683 1274 6717 1308
rect 2195 1210 2229 1244
rect 2195 1142 2229 1176
rect 2195 1074 2229 1108
rect 2195 1006 2229 1040
rect 2195 938 2229 972
rect 2195 870 2229 904
rect 2195 802 2229 836
rect 2195 734 2229 768
rect 2195 666 2229 700
rect 2195 598 2229 632
rect 2195 530 2229 564
rect 2195 462 2229 496
rect 6683 1206 6717 1240
rect 6683 1138 6717 1172
rect 6683 1070 6717 1104
rect 6683 1002 6717 1036
rect 6683 934 6717 968
rect 6683 866 6717 900
rect 6683 798 6717 832
rect 6683 730 6717 764
rect 6683 662 6717 696
rect 6683 594 6717 628
rect 6683 526 6717 560
rect 6683 458 6717 492
rect 2195 394 2229 428
rect 6683 390 6717 424
rect 2260 325 2294 359
rect 2328 325 2362 359
rect 2396 325 2430 359
rect 2464 325 2498 359
rect 2532 325 2566 359
rect 2600 325 2634 359
rect 2668 325 2702 359
rect 2736 325 2770 359
rect 2804 325 2838 359
rect 2872 325 2906 359
rect 2940 325 2974 359
rect 3008 325 3042 359
rect 3076 325 3110 359
rect 3144 325 3178 359
rect 3212 325 3246 359
rect 3280 325 3314 359
rect 3348 325 3382 359
rect 3416 325 3450 359
rect 3484 325 3518 359
rect 3552 325 3586 359
rect 3620 325 3654 359
rect 3688 325 3722 359
rect 3756 325 3790 359
rect 3824 325 3858 359
rect 3892 325 3926 359
rect 3960 325 3994 359
rect 4028 325 4062 359
rect 4096 325 4130 359
rect 4164 325 4198 359
rect 4232 325 4266 359
rect 4300 325 4334 359
rect 4368 325 4402 359
rect 4436 325 4470 359
rect 4504 325 4538 359
rect 4572 325 4606 359
rect 4640 325 4674 359
rect 4708 325 4742 359
rect 4776 325 4810 359
rect 4844 325 4878 359
rect 4912 325 4946 359
rect 4980 325 5014 359
rect 5048 325 5082 359
rect 5116 325 5150 359
rect 5184 325 5218 359
rect 5252 325 5286 359
rect 5320 325 5354 359
rect 5388 325 5422 359
rect 5456 325 5490 359
rect 5524 325 5558 359
rect 5592 325 5626 359
rect 5660 325 5694 359
rect 5728 325 5762 359
rect 5796 325 5830 359
rect 5864 325 5898 359
rect 5932 325 5966 359
rect 6000 325 6034 359
rect 6068 325 6102 359
rect 6136 325 6170 359
rect 6204 325 6238 359
rect 6272 325 6306 359
rect 6340 325 6374 359
rect 6408 325 6442 359
rect 6476 325 6510 359
rect 6544 325 6578 359
rect 6612 325 6646 359
rect 7264 1343 7298 1377
rect 7332 1343 7366 1377
rect 7400 1343 7434 1377
rect 7468 1343 7502 1377
rect 7536 1343 7570 1377
rect 7604 1343 7638 1377
rect 7672 1343 7706 1377
rect 7740 1343 7774 1377
rect 7808 1343 7842 1377
rect 7876 1343 7910 1377
rect 7944 1343 7978 1377
rect 8012 1343 8046 1377
rect 8080 1343 8114 1377
rect 8148 1343 8182 1377
rect 8216 1343 8250 1377
rect 8284 1343 8318 1377
rect 8352 1343 8386 1377
rect 8420 1343 8454 1377
rect 8488 1343 8522 1377
rect 8556 1343 8590 1377
rect 8624 1343 8658 1377
rect 8692 1343 8726 1377
rect 8760 1343 8794 1377
rect 8828 1343 8862 1377
rect 8896 1343 8930 1377
rect 8964 1343 8998 1377
rect 9032 1343 9066 1377
rect 9100 1343 9134 1377
rect 9168 1343 9202 1377
rect 9236 1343 9270 1377
rect 9304 1343 9338 1377
rect 9372 1343 9406 1377
rect 9500 1343 9534 1377
rect 9568 1343 9602 1377
rect 9636 1343 9670 1377
rect 9704 1343 9738 1377
rect 9772 1343 9806 1377
rect 9840 1343 9874 1377
rect 9908 1343 9942 1377
rect 9976 1343 10010 1377
rect 10044 1343 10078 1377
rect 10112 1343 10146 1377
rect 10180 1343 10214 1377
rect 10248 1343 10282 1377
rect 10316 1343 10350 1377
rect 10384 1343 10418 1377
rect 10452 1343 10486 1377
rect 10520 1343 10554 1377
rect 10588 1343 10622 1377
rect 10656 1343 10690 1377
rect 10724 1343 10758 1377
rect 10792 1343 10826 1377
rect 10860 1343 10894 1377
rect 10928 1343 10962 1377
rect 10996 1343 11030 1377
rect 11064 1343 11098 1377
rect 11132 1343 11166 1377
rect 11200 1343 11234 1377
rect 11268 1343 11302 1377
rect 11336 1343 11370 1377
rect 11404 1343 11438 1377
rect 11472 1343 11506 1377
rect 11540 1343 11574 1377
rect 11608 1343 11642 1377
rect 7199 1274 7233 1308
rect 11681 1278 11715 1312
rect 7199 1206 7233 1240
rect 7199 1138 7233 1172
rect 7199 1070 7233 1104
rect 7199 1002 7233 1036
rect 7199 934 7233 968
rect 7199 866 7233 900
rect 7199 798 7233 832
rect 7199 730 7233 764
rect 7199 662 7233 696
rect 7199 594 7233 628
rect 7199 526 7233 560
rect 7199 458 7233 492
rect 11681 1210 11715 1244
rect 11681 1142 11715 1176
rect 11681 1074 11715 1108
rect 11681 1006 11715 1040
rect 11681 938 11715 972
rect 11681 870 11715 904
rect 11681 802 11715 836
rect 11681 734 11715 768
rect 11681 666 11715 700
rect 11681 598 11715 632
rect 11681 530 11715 564
rect 11681 462 11715 496
rect 7199 390 7233 424
rect 11681 394 11715 428
rect 7264 325 7298 359
rect 7332 325 7366 359
rect 7400 325 7434 359
rect 7468 325 7502 359
rect 7536 325 7570 359
rect 7604 325 7638 359
rect 7672 325 7706 359
rect 7740 325 7774 359
rect 7808 325 7842 359
rect 7876 325 7910 359
rect 7944 325 7978 359
rect 8012 325 8046 359
rect 8080 325 8114 359
rect 8148 325 8182 359
rect 8216 325 8250 359
rect 8284 325 8318 359
rect 8352 325 8386 359
rect 8420 325 8454 359
rect 8488 325 8522 359
rect 8556 325 8590 359
rect 8624 325 8658 359
rect 8692 325 8726 359
rect 8760 325 8794 359
rect 8828 325 8862 359
rect 8896 325 8930 359
rect 8964 325 8998 359
rect 9032 325 9066 359
rect 9100 325 9134 359
rect 9168 325 9202 359
rect 9236 325 9270 359
rect 9304 325 9338 359
rect 9372 325 9406 359
rect 9440 325 9474 359
rect 9508 325 9542 359
rect 9576 325 9610 359
rect 9644 325 9678 359
rect 9712 325 9746 359
rect 9780 325 9814 359
rect 9848 325 9882 359
rect 9916 325 9950 359
rect 9984 325 10018 359
rect 10052 325 10086 359
rect 10120 325 10154 359
rect 10188 325 10222 359
rect 10256 325 10290 359
rect 10324 325 10358 359
rect 10392 325 10426 359
rect 10460 325 10494 359
rect 10528 325 10562 359
rect 10596 325 10630 359
rect 10664 325 10698 359
rect 10732 325 10766 359
rect 10800 325 10834 359
rect 10868 325 10902 359
rect 10936 325 10970 359
rect 11004 325 11038 359
rect 11072 325 11106 359
rect 11140 325 11174 359
rect 11208 325 11242 359
rect 11276 325 11310 359
rect 11344 325 11378 359
rect 11412 325 11446 359
rect 11480 325 11514 359
rect 11548 325 11582 359
rect 11616 325 11650 359
<< mvnsubdiffcont >>
rect 63 135 165 1461
rect 138 67 172 101
rect 206 67 1872 169
rect 1906 135 2008 1461
rect 6884 312 6986 1434
rect 2035 67 2069 101
rect 2103 67 6897 169
rect 7020 67 11814 169
rect 11902 135 12004 1393
rect 11848 67 11882 101
rect 6498 -1188 6532 -1154
rect 6566 -1188 6600 -1154
rect 6634 -1188 6668 -1154
rect 6702 -1188 6736 -1154
rect 6770 -1188 6804 -1154
rect 6838 -1188 6872 -1154
rect 6906 -1188 6940 -1154
rect 6974 -1188 7008 -1154
rect 7042 -1188 7076 -1154
rect 7110 -1188 7144 -1154
rect 7178 -1188 7212 -1154
rect 7246 -1188 7280 -1154
rect 7314 -1188 7348 -1154
rect 7382 -1188 7416 -1154
rect 7450 -1188 7484 -1154
rect 7518 -1188 7552 -1154
rect 7586 -1188 7620 -1154
rect 7654 -1188 7688 -1154
rect 7722 -1188 7756 -1154
rect 7790 -1188 7824 -1154
rect 7858 -1188 7892 -1154
rect 7926 -1188 7960 -1154
rect 7994 -1188 8028 -1154
rect 8062 -1188 8096 -1154
rect 8130 -1188 8164 -1154
rect 8198 -1188 8232 -1154
rect 8266 -1188 8300 -1154
rect 8334 -1188 8368 -1154
rect 8402 -1188 8436 -1154
rect 8470 -1188 8504 -1154
rect 8538 -1188 8572 -1154
rect 8606 -1188 8640 -1154
rect 8674 -1188 8708 -1154
rect 6417 -1256 6451 -1222
rect 6417 -1324 6451 -1290
rect 8742 -1296 8776 -1262
rect 6417 -1392 6451 -1358
rect 6417 -1460 6451 -1426
rect 6417 -1528 6451 -1494
rect 6417 -1596 6451 -1562
rect 6417 -1758 6451 -1724
rect 6417 -1826 6451 -1792
rect 6417 -1894 6451 -1860
rect 8742 -1364 8776 -1330
rect 8742 -1432 8776 -1398
rect 8742 -1500 8776 -1466
rect 8742 -1568 8776 -1534
rect 8742 -1636 8776 -1602
rect 8742 -1704 8776 -1670
rect 8742 -1772 8776 -1738
rect 8742 -1840 8776 -1806
rect 6417 -1962 6451 -1928
rect 8742 -1908 8776 -1874
rect 8742 -1976 8776 -1942
rect 6485 -2044 6519 -2010
rect 6553 -2044 6587 -2010
rect 6621 -2044 6655 -2010
rect 6689 -2044 6723 -2010
rect 6757 -2044 6791 -2010
rect 6825 -2044 6859 -2010
rect 6893 -2044 6927 -2010
rect 6961 -2044 6995 -2010
rect 7029 -2044 7063 -2010
rect 7097 -2044 7131 -2010
rect 7165 -2044 7199 -2010
rect 7233 -2044 7267 -2010
rect 7301 -2044 7335 -2010
rect 7369 -2044 7403 -2010
rect 7437 -2044 7471 -2010
rect 7505 -2044 7539 -2010
rect 7573 -2044 7607 -2010
rect 7641 -2044 7675 -2010
rect 7709 -2044 7743 -2010
rect 7777 -2044 7811 -2010
rect 7845 -2044 7879 -2010
rect 7913 -2044 7947 -2010
rect 7981 -2044 8015 -2010
rect 8049 -2044 8083 -2010
rect 8117 -2044 8151 -2010
rect 8185 -2044 8219 -2010
rect 8253 -2044 8287 -2010
rect 8321 -2044 8355 -2010
rect 8389 -2044 8423 -2010
rect 8457 -2044 8491 -2010
rect 8525 -2044 8559 -2010
rect 8593 -2044 8627 -2010
rect 8661 -2044 8695 -2010
<< poly >>
rect 460 1171 558 1187
rect 460 1137 476 1171
rect 510 1137 558 1171
rect 460 1101 558 1137
rect 460 1067 476 1101
rect 510 1087 558 1101
rect 1558 1087 1590 1187
rect 510 1067 526 1087
rect 460 1031 526 1067
rect 460 997 476 1031
rect 510 997 558 1031
rect 460 961 558 997
rect 460 927 476 961
rect 510 931 558 961
rect 1558 931 1590 1031
rect 510 927 526 931
rect 460 891 526 927
rect 460 857 476 891
rect 510 857 526 891
rect 460 821 526 857
rect 460 787 476 821
rect 510 787 526 821
rect 460 751 526 787
rect 460 717 476 751
rect 510 745 526 751
rect 510 717 558 745
rect 460 681 558 717
rect 460 647 476 681
rect 510 647 558 681
rect 460 645 558 647
rect 1558 645 1590 745
rect 460 610 526 645
rect 460 576 476 610
rect 510 589 526 610
rect 510 576 558 589
rect 460 539 558 576
rect 460 505 476 539
rect 510 505 558 539
rect 460 489 558 505
rect 1558 489 1590 589
rect 2295 1197 2393 1213
rect 2295 1163 2311 1197
rect 2345 1163 2393 1197
rect 2295 1124 2393 1163
rect 2295 1090 2311 1124
rect 2345 1113 2393 1124
rect 4393 1113 4425 1213
rect 4467 1113 4499 1213
rect 6499 1197 6597 1213
rect 6499 1163 6547 1197
rect 6581 1163 6597 1197
rect 6499 1124 6597 1163
rect 6499 1113 6547 1124
rect 2345 1090 2361 1113
rect 2295 1057 2361 1090
rect 6531 1090 6547 1113
rect 6581 1090 6597 1124
rect 6531 1057 6597 1090
rect 2295 1051 2393 1057
rect 2295 1017 2311 1051
rect 2345 1017 2393 1051
rect 2295 978 2393 1017
rect 2295 944 2311 978
rect 2345 957 2393 978
rect 4393 957 4425 1057
rect 4467 957 4499 1057
rect 6499 1051 6597 1057
rect 6499 1017 6547 1051
rect 6581 1017 6597 1051
rect 6499 978 6597 1017
rect 6499 957 6547 978
rect 2345 944 2361 957
rect 2295 905 2361 944
rect 2295 871 2311 905
rect 2345 901 2361 905
rect 6531 944 6547 957
rect 6581 944 6597 978
rect 6531 905 6597 944
rect 6531 901 6547 905
rect 2345 871 2393 901
rect 2295 832 2393 871
rect 2295 798 2311 832
rect 2345 801 2393 832
rect 4393 801 4425 901
rect 4467 801 4499 901
rect 6499 871 6547 901
rect 6581 871 6597 905
rect 6499 832 6597 871
rect 6499 801 6547 832
rect 2345 798 2361 801
rect 2295 759 2361 798
rect 2295 725 2311 759
rect 2345 745 2361 759
rect 6531 798 6547 801
rect 6581 798 6597 832
rect 6531 759 6597 798
rect 6531 745 6547 759
rect 2345 725 2393 745
rect 2295 686 2393 725
rect 2295 652 2311 686
rect 2345 652 2393 686
rect 2295 645 2393 652
rect 4393 645 4425 745
rect 4467 645 4499 745
rect 6499 725 6547 745
rect 6581 725 6597 759
rect 6499 686 6597 725
rect 6499 652 6547 686
rect 6581 652 6597 686
rect 6499 645 6597 652
rect 2295 613 2361 645
rect 2295 579 2311 613
rect 2345 589 2361 613
rect 6531 613 6597 645
rect 6531 589 6547 613
rect 2345 579 2393 589
rect 2295 539 2393 579
rect 2295 505 2311 539
rect 2345 505 2393 539
rect 2295 489 2393 505
rect 4393 489 4425 589
rect 4467 489 4499 589
rect 6499 579 6547 589
rect 6581 579 6597 613
rect 6499 539 6597 579
rect 6499 505 6547 539
rect 6581 505 6597 539
rect 6499 489 6597 505
rect 7314 1197 7412 1213
rect 7314 1163 7330 1197
rect 7364 1163 7412 1197
rect 7314 1123 7412 1163
rect 7314 1089 7330 1123
rect 7364 1113 7412 1123
rect 9412 1113 9444 1213
rect 9486 1113 9518 1213
rect 11518 1197 11615 1213
rect 11518 1163 11565 1197
rect 11599 1163 11615 1197
rect 11518 1123 11615 1163
rect 11518 1113 11565 1123
rect 7364 1089 7380 1113
rect 7314 1057 7380 1089
rect 11549 1089 11565 1113
rect 11599 1089 11615 1123
rect 11549 1057 11615 1089
rect 7314 1050 7412 1057
rect 7314 1016 7330 1050
rect 7364 1016 7412 1050
rect 7314 977 7412 1016
rect 7314 943 7330 977
rect 7364 957 7412 977
rect 9412 957 9444 1057
rect 9486 957 9518 1057
rect 11518 1050 11615 1057
rect 11518 1016 11565 1050
rect 11599 1016 11615 1050
rect 11518 977 11615 1016
rect 11518 957 11565 977
rect 7364 943 7380 957
rect 7314 904 7380 943
rect 7314 870 7330 904
rect 7364 901 7380 904
rect 11549 943 11565 957
rect 11599 943 11615 977
rect 11549 904 11615 943
rect 11549 901 11565 904
rect 7364 870 7412 901
rect 7314 831 7412 870
rect 7314 797 7330 831
rect 7364 801 7412 831
rect 9412 801 9444 901
rect 9486 801 9518 901
rect 11518 870 11565 901
rect 11599 870 11615 904
rect 11518 831 11615 870
rect 11518 801 11565 831
rect 7364 797 7380 801
rect 7314 758 7380 797
rect 7314 724 7330 758
rect 7364 745 7380 758
rect 11549 797 11565 801
rect 11599 797 11615 831
rect 11549 758 11615 797
rect 11549 745 11565 758
rect 7364 724 7412 745
rect 7314 685 7412 724
rect 7314 651 7330 685
rect 7364 651 7412 685
rect 7314 645 7412 651
rect 9412 645 9444 745
rect 9486 645 9518 745
rect 11518 724 11565 745
rect 11599 724 11615 758
rect 11518 685 11615 724
rect 11518 651 11565 685
rect 11599 651 11615 685
rect 11518 645 11615 651
rect 7314 612 7380 645
rect 7314 578 7330 612
rect 7364 589 7380 612
rect 11549 612 11615 645
rect 11549 589 11565 612
rect 7364 578 7412 589
rect 7314 539 7412 578
rect 7314 505 7330 539
rect 7364 505 7412 539
rect 7314 489 7412 505
rect 9412 489 9444 589
rect 9486 489 9518 589
rect 11518 578 11565 589
rect 11599 578 11615 612
rect 11518 539 11615 578
rect 11518 505 11565 539
rect 11599 505 11615 539
rect 11518 489 11615 505
rect 6518 -1331 6616 -1315
rect 6518 -1365 6534 -1331
rect 6568 -1365 6616 -1331
rect 6518 -1402 6616 -1365
rect 6518 -1436 6534 -1402
rect 6568 -1415 6616 -1402
rect 8616 -1415 8648 -1315
rect 6568 -1436 6584 -1415
rect 6518 -1471 6584 -1436
rect 6518 -1473 6616 -1471
rect 6518 -1507 6534 -1473
rect 6568 -1507 6616 -1473
rect 6518 -1545 6616 -1507
rect 6518 -1579 6534 -1545
rect 6568 -1571 6616 -1545
rect 8616 -1571 8648 -1471
rect 6568 -1579 6584 -1571
rect 6518 -1617 6584 -1579
rect 6518 -1651 6534 -1617
rect 6568 -1627 6584 -1617
rect 6568 -1651 6616 -1627
rect 6518 -1689 6616 -1651
rect 6518 -1723 6534 -1689
rect 6568 -1723 6616 -1689
rect 6518 -1727 6616 -1723
rect 8616 -1727 8648 -1627
rect 6518 -1761 6584 -1727
rect 6518 -1795 6534 -1761
rect 6568 -1783 6584 -1761
rect 6568 -1795 6616 -1783
rect 6518 -1833 6616 -1795
rect 6518 -1867 6534 -1833
rect 6568 -1867 6616 -1833
rect 6518 -1883 6616 -1867
rect 8616 -1883 8648 -1783
<< polycont >>
rect 476 1137 510 1171
rect 476 1067 510 1101
rect 476 997 510 1031
rect 476 927 510 961
rect 476 857 510 891
rect 476 787 510 821
rect 476 717 510 751
rect 476 647 510 681
rect 476 576 510 610
rect 476 505 510 539
rect 2311 1163 2345 1197
rect 2311 1090 2345 1124
rect 6547 1163 6581 1197
rect 6547 1090 6581 1124
rect 2311 1017 2345 1051
rect 2311 944 2345 978
rect 6547 1017 6581 1051
rect 2311 871 2345 905
rect 6547 944 6581 978
rect 2311 798 2345 832
rect 6547 871 6581 905
rect 2311 725 2345 759
rect 6547 798 6581 832
rect 2311 652 2345 686
rect 6547 725 6581 759
rect 6547 652 6581 686
rect 2311 579 2345 613
rect 2311 505 2345 539
rect 6547 579 6581 613
rect 6547 505 6581 539
rect 7330 1163 7364 1197
rect 7330 1089 7364 1123
rect 11565 1163 11599 1197
rect 11565 1089 11599 1123
rect 7330 1016 7364 1050
rect 7330 943 7364 977
rect 11565 1016 11599 1050
rect 7330 870 7364 904
rect 11565 943 11599 977
rect 7330 797 7364 831
rect 11565 870 11599 904
rect 7330 724 7364 758
rect 11565 797 11599 831
rect 7330 651 7364 685
rect 11565 724 11599 758
rect 11565 651 11599 685
rect 7330 578 7364 612
rect 7330 505 7364 539
rect 11565 578 11599 612
rect 11565 505 11599 539
rect 6534 -1365 6568 -1331
rect 6534 -1436 6568 -1402
rect 6534 -1507 6568 -1473
rect 6534 -1579 6568 -1545
rect 6534 -1651 6568 -1617
rect 6534 -1723 6568 -1689
rect 6534 -1795 6568 -1761
rect 6534 -1867 6568 -1833
<< locali >>
rect 63 1535 12004 1637
rect 63 1461 165 1535
rect -462 1395 -409 1429
rect -375 1395 -322 1429
rect -288 1395 -236 1429
rect -202 1395 -150 1429
rect -496 1319 -116 1395
rect -462 1285 -409 1319
rect -375 1285 -322 1319
rect -288 1285 -236 1319
rect -202 1285 -150 1319
rect 55 1412 63 1444
rect 1906 1461 2008 1535
rect 165 1412 173 1444
rect 55 1378 61 1412
rect 167 1378 173 1412
rect 55 1339 63 1378
rect 165 1339 173 1378
rect 55 1305 61 1339
rect 167 1305 173 1339
rect 55 1266 63 1305
rect 165 1266 173 1305
rect 55 1232 61 1266
rect 167 1232 173 1266
rect 55 1193 63 1232
rect 165 1193 173 1232
rect 55 1159 61 1193
rect 167 1159 173 1193
rect 55 1120 63 1159
rect 165 1120 173 1159
rect 55 1086 61 1120
rect 167 1086 173 1120
rect 55 1047 63 1086
rect 165 1047 173 1086
rect 55 1013 61 1047
rect 167 1013 173 1047
rect 55 974 63 1013
rect 165 974 173 1013
rect 55 940 61 974
rect 167 940 173 974
rect 55 901 63 940
rect 165 901 173 940
rect 55 867 61 901
rect 167 867 173 901
rect 55 828 63 867
rect 165 828 173 867
rect 55 794 61 828
rect 167 794 173 828
rect 55 755 63 794
rect 165 755 173 794
rect 55 721 61 755
rect 167 721 173 755
rect 55 682 63 721
rect 165 682 173 721
rect -463 623 -410 657
rect -376 623 -323 657
rect -289 623 -236 657
rect -202 623 -150 657
rect -497 579 -116 623
rect -463 545 -410 579
rect -376 545 -323 579
rect -289 545 -236 579
rect -202 545 -150 579
rect -497 501 -116 545
rect -463 467 -410 501
rect -376 467 -323 501
rect -289 467 -236 501
rect -202 467 -150 501
rect 55 648 61 682
rect 167 648 173 682
rect 55 609 63 648
rect 165 609 173 648
rect 55 575 61 609
rect 167 575 173 609
rect 55 536 63 575
rect 165 536 173 575
rect 55 502 61 536
rect 167 502 173 536
rect 55 463 63 502
rect 165 463 173 502
rect 55 429 61 463
rect 167 429 173 463
rect 55 390 63 429
rect 165 390 173 429
rect 55 356 61 390
rect 167 356 173 390
rect 55 317 63 356
rect 165 317 173 356
rect 55 283 61 317
rect 167 283 173 317
rect 318 1437 1748 1443
rect 318 1403 402 1437
rect 436 1403 480 1437
rect 514 1403 558 1437
rect 592 1403 636 1437
rect 670 1403 714 1437
rect 748 1403 792 1437
rect 826 1403 870 1437
rect 904 1403 949 1437
rect 983 1403 1059 1437
rect 318 1365 1059 1403
rect 318 1331 324 1365
rect 358 1331 396 1365
rect 430 1351 480 1365
rect 514 1351 558 1365
rect 592 1351 636 1365
rect 670 1351 714 1365
rect 748 1351 792 1365
rect 826 1351 870 1365
rect 904 1351 949 1365
rect 983 1351 1059 1365
rect 1597 1403 1636 1437
rect 1670 1403 1748 1437
rect 1597 1365 1748 1403
rect 1597 1351 1636 1365
rect 1670 1363 1748 1365
rect 430 1331 458 1351
rect 514 1331 526 1351
rect 592 1331 594 1351
rect 318 1317 458 1331
rect 492 1317 526 1331
rect 560 1317 594 1331
rect 628 1331 636 1351
rect 696 1331 714 1351
rect 764 1331 792 1351
rect 628 1317 662 1331
rect 696 1317 730 1331
rect 764 1317 798 1331
rect 832 1317 866 1351
rect 904 1331 934 1351
rect 983 1331 1002 1351
rect 900 1317 934 1331
rect 968 1317 1002 1331
rect 1036 1331 1059 1351
rect 1597 1331 1607 1351
rect 1670 1331 1708 1363
rect 1036 1317 1131 1331
rect 1165 1317 1199 1331
rect 1233 1317 1267 1331
rect 1301 1317 1335 1331
rect 1369 1317 1403 1331
rect 1437 1317 1471 1331
rect 1505 1317 1539 1331
rect 1573 1317 1607 1331
rect 1641 1329 1708 1331
rect 1742 1329 1748 1363
rect 1641 1317 1748 1329
rect 318 1314 1748 1317
rect 318 1290 436 1314
rect 318 1256 324 1290
rect 358 1286 396 1290
rect 358 1256 360 1286
rect 318 1252 360 1256
rect 394 1256 396 1286
rect 430 1256 436 1290
rect 394 1252 436 1256
rect 318 1218 436 1252
rect 1630 1289 1748 1314
rect 1630 1255 1636 1289
rect 1670 1255 1708 1289
rect 1742 1255 1748 1289
rect 1630 1240 1748 1255
rect 600 1232 641 1235
rect 675 1232 716 1235
rect 750 1232 791 1235
rect 825 1232 866 1235
rect 900 1232 940 1235
rect 974 1232 1014 1235
rect 1048 1232 1088 1235
rect 1122 1232 1162 1235
rect 1196 1232 1236 1235
rect 1270 1232 1310 1235
rect 1344 1232 1384 1235
rect 1418 1232 1458 1235
rect 318 1215 360 1218
rect 318 1181 324 1215
rect 358 1184 360 1215
rect 394 1215 436 1218
rect 394 1184 396 1215
rect 358 1181 396 1184
rect 430 1181 436 1215
rect 554 1201 566 1232
rect 554 1198 570 1201
rect 604 1198 638 1232
rect 675 1201 706 1232
rect 750 1201 774 1232
rect 825 1201 842 1232
rect 900 1201 910 1232
rect 974 1201 978 1232
rect 672 1198 706 1201
rect 740 1198 774 1201
rect 808 1198 842 1201
rect 876 1198 910 1201
rect 944 1198 978 1201
rect 1012 1201 1014 1232
rect 1080 1201 1088 1232
rect 1148 1201 1162 1232
rect 1216 1201 1236 1232
rect 1284 1201 1310 1232
rect 1352 1201 1384 1232
rect 1012 1198 1046 1201
rect 1080 1198 1114 1201
rect 1148 1198 1182 1201
rect 1216 1198 1250 1201
rect 1284 1198 1318 1201
rect 1352 1198 1386 1201
rect 1420 1198 1454 1232
rect 1492 1201 1504 1232
rect 1488 1198 1504 1201
rect 1630 1215 1672 1240
rect 318 1150 436 1181
rect 318 1140 360 1150
rect 318 1106 324 1140
rect 358 1116 360 1140
rect 394 1140 436 1150
rect 394 1116 396 1140
rect 358 1106 396 1116
rect 430 1106 436 1140
rect 318 1082 436 1106
rect 318 1065 360 1082
rect 318 1031 324 1065
rect 358 1048 360 1065
rect 394 1065 436 1082
rect 394 1048 396 1065
rect 358 1031 396 1048
rect 430 1031 436 1065
rect 318 1014 436 1031
rect 318 990 360 1014
rect 318 956 324 990
rect 358 980 360 990
rect 394 990 436 1014
rect 394 980 396 990
rect 358 956 396 980
rect 430 956 436 990
rect 318 946 436 956
rect 318 915 360 946
rect 318 881 324 915
rect 358 912 360 915
rect 394 915 436 946
rect 394 912 396 915
rect 358 881 396 912
rect 430 881 436 915
rect 318 878 436 881
rect 318 844 360 878
rect 394 844 436 878
rect 318 841 436 844
rect 318 807 324 841
rect 358 810 396 841
rect 358 807 360 810
rect 318 776 360 807
rect 394 807 396 810
rect 430 807 436 841
rect 394 776 436 807
rect 318 767 436 776
rect 318 733 324 767
rect 358 742 396 767
rect 358 733 360 742
rect 318 708 360 733
rect 394 733 396 742
rect 430 733 436 767
rect 394 708 436 733
rect 318 693 436 708
rect 318 659 324 693
rect 358 674 396 693
rect 358 659 360 674
rect 318 640 360 659
rect 394 659 396 674
rect 430 659 436 693
rect 394 640 436 659
rect 318 619 436 640
rect 318 585 324 619
rect 358 606 396 619
rect 358 585 360 606
rect 318 572 360 585
rect 394 585 396 606
rect 430 585 436 619
rect 394 572 436 585
rect 318 545 436 572
rect 318 511 324 545
rect 358 538 396 545
rect 358 511 360 538
rect 318 504 360 511
rect 394 511 396 538
rect 430 511 436 545
rect 394 504 436 511
rect 318 471 436 504
rect 476 1175 510 1187
rect 476 1102 510 1137
rect 1630 1181 1636 1215
rect 1670 1206 1672 1215
rect 1706 1215 1748 1240
rect 1706 1206 1708 1215
rect 1670 1181 1708 1206
rect 1742 1181 1748 1215
rect 1630 1172 1748 1181
rect 1630 1141 1672 1172
rect 1630 1107 1636 1141
rect 1670 1138 1672 1141
rect 1706 1141 1748 1172
rect 1706 1138 1708 1141
rect 1670 1107 1708 1138
rect 1742 1107 1748 1141
rect 1630 1104 1748 1107
rect 476 1031 510 1067
rect 554 1042 570 1076
rect 604 1042 638 1076
rect 672 1042 706 1076
rect 740 1042 774 1076
rect 808 1042 842 1076
rect 876 1042 910 1076
rect 944 1042 978 1076
rect 1012 1042 1046 1076
rect 1080 1042 1114 1076
rect 1158 1042 1182 1076
rect 1236 1042 1250 1076
rect 1314 1042 1318 1076
rect 1352 1042 1358 1076
rect 1420 1042 1435 1076
rect 1488 1042 1512 1076
rect 1630 1070 1672 1104
rect 1706 1070 1748 1104
rect 1630 1067 1748 1070
rect 476 961 510 995
rect 476 891 510 922
rect 1630 1033 1636 1067
rect 1670 1036 1708 1067
rect 1670 1033 1672 1036
rect 1630 1002 1672 1033
rect 1706 1033 1708 1036
rect 1742 1033 1748 1067
rect 1706 1002 1748 1033
rect 1630 993 1748 1002
rect 1630 959 1636 993
rect 1670 968 1708 993
rect 1670 959 1672 968
rect 1630 934 1672 959
rect 1706 959 1708 968
rect 1742 959 1748 993
rect 1706 934 1748 959
rect 600 920 641 921
rect 675 920 716 921
rect 750 920 791 921
rect 825 920 866 921
rect 900 920 940 921
rect 974 920 1014 921
rect 1048 920 1088 921
rect 1122 920 1162 921
rect 1196 920 1236 921
rect 1270 920 1310 921
rect 1344 920 1384 921
rect 1418 920 1458 921
rect 554 887 566 920
rect 554 886 570 887
rect 604 886 638 920
rect 675 887 706 920
rect 750 887 774 920
rect 825 887 842 920
rect 900 887 910 920
rect 974 887 978 920
rect 672 886 706 887
rect 740 886 774 887
rect 808 886 842 887
rect 876 886 910 887
rect 944 886 978 887
rect 1012 887 1014 920
rect 1080 887 1088 920
rect 1148 887 1162 920
rect 1216 887 1236 920
rect 1284 887 1310 920
rect 1352 887 1384 920
rect 1012 886 1046 887
rect 1080 886 1114 887
rect 1148 886 1182 887
rect 1216 886 1250 887
rect 1284 886 1318 887
rect 1352 886 1386 887
rect 1420 886 1454 920
rect 1492 887 1504 920
rect 1488 886 1504 887
rect 1630 919 1748 934
rect 476 821 510 849
rect 1630 885 1636 919
rect 1670 900 1708 919
rect 1670 885 1672 900
rect 1630 866 1672 885
rect 1706 885 1708 900
rect 1742 885 1748 919
rect 1706 866 1748 885
rect 1630 845 1748 866
rect 1630 811 1636 845
rect 1670 832 1708 845
rect 1670 811 1672 832
rect 1630 798 1672 811
rect 1706 811 1708 832
rect 1742 811 1748 845
rect 1706 798 1748 811
rect 476 751 510 776
rect 554 756 566 790
rect 604 756 638 790
rect 675 756 706 790
rect 750 756 774 790
rect 825 756 842 790
rect 900 756 910 790
rect 974 756 978 790
rect 1012 756 1014 790
rect 1080 756 1088 790
rect 1148 756 1162 790
rect 1216 756 1236 790
rect 1284 756 1310 790
rect 1352 756 1384 790
rect 1420 756 1454 790
rect 1492 756 1504 790
rect 1630 770 1748 798
rect 476 681 510 704
rect 1630 736 1636 770
rect 1670 764 1708 770
rect 1670 736 1672 764
rect 1630 730 1672 736
rect 1706 736 1708 764
rect 1742 736 1748 770
rect 1706 730 1748 736
rect 1630 696 1748 730
rect 1630 695 1672 696
rect 1630 661 1636 695
rect 1670 662 1672 695
rect 1706 695 1748 696
rect 1706 662 1708 695
rect 1670 661 1708 662
rect 1742 661 1748 695
rect 476 610 510 632
rect 554 600 570 634
rect 604 600 638 634
rect 672 600 706 634
rect 740 600 774 634
rect 808 600 842 634
rect 876 600 910 634
rect 944 600 978 634
rect 1012 600 1046 634
rect 1080 600 1114 634
rect 1157 600 1182 634
rect 1235 600 1250 634
rect 1313 600 1318 634
rect 1352 600 1357 634
rect 1420 600 1435 634
rect 1488 600 1512 634
rect 1630 628 1748 661
rect 1630 620 1672 628
rect 476 539 510 560
rect 1630 586 1636 620
rect 1670 594 1672 620
rect 1706 620 1748 628
rect 1706 594 1708 620
rect 1670 586 1708 594
rect 1742 586 1748 620
rect 1630 560 1748 586
rect 1630 545 1672 560
rect 1630 511 1636 545
rect 1670 526 1672 545
rect 1706 545 1748 560
rect 1706 526 1708 545
rect 1670 511 1708 526
rect 1742 511 1748 545
rect 1630 492 1748 511
rect 318 437 324 471
rect 358 470 396 471
rect 358 437 360 470
rect 318 436 360 437
rect 394 437 396 470
rect 430 437 436 471
rect 554 444 570 478
rect 604 444 638 478
rect 675 444 706 478
rect 750 444 774 478
rect 825 444 842 478
rect 900 444 910 478
rect 974 444 978 478
rect 1012 444 1014 478
rect 1080 444 1088 478
rect 1148 444 1162 478
rect 1216 444 1236 478
rect 1284 444 1310 478
rect 1352 444 1384 478
rect 1420 444 1454 478
rect 1492 444 1504 478
rect 1630 470 1672 492
rect 394 436 436 437
rect 318 401 436 436
rect 1630 436 1636 470
rect 1670 458 1672 470
rect 1706 470 1748 492
rect 1706 458 1708 470
rect 1670 436 1708 458
rect 1742 436 1748 470
rect 1630 424 1748 436
rect 1630 401 1672 424
rect 318 397 1672 401
rect 318 363 324 397
rect 358 395 1672 397
rect 358 363 396 395
rect 318 361 396 363
rect 430 361 469 395
rect 503 361 542 395
rect 576 361 615 395
rect 649 361 688 395
rect 722 361 761 395
rect 795 361 834 395
rect 868 361 907 395
rect 941 361 980 395
rect 1014 361 1053 395
rect 1087 361 1126 395
rect 1160 361 1199 395
rect 1233 361 1272 395
rect 1306 361 1345 395
rect 1379 361 1418 395
rect 1452 361 1491 395
rect 1525 361 1564 395
rect 318 359 1564 361
rect 1670 390 1672 395
rect 1706 395 1748 424
rect 1706 390 1708 395
rect 1670 361 1708 390
rect 1742 361 1748 395
rect 318 325 425 359
rect 459 325 493 359
rect 527 325 561 359
rect 595 325 629 359
rect 663 325 697 359
rect 731 325 765 359
rect 799 325 833 359
rect 867 325 901 359
rect 935 325 969 359
rect 1003 325 1037 359
rect 1071 325 1105 359
rect 1139 325 1173 359
rect 1207 325 1241 359
rect 1275 325 1309 359
rect 1343 325 1377 359
rect 1411 325 1445 359
rect 1479 325 1513 359
rect 1547 325 1564 359
rect 318 323 1564 325
rect 318 289 396 323
rect 430 289 469 323
rect 503 289 542 323
rect 576 289 615 323
rect 649 289 688 323
rect 722 289 761 323
rect 795 289 834 323
rect 868 289 907 323
rect 941 289 980 323
rect 1014 289 1053 323
rect 1087 289 1126 323
rect 1160 289 1199 323
rect 1233 289 1272 323
rect 1306 289 1345 323
rect 1379 289 1418 323
rect 1452 289 1491 323
rect 1525 289 1564 323
rect 1670 289 1748 361
rect 318 283 1748 289
rect 1898 1423 1906 1455
rect 6884 1456 6986 1535
rect 2008 1423 2016 1455
rect 1898 1389 1904 1423
rect 2010 1389 2016 1423
rect 1898 1349 1906 1389
rect 2008 1349 2016 1389
rect 1898 1315 1904 1349
rect 2010 1315 2016 1349
rect 1898 1275 1906 1315
rect 2008 1275 2016 1315
rect 1898 1241 1904 1275
rect 2010 1241 2016 1275
rect 1898 1201 1906 1241
rect 2008 1201 2016 1241
rect 1898 1167 1904 1201
rect 2010 1167 2016 1201
rect 1898 1127 1906 1167
rect 2008 1127 2016 1167
rect 1898 1093 1904 1127
rect 2010 1093 2016 1127
rect 1898 1053 1906 1093
rect 2008 1053 2016 1093
rect 1898 1019 1904 1053
rect 2010 1019 2016 1053
rect 1898 979 1906 1019
rect 2008 979 2016 1019
rect 1898 945 1904 979
rect 2010 945 2016 979
rect 1898 905 1906 945
rect 2008 905 2016 945
rect 1898 871 1904 905
rect 2010 871 2016 905
rect 1898 831 1906 871
rect 2008 831 2016 871
rect 1898 797 1904 831
rect 2010 797 2016 831
rect 1898 757 1906 797
rect 2008 757 2016 797
rect 1898 723 1904 757
rect 2010 723 2016 757
rect 1898 683 1906 723
rect 2008 683 2016 723
rect 1898 649 1904 683
rect 2010 649 2016 683
rect 1898 609 1906 649
rect 2008 609 2016 649
rect 1898 575 1904 609
rect 2010 575 2016 609
rect 1898 535 1906 575
rect 2008 535 2016 575
rect 1898 501 1904 535
rect 2010 501 2016 535
rect 1898 462 1906 501
rect 2008 462 2016 501
rect 1898 428 1904 462
rect 2010 428 2016 462
rect 1898 389 1906 428
rect 2008 389 2016 428
rect 1898 355 1904 389
rect 2010 355 2016 389
rect 1898 316 1906 355
rect 2008 316 2016 355
rect 55 244 63 283
rect 165 244 173 283
rect 55 210 61 244
rect 167 210 173 244
rect 55 171 63 210
rect 165 177 173 210
rect 1898 282 1904 316
rect 2010 282 2016 316
rect 1898 243 1906 282
rect 2008 243 2016 282
rect 2153 1450 6739 1456
rect 2153 1416 2237 1450
rect 2271 1416 2315 1450
rect 2349 1416 2393 1450
rect 2427 1416 2471 1450
rect 2505 1416 2549 1450
rect 2583 1416 2627 1450
rect 2661 1416 2705 1450
rect 2739 1416 2784 1450
rect 2818 1416 2894 1450
rect 2928 1416 2967 1450
rect 3001 1416 3040 1450
rect 3074 1416 3113 1450
rect 3147 1416 3186 1450
rect 3220 1416 3259 1450
rect 3293 1416 3332 1450
rect 3366 1416 3405 1450
rect 3439 1416 3478 1450
rect 3512 1416 3551 1450
rect 3585 1416 3624 1450
rect 3658 1416 3697 1450
rect 3731 1416 3770 1450
rect 3804 1416 3843 1450
rect 3877 1416 3916 1450
rect 3950 1416 3989 1450
rect 4023 1416 4062 1450
rect 4096 1416 4135 1450
rect 4169 1416 4208 1450
rect 4242 1416 4281 1450
rect 4315 1416 4354 1450
rect 4388 1416 4427 1450
rect 4461 1416 4500 1450
rect 4534 1416 4573 1450
rect 4607 1416 4646 1450
rect 4680 1416 4719 1450
rect 4753 1416 4792 1450
rect 4826 1416 4865 1450
rect 4899 1416 4938 1450
rect 4972 1416 5011 1450
rect 5045 1416 5084 1450
rect 5118 1416 5157 1450
rect 5191 1416 5230 1450
rect 5264 1416 5303 1450
rect 5337 1416 5376 1450
rect 5410 1416 5449 1450
rect 5483 1416 5522 1450
rect 5556 1416 5595 1450
rect 5629 1416 5668 1450
rect 5702 1416 5741 1450
rect 5775 1416 5814 1450
rect 5848 1416 5887 1450
rect 5921 1416 5961 1450
rect 5995 1416 6035 1450
rect 6069 1416 6109 1450
rect 6143 1416 6183 1450
rect 6217 1416 6257 1450
rect 6291 1416 6331 1450
rect 6365 1416 6405 1450
rect 6439 1416 6479 1450
rect 6513 1416 6553 1450
rect 6587 1416 6627 1450
rect 6661 1416 6739 1450
rect 2153 1378 6739 1416
rect 2153 1344 2159 1378
rect 2193 1344 2231 1378
rect 2265 1377 2315 1378
rect 2349 1377 2393 1378
rect 2427 1377 2471 1378
rect 2505 1377 2549 1378
rect 2583 1377 2627 1378
rect 2661 1377 2705 1378
rect 2739 1377 2784 1378
rect 2818 1377 2894 1378
rect 2928 1377 2967 1378
rect 3001 1377 3040 1378
rect 3074 1377 3113 1378
rect 3147 1377 3186 1378
rect 3220 1377 3259 1378
rect 3293 1377 3332 1378
rect 3366 1377 3405 1378
rect 3439 1377 3478 1378
rect 3512 1377 3551 1378
rect 3585 1377 3624 1378
rect 3658 1377 3697 1378
rect 3731 1377 3770 1378
rect 3804 1377 3843 1378
rect 3877 1377 3916 1378
rect 3950 1377 3989 1378
rect 4023 1377 4062 1378
rect 4096 1377 4135 1378
rect 4169 1377 4208 1378
rect 4242 1377 4281 1378
rect 4315 1377 4354 1378
rect 4388 1377 4427 1378
rect 2265 1344 2287 1377
rect 2349 1344 2355 1377
rect 2153 1343 2287 1344
rect 2321 1343 2355 1344
rect 2389 1344 2393 1377
rect 2457 1344 2471 1377
rect 2525 1344 2549 1377
rect 2389 1343 2423 1344
rect 2457 1343 2491 1344
rect 2525 1343 2559 1344
rect 2593 1343 2627 1377
rect 2661 1343 2695 1377
rect 2739 1344 2763 1377
rect 2818 1344 2831 1377
rect 2729 1343 2763 1344
rect 2797 1343 2831 1344
rect 2865 1344 2894 1377
rect 2865 1343 2899 1344
rect 2933 1343 2967 1377
rect 3001 1343 3035 1377
rect 3074 1344 3103 1377
rect 3147 1344 3171 1377
rect 3220 1344 3239 1377
rect 3293 1344 3307 1377
rect 3366 1344 3375 1377
rect 3439 1344 3443 1377
rect 3069 1343 3103 1344
rect 3137 1343 3171 1344
rect 3205 1343 3239 1344
rect 3273 1343 3307 1344
rect 3341 1343 3375 1344
rect 3409 1343 3443 1344
rect 3477 1344 3478 1377
rect 3545 1344 3551 1377
rect 3613 1344 3624 1377
rect 3681 1344 3697 1377
rect 3749 1344 3770 1377
rect 3817 1344 3843 1377
rect 3885 1344 3916 1377
rect 3477 1343 3511 1344
rect 3545 1343 3579 1344
rect 3613 1343 3647 1344
rect 3681 1343 3715 1344
rect 3749 1343 3783 1344
rect 3817 1343 3851 1344
rect 3885 1343 3919 1344
rect 3953 1343 3987 1377
rect 4023 1344 4055 1377
rect 4096 1344 4123 1377
rect 4169 1344 4191 1377
rect 4242 1344 4259 1377
rect 4315 1344 4327 1377
rect 4388 1344 4395 1377
rect 4461 1344 4500 1378
rect 4534 1377 4573 1378
rect 4607 1377 4646 1378
rect 4680 1377 4719 1378
rect 4753 1377 4792 1378
rect 4826 1377 4865 1378
rect 4899 1377 4938 1378
rect 4972 1377 5011 1378
rect 5045 1377 5084 1378
rect 5118 1377 5157 1378
rect 5191 1377 5230 1378
rect 5264 1377 5303 1378
rect 5337 1377 5376 1378
rect 5410 1377 5449 1378
rect 5483 1377 5522 1378
rect 5556 1377 5595 1378
rect 5629 1377 5668 1378
rect 5702 1377 5741 1378
rect 5775 1377 5814 1378
rect 5848 1377 5887 1378
rect 5921 1377 5961 1378
rect 5995 1377 6035 1378
rect 6069 1377 6109 1378
rect 6143 1377 6183 1378
rect 6217 1377 6257 1378
rect 6291 1377 6331 1378
rect 6365 1377 6405 1378
rect 6439 1377 6479 1378
rect 6513 1377 6553 1378
rect 6587 1377 6627 1378
rect 4544 1344 4573 1377
rect 4021 1343 4055 1344
rect 4089 1343 4123 1344
rect 4157 1343 4191 1344
rect 4225 1343 4259 1344
rect 4293 1343 4327 1344
rect 4361 1343 4395 1344
rect 4429 1343 4510 1344
rect 4544 1343 4578 1344
rect 4612 1343 4646 1377
rect 4680 1343 4714 1377
rect 4753 1344 4782 1377
rect 4826 1344 4850 1377
rect 4899 1344 4918 1377
rect 4972 1344 4986 1377
rect 5045 1344 5054 1377
rect 5118 1344 5122 1377
rect 4748 1343 4782 1344
rect 4816 1343 4850 1344
rect 4884 1343 4918 1344
rect 4952 1343 4986 1344
rect 5020 1343 5054 1344
rect 5088 1343 5122 1344
rect 5156 1344 5157 1377
rect 5224 1344 5230 1377
rect 5292 1344 5303 1377
rect 5360 1344 5376 1377
rect 5428 1344 5449 1377
rect 5496 1344 5522 1377
rect 5564 1344 5595 1377
rect 5156 1343 5190 1344
rect 5224 1343 5258 1344
rect 5292 1343 5326 1344
rect 5360 1343 5394 1344
rect 5428 1343 5462 1344
rect 5496 1343 5530 1344
rect 5564 1343 5598 1344
rect 5632 1343 5666 1377
rect 5702 1344 5734 1377
rect 5775 1344 5802 1377
rect 5848 1344 5870 1377
rect 5921 1344 5938 1377
rect 5995 1344 6006 1377
rect 6069 1344 6074 1377
rect 5700 1343 5734 1344
rect 5768 1343 5802 1344
rect 5836 1343 5870 1344
rect 5904 1343 5938 1344
rect 5972 1343 6006 1344
rect 6040 1343 6074 1344
rect 6108 1344 6109 1377
rect 6176 1344 6183 1377
rect 6244 1344 6257 1377
rect 6312 1344 6331 1377
rect 6380 1344 6405 1377
rect 6448 1344 6479 1377
rect 6108 1343 6142 1344
rect 6176 1343 6210 1344
rect 6244 1343 6278 1344
rect 6312 1343 6346 1344
rect 6380 1343 6414 1344
rect 6448 1343 6482 1344
rect 6516 1343 6550 1377
rect 6587 1344 6618 1377
rect 6584 1343 6618 1344
rect 2153 1338 6627 1343
rect 2153 1312 2271 1338
rect 2153 1305 2195 1312
rect 2153 1271 2159 1305
rect 2193 1278 2195 1305
rect 2229 1305 2271 1312
rect 2229 1278 2231 1305
rect 2193 1271 2231 1278
rect 2265 1271 2271 1305
rect 2153 1244 2271 1271
rect 2153 1232 2195 1244
rect 2153 1198 2159 1232
rect 2193 1210 2195 1232
rect 2229 1232 2271 1244
rect 2229 1210 2231 1232
rect 2193 1198 2231 1210
rect 2265 1198 2271 1232
rect 2389 1224 2401 1258
rect 2439 1224 2473 1258
rect 2509 1224 2541 1258
rect 2583 1224 2609 1258
rect 2657 1224 2677 1258
rect 2731 1224 2745 1258
rect 2805 1224 2813 1258
rect 2879 1224 2881 1258
rect 2915 1224 2919 1258
rect 2983 1224 2993 1258
rect 3051 1224 3067 1258
rect 3119 1224 3141 1258
rect 3187 1224 3215 1258
rect 3255 1224 3289 1258
rect 3323 1224 3357 1258
rect 3397 1224 3425 1258
rect 3471 1224 3493 1258
rect 3544 1224 3561 1258
rect 3617 1224 3629 1258
rect 3690 1224 3697 1258
rect 3763 1224 3765 1258
rect 3799 1224 3802 1258
rect 3867 1224 3875 1258
rect 3935 1224 3948 1258
rect 4003 1224 4021 1258
rect 4071 1224 4094 1258
rect 4139 1224 4167 1258
rect 4207 1224 4240 1258
rect 4275 1224 4309 1258
rect 4347 1224 4359 1258
rect 4533 1224 4545 1258
rect 4583 1224 4617 1258
rect 4652 1224 4685 1258
rect 4725 1224 4753 1258
rect 4798 1224 4821 1258
rect 4871 1224 4889 1258
rect 4944 1224 4957 1258
rect 5017 1224 5025 1258
rect 5090 1224 5093 1258
rect 5127 1224 5129 1258
rect 5195 1224 5202 1258
rect 5263 1224 5275 1258
rect 5331 1224 5348 1258
rect 5399 1224 5421 1258
rect 5467 1224 5495 1258
rect 5535 1224 5569 1258
rect 5603 1224 5637 1258
rect 5677 1224 5705 1258
rect 5751 1224 5773 1258
rect 5825 1224 5841 1258
rect 5899 1224 5909 1258
rect 5973 1224 5977 1258
rect 6011 1224 6013 1258
rect 6079 1224 6087 1258
rect 6147 1224 6161 1258
rect 6215 1224 6235 1258
rect 6283 1224 6309 1258
rect 6351 1224 6383 1258
rect 6419 1224 6453 1258
rect 6491 1224 6503 1258
rect 2153 1176 2271 1198
rect 2153 1159 2195 1176
rect 2153 1125 2159 1159
rect 2193 1142 2195 1159
rect 2229 1159 2271 1176
rect 2229 1142 2231 1159
rect 2193 1125 2231 1142
rect 2265 1125 2271 1159
rect 2153 1108 2271 1125
rect 2153 1086 2195 1108
rect 2153 1052 2159 1086
rect 2193 1074 2195 1086
rect 2229 1086 2271 1108
rect 2229 1074 2231 1086
rect 2193 1052 2231 1074
rect 2265 1052 2271 1086
rect 2153 1040 2271 1052
rect 2153 1013 2195 1040
rect 2153 979 2159 1013
rect 2193 1006 2195 1013
rect 2229 1013 2271 1040
rect 2229 1006 2231 1013
rect 2193 979 2231 1006
rect 2265 979 2271 1013
rect 2153 972 2271 979
rect 2153 940 2195 972
rect 2153 906 2159 940
rect 2193 938 2195 940
rect 2229 940 2271 972
rect 2229 938 2231 940
rect 2193 906 2231 938
rect 2265 906 2271 940
rect 2153 904 2271 906
rect 2153 870 2195 904
rect 2229 870 2271 904
rect 2153 867 2271 870
rect 2153 833 2159 867
rect 2193 836 2231 867
rect 2193 833 2195 836
rect 2153 802 2195 833
rect 2229 833 2231 836
rect 2265 833 2271 867
rect 2229 802 2271 833
rect 2153 794 2271 802
rect 2153 760 2159 794
rect 2193 768 2231 794
rect 2193 760 2195 768
rect 2153 734 2195 760
rect 2229 760 2231 768
rect 2265 760 2271 794
rect 2229 734 2271 760
rect 2153 721 2271 734
rect 2153 687 2159 721
rect 2193 700 2231 721
rect 2193 687 2195 700
rect 2153 666 2195 687
rect 2229 687 2231 700
rect 2265 687 2271 721
rect 2229 666 2271 687
rect 2153 648 2271 666
rect 2153 614 2159 648
rect 2193 632 2231 648
rect 2193 614 2195 632
rect 2153 598 2195 614
rect 2229 614 2231 632
rect 2265 614 2271 648
rect 2229 598 2271 614
rect 2153 575 2271 598
rect 2153 541 2159 575
rect 2193 564 2231 575
rect 2193 541 2195 564
rect 2153 530 2195 541
rect 2229 541 2231 564
rect 2265 541 2271 575
rect 2229 530 2271 541
rect 2153 502 2271 530
rect 2153 324 2159 502
rect 2265 364 2271 502
rect 2311 1201 2345 1213
rect 2311 1124 2345 1163
rect 6547 1201 6581 1213
rect 6547 1124 6581 1163
rect 2311 1051 2345 1086
rect 2389 1068 2401 1102
rect 2439 1068 2473 1102
rect 2509 1068 2541 1102
rect 2583 1068 2609 1102
rect 2657 1068 2677 1102
rect 2731 1068 2745 1102
rect 2805 1068 2813 1102
rect 2879 1068 2881 1102
rect 2915 1068 2919 1102
rect 2983 1068 2993 1102
rect 3051 1068 3067 1102
rect 3119 1068 3141 1102
rect 3187 1068 3215 1102
rect 3255 1068 3289 1102
rect 3323 1068 3357 1102
rect 3397 1068 3425 1102
rect 3471 1068 3493 1102
rect 3544 1068 3561 1102
rect 3617 1068 3629 1102
rect 3690 1068 3697 1102
rect 3763 1068 3765 1102
rect 3799 1068 3802 1102
rect 3867 1068 3875 1102
rect 3935 1068 3948 1102
rect 4003 1068 4021 1102
rect 4071 1068 4094 1102
rect 4139 1068 4167 1102
rect 4207 1068 4240 1102
rect 4275 1068 4309 1102
rect 4347 1068 4359 1102
rect 4533 1068 4545 1102
rect 4583 1068 4617 1102
rect 4652 1068 4685 1102
rect 4725 1068 4753 1102
rect 4798 1068 4821 1102
rect 4871 1068 4889 1102
rect 4944 1068 4957 1102
rect 5017 1068 5025 1102
rect 5090 1068 5093 1102
rect 5127 1068 5129 1102
rect 5195 1068 5202 1102
rect 5263 1068 5275 1102
rect 5331 1068 5348 1102
rect 5399 1068 5421 1102
rect 5467 1068 5495 1102
rect 5535 1068 5569 1102
rect 5603 1068 5637 1102
rect 5677 1068 5705 1102
rect 5751 1068 5773 1102
rect 5825 1068 5841 1102
rect 5899 1068 5909 1102
rect 5973 1068 5977 1102
rect 6011 1068 6013 1102
rect 6079 1068 6087 1102
rect 6147 1068 6161 1102
rect 6215 1068 6235 1102
rect 6283 1068 6309 1102
rect 6351 1068 6383 1102
rect 6419 1068 6453 1102
rect 6491 1068 6503 1102
rect 2311 978 2345 1004
rect 6547 1051 6581 1084
rect 6547 978 6581 1001
rect 2311 905 2345 922
rect 2389 912 2401 946
rect 2439 912 2473 946
rect 2509 912 2541 946
rect 2583 912 2609 946
rect 2657 912 2677 946
rect 2731 912 2745 946
rect 2805 912 2813 946
rect 2879 912 2881 946
rect 2915 912 2919 946
rect 2983 912 2993 946
rect 3051 912 3067 946
rect 3119 912 3141 946
rect 3187 912 3215 946
rect 3255 912 3289 946
rect 3323 912 3357 946
rect 3397 912 3425 946
rect 3471 912 3493 946
rect 3544 912 3561 946
rect 3617 912 3629 946
rect 3690 912 3697 946
rect 3763 912 3765 946
rect 3799 912 3802 946
rect 3867 912 3875 946
rect 3935 912 3948 946
rect 4003 912 4021 946
rect 4071 912 4094 946
rect 4139 912 4167 946
rect 4207 912 4240 946
rect 4275 912 4309 946
rect 4347 912 4359 946
rect 4533 912 4545 946
rect 4583 912 4617 946
rect 4652 912 4685 946
rect 4725 912 4753 946
rect 4798 912 4821 946
rect 4871 912 4889 946
rect 4944 912 4957 946
rect 5017 912 5025 946
rect 5090 912 5093 946
rect 5127 912 5129 946
rect 5195 912 5202 946
rect 5263 912 5275 946
rect 5331 912 5348 946
rect 5399 912 5421 946
rect 5467 912 5495 946
rect 5535 912 5569 946
rect 5603 912 5637 946
rect 5677 912 5705 946
rect 5751 912 5773 946
rect 5825 912 5841 946
rect 5899 912 5909 946
rect 5973 912 5977 946
rect 6011 912 6013 946
rect 6079 912 6087 946
rect 6147 912 6161 946
rect 6215 912 6235 946
rect 6283 912 6309 946
rect 6351 912 6383 946
rect 6419 912 6453 946
rect 6491 912 6503 946
rect 2311 832 2345 840
rect 2311 792 2345 798
rect 6547 905 6581 918
rect 6547 868 6581 871
rect 6547 832 6581 834
rect 2389 756 2401 790
rect 2439 756 2473 790
rect 2509 756 2541 790
rect 2583 756 2609 790
rect 2657 756 2677 790
rect 2731 756 2745 790
rect 2805 756 2813 790
rect 2879 756 2881 790
rect 2915 756 2919 790
rect 2983 756 2993 790
rect 3051 756 3067 790
rect 3119 756 3141 790
rect 3187 756 3215 790
rect 3255 756 3289 790
rect 3323 756 3357 790
rect 3397 756 3425 790
rect 3471 756 3493 790
rect 3544 756 3561 790
rect 3617 756 3629 790
rect 3690 756 3697 790
rect 3763 756 3765 790
rect 3799 756 3802 790
rect 3867 756 3875 790
rect 3935 756 3948 790
rect 4003 756 4021 790
rect 4071 756 4094 790
rect 4139 756 4167 790
rect 4207 756 4240 790
rect 4275 756 4309 790
rect 4347 756 4359 790
rect 4533 756 4545 790
rect 4583 756 4617 790
rect 4652 756 4685 790
rect 4725 756 4753 790
rect 4798 756 4821 790
rect 4871 756 4889 790
rect 4944 756 4957 790
rect 5017 756 5025 790
rect 5090 756 5093 790
rect 5127 756 5129 790
rect 5195 756 5202 790
rect 5263 756 5275 790
rect 5331 756 5348 790
rect 5399 756 5421 790
rect 5467 756 5495 790
rect 5535 756 5569 790
rect 5603 756 5637 790
rect 5677 756 5705 790
rect 5751 756 5773 790
rect 5825 756 5841 790
rect 5899 756 5909 790
rect 5973 756 5977 790
rect 6011 756 6013 790
rect 6079 756 6087 790
rect 6147 756 6161 790
rect 6215 756 6235 790
rect 6283 756 6309 790
rect 6351 756 6383 790
rect 6419 756 6453 790
rect 6491 756 6503 790
rect 6547 784 6581 798
rect 2311 710 2345 725
rect 2311 613 2345 652
rect 6547 700 6581 725
rect 2389 600 2401 634
rect 2439 600 2473 634
rect 2509 600 2541 634
rect 2583 600 2609 634
rect 2657 600 2677 634
rect 2731 600 2745 634
rect 2805 600 2813 634
rect 2879 600 2881 634
rect 2915 600 2919 634
rect 2983 600 2993 634
rect 3051 600 3067 634
rect 3119 600 3141 634
rect 3187 600 3215 634
rect 3255 600 3289 634
rect 3323 600 3357 634
rect 3397 600 3425 634
rect 3471 600 3493 634
rect 3544 600 3561 634
rect 3617 600 3629 634
rect 3690 600 3697 634
rect 3763 600 3765 634
rect 3799 600 3802 634
rect 3867 600 3875 634
rect 3935 600 3948 634
rect 4003 600 4021 634
rect 4071 600 4094 634
rect 4139 600 4167 634
rect 4207 600 4240 634
rect 4275 600 4309 634
rect 4347 600 4359 634
rect 4533 600 4545 634
rect 4583 600 4617 634
rect 4652 600 4685 634
rect 4725 600 4753 634
rect 4798 600 4821 634
rect 4871 600 4889 634
rect 4944 600 4957 634
rect 5017 600 5025 634
rect 5090 600 5093 634
rect 5127 600 5129 634
rect 5195 600 5202 634
rect 5263 600 5275 634
rect 5331 600 5348 634
rect 5399 600 5421 634
rect 5467 600 5495 634
rect 5535 600 5569 634
rect 5603 600 5637 634
rect 5677 600 5705 634
rect 5751 600 5773 634
rect 5825 600 5841 634
rect 5899 600 5909 634
rect 5973 600 5977 634
rect 6011 600 6013 634
rect 6079 600 6087 634
rect 6147 600 6161 634
rect 6215 600 6235 634
rect 6283 600 6309 634
rect 6351 600 6383 634
rect 6419 600 6453 634
rect 6491 600 6503 634
rect 6547 613 6581 652
rect 2311 539 2345 579
rect 2311 489 2345 505
rect 6547 539 6581 579
rect 6547 489 6581 505
rect 6621 1200 6627 1338
rect 6733 1200 6739 1378
rect 6621 1172 6739 1200
rect 6621 1161 6683 1172
rect 6717 1161 6739 1172
rect 6621 1127 6627 1161
rect 6661 1138 6683 1161
rect 6661 1127 6699 1138
rect 6733 1127 6739 1161
rect 6621 1104 6739 1127
rect 6621 1088 6683 1104
rect 6717 1088 6739 1104
rect 6621 1054 6627 1088
rect 6661 1070 6683 1088
rect 6661 1054 6699 1070
rect 6733 1054 6739 1088
rect 6621 1036 6739 1054
rect 6621 1015 6683 1036
rect 6717 1015 6739 1036
rect 6621 981 6627 1015
rect 6661 1002 6683 1015
rect 6661 981 6699 1002
rect 6733 981 6739 1015
rect 6621 968 6739 981
rect 6621 942 6683 968
rect 6717 942 6739 968
rect 6621 908 6627 942
rect 6661 934 6683 942
rect 6661 908 6699 934
rect 6733 908 6739 942
rect 6621 900 6739 908
rect 6621 869 6683 900
rect 6717 869 6739 900
rect 6621 835 6627 869
rect 6661 866 6683 869
rect 6661 835 6699 866
rect 6733 835 6739 869
rect 6621 832 6739 835
rect 6621 798 6683 832
rect 6717 798 6739 832
rect 6621 796 6739 798
rect 6621 762 6627 796
rect 6661 764 6699 796
rect 6661 762 6683 764
rect 6733 762 6739 796
rect 6621 730 6683 762
rect 6717 730 6739 762
rect 6621 723 6739 730
rect 6621 689 6627 723
rect 6661 696 6699 723
rect 6661 689 6683 696
rect 6733 689 6739 723
rect 6621 662 6683 689
rect 6717 662 6739 689
rect 6621 650 6739 662
rect 6621 616 6627 650
rect 6661 628 6699 650
rect 6661 616 6683 628
rect 6733 616 6739 650
rect 6621 594 6683 616
rect 6717 594 6739 616
rect 6621 577 6739 594
rect 6621 543 6627 577
rect 6661 560 6699 577
rect 6661 543 6683 560
rect 6733 543 6739 577
rect 6621 526 6683 543
rect 6717 526 6739 543
rect 6621 504 6739 526
rect 2389 444 2401 478
rect 2439 444 2473 478
rect 2509 444 2541 478
rect 2583 444 2609 478
rect 2657 444 2677 478
rect 2731 444 2745 478
rect 2805 444 2813 478
rect 2879 444 2881 478
rect 2915 444 2919 478
rect 2983 444 2993 478
rect 3051 444 3067 478
rect 3119 444 3141 478
rect 3187 444 3215 478
rect 3255 444 3289 478
rect 3323 444 3357 478
rect 3397 444 3425 478
rect 3471 444 3493 478
rect 3544 444 3561 478
rect 3617 444 3629 478
rect 3690 444 3697 478
rect 3763 444 3765 478
rect 3799 444 3802 478
rect 3867 444 3875 478
rect 3935 444 3948 478
rect 4003 444 4021 478
rect 4071 444 4094 478
rect 4139 444 4167 478
rect 4207 444 4240 478
rect 4275 444 4309 478
rect 4347 444 4359 478
rect 4533 444 4545 478
rect 4583 444 4617 478
rect 4652 444 4685 478
rect 4725 444 4753 478
rect 4798 444 4821 478
rect 4871 444 4889 478
rect 4944 444 4957 478
rect 5017 444 5025 478
rect 5090 444 5093 478
rect 5127 444 5129 478
rect 5195 444 5202 478
rect 5263 444 5275 478
rect 5331 444 5348 478
rect 5399 444 5421 478
rect 5467 444 5495 478
rect 5535 444 5569 478
rect 5603 444 5637 478
rect 5677 444 5705 478
rect 5751 444 5773 478
rect 5825 444 5841 478
rect 5899 444 5909 478
rect 5973 444 5977 478
rect 6011 444 6013 478
rect 6079 444 6087 478
rect 6147 444 6161 478
rect 6215 444 6235 478
rect 6283 444 6309 478
rect 6351 444 6383 478
rect 6419 444 6453 478
rect 6491 444 6503 478
rect 6621 470 6627 504
rect 6661 492 6699 504
rect 6661 470 6683 492
rect 6733 470 6739 504
rect 6621 458 6683 470
rect 6717 458 6739 470
rect 6621 431 6739 458
rect 6621 397 6627 431
rect 6661 424 6699 431
rect 6661 397 6683 424
rect 6733 397 6739 431
rect 6621 390 6683 397
rect 6717 390 6739 397
rect 6621 364 6739 390
rect 2265 359 6739 364
rect 2294 358 2328 359
rect 2362 358 2396 359
rect 2430 358 2464 359
rect 2498 358 2532 359
rect 2566 358 2600 359
rect 2634 358 2668 359
rect 2702 358 2736 359
rect 2770 358 2804 359
rect 2838 358 2872 359
rect 2906 358 2940 359
rect 2974 358 3008 359
rect 3042 358 3076 359
rect 3110 358 3144 359
rect 3178 358 3212 359
rect 3246 358 3280 359
rect 3314 358 3348 359
rect 3382 358 3416 359
rect 3450 358 3484 359
rect 3518 358 3552 359
rect 3586 358 3620 359
rect 3654 358 3688 359
rect 3722 358 3756 359
rect 3790 358 3824 359
rect 3858 358 3892 359
rect 3926 358 3960 359
rect 3994 358 4028 359
rect 4062 358 4096 359
rect 4130 358 4164 359
rect 4198 358 4232 359
rect 4266 358 4300 359
rect 4334 358 4368 359
rect 4402 358 4436 359
rect 4470 358 4504 359
rect 4538 358 4572 359
rect 4606 358 4640 359
rect 4674 358 4708 359
rect 4742 358 4776 359
rect 4810 358 4844 359
rect 4878 358 4912 359
rect 4946 358 4980 359
rect 5014 358 5048 359
rect 5082 358 5116 359
rect 5150 358 5184 359
rect 5218 358 5252 359
rect 5286 358 5320 359
rect 5354 358 5388 359
rect 5422 358 5456 359
rect 5490 358 5524 359
rect 5558 358 5592 359
rect 5626 358 5660 359
rect 5694 358 5728 359
rect 5762 358 5796 359
rect 5830 358 5864 359
rect 5898 358 5932 359
rect 5966 358 6000 359
rect 6034 358 6068 359
rect 6102 358 6136 359
rect 6170 358 6204 359
rect 6238 358 6272 359
rect 6306 358 6340 359
rect 6374 358 6408 359
rect 6442 358 6476 359
rect 6510 358 6544 359
rect 6578 358 6612 359
rect 6646 358 6739 359
rect 2294 325 2304 358
rect 2362 325 2377 358
rect 2430 325 2450 358
rect 2498 325 2523 358
rect 2265 324 2304 325
rect 2338 324 2377 325
rect 2411 324 2450 325
rect 2484 324 2523 325
rect 2153 286 2523 324
rect 2153 252 2231 286
rect 2265 252 2304 286
rect 2338 252 2377 286
rect 2411 252 2450 286
rect 2484 252 2523 286
rect 6661 324 6699 358
rect 6733 324 6739 358
rect 6661 252 6739 324
rect 2153 246 6739 252
rect 6876 1434 6994 1456
rect 6876 1424 6884 1434
rect 6986 1424 6994 1434
rect 6876 1390 6882 1424
rect 6988 1390 6994 1424
rect 6876 1351 6884 1390
rect 6986 1351 6994 1390
rect 6876 1317 6882 1351
rect 6988 1317 6994 1351
rect 6876 1278 6884 1317
rect 6986 1278 6994 1317
rect 6876 1244 6882 1278
rect 6988 1244 6994 1278
rect 6876 1205 6884 1244
rect 6986 1205 6994 1244
rect 6876 1171 6882 1205
rect 6988 1171 6994 1205
rect 6876 1131 6884 1171
rect 6986 1131 6994 1171
rect 6876 1097 6882 1131
rect 6988 1097 6994 1131
rect 6876 1057 6884 1097
rect 6986 1057 6994 1097
rect 6876 1023 6882 1057
rect 6988 1023 6994 1057
rect 6876 983 6884 1023
rect 6986 983 6994 1023
rect 6876 949 6882 983
rect 6988 949 6994 983
rect 6876 909 6884 949
rect 6986 909 6994 949
rect 6876 875 6882 909
rect 6988 875 6994 909
rect 6876 835 6884 875
rect 6986 835 6994 875
rect 6876 801 6882 835
rect 6988 801 6994 835
rect 6876 761 6884 801
rect 6986 761 6994 801
rect 6876 727 6882 761
rect 6988 727 6994 761
rect 6876 687 6884 727
rect 6986 687 6994 727
rect 6876 653 6882 687
rect 6988 653 6994 687
rect 6876 613 6884 653
rect 6986 613 6994 653
rect 6876 579 6882 613
rect 6988 579 6994 613
rect 6876 539 6884 579
rect 6986 539 6994 579
rect 6876 505 6882 539
rect 6988 505 6994 539
rect 6876 465 6884 505
rect 6986 465 6994 505
rect 6876 431 6882 465
rect 6988 431 6994 465
rect 6876 391 6884 431
rect 6986 391 6994 431
rect 6876 357 6882 391
rect 6988 357 6994 391
rect 6876 317 6884 357
rect 6986 317 6994 357
rect 6876 283 6882 317
rect 6916 283 6954 312
rect 6988 283 6994 317
rect 1898 209 1904 243
rect 2010 209 2016 243
rect 1898 177 1906 209
rect 165 171 1906 177
rect 2008 177 2016 209
rect 6876 243 6994 283
rect 7157 1440 11757 1446
rect 7157 1406 7241 1440
rect 7275 1406 7319 1440
rect 7353 1406 7397 1440
rect 7431 1406 7475 1440
rect 7509 1406 7553 1440
rect 7587 1406 7631 1440
rect 7665 1406 7709 1440
rect 7743 1406 7788 1440
rect 7822 1406 7898 1440
rect 7157 1377 7898 1406
rect 11460 1406 11499 1440
rect 11533 1406 11572 1440
rect 11606 1406 11645 1440
rect 11679 1406 11757 1440
rect 11460 1377 11757 1406
rect 7157 1368 7264 1377
rect 7298 1368 7332 1377
rect 7366 1368 7400 1377
rect 7157 1334 7163 1368
rect 7197 1334 7235 1368
rect 7298 1343 7319 1368
rect 7366 1343 7397 1368
rect 7434 1343 7468 1377
rect 7502 1368 7536 1377
rect 7570 1368 7604 1377
rect 7638 1368 7672 1377
rect 7509 1343 7536 1368
rect 7587 1343 7604 1368
rect 7665 1343 7672 1368
rect 7706 1368 7740 1377
rect 7774 1368 7808 1377
rect 7706 1343 7709 1368
rect 7774 1343 7788 1368
rect 7842 1343 7876 1377
rect 11460 1343 11472 1377
rect 11506 1368 11540 1377
rect 11574 1368 11608 1377
rect 11533 1343 11540 1368
rect 11606 1343 11608 1368
rect 11642 1368 11757 1377
rect 11642 1343 11645 1368
rect 7269 1334 7319 1343
rect 7353 1334 7397 1343
rect 7431 1334 7475 1343
rect 7509 1334 7553 1343
rect 7587 1334 7631 1343
rect 7665 1334 7709 1343
rect 7743 1334 7788 1343
rect 7822 1334 7898 1343
rect 11460 1334 11499 1343
rect 11533 1334 11572 1343
rect 11606 1334 11645 1343
rect 7157 1328 11645 1334
rect 7157 1308 7275 1328
rect 7157 1295 7199 1308
rect 7157 1261 7163 1295
rect 7197 1274 7199 1295
rect 7233 1295 7275 1308
rect 7233 1274 7235 1295
rect 7197 1261 7235 1274
rect 7269 1261 7275 1295
rect 7157 1240 7275 1261
rect 7157 1222 7199 1240
rect 7233 1222 7275 1240
rect 7454 1224 7462 1258
rect 7528 1224 7530 1258
rect 7564 1224 7568 1258
rect 7632 1224 7642 1258
rect 7700 1224 7716 1258
rect 7768 1224 7790 1258
rect 7836 1224 7864 1258
rect 7904 1224 7938 1258
rect 7972 1224 8006 1258
rect 8046 1224 8074 1258
rect 8120 1224 8142 1258
rect 8194 1224 8210 1258
rect 8268 1224 8278 1258
rect 8342 1224 8346 1258
rect 8380 1224 8382 1258
rect 8448 1224 8456 1258
rect 8516 1224 8529 1258
rect 8584 1224 8602 1258
rect 8652 1224 8675 1258
rect 8720 1224 8748 1258
rect 8788 1224 8821 1258
rect 8856 1224 8890 1258
rect 8928 1224 8958 1258
rect 9001 1224 9026 1258
rect 9074 1224 9094 1258
rect 9147 1224 9162 1258
rect 9220 1224 9230 1258
rect 9293 1224 9298 1258
rect 9400 1224 9416 1258
rect 9552 1224 9564 1258
rect 9602 1224 9636 1258
rect 9671 1224 9704 1258
rect 9744 1224 9772 1258
rect 9817 1224 9840 1258
rect 9890 1224 9908 1258
rect 9963 1224 9976 1258
rect 10036 1224 10044 1258
rect 10109 1224 10112 1258
rect 10146 1224 10148 1258
rect 10214 1224 10221 1258
rect 10282 1224 10294 1258
rect 10350 1224 10367 1258
rect 10418 1224 10440 1258
rect 10486 1224 10514 1258
rect 10554 1224 10588 1258
rect 10622 1224 10656 1258
rect 10696 1224 10724 1258
rect 10770 1224 10792 1258
rect 10844 1224 10860 1258
rect 10918 1224 10928 1258
rect 10992 1224 10996 1258
rect 11030 1224 11032 1258
rect 11098 1224 11106 1258
rect 11166 1224 11180 1258
rect 11234 1224 11254 1258
rect 11302 1224 11328 1258
rect 11370 1224 11402 1258
rect 11438 1224 11472 1258
rect 11510 1224 11522 1258
rect 7157 324 7163 1222
rect 7269 364 7275 1222
rect 7330 1201 7364 1213
rect 7330 1127 7364 1163
rect 11565 1201 11599 1213
rect 11565 1197 11566 1201
rect 11599 1163 11600 1167
rect 11565 1127 11600 1163
rect 11565 1123 11566 1127
rect 7330 1053 7364 1089
rect 7454 1068 7462 1102
rect 7528 1068 7530 1102
rect 7564 1068 7568 1102
rect 7632 1068 7642 1102
rect 7700 1068 7716 1102
rect 7768 1068 7790 1102
rect 7836 1068 7864 1102
rect 7904 1068 7938 1102
rect 7972 1068 8006 1102
rect 8046 1068 8074 1102
rect 8120 1068 8142 1102
rect 8194 1068 8210 1102
rect 8268 1068 8278 1102
rect 8342 1068 8346 1102
rect 8380 1068 8382 1102
rect 8448 1068 8456 1102
rect 8516 1068 8529 1102
rect 8584 1068 8602 1102
rect 8652 1068 8675 1102
rect 8720 1068 8748 1102
rect 8788 1068 8821 1102
rect 8856 1068 8890 1102
rect 8928 1068 8958 1102
rect 9001 1068 9026 1102
rect 9074 1068 9094 1102
rect 9147 1068 9162 1102
rect 9220 1068 9230 1102
rect 9293 1068 9298 1102
rect 9400 1068 9416 1102
rect 9552 1068 9564 1102
rect 9602 1068 9636 1102
rect 9671 1068 9704 1102
rect 9744 1068 9772 1102
rect 9817 1068 9840 1102
rect 9890 1068 9908 1102
rect 9963 1068 9976 1102
rect 10036 1068 10044 1102
rect 10109 1068 10112 1102
rect 10146 1068 10148 1102
rect 10214 1068 10221 1102
rect 10282 1068 10294 1102
rect 10350 1068 10367 1102
rect 10418 1068 10440 1102
rect 10486 1068 10514 1102
rect 10554 1068 10588 1102
rect 10622 1068 10656 1102
rect 10696 1068 10724 1102
rect 10770 1068 10792 1102
rect 10844 1068 10860 1102
rect 10918 1068 10928 1102
rect 10992 1068 10996 1102
rect 11030 1068 11032 1102
rect 11098 1068 11106 1102
rect 11166 1068 11180 1102
rect 11234 1068 11254 1102
rect 11302 1068 11328 1102
rect 11370 1068 11402 1102
rect 11438 1068 11472 1102
rect 11510 1068 11522 1102
rect 11599 1089 11600 1093
rect 7330 979 7364 1016
rect 11565 1053 11600 1089
rect 11565 1050 11566 1053
rect 11599 1016 11600 1019
rect 11565 979 11600 1016
rect 11565 977 11566 979
rect 7330 905 7364 943
rect 7454 912 7462 946
rect 7528 912 7530 946
rect 7564 912 7568 946
rect 7632 912 7642 946
rect 7700 912 7716 946
rect 7768 912 7790 946
rect 7836 912 7864 946
rect 7904 912 7938 946
rect 7972 912 8006 946
rect 8046 912 8074 946
rect 8120 912 8142 946
rect 8194 912 8210 946
rect 8268 912 8278 946
rect 8342 912 8346 946
rect 8380 912 8382 946
rect 8448 912 8456 946
rect 8516 912 8529 946
rect 8584 912 8602 946
rect 8652 912 8675 946
rect 8720 912 8748 946
rect 8788 912 8821 946
rect 8856 912 8890 946
rect 8928 912 8958 946
rect 9001 912 9026 946
rect 9074 912 9094 946
rect 9147 912 9162 946
rect 9220 912 9230 946
rect 9293 912 9298 946
rect 9400 912 9416 946
rect 9552 912 9564 946
rect 9602 912 9636 946
rect 9671 912 9704 946
rect 9744 912 9772 946
rect 9817 912 9840 946
rect 9890 912 9908 946
rect 9963 912 9976 946
rect 10036 912 10044 946
rect 10109 912 10112 946
rect 10146 912 10148 946
rect 10214 912 10221 946
rect 10282 912 10294 946
rect 10350 912 10367 946
rect 10418 912 10440 946
rect 10486 912 10514 946
rect 10554 912 10588 946
rect 10622 912 10656 946
rect 10696 912 10724 946
rect 10770 912 10792 946
rect 10844 912 10860 946
rect 10918 912 10928 946
rect 10992 912 10996 946
rect 11030 912 11032 946
rect 11098 912 11106 946
rect 11166 912 11180 946
rect 11234 912 11254 946
rect 11302 912 11328 946
rect 11370 912 11402 946
rect 11438 912 11472 946
rect 11510 912 11522 946
rect 11599 943 11600 945
rect 7330 831 7364 870
rect 7330 758 7364 797
rect 11565 905 11600 943
rect 11565 904 11566 905
rect 11599 870 11600 871
rect 11565 831 11600 870
rect 7454 756 7462 790
rect 7528 756 7530 790
rect 7564 756 7568 790
rect 7632 756 7642 790
rect 7700 756 7716 790
rect 7768 756 7790 790
rect 7836 756 7864 790
rect 7904 756 7938 790
rect 7972 756 8006 790
rect 8046 756 8074 790
rect 8120 756 8142 790
rect 8194 756 8210 790
rect 8268 756 8278 790
rect 8342 756 8346 790
rect 8380 756 8382 790
rect 8448 756 8456 790
rect 8516 756 8529 790
rect 8584 756 8602 790
rect 8652 756 8675 790
rect 8720 756 8748 790
rect 8788 756 8821 790
rect 8856 756 8890 790
rect 8928 756 8958 790
rect 9001 756 9026 790
rect 9074 756 9094 790
rect 9147 756 9162 790
rect 9220 756 9230 790
rect 9293 756 9298 790
rect 9400 756 9416 790
rect 9552 756 9564 790
rect 9602 756 9636 790
rect 9671 756 9704 790
rect 9744 756 9772 790
rect 9817 756 9840 790
rect 9890 756 9908 790
rect 9963 756 9976 790
rect 10036 756 10044 790
rect 10109 756 10112 790
rect 10146 756 10148 790
rect 10214 756 10221 790
rect 10282 756 10294 790
rect 10350 756 10367 790
rect 10418 756 10440 790
rect 10486 756 10514 790
rect 10554 756 10588 790
rect 10622 756 10656 790
rect 10696 756 10724 790
rect 10770 756 10792 790
rect 10844 756 10860 790
rect 10918 756 10928 790
rect 10992 756 10996 790
rect 11030 756 11032 790
rect 11098 756 11106 790
rect 11166 756 11180 790
rect 11234 756 11254 790
rect 11302 756 11328 790
rect 11370 756 11402 790
rect 11438 756 11472 790
rect 11510 756 11522 790
rect 11565 758 11600 797
rect 11599 757 11600 758
rect 7330 685 7364 723
rect 7330 612 7364 649
rect 11565 723 11566 724
rect 11565 685 11600 723
rect 11599 683 11600 685
rect 11565 649 11566 651
rect 7454 600 7462 634
rect 7528 600 7530 634
rect 7564 600 7568 634
rect 7632 600 7642 634
rect 7700 600 7716 634
rect 7768 600 7790 634
rect 7836 600 7864 634
rect 7904 600 7938 634
rect 7972 600 8006 634
rect 8046 600 8074 634
rect 8120 600 8142 634
rect 8194 600 8210 634
rect 8268 600 8278 634
rect 8342 600 8346 634
rect 8380 600 8382 634
rect 8448 600 8456 634
rect 8516 600 8529 634
rect 8584 600 8602 634
rect 8652 600 8675 634
rect 8720 600 8748 634
rect 8788 600 8821 634
rect 8856 600 8890 634
rect 8928 600 8958 634
rect 9001 600 9026 634
rect 9074 600 9094 634
rect 9147 600 9162 634
rect 9220 600 9230 634
rect 9293 600 9298 634
rect 9400 600 9416 634
rect 9552 600 9564 634
rect 9602 600 9636 634
rect 9671 600 9704 634
rect 9744 600 9772 634
rect 9817 600 9840 634
rect 9890 600 9908 634
rect 9963 600 9976 634
rect 10036 600 10044 634
rect 10109 600 10112 634
rect 10146 600 10148 634
rect 10214 600 10221 634
rect 10282 600 10294 634
rect 10350 600 10367 634
rect 10418 600 10440 634
rect 10486 600 10514 634
rect 10554 600 10588 634
rect 10622 600 10656 634
rect 10696 600 10724 634
rect 10770 600 10792 634
rect 10844 600 10860 634
rect 10918 600 10928 634
rect 10992 600 10996 634
rect 11030 600 11032 634
rect 11098 600 11106 634
rect 11166 600 11180 634
rect 11234 600 11254 634
rect 11302 600 11328 634
rect 11370 600 11402 634
rect 11438 600 11472 634
rect 11510 600 11522 634
rect 11565 612 11600 649
rect 11599 609 11600 612
rect 7330 539 7364 575
rect 7330 489 7364 501
rect 11565 575 11566 578
rect 11565 539 11600 575
rect 11599 535 11600 539
rect 11565 501 11566 505
rect 11565 489 11599 501
rect 7454 444 7462 478
rect 7528 444 7530 478
rect 7564 444 7568 478
rect 7632 444 7642 478
rect 7700 444 7716 478
rect 7768 444 7790 478
rect 7836 444 7864 478
rect 7904 444 7938 478
rect 7972 444 8006 478
rect 8046 444 8074 478
rect 8120 444 8142 478
rect 8194 444 8210 478
rect 8268 444 8278 478
rect 8342 444 8346 478
rect 8380 444 8382 478
rect 8448 444 8456 478
rect 8516 444 8529 478
rect 8584 444 8602 478
rect 8652 444 8675 478
rect 8720 444 8748 478
rect 8788 444 8821 478
rect 8856 444 8890 478
rect 8928 444 8958 478
rect 9001 444 9026 478
rect 9074 444 9094 478
rect 9147 444 9162 478
rect 9220 444 9230 478
rect 9293 444 9298 478
rect 9400 444 9416 478
rect 9552 444 9564 478
rect 9602 444 9636 478
rect 9671 444 9704 478
rect 9744 444 9772 478
rect 9817 444 9840 478
rect 9890 444 9908 478
rect 9963 444 9976 478
rect 10036 444 10044 478
rect 10109 444 10112 478
rect 10146 444 10148 478
rect 10214 444 10221 478
rect 10282 444 10294 478
rect 10350 444 10367 478
rect 10418 444 10440 478
rect 10486 444 10514 478
rect 10554 444 10588 478
rect 10622 444 10656 478
rect 10696 444 10724 478
rect 10770 444 10792 478
rect 10844 444 10860 478
rect 10918 444 10928 478
rect 10992 444 10996 478
rect 11030 444 11032 478
rect 11098 444 11106 478
rect 11166 444 11180 478
rect 11234 444 11254 478
rect 11302 444 11328 478
rect 11370 444 11402 478
rect 11438 444 11472 478
rect 11510 444 11522 478
rect 11639 470 11645 1328
rect 11751 470 11757 1368
rect 11639 462 11681 470
rect 11715 462 11757 470
rect 11639 431 11757 462
rect 11639 397 11645 431
rect 11679 428 11717 431
rect 11679 397 11681 428
rect 11639 394 11681 397
rect 11715 397 11717 428
rect 11751 397 11757 431
rect 11715 394 11757 397
rect 11639 364 11757 394
rect 7269 359 11757 364
rect 7298 358 7332 359
rect 7366 358 7400 359
rect 7434 358 7468 359
rect 7502 358 7536 359
rect 7570 358 7604 359
rect 7298 325 7308 358
rect 7366 325 7381 358
rect 7434 325 7454 358
rect 7502 325 7527 358
rect 7570 325 7600 358
rect 7638 325 7672 359
rect 7706 358 7740 359
rect 7774 358 7808 359
rect 7842 358 7876 359
rect 7910 358 7944 359
rect 7978 358 8012 359
rect 8046 358 8080 359
rect 8114 358 8148 359
rect 7707 325 7740 358
rect 7780 325 7808 358
rect 7853 325 7876 358
rect 7926 325 7944 358
rect 7999 325 8012 358
rect 8072 325 8080 358
rect 8145 325 8148 358
rect 8182 358 8216 359
rect 8250 358 8284 359
rect 8318 358 8352 359
rect 8386 358 8420 359
rect 8454 358 8488 359
rect 8522 358 8556 359
rect 8590 358 8624 359
rect 8658 358 8692 359
rect 8726 358 8760 359
rect 8794 358 8828 359
rect 8862 358 8896 359
rect 8930 358 8964 359
rect 8998 358 9032 359
rect 9066 358 9100 359
rect 9134 358 9168 359
rect 9202 358 9236 359
rect 9270 358 9304 359
rect 9338 358 9372 359
rect 9406 358 9440 359
rect 9474 358 9508 359
rect 9542 358 9576 359
rect 9610 358 9644 359
rect 9678 358 9712 359
rect 9746 358 9780 359
rect 9814 358 9848 359
rect 9882 358 9916 359
rect 9950 358 9984 359
rect 10018 358 10052 359
rect 10086 358 10120 359
rect 10154 358 10188 359
rect 10222 358 10256 359
rect 10290 358 10324 359
rect 10358 358 10392 359
rect 10426 358 10460 359
rect 10494 358 10528 359
rect 10562 358 10596 359
rect 10630 358 10664 359
rect 10698 358 10732 359
rect 10766 358 10800 359
rect 10834 358 10868 359
rect 10902 358 10936 359
rect 10970 358 11004 359
rect 11038 358 11072 359
rect 11106 358 11140 359
rect 11174 358 11208 359
rect 11242 358 11276 359
rect 11310 358 11344 359
rect 11378 358 11412 359
rect 11446 358 11480 359
rect 11514 358 11548 359
rect 11582 358 11616 359
rect 11650 358 11757 359
rect 8182 325 8184 358
rect 8250 325 8257 358
rect 8318 325 8330 358
rect 8386 325 8403 358
rect 8454 325 8476 358
rect 8522 325 8549 358
rect 7269 324 7308 325
rect 7342 324 7381 325
rect 7415 324 7454 325
rect 7488 324 7527 325
rect 7561 324 7600 325
rect 7634 324 7673 325
rect 7707 324 7746 325
rect 7780 324 7819 325
rect 7853 324 7892 325
rect 7926 324 7965 325
rect 7999 324 8038 325
rect 8072 324 8111 325
rect 8145 324 8184 325
rect 8218 324 8257 325
rect 8291 324 8330 325
rect 8364 324 8403 325
rect 8437 324 8476 325
rect 8510 324 8549 325
rect 7157 286 8549 324
rect 7157 252 7235 286
rect 7269 252 7308 286
rect 7342 252 7381 286
rect 7415 252 7454 286
rect 7488 252 7527 286
rect 7561 252 7600 286
rect 7634 252 7673 286
rect 7707 252 7746 286
rect 7780 252 7819 286
rect 7853 252 7892 286
rect 7926 252 7965 286
rect 7999 252 8038 286
rect 8072 252 8111 286
rect 8145 252 8184 286
rect 8218 252 8257 286
rect 8291 252 8330 286
rect 8364 252 8403 286
rect 8437 252 8476 286
rect 8510 252 8549 286
rect 11679 324 11717 358
rect 11751 324 11757 358
rect 11679 252 11757 324
rect 7157 246 11757 252
rect 11902 1393 12004 1535
rect 6876 177 6882 243
rect 2008 171 6882 177
rect 6988 177 6994 243
rect 6988 171 11893 177
rect 55 137 61 171
rect 167 137 206 171
rect 240 169 279 171
rect 313 169 352 171
rect 386 169 425 171
rect 459 169 498 171
rect 532 169 571 171
rect 605 169 644 171
rect 678 169 717 171
rect 751 169 790 171
rect 824 169 863 171
rect 897 169 936 171
rect 970 169 1009 171
rect 1043 169 1082 171
rect 1116 169 1155 171
rect 1189 169 1228 171
rect 1262 169 1301 171
rect 1335 169 1374 171
rect 1408 169 1447 171
rect 1481 169 1520 171
rect 1554 169 1593 171
rect 1627 169 1666 171
rect 1700 169 1739 171
rect 1773 169 1812 171
rect 1846 169 1885 171
rect 1872 137 1885 169
rect 2008 137 2031 171
rect 2065 169 2104 171
rect 2138 169 2177 171
rect 2211 169 2250 171
rect 2284 169 2323 171
rect 11861 169 11893 171
rect 2065 137 2103 169
rect 55 135 63 137
rect 165 135 206 137
rect 55 101 206 135
rect 55 99 138 101
rect 55 65 133 99
rect 172 67 206 101
rect 1872 135 1906 137
rect 2008 135 2103 137
rect 1872 101 2103 135
rect 1872 99 2035 101
rect 1872 67 1885 99
rect 167 65 206 67
rect 240 65 279 67
rect 313 65 352 67
rect 386 65 425 67
rect 459 65 498 67
rect 532 65 571 67
rect 605 65 644 67
rect 678 65 717 67
rect 751 65 790 67
rect 824 65 863 67
rect 897 65 936 67
rect 970 65 1009 67
rect 1043 65 1082 67
rect 1116 65 1155 67
rect 1189 65 1228 67
rect 1262 65 1301 67
rect 1335 65 1374 67
rect 1408 65 1447 67
rect 1481 65 1520 67
rect 1554 65 1593 67
rect 1627 65 1666 67
rect 1700 65 1739 67
rect 1773 65 1812 67
rect 1846 65 1885 67
rect 1919 65 1958 99
rect 1992 65 2031 99
rect 2069 67 2103 101
rect 11861 135 11902 169
rect 11861 101 12004 135
rect 11882 67 12004 101
rect 2065 65 2104 67
rect 2138 65 2177 67
rect 2211 65 2250 67
rect 2284 65 2323 67
rect 11861 65 11893 67
rect 55 59 11893 65
rect -462 -217 -409 -183
rect -375 -217 -322 -183
rect -288 -217 -236 -183
rect -202 -217 -150 -183
rect -496 -293 -116 -217
rect -462 -327 -409 -293
rect -375 -327 -322 -293
rect -288 -327 -236 -293
rect -202 -327 -150 -293
rect 6402 -1153 8791 -1138
rect 6402 -1187 6483 -1153
rect 6517 -1154 6558 -1153
rect 6592 -1154 6633 -1153
rect 6667 -1154 6708 -1153
rect 6742 -1154 6783 -1153
rect 6817 -1154 6859 -1153
rect 6893 -1154 6935 -1153
rect 6969 -1154 7011 -1153
rect 7045 -1154 7087 -1153
rect 7121 -1154 7197 -1153
rect 7231 -1154 7271 -1153
rect 7305 -1154 7345 -1153
rect 7379 -1154 7419 -1153
rect 7453 -1154 7493 -1153
rect 7527 -1154 7567 -1153
rect 7601 -1154 7641 -1153
rect 7675 -1154 7715 -1153
rect 7749 -1154 7789 -1153
rect 7823 -1154 7863 -1153
rect 7897 -1154 7937 -1153
rect 7971 -1154 8011 -1153
rect 8045 -1154 8085 -1153
rect 8119 -1154 8159 -1153
rect 8193 -1154 8233 -1153
rect 8267 -1154 8307 -1153
rect 8341 -1154 8381 -1153
rect 8415 -1154 8455 -1153
rect 8489 -1154 8529 -1153
rect 8563 -1154 8604 -1153
rect 8638 -1154 8679 -1153
rect 6532 -1187 6558 -1154
rect 6600 -1187 6633 -1154
rect 6402 -1188 6498 -1187
rect 6532 -1188 6566 -1187
rect 6600 -1188 6634 -1187
rect 6668 -1188 6702 -1154
rect 6742 -1187 6770 -1154
rect 6817 -1187 6838 -1154
rect 6893 -1187 6906 -1154
rect 6969 -1187 6974 -1154
rect 6736 -1188 6770 -1187
rect 6804 -1188 6838 -1187
rect 6872 -1188 6906 -1187
rect 6940 -1188 6974 -1187
rect 7008 -1187 7011 -1154
rect 7076 -1187 7087 -1154
rect 7008 -1188 7042 -1187
rect 7076 -1188 7110 -1187
rect 7144 -1188 7178 -1154
rect 7231 -1187 7246 -1154
rect 7305 -1187 7314 -1154
rect 7379 -1187 7382 -1154
rect 7212 -1188 7246 -1187
rect 7280 -1188 7314 -1187
rect 7348 -1188 7382 -1187
rect 7416 -1187 7419 -1154
rect 7484 -1187 7493 -1154
rect 7552 -1187 7567 -1154
rect 7620 -1187 7641 -1154
rect 7688 -1187 7715 -1154
rect 7756 -1187 7789 -1154
rect 7416 -1188 7450 -1187
rect 7484 -1188 7518 -1187
rect 7552 -1188 7586 -1187
rect 7620 -1188 7654 -1187
rect 7688 -1188 7722 -1187
rect 7756 -1188 7790 -1187
rect 7824 -1188 7858 -1154
rect 7897 -1187 7926 -1154
rect 7971 -1187 7994 -1154
rect 8045 -1187 8062 -1154
rect 8119 -1187 8130 -1154
rect 8193 -1187 8198 -1154
rect 7892 -1188 7926 -1187
rect 7960 -1188 7994 -1187
rect 8028 -1188 8062 -1187
rect 8096 -1188 8130 -1187
rect 8164 -1188 8198 -1187
rect 8232 -1187 8233 -1154
rect 8300 -1187 8307 -1154
rect 8368 -1187 8381 -1154
rect 8436 -1187 8455 -1154
rect 8504 -1187 8529 -1154
rect 8572 -1187 8604 -1154
rect 8232 -1188 8266 -1187
rect 8300 -1188 8334 -1187
rect 8368 -1188 8402 -1187
rect 8436 -1188 8470 -1187
rect 8504 -1188 8538 -1187
rect 8572 -1188 8606 -1187
rect 8640 -1188 8674 -1154
rect 8713 -1187 8791 -1153
rect 8708 -1188 8791 -1187
rect 6402 -1202 8791 -1188
rect 6402 -1216 6466 -1202
rect 6402 -1256 6417 -1216
rect 6451 -1256 6466 -1216
rect 6402 -1290 6466 -1256
rect 8727 -1217 8791 -1202
rect 8727 -1251 8742 -1217
rect 8776 -1251 8791 -1217
rect 8727 -1262 8791 -1251
rect 6402 -1328 6417 -1290
rect 6451 -1328 6466 -1290
rect 6650 -1304 6652 -1270
rect 6700 -1304 6727 -1270
rect 6768 -1304 6802 -1270
rect 6836 -1304 6870 -1270
rect 6911 -1304 6938 -1270
rect 6986 -1304 7006 -1270
rect 7061 -1304 7074 -1270
rect 7136 -1304 7142 -1270
rect 7176 -1304 7177 -1270
rect 7244 -1304 7252 -1270
rect 7312 -1304 7327 -1270
rect 7380 -1304 7402 -1270
rect 7448 -1304 7476 -1270
rect 7516 -1304 7550 -1270
rect 7584 -1304 7618 -1270
rect 7658 -1304 7686 -1270
rect 7732 -1304 7754 -1270
rect 7806 -1304 7822 -1270
rect 7880 -1304 7890 -1270
rect 7954 -1304 7958 -1270
rect 7992 -1304 7994 -1270
rect 8060 -1304 8068 -1270
rect 8128 -1304 8142 -1270
rect 8196 -1304 8216 -1270
rect 8264 -1304 8290 -1270
rect 8332 -1304 8364 -1270
rect 8400 -1304 8434 -1270
rect 8472 -1304 8502 -1270
rect 8546 -1304 8570 -1270
rect 6402 -1358 6466 -1328
rect 6402 -1406 6417 -1358
rect 6451 -1406 6466 -1358
rect 6402 -1426 6466 -1406
rect 6402 -1484 6417 -1426
rect 6451 -1484 6466 -1426
rect 6402 -1494 6466 -1484
rect 6402 -1596 6417 -1494
rect 6451 -1596 6466 -1494
rect 6402 -1606 6466 -1596
rect 6402 -1640 6417 -1606
rect 6451 -1640 6466 -1606
rect 6402 -1684 6466 -1640
rect 6402 -1718 6417 -1684
rect 6451 -1718 6466 -1684
rect 6402 -1724 6466 -1718
rect 6402 -1758 6417 -1724
rect 6451 -1758 6466 -1724
rect 6402 -1762 6466 -1758
rect 6402 -1826 6417 -1762
rect 6451 -1826 6466 -1762
rect 6402 -1840 6466 -1826
rect 6402 -1894 6417 -1840
rect 6451 -1894 6466 -1840
rect 6534 -1327 6568 -1315
rect 6534 -1399 6568 -1365
rect 8727 -1324 8742 -1262
rect 8776 -1324 8791 -1262
rect 8727 -1330 8791 -1324
rect 8727 -1397 8742 -1330
rect 8776 -1397 8791 -1330
rect 8727 -1398 8791 -1397
rect 6534 -1472 6568 -1436
rect 6650 -1460 6652 -1426
rect 6700 -1460 6727 -1426
rect 6768 -1460 6802 -1426
rect 6836 -1460 6870 -1426
rect 6911 -1460 6938 -1426
rect 6986 -1460 7006 -1426
rect 7061 -1460 7074 -1426
rect 7136 -1460 7142 -1426
rect 7176 -1460 7177 -1426
rect 7244 -1460 7252 -1426
rect 7312 -1460 7327 -1426
rect 7380 -1460 7402 -1426
rect 7448 -1460 7476 -1426
rect 7516 -1460 7550 -1426
rect 7584 -1460 7618 -1426
rect 7658 -1460 7686 -1426
rect 7732 -1460 7754 -1426
rect 7806 -1460 7822 -1426
rect 7880 -1460 7890 -1426
rect 7954 -1460 7958 -1426
rect 7992 -1460 7994 -1426
rect 8060 -1460 8068 -1426
rect 8128 -1460 8142 -1426
rect 8196 -1460 8216 -1426
rect 8264 -1460 8290 -1426
rect 8332 -1460 8364 -1426
rect 8400 -1460 8434 -1426
rect 8472 -1460 8502 -1426
rect 8546 -1460 8570 -1426
rect 8727 -1432 8742 -1398
rect 8776 -1432 8791 -1398
rect 8727 -1436 8791 -1432
rect 6534 -1545 6568 -1507
rect 6534 -1617 6568 -1579
rect 8727 -1500 8742 -1436
rect 8776 -1500 8791 -1436
rect 8727 -1509 8791 -1500
rect 8727 -1568 8742 -1509
rect 8776 -1568 8791 -1509
rect 8727 -1582 8791 -1568
rect 6650 -1616 6652 -1582
rect 6700 -1616 6727 -1582
rect 6768 -1616 6802 -1582
rect 6836 -1616 6870 -1582
rect 6911 -1616 6938 -1582
rect 6986 -1616 7006 -1582
rect 7061 -1616 7074 -1582
rect 7136 -1616 7142 -1582
rect 7176 -1616 7177 -1582
rect 7244 -1616 7252 -1582
rect 7312 -1616 7327 -1582
rect 7380 -1616 7402 -1582
rect 7448 -1616 7476 -1582
rect 7516 -1616 7550 -1582
rect 7584 -1616 7618 -1582
rect 7658 -1616 7686 -1582
rect 7732 -1616 7754 -1582
rect 7806 -1616 7822 -1582
rect 7880 -1616 7890 -1582
rect 7954 -1616 7958 -1582
rect 7992 -1616 7994 -1582
rect 8060 -1616 8068 -1582
rect 8128 -1616 8142 -1582
rect 8196 -1616 8216 -1582
rect 8264 -1616 8290 -1582
rect 8332 -1616 8364 -1582
rect 8400 -1616 8434 -1582
rect 8472 -1616 8502 -1582
rect 8546 -1616 8570 -1582
rect 6534 -1689 6568 -1652
rect 6534 -1761 6568 -1725
rect 8727 -1636 8742 -1582
rect 8776 -1636 8791 -1582
rect 8727 -1655 8791 -1636
rect 8727 -1704 8742 -1655
rect 8776 -1704 8791 -1655
rect 8727 -1728 8791 -1704
rect 6650 -1772 6652 -1738
rect 6700 -1772 6727 -1738
rect 6768 -1772 6802 -1738
rect 6836 -1772 6870 -1738
rect 6911 -1772 6938 -1738
rect 6986 -1772 7006 -1738
rect 7061 -1772 7074 -1738
rect 7136 -1772 7142 -1738
rect 7176 -1772 7177 -1738
rect 7244 -1772 7252 -1738
rect 7312 -1772 7327 -1738
rect 7380 -1772 7402 -1738
rect 7448 -1772 7476 -1738
rect 7516 -1772 7550 -1738
rect 7584 -1772 7618 -1738
rect 7658 -1772 7686 -1738
rect 7732 -1772 7754 -1738
rect 7806 -1772 7822 -1738
rect 7880 -1772 7890 -1738
rect 7954 -1772 7958 -1738
rect 7992 -1772 7994 -1738
rect 8060 -1772 8068 -1738
rect 8128 -1772 8142 -1738
rect 8196 -1772 8216 -1738
rect 8264 -1772 8290 -1738
rect 8332 -1772 8364 -1738
rect 8400 -1772 8434 -1738
rect 8472 -1772 8502 -1738
rect 8546 -1772 8570 -1738
rect 8727 -1772 8742 -1728
rect 8776 -1772 8791 -1728
rect 6534 -1833 6568 -1798
rect 6534 -1883 6568 -1871
rect 8727 -1801 8791 -1772
rect 8727 -1840 8742 -1801
rect 8776 -1840 8791 -1801
rect 8727 -1874 8791 -1840
rect 6402 -1918 6466 -1894
rect 6402 -1962 6417 -1918
rect 6451 -1962 6466 -1918
rect 6650 -1928 6652 -1894
rect 6700 -1928 6727 -1894
rect 6768 -1928 6802 -1894
rect 6836 -1928 6870 -1894
rect 6911 -1928 6938 -1894
rect 6986 -1928 7006 -1894
rect 7061 -1928 7074 -1894
rect 7136 -1928 7142 -1894
rect 7176 -1928 7177 -1894
rect 7244 -1928 7252 -1894
rect 7312 -1928 7327 -1894
rect 7380 -1928 7402 -1894
rect 7448 -1928 7476 -1894
rect 7516 -1928 7550 -1894
rect 7584 -1928 7618 -1894
rect 7658 -1928 7686 -1894
rect 7732 -1928 7754 -1894
rect 7806 -1928 7822 -1894
rect 7880 -1928 7890 -1894
rect 7954 -1928 7958 -1894
rect 7992 -1928 7994 -1894
rect 8060 -1928 8068 -1894
rect 8128 -1928 8142 -1894
rect 8196 -1928 8216 -1894
rect 8264 -1928 8290 -1894
rect 8332 -1928 8364 -1894
rect 8400 -1928 8434 -1894
rect 8472 -1928 8502 -1894
rect 8546 -1928 8570 -1894
rect 8727 -1908 8742 -1874
rect 8776 -1908 8791 -1874
rect 6402 -1971 6466 -1962
rect 8727 -1942 8791 -1908
rect 6402 -1986 6721 -1971
rect 6402 -2020 6480 -1986
rect 6514 -2010 6581 -1986
rect 6615 -1995 6721 -1986
rect 8727 -1981 8742 -1942
rect 8776 -1981 8791 -1942
rect 8727 -1995 8791 -1981
rect 6615 -2010 8791 -1995
rect 6402 -2035 6485 -2020
rect 6417 -2044 6485 -2035
rect 6519 -2044 6553 -2010
rect 6615 -2020 6621 -2010
rect 6587 -2044 6621 -2020
rect 6655 -2044 6689 -2010
rect 6723 -2044 6735 -2010
rect 6791 -2044 6807 -2010
rect 6859 -2044 6879 -2010
rect 6927 -2044 6951 -2010
rect 6995 -2044 7023 -2010
rect 7063 -2044 7095 -2010
rect 7131 -2044 7165 -2010
rect 7201 -2044 7233 -2010
rect 7273 -2044 7301 -2010
rect 7345 -2044 7369 -2010
rect 7417 -2044 7437 -2010
rect 7489 -2044 7505 -2010
rect 7561 -2044 7573 -2010
rect 7633 -2044 7641 -2010
rect 7705 -2044 7709 -2010
rect 7811 -2044 7815 -2010
rect 7879 -2044 7887 -2010
rect 7947 -2044 7959 -2010
rect 8015 -2044 8031 -2010
rect 8083 -2044 8103 -2010
rect 8151 -2044 8175 -2010
rect 8219 -2044 8247 -2010
rect 8287 -2044 8319 -2010
rect 8355 -2044 8389 -2010
rect 8425 -2044 8457 -2010
rect 8497 -2044 8525 -2010
rect 8569 -2044 8593 -2010
rect 8641 -2044 8661 -2010
rect 8713 -2044 8791 -2010
rect 6657 -2059 8791 -2044
<< viali >>
rect -496 1395 -462 1429
rect -409 1395 -375 1429
rect -322 1395 -288 1429
rect -236 1395 -202 1429
rect -150 1395 -116 1429
rect -496 1285 -462 1319
rect -409 1285 -375 1319
rect -322 1285 -288 1319
rect -236 1285 -202 1319
rect -150 1285 -116 1319
rect 61 1378 63 1412
rect 63 1378 95 1412
rect 133 1378 165 1412
rect 165 1378 167 1412
rect 61 1305 63 1339
rect 63 1305 95 1339
rect 133 1305 165 1339
rect 165 1305 167 1339
rect 61 1232 63 1266
rect 63 1232 95 1266
rect 133 1232 165 1266
rect 165 1232 167 1266
rect 61 1159 63 1193
rect 63 1159 95 1193
rect 133 1159 165 1193
rect 165 1159 167 1193
rect 61 1086 63 1120
rect 63 1086 95 1120
rect 133 1086 165 1120
rect 165 1086 167 1120
rect 61 1013 63 1047
rect 63 1013 95 1047
rect 133 1013 165 1047
rect 165 1013 167 1047
rect 61 940 63 974
rect 63 940 95 974
rect 133 940 165 974
rect 165 940 167 974
rect 61 867 63 901
rect 63 867 95 901
rect 133 867 165 901
rect 165 867 167 901
rect 61 794 63 828
rect 63 794 95 828
rect 133 794 165 828
rect 165 794 167 828
rect 61 721 63 755
rect 63 721 95 755
rect 133 721 165 755
rect 165 721 167 755
rect -497 623 -463 657
rect -410 623 -376 657
rect -323 623 -289 657
rect -236 623 -202 657
rect -150 623 -116 657
rect -497 545 -463 579
rect -410 545 -376 579
rect -323 545 -289 579
rect -236 545 -202 579
rect -150 545 -116 579
rect -497 467 -463 501
rect -410 467 -376 501
rect -323 467 -289 501
rect -236 467 -202 501
rect -150 467 -116 501
rect 61 648 63 682
rect 63 648 95 682
rect 133 648 165 682
rect 165 648 167 682
rect 61 575 63 609
rect 63 575 95 609
rect 133 575 165 609
rect 165 575 167 609
rect 61 502 63 536
rect 63 502 95 536
rect 133 502 165 536
rect 165 502 167 536
rect 61 429 63 463
rect 63 429 95 463
rect 133 429 165 463
rect 165 429 167 463
rect 61 356 63 390
rect 63 356 95 390
rect 133 356 165 390
rect 165 356 167 390
rect 61 283 63 317
rect 63 283 95 317
rect 133 283 165 317
rect 165 283 167 317
rect 402 1403 436 1437
rect 480 1403 514 1437
rect 558 1403 592 1437
rect 636 1403 670 1437
rect 714 1403 748 1437
rect 792 1403 826 1437
rect 870 1403 904 1437
rect 949 1403 983 1437
rect 324 1331 358 1365
rect 396 1331 430 1365
rect 480 1351 514 1365
rect 558 1351 592 1365
rect 636 1351 670 1365
rect 714 1351 748 1365
rect 792 1351 826 1365
rect 870 1351 904 1365
rect 949 1351 983 1365
rect 1059 1351 1597 1437
rect 1636 1403 1670 1437
rect 1636 1351 1670 1365
rect 480 1331 492 1351
rect 492 1331 514 1351
rect 558 1331 560 1351
rect 560 1331 592 1351
rect 636 1331 662 1351
rect 662 1331 670 1351
rect 714 1331 730 1351
rect 730 1331 748 1351
rect 792 1331 798 1351
rect 798 1331 826 1351
rect 870 1331 900 1351
rect 900 1331 904 1351
rect 949 1331 968 1351
rect 968 1331 983 1351
rect 1059 1331 1131 1351
rect 1131 1331 1165 1351
rect 1165 1331 1199 1351
rect 1199 1331 1233 1351
rect 1233 1331 1267 1351
rect 1267 1331 1301 1351
rect 1301 1331 1335 1351
rect 1335 1331 1369 1351
rect 1369 1331 1403 1351
rect 1403 1331 1437 1351
rect 1437 1331 1471 1351
rect 1471 1331 1505 1351
rect 1505 1331 1539 1351
rect 1539 1331 1573 1351
rect 1573 1331 1597 1351
rect 1636 1331 1641 1351
rect 1641 1331 1670 1351
rect 1708 1329 1742 1363
rect 324 1256 358 1290
rect 396 1256 430 1290
rect 1636 1255 1670 1289
rect 1708 1255 1742 1289
rect 566 1232 600 1235
rect 641 1232 675 1235
rect 716 1232 750 1235
rect 791 1232 825 1235
rect 866 1232 900 1235
rect 940 1232 974 1235
rect 1014 1232 1048 1235
rect 1088 1232 1122 1235
rect 1162 1232 1196 1235
rect 1236 1232 1270 1235
rect 1310 1232 1344 1235
rect 1384 1232 1418 1235
rect 1458 1232 1492 1235
rect 324 1181 358 1215
rect 396 1181 430 1215
rect 566 1201 570 1232
rect 570 1201 600 1232
rect 641 1201 672 1232
rect 672 1201 675 1232
rect 716 1201 740 1232
rect 740 1201 750 1232
rect 791 1201 808 1232
rect 808 1201 825 1232
rect 866 1201 876 1232
rect 876 1201 900 1232
rect 940 1201 944 1232
rect 944 1201 974 1232
rect 1014 1201 1046 1232
rect 1046 1201 1048 1232
rect 1088 1201 1114 1232
rect 1114 1201 1122 1232
rect 1162 1201 1182 1232
rect 1182 1201 1196 1232
rect 1236 1201 1250 1232
rect 1250 1201 1270 1232
rect 1310 1201 1318 1232
rect 1318 1201 1344 1232
rect 1384 1201 1386 1232
rect 1386 1201 1418 1232
rect 1458 1201 1488 1232
rect 1488 1201 1492 1232
rect 324 1106 358 1140
rect 396 1106 430 1140
rect 324 1031 358 1065
rect 396 1031 430 1065
rect 324 956 358 990
rect 396 956 430 990
rect 324 881 358 915
rect 396 881 430 915
rect 324 807 358 841
rect 396 807 430 841
rect 324 733 358 767
rect 396 733 430 767
rect 324 659 358 693
rect 396 659 430 693
rect 324 585 358 619
rect 396 585 430 619
rect 324 511 358 545
rect 396 511 430 545
rect 476 1171 510 1175
rect 476 1141 510 1171
rect 476 1101 510 1102
rect 476 1068 510 1101
rect 1636 1181 1670 1215
rect 1708 1181 1742 1215
rect 1636 1107 1670 1141
rect 1708 1107 1742 1141
rect 1124 1042 1148 1076
rect 1148 1042 1158 1076
rect 1202 1042 1216 1076
rect 1216 1042 1236 1076
rect 1280 1042 1284 1076
rect 1284 1042 1314 1076
rect 1358 1042 1386 1076
rect 1386 1042 1392 1076
rect 1435 1042 1454 1076
rect 1454 1042 1469 1076
rect 1512 1042 1546 1076
rect 476 997 510 1029
rect 476 995 510 997
rect 476 927 510 956
rect 476 922 510 927
rect 1636 1033 1670 1067
rect 1708 1033 1742 1067
rect 1636 959 1670 993
rect 1708 959 1742 993
rect 566 920 600 921
rect 641 920 675 921
rect 716 920 750 921
rect 791 920 825 921
rect 866 920 900 921
rect 940 920 974 921
rect 1014 920 1048 921
rect 1088 920 1122 921
rect 1162 920 1196 921
rect 1236 920 1270 921
rect 1310 920 1344 921
rect 1384 920 1418 921
rect 1458 920 1492 921
rect 566 887 570 920
rect 570 887 600 920
rect 641 887 672 920
rect 672 887 675 920
rect 716 887 740 920
rect 740 887 750 920
rect 791 887 808 920
rect 808 887 825 920
rect 866 887 876 920
rect 876 887 900 920
rect 940 887 944 920
rect 944 887 974 920
rect 1014 887 1046 920
rect 1046 887 1048 920
rect 1088 887 1114 920
rect 1114 887 1122 920
rect 1162 887 1182 920
rect 1182 887 1196 920
rect 1236 887 1250 920
rect 1250 887 1270 920
rect 1310 887 1318 920
rect 1318 887 1344 920
rect 1384 887 1386 920
rect 1386 887 1418 920
rect 1458 887 1488 920
rect 1488 887 1492 920
rect 476 857 510 883
rect 476 849 510 857
rect 476 787 510 810
rect 1636 885 1670 919
rect 1708 885 1742 919
rect 1636 811 1670 845
rect 1708 811 1742 845
rect 476 776 510 787
rect 566 756 570 790
rect 570 756 600 790
rect 641 756 672 790
rect 672 756 675 790
rect 716 756 740 790
rect 740 756 750 790
rect 791 756 808 790
rect 808 756 825 790
rect 866 756 876 790
rect 876 756 900 790
rect 940 756 944 790
rect 944 756 974 790
rect 1014 756 1046 790
rect 1046 756 1048 790
rect 1088 756 1114 790
rect 1114 756 1122 790
rect 1162 756 1182 790
rect 1182 756 1196 790
rect 1236 756 1250 790
rect 1250 756 1270 790
rect 1310 756 1318 790
rect 1318 756 1344 790
rect 1384 756 1386 790
rect 1386 756 1418 790
rect 1458 756 1488 790
rect 1488 756 1492 790
rect 476 717 510 738
rect 476 704 510 717
rect 476 647 510 666
rect 476 632 510 647
rect 1636 736 1670 770
rect 1708 736 1742 770
rect 1636 661 1670 695
rect 1708 661 1742 695
rect 1123 600 1148 634
rect 1148 600 1157 634
rect 1201 600 1216 634
rect 1216 600 1235 634
rect 1279 600 1284 634
rect 1284 600 1313 634
rect 1357 600 1386 634
rect 1386 600 1391 634
rect 1435 600 1454 634
rect 1454 600 1469 634
rect 1512 600 1546 634
rect 476 576 510 594
rect 476 560 510 576
rect 476 505 510 522
rect 476 488 510 505
rect 1636 586 1670 620
rect 1708 586 1742 620
rect 1636 511 1670 545
rect 1708 511 1742 545
rect 324 437 358 471
rect 396 437 430 471
rect 641 444 672 478
rect 672 444 675 478
rect 716 444 740 478
rect 740 444 750 478
rect 791 444 808 478
rect 808 444 825 478
rect 866 444 876 478
rect 876 444 900 478
rect 940 444 944 478
rect 944 444 974 478
rect 1014 444 1046 478
rect 1046 444 1048 478
rect 1088 444 1114 478
rect 1114 444 1122 478
rect 1162 444 1182 478
rect 1182 444 1196 478
rect 1236 444 1250 478
rect 1250 444 1270 478
rect 1310 444 1318 478
rect 1318 444 1344 478
rect 1384 444 1386 478
rect 1386 444 1418 478
rect 1458 444 1488 478
rect 1488 444 1492 478
rect 1636 436 1670 470
rect 1708 436 1742 470
rect 324 363 358 397
rect 396 361 430 395
rect 469 361 503 395
rect 542 361 576 395
rect 615 361 649 395
rect 688 361 722 395
rect 761 361 795 395
rect 834 361 868 395
rect 907 361 941 395
rect 980 361 1014 395
rect 1053 361 1087 395
rect 1126 361 1160 395
rect 1199 361 1233 395
rect 1272 361 1306 395
rect 1345 361 1379 395
rect 1418 361 1452 395
rect 1491 361 1525 395
rect 1564 359 1670 395
rect 1708 361 1742 395
rect 1564 325 1581 359
rect 1581 325 1615 359
rect 1615 325 1670 359
rect 396 289 430 323
rect 469 289 503 323
rect 542 289 576 323
rect 615 289 649 323
rect 688 289 722 323
rect 761 289 795 323
rect 834 289 868 323
rect 907 289 941 323
rect 980 289 1014 323
rect 1053 289 1087 323
rect 1126 289 1160 323
rect 1199 289 1233 323
rect 1272 289 1306 323
rect 1345 289 1379 323
rect 1418 289 1452 323
rect 1491 289 1525 323
rect 1564 289 1670 325
rect 1904 1389 1906 1423
rect 1906 1389 1938 1423
rect 1976 1389 2008 1423
rect 2008 1389 2010 1423
rect 1904 1315 1906 1349
rect 1906 1315 1938 1349
rect 1976 1315 2008 1349
rect 2008 1315 2010 1349
rect 1904 1241 1906 1275
rect 1906 1241 1938 1275
rect 1976 1241 2008 1275
rect 2008 1241 2010 1275
rect 1904 1167 1906 1201
rect 1906 1167 1938 1201
rect 1976 1167 2008 1201
rect 2008 1167 2010 1201
rect 1904 1093 1906 1127
rect 1906 1093 1938 1127
rect 1976 1093 2008 1127
rect 2008 1093 2010 1127
rect 1904 1019 1906 1053
rect 1906 1019 1938 1053
rect 1976 1019 2008 1053
rect 2008 1019 2010 1053
rect 1904 945 1906 979
rect 1906 945 1938 979
rect 1976 945 2008 979
rect 2008 945 2010 979
rect 1904 871 1906 905
rect 1906 871 1938 905
rect 1976 871 2008 905
rect 2008 871 2010 905
rect 1904 797 1906 831
rect 1906 797 1938 831
rect 1976 797 2008 831
rect 2008 797 2010 831
rect 1904 723 1906 757
rect 1906 723 1938 757
rect 1976 723 2008 757
rect 2008 723 2010 757
rect 1904 649 1906 683
rect 1906 649 1938 683
rect 1976 649 2008 683
rect 2008 649 2010 683
rect 1904 575 1906 609
rect 1906 575 1938 609
rect 1976 575 2008 609
rect 2008 575 2010 609
rect 1904 501 1906 535
rect 1906 501 1938 535
rect 1976 501 2008 535
rect 2008 501 2010 535
rect 1904 428 1906 462
rect 1906 428 1938 462
rect 1976 428 2008 462
rect 2008 428 2010 462
rect 1904 355 1906 389
rect 1906 355 1938 389
rect 1976 355 2008 389
rect 2008 355 2010 389
rect 61 210 63 244
rect 63 210 95 244
rect 133 210 165 244
rect 165 210 167 244
rect 1904 282 1906 316
rect 1906 282 1938 316
rect 1976 282 2008 316
rect 2008 282 2010 316
rect 2237 1416 2271 1450
rect 2315 1416 2349 1450
rect 2393 1416 2427 1450
rect 2471 1416 2505 1450
rect 2549 1416 2583 1450
rect 2627 1416 2661 1450
rect 2705 1416 2739 1450
rect 2784 1416 2818 1450
rect 2894 1416 2928 1450
rect 2967 1416 3001 1450
rect 3040 1416 3074 1450
rect 3113 1416 3147 1450
rect 3186 1416 3220 1450
rect 3259 1416 3293 1450
rect 3332 1416 3366 1450
rect 3405 1416 3439 1450
rect 3478 1416 3512 1450
rect 3551 1416 3585 1450
rect 3624 1416 3658 1450
rect 3697 1416 3731 1450
rect 3770 1416 3804 1450
rect 3843 1416 3877 1450
rect 3916 1416 3950 1450
rect 3989 1416 4023 1450
rect 4062 1416 4096 1450
rect 4135 1416 4169 1450
rect 4208 1416 4242 1450
rect 4281 1416 4315 1450
rect 4354 1416 4388 1450
rect 4427 1416 4461 1450
rect 4500 1416 4534 1450
rect 4573 1416 4607 1450
rect 4646 1416 4680 1450
rect 4719 1416 4753 1450
rect 4792 1416 4826 1450
rect 4865 1416 4899 1450
rect 4938 1416 4972 1450
rect 5011 1416 5045 1450
rect 5084 1416 5118 1450
rect 5157 1416 5191 1450
rect 5230 1416 5264 1450
rect 5303 1416 5337 1450
rect 5376 1416 5410 1450
rect 5449 1416 5483 1450
rect 5522 1416 5556 1450
rect 5595 1416 5629 1450
rect 5668 1416 5702 1450
rect 5741 1416 5775 1450
rect 5814 1416 5848 1450
rect 5887 1416 5921 1450
rect 5961 1416 5995 1450
rect 6035 1416 6069 1450
rect 6109 1416 6143 1450
rect 6183 1416 6217 1450
rect 6257 1416 6291 1450
rect 6331 1416 6365 1450
rect 6405 1416 6439 1450
rect 6479 1416 6513 1450
rect 6553 1416 6587 1450
rect 6627 1416 6661 1450
rect 2159 1344 2193 1378
rect 2231 1344 2265 1378
rect 2315 1377 2349 1378
rect 2393 1377 2427 1378
rect 2471 1377 2505 1378
rect 2549 1377 2583 1378
rect 2627 1377 2661 1378
rect 2705 1377 2739 1378
rect 2784 1377 2818 1378
rect 2894 1377 2928 1378
rect 2967 1377 3001 1378
rect 3040 1377 3074 1378
rect 3113 1377 3147 1378
rect 3186 1377 3220 1378
rect 3259 1377 3293 1378
rect 3332 1377 3366 1378
rect 3405 1377 3439 1378
rect 3478 1377 3512 1378
rect 3551 1377 3585 1378
rect 3624 1377 3658 1378
rect 3697 1377 3731 1378
rect 3770 1377 3804 1378
rect 3843 1377 3877 1378
rect 3916 1377 3950 1378
rect 3989 1377 4023 1378
rect 4062 1377 4096 1378
rect 4135 1377 4169 1378
rect 4208 1377 4242 1378
rect 4281 1377 4315 1378
rect 4354 1377 4388 1378
rect 4427 1377 4461 1378
rect 2315 1344 2321 1377
rect 2321 1344 2349 1377
rect 2393 1344 2423 1377
rect 2423 1344 2427 1377
rect 2471 1344 2491 1377
rect 2491 1344 2505 1377
rect 2549 1344 2559 1377
rect 2559 1344 2583 1377
rect 2627 1344 2661 1377
rect 2705 1344 2729 1377
rect 2729 1344 2739 1377
rect 2784 1344 2797 1377
rect 2797 1344 2818 1377
rect 2894 1344 2899 1377
rect 2899 1344 2928 1377
rect 2967 1344 3001 1377
rect 3040 1344 3069 1377
rect 3069 1344 3074 1377
rect 3113 1344 3137 1377
rect 3137 1344 3147 1377
rect 3186 1344 3205 1377
rect 3205 1344 3220 1377
rect 3259 1344 3273 1377
rect 3273 1344 3293 1377
rect 3332 1344 3341 1377
rect 3341 1344 3366 1377
rect 3405 1344 3409 1377
rect 3409 1344 3439 1377
rect 3478 1344 3511 1377
rect 3511 1344 3512 1377
rect 3551 1344 3579 1377
rect 3579 1344 3585 1377
rect 3624 1344 3647 1377
rect 3647 1344 3658 1377
rect 3697 1344 3715 1377
rect 3715 1344 3731 1377
rect 3770 1344 3783 1377
rect 3783 1344 3804 1377
rect 3843 1344 3851 1377
rect 3851 1344 3877 1377
rect 3916 1344 3919 1377
rect 3919 1344 3950 1377
rect 3989 1344 4021 1377
rect 4021 1344 4023 1377
rect 4062 1344 4089 1377
rect 4089 1344 4096 1377
rect 4135 1344 4157 1377
rect 4157 1344 4169 1377
rect 4208 1344 4225 1377
rect 4225 1344 4242 1377
rect 4281 1344 4293 1377
rect 4293 1344 4315 1377
rect 4354 1344 4361 1377
rect 4361 1344 4388 1377
rect 4427 1344 4429 1377
rect 4429 1344 4461 1377
rect 4500 1377 4534 1378
rect 4573 1377 4607 1378
rect 4646 1377 4680 1378
rect 4719 1377 4753 1378
rect 4792 1377 4826 1378
rect 4865 1377 4899 1378
rect 4938 1377 4972 1378
rect 5011 1377 5045 1378
rect 5084 1377 5118 1378
rect 5157 1377 5191 1378
rect 5230 1377 5264 1378
rect 5303 1377 5337 1378
rect 5376 1377 5410 1378
rect 5449 1377 5483 1378
rect 5522 1377 5556 1378
rect 5595 1377 5629 1378
rect 5668 1377 5702 1378
rect 5741 1377 5775 1378
rect 5814 1377 5848 1378
rect 5887 1377 5921 1378
rect 5961 1377 5995 1378
rect 6035 1377 6069 1378
rect 6109 1377 6143 1378
rect 6183 1377 6217 1378
rect 6257 1377 6291 1378
rect 6331 1377 6365 1378
rect 6405 1377 6439 1378
rect 6479 1377 6513 1378
rect 6553 1377 6587 1378
rect 6627 1377 6733 1378
rect 4500 1344 4510 1377
rect 4510 1344 4534 1377
rect 4573 1344 4578 1377
rect 4578 1344 4607 1377
rect 4646 1344 4680 1377
rect 4719 1344 4748 1377
rect 4748 1344 4753 1377
rect 4792 1344 4816 1377
rect 4816 1344 4826 1377
rect 4865 1344 4884 1377
rect 4884 1344 4899 1377
rect 4938 1344 4952 1377
rect 4952 1344 4972 1377
rect 5011 1344 5020 1377
rect 5020 1344 5045 1377
rect 5084 1344 5088 1377
rect 5088 1344 5118 1377
rect 5157 1344 5190 1377
rect 5190 1344 5191 1377
rect 5230 1344 5258 1377
rect 5258 1344 5264 1377
rect 5303 1344 5326 1377
rect 5326 1344 5337 1377
rect 5376 1344 5394 1377
rect 5394 1344 5410 1377
rect 5449 1344 5462 1377
rect 5462 1344 5483 1377
rect 5522 1344 5530 1377
rect 5530 1344 5556 1377
rect 5595 1344 5598 1377
rect 5598 1344 5629 1377
rect 5668 1344 5700 1377
rect 5700 1344 5702 1377
rect 5741 1344 5768 1377
rect 5768 1344 5775 1377
rect 5814 1344 5836 1377
rect 5836 1344 5848 1377
rect 5887 1344 5904 1377
rect 5904 1344 5921 1377
rect 5961 1344 5972 1377
rect 5972 1344 5995 1377
rect 6035 1344 6040 1377
rect 6040 1344 6069 1377
rect 6109 1344 6142 1377
rect 6142 1344 6143 1377
rect 6183 1344 6210 1377
rect 6210 1344 6217 1377
rect 6257 1344 6278 1377
rect 6278 1344 6291 1377
rect 6331 1344 6346 1377
rect 6346 1344 6365 1377
rect 6405 1344 6414 1377
rect 6414 1344 6439 1377
rect 6479 1344 6482 1377
rect 6482 1344 6513 1377
rect 6553 1344 6584 1377
rect 6584 1344 6587 1377
rect 6627 1343 6652 1377
rect 6652 1343 6733 1377
rect 2159 1271 2193 1305
rect 2231 1271 2265 1305
rect 2159 1198 2193 1232
rect 2231 1198 2265 1232
rect 2401 1224 2405 1258
rect 2405 1224 2435 1258
rect 2475 1224 2507 1258
rect 2507 1224 2509 1258
rect 2549 1224 2575 1258
rect 2575 1224 2583 1258
rect 2623 1224 2643 1258
rect 2643 1224 2657 1258
rect 2697 1224 2711 1258
rect 2711 1224 2731 1258
rect 2771 1224 2779 1258
rect 2779 1224 2805 1258
rect 2845 1224 2847 1258
rect 2847 1224 2879 1258
rect 2919 1224 2949 1258
rect 2949 1224 2953 1258
rect 2993 1224 3017 1258
rect 3017 1224 3027 1258
rect 3067 1224 3085 1258
rect 3085 1224 3101 1258
rect 3141 1224 3153 1258
rect 3153 1224 3175 1258
rect 3215 1224 3221 1258
rect 3221 1224 3249 1258
rect 3289 1224 3323 1258
rect 3363 1224 3391 1258
rect 3391 1224 3397 1258
rect 3437 1224 3459 1258
rect 3459 1224 3471 1258
rect 3510 1224 3527 1258
rect 3527 1224 3544 1258
rect 3583 1224 3595 1258
rect 3595 1224 3617 1258
rect 3656 1224 3663 1258
rect 3663 1224 3690 1258
rect 3729 1224 3731 1258
rect 3731 1224 3763 1258
rect 3802 1224 3833 1258
rect 3833 1224 3836 1258
rect 3875 1224 3901 1258
rect 3901 1224 3909 1258
rect 3948 1224 3969 1258
rect 3969 1224 3982 1258
rect 4021 1224 4037 1258
rect 4037 1224 4055 1258
rect 4094 1224 4105 1258
rect 4105 1224 4128 1258
rect 4167 1224 4173 1258
rect 4173 1224 4201 1258
rect 4240 1224 4241 1258
rect 4241 1224 4274 1258
rect 4313 1224 4343 1258
rect 4343 1224 4347 1258
rect 4545 1224 4549 1258
rect 4549 1224 4579 1258
rect 4618 1224 4651 1258
rect 4651 1224 4652 1258
rect 4691 1224 4719 1258
rect 4719 1224 4725 1258
rect 4764 1224 4787 1258
rect 4787 1224 4798 1258
rect 4837 1224 4855 1258
rect 4855 1224 4871 1258
rect 4910 1224 4923 1258
rect 4923 1224 4944 1258
rect 4983 1224 4991 1258
rect 4991 1224 5017 1258
rect 5056 1224 5059 1258
rect 5059 1224 5090 1258
rect 5129 1224 5161 1258
rect 5161 1224 5163 1258
rect 5202 1224 5229 1258
rect 5229 1224 5236 1258
rect 5275 1224 5297 1258
rect 5297 1224 5309 1258
rect 5348 1224 5365 1258
rect 5365 1224 5382 1258
rect 5421 1224 5433 1258
rect 5433 1224 5455 1258
rect 5495 1224 5501 1258
rect 5501 1224 5529 1258
rect 5569 1224 5603 1258
rect 5643 1224 5671 1258
rect 5671 1224 5677 1258
rect 5717 1224 5739 1258
rect 5739 1224 5751 1258
rect 5791 1224 5807 1258
rect 5807 1224 5825 1258
rect 5865 1224 5875 1258
rect 5875 1224 5899 1258
rect 5939 1224 5943 1258
rect 5943 1224 5973 1258
rect 6013 1224 6045 1258
rect 6045 1224 6047 1258
rect 6087 1224 6113 1258
rect 6113 1224 6121 1258
rect 6161 1224 6181 1258
rect 6181 1224 6195 1258
rect 6235 1224 6249 1258
rect 6249 1224 6269 1258
rect 6309 1224 6317 1258
rect 6317 1224 6343 1258
rect 6383 1224 6385 1258
rect 6385 1224 6417 1258
rect 6457 1224 6487 1258
rect 6487 1224 6491 1258
rect 2159 1125 2193 1159
rect 2231 1125 2265 1159
rect 2159 1052 2193 1086
rect 2231 1052 2265 1086
rect 2159 979 2193 1013
rect 2231 979 2265 1013
rect 2159 906 2193 940
rect 2231 906 2265 940
rect 2159 833 2193 867
rect 2231 833 2265 867
rect 2159 760 2193 794
rect 2231 760 2265 794
rect 2159 687 2193 721
rect 2231 687 2265 721
rect 2159 614 2193 648
rect 2231 614 2265 648
rect 2159 541 2193 575
rect 2231 541 2265 575
rect 2159 496 2265 502
rect 2159 462 2195 496
rect 2195 462 2229 496
rect 2229 462 2265 496
rect 2159 428 2265 462
rect 2159 394 2195 428
rect 2195 394 2229 428
rect 2229 394 2265 428
rect 2159 359 2265 394
rect 2311 1197 2345 1201
rect 2311 1167 2345 1197
rect 2311 1090 2345 1120
rect 6547 1197 6581 1201
rect 6547 1167 6581 1197
rect 2311 1086 2345 1090
rect 2401 1068 2405 1102
rect 2405 1068 2435 1102
rect 2475 1068 2507 1102
rect 2507 1068 2509 1102
rect 2549 1068 2575 1102
rect 2575 1068 2583 1102
rect 2623 1068 2643 1102
rect 2643 1068 2657 1102
rect 2697 1068 2711 1102
rect 2711 1068 2731 1102
rect 2771 1068 2779 1102
rect 2779 1068 2805 1102
rect 2845 1068 2847 1102
rect 2847 1068 2879 1102
rect 2919 1068 2949 1102
rect 2949 1068 2953 1102
rect 2993 1068 3017 1102
rect 3017 1068 3027 1102
rect 3067 1068 3085 1102
rect 3085 1068 3101 1102
rect 3141 1068 3153 1102
rect 3153 1068 3175 1102
rect 3215 1068 3221 1102
rect 3221 1068 3249 1102
rect 3289 1068 3323 1102
rect 3363 1068 3391 1102
rect 3391 1068 3397 1102
rect 3437 1068 3459 1102
rect 3459 1068 3471 1102
rect 3510 1068 3527 1102
rect 3527 1068 3544 1102
rect 3583 1068 3595 1102
rect 3595 1068 3617 1102
rect 3656 1068 3663 1102
rect 3663 1068 3690 1102
rect 3729 1068 3731 1102
rect 3731 1068 3763 1102
rect 3802 1068 3833 1102
rect 3833 1068 3836 1102
rect 3875 1068 3901 1102
rect 3901 1068 3909 1102
rect 3948 1068 3969 1102
rect 3969 1068 3982 1102
rect 4021 1068 4037 1102
rect 4037 1068 4055 1102
rect 4094 1068 4105 1102
rect 4105 1068 4128 1102
rect 4167 1068 4173 1102
rect 4173 1068 4201 1102
rect 4240 1068 4241 1102
rect 4241 1068 4274 1102
rect 4313 1068 4343 1102
rect 4343 1068 4347 1102
rect 4545 1068 4549 1102
rect 4549 1068 4579 1102
rect 4618 1068 4651 1102
rect 4651 1068 4652 1102
rect 4691 1068 4719 1102
rect 4719 1068 4725 1102
rect 4764 1068 4787 1102
rect 4787 1068 4798 1102
rect 4837 1068 4855 1102
rect 4855 1068 4871 1102
rect 4910 1068 4923 1102
rect 4923 1068 4944 1102
rect 4983 1068 4991 1102
rect 4991 1068 5017 1102
rect 5056 1068 5059 1102
rect 5059 1068 5090 1102
rect 5129 1068 5161 1102
rect 5161 1068 5163 1102
rect 5202 1068 5229 1102
rect 5229 1068 5236 1102
rect 5275 1068 5297 1102
rect 5297 1068 5309 1102
rect 5348 1068 5365 1102
rect 5365 1068 5382 1102
rect 5421 1068 5433 1102
rect 5433 1068 5455 1102
rect 5495 1068 5501 1102
rect 5501 1068 5529 1102
rect 5569 1068 5603 1102
rect 5643 1068 5671 1102
rect 5671 1068 5677 1102
rect 5717 1068 5739 1102
rect 5739 1068 5751 1102
rect 5791 1068 5807 1102
rect 5807 1068 5825 1102
rect 5865 1068 5875 1102
rect 5875 1068 5899 1102
rect 5939 1068 5943 1102
rect 5943 1068 5973 1102
rect 6013 1068 6045 1102
rect 6045 1068 6047 1102
rect 6087 1068 6113 1102
rect 6113 1068 6121 1102
rect 6161 1068 6181 1102
rect 6181 1068 6195 1102
rect 6235 1068 6249 1102
rect 6249 1068 6269 1102
rect 6309 1068 6317 1102
rect 6317 1068 6343 1102
rect 6383 1068 6385 1102
rect 6385 1068 6417 1102
rect 6457 1068 6487 1102
rect 6487 1068 6491 1102
rect 6547 1090 6581 1118
rect 6547 1084 6581 1090
rect 2311 1017 2345 1038
rect 2311 1004 2345 1017
rect 2311 944 2345 956
rect 6547 1017 6581 1035
rect 6547 1001 6581 1017
rect 2311 922 2345 944
rect 2401 912 2405 946
rect 2405 912 2435 946
rect 2475 912 2507 946
rect 2507 912 2509 946
rect 2549 912 2575 946
rect 2575 912 2583 946
rect 2623 912 2643 946
rect 2643 912 2657 946
rect 2697 912 2711 946
rect 2711 912 2731 946
rect 2771 912 2779 946
rect 2779 912 2805 946
rect 2845 912 2847 946
rect 2847 912 2879 946
rect 2919 912 2949 946
rect 2949 912 2953 946
rect 2993 912 3017 946
rect 3017 912 3027 946
rect 3067 912 3085 946
rect 3085 912 3101 946
rect 3141 912 3153 946
rect 3153 912 3175 946
rect 3215 912 3221 946
rect 3221 912 3249 946
rect 3289 912 3323 946
rect 3363 912 3391 946
rect 3391 912 3397 946
rect 3437 912 3459 946
rect 3459 912 3471 946
rect 3510 912 3527 946
rect 3527 912 3544 946
rect 3583 912 3595 946
rect 3595 912 3617 946
rect 3656 912 3663 946
rect 3663 912 3690 946
rect 3729 912 3731 946
rect 3731 912 3763 946
rect 3802 912 3833 946
rect 3833 912 3836 946
rect 3875 912 3901 946
rect 3901 912 3909 946
rect 3948 912 3969 946
rect 3969 912 3982 946
rect 4021 912 4037 946
rect 4037 912 4055 946
rect 4094 912 4105 946
rect 4105 912 4128 946
rect 4167 912 4173 946
rect 4173 912 4201 946
rect 4240 912 4241 946
rect 4241 912 4274 946
rect 4313 912 4343 946
rect 4343 912 4347 946
rect 4545 912 4549 946
rect 4549 912 4579 946
rect 4618 912 4651 946
rect 4651 912 4652 946
rect 4691 912 4719 946
rect 4719 912 4725 946
rect 4764 912 4787 946
rect 4787 912 4798 946
rect 4837 912 4855 946
rect 4855 912 4871 946
rect 4910 912 4923 946
rect 4923 912 4944 946
rect 4983 912 4991 946
rect 4991 912 5017 946
rect 5056 912 5059 946
rect 5059 912 5090 946
rect 5129 912 5161 946
rect 5161 912 5163 946
rect 5202 912 5229 946
rect 5229 912 5236 946
rect 5275 912 5297 946
rect 5297 912 5309 946
rect 5348 912 5365 946
rect 5365 912 5382 946
rect 5421 912 5433 946
rect 5433 912 5455 946
rect 5495 912 5501 946
rect 5501 912 5529 946
rect 5569 912 5603 946
rect 5643 912 5671 946
rect 5671 912 5677 946
rect 5717 912 5739 946
rect 5739 912 5751 946
rect 5791 912 5807 946
rect 5807 912 5825 946
rect 5865 912 5875 946
rect 5875 912 5899 946
rect 5939 912 5943 946
rect 5943 912 5973 946
rect 6013 912 6045 946
rect 6045 912 6047 946
rect 6087 912 6113 946
rect 6113 912 6121 946
rect 6161 912 6181 946
rect 6181 912 6195 946
rect 6235 912 6249 946
rect 6249 912 6269 946
rect 6309 912 6317 946
rect 6317 912 6343 946
rect 6383 912 6385 946
rect 6385 912 6417 946
rect 6457 912 6487 946
rect 6487 912 6491 946
rect 6547 944 6581 952
rect 6547 918 6581 944
rect 2311 871 2345 874
rect 2311 840 2345 871
rect 2311 759 2345 792
rect 6547 834 6581 868
rect 2311 758 2345 759
rect 2401 756 2405 790
rect 2405 756 2435 790
rect 2475 756 2507 790
rect 2507 756 2509 790
rect 2549 756 2575 790
rect 2575 756 2583 790
rect 2623 756 2643 790
rect 2643 756 2657 790
rect 2697 756 2711 790
rect 2711 756 2731 790
rect 2771 756 2779 790
rect 2779 756 2805 790
rect 2845 756 2847 790
rect 2847 756 2879 790
rect 2919 756 2949 790
rect 2949 756 2953 790
rect 2993 756 3017 790
rect 3017 756 3027 790
rect 3067 756 3085 790
rect 3085 756 3101 790
rect 3141 756 3153 790
rect 3153 756 3175 790
rect 3215 756 3221 790
rect 3221 756 3249 790
rect 3289 756 3323 790
rect 3363 756 3391 790
rect 3391 756 3397 790
rect 3437 756 3459 790
rect 3459 756 3471 790
rect 3510 756 3527 790
rect 3527 756 3544 790
rect 3583 756 3595 790
rect 3595 756 3617 790
rect 3656 756 3663 790
rect 3663 756 3690 790
rect 3729 756 3731 790
rect 3731 756 3763 790
rect 3802 756 3833 790
rect 3833 756 3836 790
rect 3875 756 3901 790
rect 3901 756 3909 790
rect 3948 756 3969 790
rect 3969 756 3982 790
rect 4021 756 4037 790
rect 4037 756 4055 790
rect 4094 756 4105 790
rect 4105 756 4128 790
rect 4167 756 4173 790
rect 4173 756 4201 790
rect 4240 756 4241 790
rect 4241 756 4274 790
rect 4313 756 4343 790
rect 4343 756 4347 790
rect 4545 756 4549 790
rect 4549 756 4579 790
rect 4618 756 4651 790
rect 4651 756 4652 790
rect 4691 756 4719 790
rect 4719 756 4725 790
rect 4764 756 4787 790
rect 4787 756 4798 790
rect 4837 756 4855 790
rect 4855 756 4871 790
rect 4910 756 4923 790
rect 4923 756 4944 790
rect 4983 756 4991 790
rect 4991 756 5017 790
rect 5056 756 5059 790
rect 5059 756 5090 790
rect 5129 756 5161 790
rect 5161 756 5163 790
rect 5202 756 5229 790
rect 5229 756 5236 790
rect 5275 756 5297 790
rect 5297 756 5309 790
rect 5348 756 5365 790
rect 5365 756 5382 790
rect 5421 756 5433 790
rect 5433 756 5455 790
rect 5495 756 5501 790
rect 5501 756 5529 790
rect 5569 756 5603 790
rect 5643 756 5671 790
rect 5671 756 5677 790
rect 5717 756 5739 790
rect 5739 756 5751 790
rect 5791 756 5807 790
rect 5807 756 5825 790
rect 5865 756 5875 790
rect 5875 756 5899 790
rect 5939 756 5943 790
rect 5943 756 5973 790
rect 6013 756 6045 790
rect 6045 756 6047 790
rect 6087 756 6113 790
rect 6113 756 6121 790
rect 6161 756 6181 790
rect 6181 756 6195 790
rect 6235 756 6249 790
rect 6249 756 6269 790
rect 6309 756 6317 790
rect 6317 756 6343 790
rect 6383 756 6385 790
rect 6385 756 6417 790
rect 6457 756 6487 790
rect 6487 756 6491 790
rect 6547 759 6581 784
rect 2311 686 2345 710
rect 2311 676 2345 686
rect 6547 750 6581 759
rect 6547 686 6581 700
rect 6547 666 6581 686
rect 2401 600 2405 634
rect 2405 600 2435 634
rect 2475 600 2507 634
rect 2507 600 2509 634
rect 2549 600 2575 634
rect 2575 600 2583 634
rect 2623 600 2643 634
rect 2643 600 2657 634
rect 2697 600 2711 634
rect 2711 600 2731 634
rect 2771 600 2779 634
rect 2779 600 2805 634
rect 2845 600 2847 634
rect 2847 600 2879 634
rect 2919 600 2949 634
rect 2949 600 2953 634
rect 2993 600 3017 634
rect 3017 600 3027 634
rect 3067 600 3085 634
rect 3085 600 3101 634
rect 3141 600 3153 634
rect 3153 600 3175 634
rect 3215 600 3221 634
rect 3221 600 3249 634
rect 3289 600 3323 634
rect 3363 600 3391 634
rect 3391 600 3397 634
rect 3437 600 3459 634
rect 3459 600 3471 634
rect 3510 600 3527 634
rect 3527 600 3544 634
rect 3583 600 3595 634
rect 3595 600 3617 634
rect 3656 600 3663 634
rect 3663 600 3690 634
rect 3729 600 3731 634
rect 3731 600 3763 634
rect 3802 600 3833 634
rect 3833 600 3836 634
rect 3875 600 3901 634
rect 3901 600 3909 634
rect 3948 600 3969 634
rect 3969 600 3982 634
rect 4021 600 4037 634
rect 4037 600 4055 634
rect 4094 600 4105 634
rect 4105 600 4128 634
rect 4167 600 4173 634
rect 4173 600 4201 634
rect 4240 600 4241 634
rect 4241 600 4274 634
rect 4313 600 4343 634
rect 4343 600 4347 634
rect 4545 600 4549 634
rect 4549 600 4579 634
rect 4618 600 4651 634
rect 4651 600 4652 634
rect 4691 600 4719 634
rect 4719 600 4725 634
rect 4764 600 4787 634
rect 4787 600 4798 634
rect 4837 600 4855 634
rect 4855 600 4871 634
rect 4910 600 4923 634
rect 4923 600 4944 634
rect 4983 600 4991 634
rect 4991 600 5017 634
rect 5056 600 5059 634
rect 5059 600 5090 634
rect 5129 600 5161 634
rect 5161 600 5163 634
rect 5202 600 5229 634
rect 5229 600 5236 634
rect 5275 600 5297 634
rect 5297 600 5309 634
rect 5348 600 5365 634
rect 5365 600 5382 634
rect 5421 600 5433 634
rect 5433 600 5455 634
rect 5495 600 5501 634
rect 5501 600 5529 634
rect 5569 600 5603 634
rect 5643 600 5671 634
rect 5671 600 5677 634
rect 5717 600 5739 634
rect 5739 600 5751 634
rect 5791 600 5807 634
rect 5807 600 5825 634
rect 5865 600 5875 634
rect 5875 600 5899 634
rect 5939 600 5943 634
rect 5943 600 5973 634
rect 6013 600 6045 634
rect 6045 600 6047 634
rect 6087 600 6113 634
rect 6113 600 6121 634
rect 6161 600 6181 634
rect 6181 600 6195 634
rect 6235 600 6249 634
rect 6249 600 6269 634
rect 6309 600 6317 634
rect 6317 600 6343 634
rect 6383 600 6385 634
rect 6385 600 6417 634
rect 6457 600 6487 634
rect 6487 600 6491 634
rect 6627 1308 6733 1343
rect 6627 1274 6683 1308
rect 6683 1274 6717 1308
rect 6717 1274 6733 1308
rect 6627 1240 6733 1274
rect 6627 1206 6683 1240
rect 6683 1206 6717 1240
rect 6717 1206 6733 1240
rect 6627 1200 6733 1206
rect 6627 1127 6661 1161
rect 6699 1138 6717 1161
rect 6717 1138 6733 1161
rect 6699 1127 6733 1138
rect 6627 1054 6661 1088
rect 6699 1070 6717 1088
rect 6717 1070 6733 1088
rect 6699 1054 6733 1070
rect 6627 981 6661 1015
rect 6699 1002 6717 1015
rect 6717 1002 6733 1015
rect 6699 981 6733 1002
rect 6627 908 6661 942
rect 6699 934 6717 942
rect 6717 934 6733 942
rect 6699 908 6733 934
rect 6627 835 6661 869
rect 6699 866 6717 869
rect 6717 866 6733 869
rect 6699 835 6733 866
rect 6627 762 6661 796
rect 6699 764 6733 796
rect 6699 762 6717 764
rect 6717 762 6733 764
rect 6627 689 6661 723
rect 6699 696 6733 723
rect 6699 689 6717 696
rect 6717 689 6733 696
rect 6627 616 6661 650
rect 6699 628 6733 650
rect 6699 616 6717 628
rect 6717 616 6733 628
rect 6627 543 6661 577
rect 6699 560 6733 577
rect 6699 543 6717 560
rect 6717 543 6733 560
rect 2401 444 2405 478
rect 2405 444 2435 478
rect 2475 444 2507 478
rect 2507 444 2509 478
rect 2549 444 2575 478
rect 2575 444 2583 478
rect 2623 444 2643 478
rect 2643 444 2657 478
rect 2697 444 2711 478
rect 2711 444 2731 478
rect 2771 444 2779 478
rect 2779 444 2805 478
rect 2845 444 2847 478
rect 2847 444 2879 478
rect 2919 444 2949 478
rect 2949 444 2953 478
rect 2993 444 3017 478
rect 3017 444 3027 478
rect 3067 444 3085 478
rect 3085 444 3101 478
rect 3141 444 3153 478
rect 3153 444 3175 478
rect 3215 444 3221 478
rect 3221 444 3249 478
rect 3289 444 3323 478
rect 3363 444 3391 478
rect 3391 444 3397 478
rect 3437 444 3459 478
rect 3459 444 3471 478
rect 3510 444 3527 478
rect 3527 444 3544 478
rect 3583 444 3595 478
rect 3595 444 3617 478
rect 3656 444 3663 478
rect 3663 444 3690 478
rect 3729 444 3731 478
rect 3731 444 3763 478
rect 3802 444 3833 478
rect 3833 444 3836 478
rect 3875 444 3901 478
rect 3901 444 3909 478
rect 3948 444 3969 478
rect 3969 444 3982 478
rect 4021 444 4037 478
rect 4037 444 4055 478
rect 4094 444 4105 478
rect 4105 444 4128 478
rect 4167 444 4173 478
rect 4173 444 4201 478
rect 4240 444 4241 478
rect 4241 444 4274 478
rect 4313 444 4343 478
rect 4343 444 4347 478
rect 4545 444 4549 478
rect 4549 444 4579 478
rect 4618 444 4651 478
rect 4651 444 4652 478
rect 4691 444 4719 478
rect 4719 444 4725 478
rect 4764 444 4787 478
rect 4787 444 4798 478
rect 4837 444 4855 478
rect 4855 444 4871 478
rect 4910 444 4923 478
rect 4923 444 4944 478
rect 4983 444 4991 478
rect 4991 444 5017 478
rect 5056 444 5059 478
rect 5059 444 5090 478
rect 5129 444 5161 478
rect 5161 444 5163 478
rect 5202 444 5229 478
rect 5229 444 5236 478
rect 5275 444 5297 478
rect 5297 444 5309 478
rect 5348 444 5365 478
rect 5365 444 5382 478
rect 5421 444 5433 478
rect 5433 444 5455 478
rect 5495 444 5501 478
rect 5501 444 5529 478
rect 5569 444 5603 478
rect 5643 444 5671 478
rect 5671 444 5677 478
rect 5717 444 5739 478
rect 5739 444 5751 478
rect 5791 444 5807 478
rect 5807 444 5825 478
rect 5865 444 5875 478
rect 5875 444 5899 478
rect 5939 444 5943 478
rect 5943 444 5973 478
rect 6013 444 6045 478
rect 6045 444 6047 478
rect 6087 444 6113 478
rect 6113 444 6121 478
rect 6161 444 6181 478
rect 6181 444 6195 478
rect 6235 444 6249 478
rect 6249 444 6269 478
rect 6309 444 6317 478
rect 6317 444 6343 478
rect 6383 444 6385 478
rect 6385 444 6417 478
rect 6457 444 6487 478
rect 6487 444 6491 478
rect 6627 470 6661 504
rect 6699 492 6733 504
rect 6699 470 6717 492
rect 6717 470 6733 492
rect 6627 397 6661 431
rect 6699 424 6733 431
rect 6699 397 6717 424
rect 6717 397 6733 424
rect 2159 325 2260 359
rect 2260 325 2265 359
rect 2304 325 2328 358
rect 2328 325 2338 358
rect 2377 325 2396 358
rect 2396 325 2411 358
rect 2450 325 2464 358
rect 2464 325 2484 358
rect 2523 325 2532 358
rect 2532 325 2566 358
rect 2566 325 2600 358
rect 2600 325 2634 358
rect 2634 325 2668 358
rect 2668 325 2702 358
rect 2702 325 2736 358
rect 2736 325 2770 358
rect 2770 325 2804 358
rect 2804 325 2838 358
rect 2838 325 2872 358
rect 2872 325 2906 358
rect 2906 325 2940 358
rect 2940 325 2974 358
rect 2974 325 3008 358
rect 3008 325 3042 358
rect 3042 325 3076 358
rect 3076 325 3110 358
rect 3110 325 3144 358
rect 3144 325 3178 358
rect 3178 325 3212 358
rect 3212 325 3246 358
rect 3246 325 3280 358
rect 3280 325 3314 358
rect 3314 325 3348 358
rect 3348 325 3382 358
rect 3382 325 3416 358
rect 3416 325 3450 358
rect 3450 325 3484 358
rect 3484 325 3518 358
rect 3518 325 3552 358
rect 3552 325 3586 358
rect 3586 325 3620 358
rect 3620 325 3654 358
rect 3654 325 3688 358
rect 3688 325 3722 358
rect 3722 325 3756 358
rect 3756 325 3790 358
rect 3790 325 3824 358
rect 3824 325 3858 358
rect 3858 325 3892 358
rect 3892 325 3926 358
rect 3926 325 3960 358
rect 3960 325 3994 358
rect 3994 325 4028 358
rect 4028 325 4062 358
rect 4062 325 4096 358
rect 4096 325 4130 358
rect 4130 325 4164 358
rect 4164 325 4198 358
rect 4198 325 4232 358
rect 4232 325 4266 358
rect 4266 325 4300 358
rect 4300 325 4334 358
rect 4334 325 4368 358
rect 4368 325 4402 358
rect 4402 325 4436 358
rect 4436 325 4470 358
rect 4470 325 4504 358
rect 4504 325 4538 358
rect 4538 325 4572 358
rect 4572 325 4606 358
rect 4606 325 4640 358
rect 4640 325 4674 358
rect 4674 325 4708 358
rect 4708 325 4742 358
rect 4742 325 4776 358
rect 4776 325 4810 358
rect 4810 325 4844 358
rect 4844 325 4878 358
rect 4878 325 4912 358
rect 4912 325 4946 358
rect 4946 325 4980 358
rect 4980 325 5014 358
rect 5014 325 5048 358
rect 5048 325 5082 358
rect 5082 325 5116 358
rect 5116 325 5150 358
rect 5150 325 5184 358
rect 5184 325 5218 358
rect 5218 325 5252 358
rect 5252 325 5286 358
rect 5286 325 5320 358
rect 5320 325 5354 358
rect 5354 325 5388 358
rect 5388 325 5422 358
rect 5422 325 5456 358
rect 5456 325 5490 358
rect 5490 325 5524 358
rect 5524 325 5558 358
rect 5558 325 5592 358
rect 5592 325 5626 358
rect 5626 325 5660 358
rect 5660 325 5694 358
rect 5694 325 5728 358
rect 5728 325 5762 358
rect 5762 325 5796 358
rect 5796 325 5830 358
rect 5830 325 5864 358
rect 5864 325 5898 358
rect 5898 325 5932 358
rect 5932 325 5966 358
rect 5966 325 6000 358
rect 6000 325 6034 358
rect 6034 325 6068 358
rect 6068 325 6102 358
rect 6102 325 6136 358
rect 6136 325 6170 358
rect 6170 325 6204 358
rect 6204 325 6238 358
rect 6238 325 6272 358
rect 6272 325 6306 358
rect 6306 325 6340 358
rect 6340 325 6374 358
rect 6374 325 6408 358
rect 6408 325 6442 358
rect 6442 325 6476 358
rect 6476 325 6510 358
rect 6510 325 6544 358
rect 6544 325 6578 358
rect 6578 325 6612 358
rect 6612 325 6646 358
rect 6646 325 6661 358
rect 2159 324 2265 325
rect 2304 324 2338 325
rect 2377 324 2411 325
rect 2450 324 2484 325
rect 2231 252 2265 286
rect 2304 252 2338 286
rect 2377 252 2411 286
rect 2450 252 2484 286
rect 2523 252 6661 325
rect 6699 324 6733 358
rect 6882 1390 6884 1424
rect 6884 1390 6916 1424
rect 6954 1390 6986 1424
rect 6986 1390 6988 1424
rect 6882 1317 6884 1351
rect 6884 1317 6916 1351
rect 6954 1317 6986 1351
rect 6986 1317 6988 1351
rect 6882 1244 6884 1278
rect 6884 1244 6916 1278
rect 6954 1244 6986 1278
rect 6986 1244 6988 1278
rect 6882 1171 6884 1205
rect 6884 1171 6916 1205
rect 6954 1171 6986 1205
rect 6986 1171 6988 1205
rect 6882 1097 6884 1131
rect 6884 1097 6916 1131
rect 6954 1097 6986 1131
rect 6986 1097 6988 1131
rect 6882 1023 6884 1057
rect 6884 1023 6916 1057
rect 6954 1023 6986 1057
rect 6986 1023 6988 1057
rect 6882 949 6884 983
rect 6884 949 6916 983
rect 6954 949 6986 983
rect 6986 949 6988 983
rect 6882 875 6884 909
rect 6884 875 6916 909
rect 6954 875 6986 909
rect 6986 875 6988 909
rect 6882 801 6884 835
rect 6884 801 6916 835
rect 6954 801 6986 835
rect 6986 801 6988 835
rect 6882 727 6884 761
rect 6884 727 6916 761
rect 6954 727 6986 761
rect 6986 727 6988 761
rect 6882 653 6884 687
rect 6884 653 6916 687
rect 6954 653 6986 687
rect 6986 653 6988 687
rect 6882 579 6884 613
rect 6884 579 6916 613
rect 6954 579 6986 613
rect 6986 579 6988 613
rect 6882 505 6884 539
rect 6884 505 6916 539
rect 6954 505 6986 539
rect 6986 505 6988 539
rect 6882 431 6884 465
rect 6884 431 6916 465
rect 6954 431 6986 465
rect 6986 431 6988 465
rect 6882 357 6884 391
rect 6884 357 6916 391
rect 6954 357 6986 391
rect 6986 357 6988 391
rect 6882 312 6884 317
rect 6884 312 6916 317
rect 6954 312 6986 317
rect 6986 312 6988 317
rect 6882 283 6916 312
rect 6954 283 6988 312
rect 1904 209 1906 243
rect 1906 209 1938 243
rect 1976 209 2008 243
rect 2008 209 2010 243
rect 7241 1406 7275 1440
rect 7319 1406 7353 1440
rect 7397 1406 7431 1440
rect 7475 1406 7509 1440
rect 7553 1406 7587 1440
rect 7631 1406 7665 1440
rect 7709 1406 7743 1440
rect 7788 1406 7822 1440
rect 7898 1377 11460 1440
rect 11499 1406 11533 1440
rect 11572 1406 11606 1440
rect 11645 1406 11679 1440
rect 7163 1334 7197 1368
rect 7235 1343 7264 1368
rect 7264 1343 7269 1368
rect 7319 1343 7332 1368
rect 7332 1343 7353 1368
rect 7397 1343 7400 1368
rect 7400 1343 7431 1368
rect 7475 1343 7502 1368
rect 7502 1343 7509 1368
rect 7553 1343 7570 1368
rect 7570 1343 7587 1368
rect 7631 1343 7638 1368
rect 7638 1343 7665 1368
rect 7709 1343 7740 1368
rect 7740 1343 7743 1368
rect 7788 1343 7808 1368
rect 7808 1343 7822 1368
rect 7898 1343 7910 1377
rect 7910 1343 7944 1377
rect 7944 1343 7978 1377
rect 7978 1343 8012 1377
rect 8012 1343 8046 1377
rect 8046 1343 8080 1377
rect 8080 1343 8114 1377
rect 8114 1343 8148 1377
rect 8148 1343 8182 1377
rect 8182 1343 8216 1377
rect 8216 1343 8250 1377
rect 8250 1343 8284 1377
rect 8284 1343 8318 1377
rect 8318 1343 8352 1377
rect 8352 1343 8386 1377
rect 8386 1343 8420 1377
rect 8420 1343 8454 1377
rect 8454 1343 8488 1377
rect 8488 1343 8522 1377
rect 8522 1343 8556 1377
rect 8556 1343 8590 1377
rect 8590 1343 8624 1377
rect 8624 1343 8658 1377
rect 8658 1343 8692 1377
rect 8692 1343 8726 1377
rect 8726 1343 8760 1377
rect 8760 1343 8794 1377
rect 8794 1343 8828 1377
rect 8828 1343 8862 1377
rect 8862 1343 8896 1377
rect 8896 1343 8930 1377
rect 8930 1343 8964 1377
rect 8964 1343 8998 1377
rect 8998 1343 9032 1377
rect 9032 1343 9066 1377
rect 9066 1343 9100 1377
rect 9100 1343 9134 1377
rect 9134 1343 9168 1377
rect 9168 1343 9202 1377
rect 9202 1343 9236 1377
rect 9236 1343 9270 1377
rect 9270 1343 9304 1377
rect 9304 1343 9338 1377
rect 9338 1343 9372 1377
rect 9372 1343 9406 1377
rect 9406 1343 9500 1377
rect 9500 1343 9534 1377
rect 9534 1343 9568 1377
rect 9568 1343 9602 1377
rect 9602 1343 9636 1377
rect 9636 1343 9670 1377
rect 9670 1343 9704 1377
rect 9704 1343 9738 1377
rect 9738 1343 9772 1377
rect 9772 1343 9806 1377
rect 9806 1343 9840 1377
rect 9840 1343 9874 1377
rect 9874 1343 9908 1377
rect 9908 1343 9942 1377
rect 9942 1343 9976 1377
rect 9976 1343 10010 1377
rect 10010 1343 10044 1377
rect 10044 1343 10078 1377
rect 10078 1343 10112 1377
rect 10112 1343 10146 1377
rect 10146 1343 10180 1377
rect 10180 1343 10214 1377
rect 10214 1343 10248 1377
rect 10248 1343 10282 1377
rect 10282 1343 10316 1377
rect 10316 1343 10350 1377
rect 10350 1343 10384 1377
rect 10384 1343 10418 1377
rect 10418 1343 10452 1377
rect 10452 1343 10486 1377
rect 10486 1343 10520 1377
rect 10520 1343 10554 1377
rect 10554 1343 10588 1377
rect 10588 1343 10622 1377
rect 10622 1343 10656 1377
rect 10656 1343 10690 1377
rect 10690 1343 10724 1377
rect 10724 1343 10758 1377
rect 10758 1343 10792 1377
rect 10792 1343 10826 1377
rect 10826 1343 10860 1377
rect 10860 1343 10894 1377
rect 10894 1343 10928 1377
rect 10928 1343 10962 1377
rect 10962 1343 10996 1377
rect 10996 1343 11030 1377
rect 11030 1343 11064 1377
rect 11064 1343 11098 1377
rect 11098 1343 11132 1377
rect 11132 1343 11166 1377
rect 11166 1343 11200 1377
rect 11200 1343 11234 1377
rect 11234 1343 11268 1377
rect 11268 1343 11302 1377
rect 11302 1343 11336 1377
rect 11336 1343 11370 1377
rect 11370 1343 11404 1377
rect 11404 1343 11438 1377
rect 11438 1343 11460 1377
rect 11499 1343 11506 1368
rect 11506 1343 11533 1368
rect 11572 1343 11574 1368
rect 11574 1343 11606 1368
rect 7235 1334 7269 1343
rect 7319 1334 7353 1343
rect 7397 1334 7431 1343
rect 7475 1334 7509 1343
rect 7553 1334 7587 1343
rect 7631 1334 7665 1343
rect 7709 1334 7743 1343
rect 7788 1334 7822 1343
rect 7898 1334 11460 1343
rect 11499 1334 11533 1343
rect 11572 1334 11606 1343
rect 7163 1261 7197 1295
rect 7235 1261 7269 1295
rect 7420 1224 7454 1258
rect 7494 1224 7496 1258
rect 7496 1224 7528 1258
rect 7568 1224 7598 1258
rect 7598 1224 7602 1258
rect 7642 1224 7666 1258
rect 7666 1224 7676 1258
rect 7716 1224 7734 1258
rect 7734 1224 7750 1258
rect 7790 1224 7802 1258
rect 7802 1224 7824 1258
rect 7864 1224 7870 1258
rect 7870 1224 7898 1258
rect 7938 1224 7972 1258
rect 8012 1224 8040 1258
rect 8040 1224 8046 1258
rect 8086 1224 8108 1258
rect 8108 1224 8120 1258
rect 8160 1224 8176 1258
rect 8176 1224 8194 1258
rect 8234 1224 8244 1258
rect 8244 1224 8268 1258
rect 8308 1224 8312 1258
rect 8312 1224 8342 1258
rect 8382 1224 8414 1258
rect 8414 1224 8416 1258
rect 8456 1224 8482 1258
rect 8482 1224 8490 1258
rect 8529 1224 8550 1258
rect 8550 1224 8563 1258
rect 8602 1224 8618 1258
rect 8618 1224 8636 1258
rect 8675 1224 8686 1258
rect 8686 1224 8709 1258
rect 8748 1224 8754 1258
rect 8754 1224 8782 1258
rect 8821 1224 8822 1258
rect 8822 1224 8855 1258
rect 8894 1224 8924 1258
rect 8924 1224 8928 1258
rect 8967 1224 8992 1258
rect 8992 1224 9001 1258
rect 9040 1224 9060 1258
rect 9060 1224 9074 1258
rect 9113 1224 9128 1258
rect 9128 1224 9147 1258
rect 9186 1224 9196 1258
rect 9196 1224 9220 1258
rect 9259 1224 9264 1258
rect 9264 1224 9293 1258
rect 9332 1224 9366 1258
rect 9564 1224 9568 1258
rect 9568 1224 9598 1258
rect 9637 1224 9670 1258
rect 9670 1224 9671 1258
rect 9710 1224 9738 1258
rect 9738 1224 9744 1258
rect 9783 1224 9806 1258
rect 9806 1224 9817 1258
rect 9856 1224 9874 1258
rect 9874 1224 9890 1258
rect 9929 1224 9942 1258
rect 9942 1224 9963 1258
rect 10002 1224 10010 1258
rect 10010 1224 10036 1258
rect 10075 1224 10078 1258
rect 10078 1224 10109 1258
rect 10148 1224 10180 1258
rect 10180 1224 10182 1258
rect 10221 1224 10248 1258
rect 10248 1224 10255 1258
rect 10294 1224 10316 1258
rect 10316 1224 10328 1258
rect 10367 1224 10384 1258
rect 10384 1224 10401 1258
rect 10440 1224 10452 1258
rect 10452 1224 10474 1258
rect 10514 1224 10520 1258
rect 10520 1224 10548 1258
rect 10588 1224 10622 1258
rect 10662 1224 10690 1258
rect 10690 1224 10696 1258
rect 10736 1224 10758 1258
rect 10758 1224 10770 1258
rect 10810 1224 10826 1258
rect 10826 1224 10844 1258
rect 10884 1224 10894 1258
rect 10894 1224 10918 1258
rect 10958 1224 10962 1258
rect 10962 1224 10992 1258
rect 11032 1224 11064 1258
rect 11064 1224 11066 1258
rect 11106 1224 11132 1258
rect 11132 1224 11140 1258
rect 11180 1224 11200 1258
rect 11200 1224 11214 1258
rect 11254 1224 11268 1258
rect 11268 1224 11288 1258
rect 11328 1224 11336 1258
rect 11336 1224 11362 1258
rect 11402 1224 11404 1258
rect 11404 1224 11436 1258
rect 11476 1224 11506 1258
rect 11506 1224 11510 1258
rect 7163 1206 7199 1222
rect 7199 1206 7233 1222
rect 7233 1206 7269 1222
rect 7163 1172 7269 1206
rect 7163 1138 7199 1172
rect 7199 1138 7233 1172
rect 7233 1138 7269 1172
rect 7163 1104 7269 1138
rect 7163 1070 7199 1104
rect 7199 1070 7233 1104
rect 7233 1070 7269 1104
rect 7163 1036 7269 1070
rect 7163 1002 7199 1036
rect 7199 1002 7233 1036
rect 7233 1002 7269 1036
rect 7163 968 7269 1002
rect 7163 934 7199 968
rect 7199 934 7233 968
rect 7233 934 7269 968
rect 7163 900 7269 934
rect 7163 866 7199 900
rect 7199 866 7233 900
rect 7233 866 7269 900
rect 7163 832 7269 866
rect 7163 798 7199 832
rect 7199 798 7233 832
rect 7233 798 7269 832
rect 7163 764 7269 798
rect 7163 730 7199 764
rect 7199 730 7233 764
rect 7233 730 7269 764
rect 7163 696 7269 730
rect 7163 662 7199 696
rect 7199 662 7233 696
rect 7233 662 7269 696
rect 7163 628 7269 662
rect 7163 594 7199 628
rect 7199 594 7233 628
rect 7233 594 7269 628
rect 7163 560 7269 594
rect 7163 526 7199 560
rect 7199 526 7233 560
rect 7233 526 7269 560
rect 7163 492 7269 526
rect 7163 458 7199 492
rect 7199 458 7233 492
rect 7233 458 7269 492
rect 7163 424 7269 458
rect 7163 390 7199 424
rect 7199 390 7233 424
rect 7233 390 7269 424
rect 7163 359 7269 390
rect 7330 1197 7364 1201
rect 7330 1167 7364 1197
rect 7330 1123 7364 1127
rect 7330 1093 7364 1123
rect 11566 1197 11600 1201
rect 11566 1167 11599 1197
rect 11599 1167 11600 1197
rect 11566 1123 11600 1127
rect 7420 1068 7454 1102
rect 7494 1068 7496 1102
rect 7496 1068 7528 1102
rect 7568 1068 7598 1102
rect 7598 1068 7602 1102
rect 7642 1068 7666 1102
rect 7666 1068 7676 1102
rect 7716 1068 7734 1102
rect 7734 1068 7750 1102
rect 7790 1068 7802 1102
rect 7802 1068 7824 1102
rect 7864 1068 7870 1102
rect 7870 1068 7898 1102
rect 7938 1068 7972 1102
rect 8012 1068 8040 1102
rect 8040 1068 8046 1102
rect 8086 1068 8108 1102
rect 8108 1068 8120 1102
rect 8160 1068 8176 1102
rect 8176 1068 8194 1102
rect 8234 1068 8244 1102
rect 8244 1068 8268 1102
rect 8308 1068 8312 1102
rect 8312 1068 8342 1102
rect 8382 1068 8414 1102
rect 8414 1068 8416 1102
rect 8456 1068 8482 1102
rect 8482 1068 8490 1102
rect 8529 1068 8550 1102
rect 8550 1068 8563 1102
rect 8602 1068 8618 1102
rect 8618 1068 8636 1102
rect 8675 1068 8686 1102
rect 8686 1068 8709 1102
rect 8748 1068 8754 1102
rect 8754 1068 8782 1102
rect 8821 1068 8822 1102
rect 8822 1068 8855 1102
rect 8894 1068 8924 1102
rect 8924 1068 8928 1102
rect 8967 1068 8992 1102
rect 8992 1068 9001 1102
rect 9040 1068 9060 1102
rect 9060 1068 9074 1102
rect 9113 1068 9128 1102
rect 9128 1068 9147 1102
rect 9186 1068 9196 1102
rect 9196 1068 9220 1102
rect 9259 1068 9264 1102
rect 9264 1068 9293 1102
rect 9332 1068 9366 1102
rect 9564 1068 9568 1102
rect 9568 1068 9598 1102
rect 9637 1068 9670 1102
rect 9670 1068 9671 1102
rect 9710 1068 9738 1102
rect 9738 1068 9744 1102
rect 9783 1068 9806 1102
rect 9806 1068 9817 1102
rect 9856 1068 9874 1102
rect 9874 1068 9890 1102
rect 9929 1068 9942 1102
rect 9942 1068 9963 1102
rect 10002 1068 10010 1102
rect 10010 1068 10036 1102
rect 10075 1068 10078 1102
rect 10078 1068 10109 1102
rect 10148 1068 10180 1102
rect 10180 1068 10182 1102
rect 10221 1068 10248 1102
rect 10248 1068 10255 1102
rect 10294 1068 10316 1102
rect 10316 1068 10328 1102
rect 10367 1068 10384 1102
rect 10384 1068 10401 1102
rect 10440 1068 10452 1102
rect 10452 1068 10474 1102
rect 10514 1068 10520 1102
rect 10520 1068 10548 1102
rect 10588 1068 10622 1102
rect 10662 1068 10690 1102
rect 10690 1068 10696 1102
rect 10736 1068 10758 1102
rect 10758 1068 10770 1102
rect 10810 1068 10826 1102
rect 10826 1068 10844 1102
rect 10884 1068 10894 1102
rect 10894 1068 10918 1102
rect 10958 1068 10962 1102
rect 10962 1068 10992 1102
rect 11032 1068 11064 1102
rect 11064 1068 11066 1102
rect 11106 1068 11132 1102
rect 11132 1068 11140 1102
rect 11180 1068 11200 1102
rect 11200 1068 11214 1102
rect 11254 1068 11268 1102
rect 11268 1068 11288 1102
rect 11328 1068 11336 1102
rect 11336 1068 11362 1102
rect 11402 1068 11404 1102
rect 11404 1068 11436 1102
rect 11476 1068 11506 1102
rect 11506 1068 11510 1102
rect 11566 1093 11599 1123
rect 11599 1093 11600 1123
rect 7330 1050 7364 1053
rect 7330 1019 7364 1050
rect 7330 977 7364 979
rect 7330 945 7364 977
rect 11566 1050 11600 1053
rect 11566 1019 11599 1050
rect 11599 1019 11600 1050
rect 11566 977 11600 979
rect 7420 912 7454 946
rect 7494 912 7496 946
rect 7496 912 7528 946
rect 7568 912 7598 946
rect 7598 912 7602 946
rect 7642 912 7666 946
rect 7666 912 7676 946
rect 7716 912 7734 946
rect 7734 912 7750 946
rect 7790 912 7802 946
rect 7802 912 7824 946
rect 7864 912 7870 946
rect 7870 912 7898 946
rect 7938 912 7972 946
rect 8012 912 8040 946
rect 8040 912 8046 946
rect 8086 912 8108 946
rect 8108 912 8120 946
rect 8160 912 8176 946
rect 8176 912 8194 946
rect 8234 912 8244 946
rect 8244 912 8268 946
rect 8308 912 8312 946
rect 8312 912 8342 946
rect 8382 912 8414 946
rect 8414 912 8416 946
rect 8456 912 8482 946
rect 8482 912 8490 946
rect 8529 912 8550 946
rect 8550 912 8563 946
rect 8602 912 8618 946
rect 8618 912 8636 946
rect 8675 912 8686 946
rect 8686 912 8709 946
rect 8748 912 8754 946
rect 8754 912 8782 946
rect 8821 912 8822 946
rect 8822 912 8855 946
rect 8894 912 8924 946
rect 8924 912 8928 946
rect 8967 912 8992 946
rect 8992 912 9001 946
rect 9040 912 9060 946
rect 9060 912 9074 946
rect 9113 912 9128 946
rect 9128 912 9147 946
rect 9186 912 9196 946
rect 9196 912 9220 946
rect 9259 912 9264 946
rect 9264 912 9293 946
rect 9332 912 9366 946
rect 9564 912 9568 946
rect 9568 912 9598 946
rect 9637 912 9670 946
rect 9670 912 9671 946
rect 9710 912 9738 946
rect 9738 912 9744 946
rect 9783 912 9806 946
rect 9806 912 9817 946
rect 9856 912 9874 946
rect 9874 912 9890 946
rect 9929 912 9942 946
rect 9942 912 9963 946
rect 10002 912 10010 946
rect 10010 912 10036 946
rect 10075 912 10078 946
rect 10078 912 10109 946
rect 10148 912 10180 946
rect 10180 912 10182 946
rect 10221 912 10248 946
rect 10248 912 10255 946
rect 10294 912 10316 946
rect 10316 912 10328 946
rect 10367 912 10384 946
rect 10384 912 10401 946
rect 10440 912 10452 946
rect 10452 912 10474 946
rect 10514 912 10520 946
rect 10520 912 10548 946
rect 10588 912 10622 946
rect 10662 912 10690 946
rect 10690 912 10696 946
rect 10736 912 10758 946
rect 10758 912 10770 946
rect 10810 912 10826 946
rect 10826 912 10844 946
rect 10884 912 10894 946
rect 10894 912 10918 946
rect 10958 912 10962 946
rect 10962 912 10992 946
rect 11032 912 11064 946
rect 11064 912 11066 946
rect 11106 912 11132 946
rect 11132 912 11140 946
rect 11180 912 11200 946
rect 11200 912 11214 946
rect 11254 912 11268 946
rect 11268 912 11288 946
rect 11328 912 11336 946
rect 11336 912 11362 946
rect 11402 912 11404 946
rect 11404 912 11436 946
rect 11476 912 11506 946
rect 11506 912 11510 946
rect 11566 945 11599 977
rect 11599 945 11600 977
rect 7330 904 7364 905
rect 7330 871 7364 904
rect 7330 797 7364 831
rect 11566 904 11600 905
rect 11566 871 11599 904
rect 11599 871 11600 904
rect 11566 797 11599 831
rect 11599 797 11600 831
rect 7330 724 7364 757
rect 7420 756 7454 790
rect 7494 756 7496 790
rect 7496 756 7528 790
rect 7568 756 7598 790
rect 7598 756 7602 790
rect 7642 756 7666 790
rect 7666 756 7676 790
rect 7716 756 7734 790
rect 7734 756 7750 790
rect 7790 756 7802 790
rect 7802 756 7824 790
rect 7864 756 7870 790
rect 7870 756 7898 790
rect 7938 756 7972 790
rect 8012 756 8040 790
rect 8040 756 8046 790
rect 8086 756 8108 790
rect 8108 756 8120 790
rect 8160 756 8176 790
rect 8176 756 8194 790
rect 8234 756 8244 790
rect 8244 756 8268 790
rect 8308 756 8312 790
rect 8312 756 8342 790
rect 8382 756 8414 790
rect 8414 756 8416 790
rect 8456 756 8482 790
rect 8482 756 8490 790
rect 8529 756 8550 790
rect 8550 756 8563 790
rect 8602 756 8618 790
rect 8618 756 8636 790
rect 8675 756 8686 790
rect 8686 756 8709 790
rect 8748 756 8754 790
rect 8754 756 8782 790
rect 8821 756 8822 790
rect 8822 756 8855 790
rect 8894 756 8924 790
rect 8924 756 8928 790
rect 8967 756 8992 790
rect 8992 756 9001 790
rect 9040 756 9060 790
rect 9060 756 9074 790
rect 9113 756 9128 790
rect 9128 756 9147 790
rect 9186 756 9196 790
rect 9196 756 9220 790
rect 9259 756 9264 790
rect 9264 756 9293 790
rect 9332 756 9366 790
rect 9564 756 9568 790
rect 9568 756 9598 790
rect 9637 756 9670 790
rect 9670 756 9671 790
rect 9710 756 9738 790
rect 9738 756 9744 790
rect 9783 756 9806 790
rect 9806 756 9817 790
rect 9856 756 9874 790
rect 9874 756 9890 790
rect 9929 756 9942 790
rect 9942 756 9963 790
rect 10002 756 10010 790
rect 10010 756 10036 790
rect 10075 756 10078 790
rect 10078 756 10109 790
rect 10148 756 10180 790
rect 10180 756 10182 790
rect 10221 756 10248 790
rect 10248 756 10255 790
rect 10294 756 10316 790
rect 10316 756 10328 790
rect 10367 756 10384 790
rect 10384 756 10401 790
rect 10440 756 10452 790
rect 10452 756 10474 790
rect 10514 756 10520 790
rect 10520 756 10548 790
rect 10588 756 10622 790
rect 10662 756 10690 790
rect 10690 756 10696 790
rect 10736 756 10758 790
rect 10758 756 10770 790
rect 10810 756 10826 790
rect 10826 756 10844 790
rect 10884 756 10894 790
rect 10894 756 10918 790
rect 10958 756 10962 790
rect 10962 756 10992 790
rect 11032 756 11064 790
rect 11064 756 11066 790
rect 11106 756 11132 790
rect 11132 756 11140 790
rect 11180 756 11200 790
rect 11200 756 11214 790
rect 11254 756 11268 790
rect 11268 756 11288 790
rect 11328 756 11336 790
rect 11336 756 11362 790
rect 11402 756 11404 790
rect 11404 756 11436 790
rect 11476 756 11506 790
rect 11506 756 11510 790
rect 7330 723 7364 724
rect 7330 651 7364 683
rect 7330 649 7364 651
rect 11566 724 11599 757
rect 11599 724 11600 757
rect 11566 723 11600 724
rect 11566 651 11599 683
rect 11599 651 11600 683
rect 11566 649 11600 651
rect 7330 578 7364 609
rect 7420 600 7454 634
rect 7494 600 7496 634
rect 7496 600 7528 634
rect 7568 600 7598 634
rect 7598 600 7602 634
rect 7642 600 7666 634
rect 7666 600 7676 634
rect 7716 600 7734 634
rect 7734 600 7750 634
rect 7790 600 7802 634
rect 7802 600 7824 634
rect 7864 600 7870 634
rect 7870 600 7898 634
rect 7938 600 7972 634
rect 8012 600 8040 634
rect 8040 600 8046 634
rect 8086 600 8108 634
rect 8108 600 8120 634
rect 8160 600 8176 634
rect 8176 600 8194 634
rect 8234 600 8244 634
rect 8244 600 8268 634
rect 8308 600 8312 634
rect 8312 600 8342 634
rect 8382 600 8414 634
rect 8414 600 8416 634
rect 8456 600 8482 634
rect 8482 600 8490 634
rect 8529 600 8550 634
rect 8550 600 8563 634
rect 8602 600 8618 634
rect 8618 600 8636 634
rect 8675 600 8686 634
rect 8686 600 8709 634
rect 8748 600 8754 634
rect 8754 600 8782 634
rect 8821 600 8822 634
rect 8822 600 8855 634
rect 8894 600 8924 634
rect 8924 600 8928 634
rect 8967 600 8992 634
rect 8992 600 9001 634
rect 9040 600 9060 634
rect 9060 600 9074 634
rect 9113 600 9128 634
rect 9128 600 9147 634
rect 9186 600 9196 634
rect 9196 600 9220 634
rect 9259 600 9264 634
rect 9264 600 9293 634
rect 9332 600 9366 634
rect 9564 600 9568 634
rect 9568 600 9598 634
rect 9637 600 9670 634
rect 9670 600 9671 634
rect 9710 600 9738 634
rect 9738 600 9744 634
rect 9783 600 9806 634
rect 9806 600 9817 634
rect 9856 600 9874 634
rect 9874 600 9890 634
rect 9929 600 9942 634
rect 9942 600 9963 634
rect 10002 600 10010 634
rect 10010 600 10036 634
rect 10075 600 10078 634
rect 10078 600 10109 634
rect 10148 600 10180 634
rect 10180 600 10182 634
rect 10221 600 10248 634
rect 10248 600 10255 634
rect 10294 600 10316 634
rect 10316 600 10328 634
rect 10367 600 10384 634
rect 10384 600 10401 634
rect 10440 600 10452 634
rect 10452 600 10474 634
rect 10514 600 10520 634
rect 10520 600 10548 634
rect 10588 600 10622 634
rect 10662 600 10690 634
rect 10690 600 10696 634
rect 10736 600 10758 634
rect 10758 600 10770 634
rect 10810 600 10826 634
rect 10826 600 10844 634
rect 10884 600 10894 634
rect 10894 600 10918 634
rect 10958 600 10962 634
rect 10962 600 10992 634
rect 11032 600 11064 634
rect 11064 600 11066 634
rect 11106 600 11132 634
rect 11132 600 11140 634
rect 11180 600 11200 634
rect 11200 600 11214 634
rect 11254 600 11268 634
rect 11268 600 11288 634
rect 11328 600 11336 634
rect 11336 600 11362 634
rect 11402 600 11404 634
rect 11404 600 11436 634
rect 11476 600 11506 634
rect 11506 600 11510 634
rect 7330 575 7364 578
rect 7330 505 7364 535
rect 7330 501 7364 505
rect 11566 578 11599 609
rect 11599 578 11600 609
rect 11566 575 11600 578
rect 11566 505 11599 535
rect 11599 505 11600 535
rect 11566 501 11600 505
rect 7420 444 7454 478
rect 7494 444 7496 478
rect 7496 444 7528 478
rect 7568 444 7598 478
rect 7598 444 7602 478
rect 7642 444 7666 478
rect 7666 444 7676 478
rect 7716 444 7734 478
rect 7734 444 7750 478
rect 7790 444 7802 478
rect 7802 444 7824 478
rect 7864 444 7870 478
rect 7870 444 7898 478
rect 7938 444 7972 478
rect 8012 444 8040 478
rect 8040 444 8046 478
rect 8086 444 8108 478
rect 8108 444 8120 478
rect 8160 444 8176 478
rect 8176 444 8194 478
rect 8234 444 8244 478
rect 8244 444 8268 478
rect 8308 444 8312 478
rect 8312 444 8342 478
rect 8382 444 8414 478
rect 8414 444 8416 478
rect 8456 444 8482 478
rect 8482 444 8490 478
rect 8529 444 8550 478
rect 8550 444 8563 478
rect 8602 444 8618 478
rect 8618 444 8636 478
rect 8675 444 8686 478
rect 8686 444 8709 478
rect 8748 444 8754 478
rect 8754 444 8782 478
rect 8821 444 8822 478
rect 8822 444 8855 478
rect 8894 444 8924 478
rect 8924 444 8928 478
rect 8967 444 8992 478
rect 8992 444 9001 478
rect 9040 444 9060 478
rect 9060 444 9074 478
rect 9113 444 9128 478
rect 9128 444 9147 478
rect 9186 444 9196 478
rect 9196 444 9220 478
rect 9259 444 9264 478
rect 9264 444 9293 478
rect 9332 444 9366 478
rect 9564 444 9568 478
rect 9568 444 9598 478
rect 9637 444 9670 478
rect 9670 444 9671 478
rect 9710 444 9738 478
rect 9738 444 9744 478
rect 9783 444 9806 478
rect 9806 444 9817 478
rect 9856 444 9874 478
rect 9874 444 9890 478
rect 9929 444 9942 478
rect 9942 444 9963 478
rect 10002 444 10010 478
rect 10010 444 10036 478
rect 10075 444 10078 478
rect 10078 444 10109 478
rect 10148 444 10180 478
rect 10180 444 10182 478
rect 10221 444 10248 478
rect 10248 444 10255 478
rect 10294 444 10316 478
rect 10316 444 10328 478
rect 10367 444 10384 478
rect 10384 444 10401 478
rect 10440 444 10452 478
rect 10452 444 10474 478
rect 10514 444 10520 478
rect 10520 444 10548 478
rect 10588 444 10622 478
rect 10662 444 10690 478
rect 10690 444 10696 478
rect 10736 444 10758 478
rect 10758 444 10770 478
rect 10810 444 10826 478
rect 10826 444 10844 478
rect 10884 444 10894 478
rect 10894 444 10918 478
rect 10958 444 10962 478
rect 10962 444 10992 478
rect 11032 444 11064 478
rect 11064 444 11066 478
rect 11106 444 11132 478
rect 11132 444 11140 478
rect 11180 444 11200 478
rect 11200 444 11214 478
rect 11254 444 11268 478
rect 11268 444 11288 478
rect 11328 444 11336 478
rect 11336 444 11362 478
rect 11402 444 11404 478
rect 11404 444 11436 478
rect 11476 444 11506 478
rect 11506 444 11510 478
rect 11645 1312 11751 1368
rect 11645 1278 11681 1312
rect 11681 1278 11715 1312
rect 11715 1278 11751 1312
rect 11645 1244 11751 1278
rect 11645 1210 11681 1244
rect 11681 1210 11715 1244
rect 11715 1210 11751 1244
rect 11645 1176 11751 1210
rect 11645 1142 11681 1176
rect 11681 1142 11715 1176
rect 11715 1142 11751 1176
rect 11645 1108 11751 1142
rect 11645 1074 11681 1108
rect 11681 1074 11715 1108
rect 11715 1074 11751 1108
rect 11645 1040 11751 1074
rect 11645 1006 11681 1040
rect 11681 1006 11715 1040
rect 11715 1006 11751 1040
rect 11645 972 11751 1006
rect 11645 938 11681 972
rect 11681 938 11715 972
rect 11715 938 11751 972
rect 11645 904 11751 938
rect 11645 870 11681 904
rect 11681 870 11715 904
rect 11715 870 11751 904
rect 11645 836 11751 870
rect 11645 802 11681 836
rect 11681 802 11715 836
rect 11715 802 11751 836
rect 11645 768 11751 802
rect 11645 734 11681 768
rect 11681 734 11715 768
rect 11715 734 11751 768
rect 11645 700 11751 734
rect 11645 666 11681 700
rect 11681 666 11715 700
rect 11715 666 11751 700
rect 11645 632 11751 666
rect 11645 598 11681 632
rect 11681 598 11715 632
rect 11715 598 11751 632
rect 11645 564 11751 598
rect 11645 530 11681 564
rect 11681 530 11715 564
rect 11715 530 11751 564
rect 11645 496 11751 530
rect 11645 470 11681 496
rect 11681 470 11715 496
rect 11715 470 11751 496
rect 11645 397 11679 431
rect 11717 397 11751 431
rect 7163 325 7264 359
rect 7264 325 7269 359
rect 7308 325 7332 358
rect 7332 325 7342 358
rect 7381 325 7400 358
rect 7400 325 7415 358
rect 7454 325 7468 358
rect 7468 325 7488 358
rect 7527 325 7536 358
rect 7536 325 7561 358
rect 7600 325 7604 358
rect 7604 325 7634 358
rect 7673 325 7706 358
rect 7706 325 7707 358
rect 7746 325 7774 358
rect 7774 325 7780 358
rect 7819 325 7842 358
rect 7842 325 7853 358
rect 7892 325 7910 358
rect 7910 325 7926 358
rect 7965 325 7978 358
rect 7978 325 7999 358
rect 8038 325 8046 358
rect 8046 325 8072 358
rect 8111 325 8114 358
rect 8114 325 8145 358
rect 8184 325 8216 358
rect 8216 325 8218 358
rect 8257 325 8284 358
rect 8284 325 8291 358
rect 8330 325 8352 358
rect 8352 325 8364 358
rect 8403 325 8420 358
rect 8420 325 8437 358
rect 8476 325 8488 358
rect 8488 325 8510 358
rect 8549 325 8556 358
rect 8556 325 8590 358
rect 8590 325 8624 358
rect 8624 325 8658 358
rect 8658 325 8692 358
rect 8692 325 8726 358
rect 8726 325 8760 358
rect 8760 325 8794 358
rect 8794 325 8828 358
rect 8828 325 8862 358
rect 8862 325 8896 358
rect 8896 325 8930 358
rect 8930 325 8964 358
rect 8964 325 8998 358
rect 8998 325 9032 358
rect 9032 325 9066 358
rect 9066 325 9100 358
rect 9100 325 9134 358
rect 9134 325 9168 358
rect 9168 325 9202 358
rect 9202 325 9236 358
rect 9236 325 9270 358
rect 9270 325 9304 358
rect 9304 325 9338 358
rect 9338 325 9372 358
rect 9372 325 9406 358
rect 9406 325 9440 358
rect 9440 325 9474 358
rect 9474 325 9508 358
rect 9508 325 9542 358
rect 9542 325 9576 358
rect 9576 325 9610 358
rect 9610 325 9644 358
rect 9644 325 9678 358
rect 9678 325 9712 358
rect 9712 325 9746 358
rect 9746 325 9780 358
rect 9780 325 9814 358
rect 9814 325 9848 358
rect 9848 325 9882 358
rect 9882 325 9916 358
rect 9916 325 9950 358
rect 9950 325 9984 358
rect 9984 325 10018 358
rect 10018 325 10052 358
rect 10052 325 10086 358
rect 10086 325 10120 358
rect 10120 325 10154 358
rect 10154 325 10188 358
rect 10188 325 10222 358
rect 10222 325 10256 358
rect 10256 325 10290 358
rect 10290 325 10324 358
rect 10324 325 10358 358
rect 10358 325 10392 358
rect 10392 325 10426 358
rect 10426 325 10460 358
rect 10460 325 10494 358
rect 10494 325 10528 358
rect 10528 325 10562 358
rect 10562 325 10596 358
rect 10596 325 10630 358
rect 10630 325 10664 358
rect 10664 325 10698 358
rect 10698 325 10732 358
rect 10732 325 10766 358
rect 10766 325 10800 358
rect 10800 325 10834 358
rect 10834 325 10868 358
rect 10868 325 10902 358
rect 10902 325 10936 358
rect 10936 325 10970 358
rect 10970 325 11004 358
rect 11004 325 11038 358
rect 11038 325 11072 358
rect 11072 325 11106 358
rect 11106 325 11140 358
rect 11140 325 11174 358
rect 11174 325 11208 358
rect 11208 325 11242 358
rect 11242 325 11276 358
rect 11276 325 11310 358
rect 11310 325 11344 358
rect 11344 325 11378 358
rect 11378 325 11412 358
rect 11412 325 11446 358
rect 11446 325 11480 358
rect 11480 325 11514 358
rect 11514 325 11548 358
rect 11548 325 11582 358
rect 11582 325 11616 358
rect 11616 325 11650 358
rect 11650 325 11679 358
rect 7163 324 7269 325
rect 7308 324 7342 325
rect 7381 324 7415 325
rect 7454 324 7488 325
rect 7527 324 7561 325
rect 7600 324 7634 325
rect 7673 324 7707 325
rect 7746 324 7780 325
rect 7819 324 7853 325
rect 7892 324 7926 325
rect 7965 324 7999 325
rect 8038 324 8072 325
rect 8111 324 8145 325
rect 8184 324 8218 325
rect 8257 324 8291 325
rect 8330 324 8364 325
rect 8403 324 8437 325
rect 8476 324 8510 325
rect 7235 252 7269 286
rect 7308 252 7342 286
rect 7381 252 7415 286
rect 7454 252 7488 286
rect 7527 252 7561 286
rect 7600 252 7634 286
rect 7673 252 7707 286
rect 7746 252 7780 286
rect 7819 252 7853 286
rect 7892 252 7926 286
rect 7965 252 7999 286
rect 8038 252 8072 286
rect 8111 252 8145 286
rect 8184 252 8218 286
rect 8257 252 8291 286
rect 8330 252 8364 286
rect 8403 252 8437 286
rect 8476 252 8510 286
rect 8549 252 11679 325
rect 11717 324 11751 358
rect 6882 171 6988 243
rect 61 137 63 171
rect 63 137 95 171
rect 133 137 165 171
rect 165 137 167 171
rect 206 169 240 171
rect 279 169 313 171
rect 352 169 386 171
rect 425 169 459 171
rect 498 169 532 171
rect 571 169 605 171
rect 644 169 678 171
rect 717 169 751 171
rect 790 169 824 171
rect 863 169 897 171
rect 936 169 970 171
rect 1009 169 1043 171
rect 1082 169 1116 171
rect 1155 169 1189 171
rect 1228 169 1262 171
rect 1301 169 1335 171
rect 1374 169 1408 171
rect 1447 169 1481 171
rect 1520 169 1554 171
rect 1593 169 1627 171
rect 1666 169 1700 171
rect 1739 169 1773 171
rect 1812 169 1846 171
rect 206 137 240 169
rect 279 137 313 169
rect 352 137 386 169
rect 425 137 459 169
rect 498 137 532 169
rect 571 137 605 169
rect 644 137 678 169
rect 717 137 751 169
rect 790 137 824 169
rect 863 137 897 169
rect 936 137 970 169
rect 1009 137 1043 169
rect 1082 137 1116 169
rect 1155 137 1189 169
rect 1228 137 1262 169
rect 1301 137 1335 169
rect 1374 137 1408 169
rect 1447 137 1481 169
rect 1520 137 1554 169
rect 1593 137 1627 169
rect 1666 137 1700 169
rect 1739 137 1773 169
rect 1812 137 1846 169
rect 1885 137 1906 171
rect 1906 137 1919 171
rect 1958 137 1992 171
rect 2031 137 2065 171
rect 2104 169 2138 171
rect 2177 169 2211 171
rect 2250 169 2284 171
rect 2323 169 11861 171
rect 2104 137 2138 169
rect 2177 137 2211 169
rect 2250 137 2284 169
rect 133 67 138 99
rect 138 67 167 99
rect 206 67 240 99
rect 279 67 313 99
rect 352 67 386 99
rect 425 67 459 99
rect 498 67 532 99
rect 571 67 605 99
rect 644 67 678 99
rect 717 67 751 99
rect 790 67 824 99
rect 863 67 897 99
rect 936 67 970 99
rect 1009 67 1043 99
rect 1082 67 1116 99
rect 1155 67 1189 99
rect 1228 67 1262 99
rect 1301 67 1335 99
rect 1374 67 1408 99
rect 1447 67 1481 99
rect 1520 67 1554 99
rect 1593 67 1627 99
rect 1666 67 1700 99
rect 1739 67 1773 99
rect 1812 67 1846 99
rect 133 65 167 67
rect 206 65 240 67
rect 279 65 313 67
rect 352 65 386 67
rect 425 65 459 67
rect 498 65 532 67
rect 571 65 605 67
rect 644 65 678 67
rect 717 65 751 67
rect 790 65 824 67
rect 863 65 897 67
rect 936 65 970 67
rect 1009 65 1043 67
rect 1082 65 1116 67
rect 1155 65 1189 67
rect 1228 65 1262 67
rect 1301 65 1335 67
rect 1374 65 1408 67
rect 1447 65 1481 67
rect 1520 65 1554 67
rect 1593 65 1627 67
rect 1666 65 1700 67
rect 1739 65 1773 67
rect 1812 65 1846 67
rect 1885 65 1919 99
rect 1958 65 1992 99
rect 2031 67 2035 99
rect 2035 67 2065 99
rect 2104 67 2138 99
rect 2177 67 2211 99
rect 2250 67 2284 99
rect 2323 67 6897 169
rect 6897 67 7020 169
rect 7020 67 11814 169
rect 11814 101 11861 169
rect 11814 67 11848 101
rect 11848 67 11861 101
rect 2031 65 2065 67
rect 2104 65 2138 67
rect 2177 65 2211 67
rect 2250 65 2284 67
rect 2323 65 11861 67
rect -496 -217 -462 -183
rect -409 -217 -375 -183
rect -322 -217 -288 -183
rect -236 -217 -202 -183
rect -150 -217 -116 -183
rect -496 -327 -462 -293
rect -409 -327 -375 -293
rect -322 -327 -288 -293
rect -236 -327 -202 -293
rect -150 -327 -116 -293
rect 6483 -1154 6517 -1153
rect 6558 -1154 6592 -1153
rect 6633 -1154 6667 -1153
rect 6708 -1154 6742 -1153
rect 6783 -1154 6817 -1153
rect 6859 -1154 6893 -1153
rect 6935 -1154 6969 -1153
rect 7011 -1154 7045 -1153
rect 7087 -1154 7121 -1153
rect 7197 -1154 7231 -1153
rect 7271 -1154 7305 -1153
rect 7345 -1154 7379 -1153
rect 7419 -1154 7453 -1153
rect 7493 -1154 7527 -1153
rect 7567 -1154 7601 -1153
rect 7641 -1154 7675 -1153
rect 7715 -1154 7749 -1153
rect 7789 -1154 7823 -1153
rect 7863 -1154 7897 -1153
rect 7937 -1154 7971 -1153
rect 8011 -1154 8045 -1153
rect 8085 -1154 8119 -1153
rect 8159 -1154 8193 -1153
rect 8233 -1154 8267 -1153
rect 8307 -1154 8341 -1153
rect 8381 -1154 8415 -1153
rect 8455 -1154 8489 -1153
rect 8529 -1154 8563 -1153
rect 8604 -1154 8638 -1153
rect 8679 -1154 8713 -1153
rect 6483 -1187 6498 -1154
rect 6498 -1187 6517 -1154
rect 6558 -1187 6566 -1154
rect 6566 -1187 6592 -1154
rect 6633 -1187 6634 -1154
rect 6634 -1187 6667 -1154
rect 6708 -1187 6736 -1154
rect 6736 -1187 6742 -1154
rect 6783 -1187 6804 -1154
rect 6804 -1187 6817 -1154
rect 6859 -1187 6872 -1154
rect 6872 -1187 6893 -1154
rect 6935 -1187 6940 -1154
rect 6940 -1187 6969 -1154
rect 7011 -1187 7042 -1154
rect 7042 -1187 7045 -1154
rect 7087 -1187 7110 -1154
rect 7110 -1187 7121 -1154
rect 7197 -1187 7212 -1154
rect 7212 -1187 7231 -1154
rect 7271 -1187 7280 -1154
rect 7280 -1187 7305 -1154
rect 7345 -1187 7348 -1154
rect 7348 -1187 7379 -1154
rect 7419 -1187 7450 -1154
rect 7450 -1187 7453 -1154
rect 7493 -1187 7518 -1154
rect 7518 -1187 7527 -1154
rect 7567 -1187 7586 -1154
rect 7586 -1187 7601 -1154
rect 7641 -1187 7654 -1154
rect 7654 -1187 7675 -1154
rect 7715 -1187 7722 -1154
rect 7722 -1187 7749 -1154
rect 7789 -1187 7790 -1154
rect 7790 -1187 7823 -1154
rect 7863 -1187 7892 -1154
rect 7892 -1187 7897 -1154
rect 7937 -1187 7960 -1154
rect 7960 -1187 7971 -1154
rect 8011 -1187 8028 -1154
rect 8028 -1187 8045 -1154
rect 8085 -1187 8096 -1154
rect 8096 -1187 8119 -1154
rect 8159 -1187 8164 -1154
rect 8164 -1187 8193 -1154
rect 8233 -1187 8266 -1154
rect 8266 -1187 8267 -1154
rect 8307 -1187 8334 -1154
rect 8334 -1187 8341 -1154
rect 8381 -1187 8402 -1154
rect 8402 -1187 8415 -1154
rect 8455 -1187 8470 -1154
rect 8470 -1187 8489 -1154
rect 8529 -1187 8538 -1154
rect 8538 -1187 8563 -1154
rect 8604 -1187 8606 -1154
rect 8606 -1187 8638 -1154
rect 8679 -1187 8708 -1154
rect 8708 -1187 8713 -1154
rect 6417 -1222 6451 -1216
rect 6417 -1250 6451 -1222
rect 8742 -1251 8776 -1217
rect 6417 -1324 6451 -1294
rect 6417 -1328 6451 -1324
rect 6652 -1304 6666 -1270
rect 6666 -1304 6686 -1270
rect 6727 -1304 6734 -1270
rect 6734 -1304 6761 -1270
rect 6802 -1304 6836 -1270
rect 6877 -1304 6904 -1270
rect 6904 -1304 6911 -1270
rect 6952 -1304 6972 -1270
rect 6972 -1304 6986 -1270
rect 7027 -1304 7040 -1270
rect 7040 -1304 7061 -1270
rect 7102 -1304 7108 -1270
rect 7108 -1304 7136 -1270
rect 7177 -1304 7210 -1270
rect 7210 -1304 7211 -1270
rect 7252 -1304 7278 -1270
rect 7278 -1304 7286 -1270
rect 7327 -1304 7346 -1270
rect 7346 -1304 7361 -1270
rect 7402 -1304 7414 -1270
rect 7414 -1304 7436 -1270
rect 7476 -1304 7482 -1270
rect 7482 -1304 7510 -1270
rect 7550 -1304 7584 -1270
rect 7624 -1304 7652 -1270
rect 7652 -1304 7658 -1270
rect 7698 -1304 7720 -1270
rect 7720 -1304 7732 -1270
rect 7772 -1304 7788 -1270
rect 7788 -1304 7806 -1270
rect 7846 -1304 7856 -1270
rect 7856 -1304 7880 -1270
rect 7920 -1304 7924 -1270
rect 7924 -1304 7954 -1270
rect 7994 -1304 8026 -1270
rect 8026 -1304 8028 -1270
rect 8068 -1304 8094 -1270
rect 8094 -1304 8102 -1270
rect 8142 -1304 8162 -1270
rect 8162 -1304 8176 -1270
rect 8216 -1304 8230 -1270
rect 8230 -1304 8250 -1270
rect 8290 -1304 8298 -1270
rect 8298 -1304 8324 -1270
rect 8364 -1304 8366 -1270
rect 8366 -1304 8398 -1270
rect 8438 -1304 8468 -1270
rect 8468 -1304 8472 -1270
rect 8512 -1304 8536 -1270
rect 8536 -1304 8546 -1270
rect 8586 -1304 8604 -1270
rect 8604 -1304 8620 -1270
rect 6417 -1392 6451 -1372
rect 6417 -1406 6451 -1392
rect 6417 -1460 6451 -1450
rect 6417 -1484 6451 -1460
rect 6417 -1562 6451 -1528
rect 6417 -1640 6451 -1606
rect 6417 -1718 6451 -1684
rect 6417 -1792 6451 -1762
rect 6417 -1796 6451 -1792
rect 6417 -1860 6451 -1840
rect 6417 -1874 6451 -1860
rect 6534 -1331 6568 -1327
rect 6534 -1361 6568 -1331
rect 6534 -1402 6568 -1399
rect 6534 -1433 6568 -1402
rect 8742 -1296 8776 -1290
rect 8742 -1324 8776 -1296
rect 8742 -1364 8776 -1363
rect 8742 -1397 8776 -1364
rect 6652 -1460 6666 -1426
rect 6666 -1460 6686 -1426
rect 6727 -1460 6734 -1426
rect 6734 -1460 6761 -1426
rect 6802 -1460 6836 -1426
rect 6877 -1460 6904 -1426
rect 6904 -1460 6911 -1426
rect 6952 -1460 6972 -1426
rect 6972 -1460 6986 -1426
rect 7027 -1460 7040 -1426
rect 7040 -1460 7061 -1426
rect 7102 -1460 7108 -1426
rect 7108 -1460 7136 -1426
rect 7177 -1460 7210 -1426
rect 7210 -1460 7211 -1426
rect 7252 -1460 7278 -1426
rect 7278 -1460 7286 -1426
rect 7327 -1460 7346 -1426
rect 7346 -1460 7361 -1426
rect 7402 -1460 7414 -1426
rect 7414 -1460 7436 -1426
rect 7476 -1460 7482 -1426
rect 7482 -1460 7510 -1426
rect 7550 -1460 7584 -1426
rect 7624 -1460 7652 -1426
rect 7652 -1460 7658 -1426
rect 7698 -1460 7720 -1426
rect 7720 -1460 7732 -1426
rect 7772 -1460 7788 -1426
rect 7788 -1460 7806 -1426
rect 7846 -1460 7856 -1426
rect 7856 -1460 7880 -1426
rect 7920 -1460 7924 -1426
rect 7924 -1460 7954 -1426
rect 7994 -1460 8026 -1426
rect 8026 -1460 8028 -1426
rect 8068 -1460 8094 -1426
rect 8094 -1460 8102 -1426
rect 8142 -1460 8162 -1426
rect 8162 -1460 8176 -1426
rect 8216 -1460 8230 -1426
rect 8230 -1460 8250 -1426
rect 8290 -1460 8298 -1426
rect 8298 -1460 8324 -1426
rect 8364 -1460 8366 -1426
rect 8366 -1460 8398 -1426
rect 8438 -1460 8468 -1426
rect 8468 -1460 8472 -1426
rect 8512 -1460 8536 -1426
rect 8536 -1460 8546 -1426
rect 8586 -1460 8604 -1426
rect 8604 -1460 8620 -1426
rect 6534 -1473 6568 -1472
rect 6534 -1506 6568 -1473
rect 6534 -1579 6568 -1545
rect 8742 -1466 8776 -1436
rect 8742 -1470 8776 -1466
rect 8742 -1534 8776 -1509
rect 8742 -1543 8776 -1534
rect 6652 -1616 6666 -1582
rect 6666 -1616 6686 -1582
rect 6727 -1616 6734 -1582
rect 6734 -1616 6761 -1582
rect 6802 -1616 6836 -1582
rect 6877 -1616 6904 -1582
rect 6904 -1616 6911 -1582
rect 6952 -1616 6972 -1582
rect 6972 -1616 6986 -1582
rect 7027 -1616 7040 -1582
rect 7040 -1616 7061 -1582
rect 7102 -1616 7108 -1582
rect 7108 -1616 7136 -1582
rect 7177 -1616 7210 -1582
rect 7210 -1616 7211 -1582
rect 7252 -1616 7278 -1582
rect 7278 -1616 7286 -1582
rect 7327 -1616 7346 -1582
rect 7346 -1616 7361 -1582
rect 7402 -1616 7414 -1582
rect 7414 -1616 7436 -1582
rect 7476 -1616 7482 -1582
rect 7482 -1616 7510 -1582
rect 7550 -1616 7584 -1582
rect 7624 -1616 7652 -1582
rect 7652 -1616 7658 -1582
rect 7698 -1616 7720 -1582
rect 7720 -1616 7732 -1582
rect 7772 -1616 7788 -1582
rect 7788 -1616 7806 -1582
rect 7846 -1616 7856 -1582
rect 7856 -1616 7880 -1582
rect 7920 -1616 7924 -1582
rect 7924 -1616 7954 -1582
rect 7994 -1616 8026 -1582
rect 8026 -1616 8028 -1582
rect 8068 -1616 8094 -1582
rect 8094 -1616 8102 -1582
rect 8142 -1616 8162 -1582
rect 8162 -1616 8176 -1582
rect 8216 -1616 8230 -1582
rect 8230 -1616 8250 -1582
rect 8290 -1616 8298 -1582
rect 8298 -1616 8324 -1582
rect 8364 -1616 8366 -1582
rect 8366 -1616 8398 -1582
rect 8438 -1616 8468 -1582
rect 8468 -1616 8472 -1582
rect 8512 -1616 8536 -1582
rect 8536 -1616 8546 -1582
rect 8586 -1616 8604 -1582
rect 8604 -1616 8620 -1582
rect 6534 -1651 6568 -1618
rect 6534 -1652 6568 -1651
rect 6534 -1723 6568 -1691
rect 6534 -1725 6568 -1723
rect 8742 -1602 8776 -1582
rect 8742 -1616 8776 -1602
rect 8742 -1670 8776 -1655
rect 8742 -1689 8776 -1670
rect 6534 -1795 6568 -1764
rect 6652 -1772 6666 -1738
rect 6666 -1772 6686 -1738
rect 6727 -1772 6734 -1738
rect 6734 -1772 6761 -1738
rect 6802 -1772 6836 -1738
rect 6877 -1772 6904 -1738
rect 6904 -1772 6911 -1738
rect 6952 -1772 6972 -1738
rect 6972 -1772 6986 -1738
rect 7027 -1772 7040 -1738
rect 7040 -1772 7061 -1738
rect 7102 -1772 7108 -1738
rect 7108 -1772 7136 -1738
rect 7177 -1772 7210 -1738
rect 7210 -1772 7211 -1738
rect 7252 -1772 7278 -1738
rect 7278 -1772 7286 -1738
rect 7327 -1772 7346 -1738
rect 7346 -1772 7361 -1738
rect 7402 -1772 7414 -1738
rect 7414 -1772 7436 -1738
rect 7476 -1772 7482 -1738
rect 7482 -1772 7510 -1738
rect 7550 -1772 7584 -1738
rect 7624 -1772 7652 -1738
rect 7652 -1772 7658 -1738
rect 7698 -1772 7720 -1738
rect 7720 -1772 7732 -1738
rect 7772 -1772 7788 -1738
rect 7788 -1772 7806 -1738
rect 7846 -1772 7856 -1738
rect 7856 -1772 7880 -1738
rect 7920 -1772 7924 -1738
rect 7924 -1772 7954 -1738
rect 7994 -1772 8026 -1738
rect 8026 -1772 8028 -1738
rect 8068 -1772 8094 -1738
rect 8094 -1772 8102 -1738
rect 8142 -1772 8162 -1738
rect 8162 -1772 8176 -1738
rect 8216 -1772 8230 -1738
rect 8230 -1772 8250 -1738
rect 8290 -1772 8298 -1738
rect 8298 -1772 8324 -1738
rect 8364 -1772 8366 -1738
rect 8366 -1772 8398 -1738
rect 8438 -1772 8468 -1738
rect 8468 -1772 8472 -1738
rect 8512 -1772 8536 -1738
rect 8536 -1772 8546 -1738
rect 8586 -1772 8604 -1738
rect 8604 -1772 8620 -1738
rect 8742 -1738 8776 -1728
rect 8742 -1762 8776 -1738
rect 6534 -1798 6568 -1795
rect 6534 -1867 6568 -1837
rect 6534 -1871 6568 -1867
rect 8742 -1806 8776 -1801
rect 8742 -1835 8776 -1806
rect 6417 -1928 6451 -1918
rect 6417 -1952 6451 -1928
rect 6652 -1928 6666 -1894
rect 6666 -1928 6686 -1894
rect 6727 -1928 6734 -1894
rect 6734 -1928 6761 -1894
rect 6802 -1928 6836 -1894
rect 6877 -1928 6904 -1894
rect 6904 -1928 6911 -1894
rect 6952 -1928 6972 -1894
rect 6972 -1928 6986 -1894
rect 7027 -1928 7040 -1894
rect 7040 -1928 7061 -1894
rect 7102 -1928 7108 -1894
rect 7108 -1928 7136 -1894
rect 7177 -1928 7210 -1894
rect 7210 -1928 7211 -1894
rect 7252 -1928 7278 -1894
rect 7278 -1928 7286 -1894
rect 7327 -1928 7346 -1894
rect 7346 -1928 7361 -1894
rect 7402 -1928 7414 -1894
rect 7414 -1928 7436 -1894
rect 7476 -1928 7482 -1894
rect 7482 -1928 7510 -1894
rect 7550 -1928 7584 -1894
rect 7624 -1928 7652 -1894
rect 7652 -1928 7658 -1894
rect 7698 -1928 7720 -1894
rect 7720 -1928 7732 -1894
rect 7772 -1928 7788 -1894
rect 7788 -1928 7806 -1894
rect 7846 -1928 7856 -1894
rect 7856 -1928 7880 -1894
rect 7920 -1928 7924 -1894
rect 7924 -1928 7954 -1894
rect 7994 -1928 8026 -1894
rect 8026 -1928 8028 -1894
rect 8068 -1928 8094 -1894
rect 8094 -1928 8102 -1894
rect 8142 -1928 8162 -1894
rect 8162 -1928 8176 -1894
rect 8216 -1928 8230 -1894
rect 8230 -1928 8250 -1894
rect 8290 -1928 8298 -1894
rect 8298 -1928 8324 -1894
rect 8364 -1928 8366 -1894
rect 8366 -1928 8398 -1894
rect 8438 -1928 8468 -1894
rect 8468 -1928 8472 -1894
rect 8512 -1928 8536 -1894
rect 8536 -1928 8546 -1894
rect 8586 -1928 8604 -1894
rect 8604 -1928 8620 -1894
rect 8742 -1908 8776 -1874
rect 6480 -2010 6514 -1986
rect 6581 -2010 6615 -1986
rect 8742 -1976 8776 -1947
rect 8742 -1981 8776 -1976
rect 6480 -2020 6485 -2010
rect 6485 -2020 6514 -2010
rect 6581 -2020 6587 -2010
rect 6587 -2020 6615 -2010
rect 6735 -2044 6757 -2010
rect 6757 -2044 6769 -2010
rect 6807 -2044 6825 -2010
rect 6825 -2044 6841 -2010
rect 6879 -2044 6893 -2010
rect 6893 -2044 6913 -2010
rect 6951 -2044 6961 -2010
rect 6961 -2044 6985 -2010
rect 7023 -2044 7029 -2010
rect 7029 -2044 7057 -2010
rect 7095 -2044 7097 -2010
rect 7097 -2044 7129 -2010
rect 7167 -2044 7199 -2010
rect 7199 -2044 7201 -2010
rect 7239 -2044 7267 -2010
rect 7267 -2044 7273 -2010
rect 7311 -2044 7335 -2010
rect 7335 -2044 7345 -2010
rect 7383 -2044 7403 -2010
rect 7403 -2044 7417 -2010
rect 7455 -2044 7471 -2010
rect 7471 -2044 7489 -2010
rect 7527 -2044 7539 -2010
rect 7539 -2044 7561 -2010
rect 7599 -2044 7607 -2010
rect 7607 -2044 7633 -2010
rect 7671 -2044 7675 -2010
rect 7675 -2044 7705 -2010
rect 7743 -2044 7777 -2010
rect 7815 -2044 7845 -2010
rect 7845 -2044 7849 -2010
rect 7887 -2044 7913 -2010
rect 7913 -2044 7921 -2010
rect 7959 -2044 7981 -2010
rect 7981 -2044 7993 -2010
rect 8031 -2044 8049 -2010
rect 8049 -2044 8065 -2010
rect 8103 -2044 8117 -2010
rect 8117 -2044 8137 -2010
rect 8175 -2044 8185 -2010
rect 8185 -2044 8209 -2010
rect 8247 -2044 8253 -2010
rect 8253 -2044 8281 -2010
rect 8319 -2044 8321 -2010
rect 8321 -2044 8353 -2010
rect 8391 -2044 8423 -2010
rect 8423 -2044 8425 -2010
rect 8463 -2044 8491 -2010
rect 8491 -2044 8497 -2010
rect 8535 -2044 8559 -2010
rect 8559 -2044 8569 -2010
rect 8607 -2044 8627 -2010
rect 8627 -2044 8641 -2010
rect 8679 -2044 8695 -2010
rect 8695 -2044 8713 -2010
<< metal1 >>
rect -508 1429 -104 1435
rect -508 1395 -496 1429
rect -462 1395 -409 1429
rect -375 1428 -322 1429
rect -288 1428 -236 1429
rect -375 1395 -358 1428
rect -242 1395 -236 1428
rect -202 1395 -150 1429
rect -116 1395 -104 1429
rect -508 1376 -358 1395
rect -306 1376 -294 1395
rect -242 1376 -104 1395
rect -508 1355 -104 1376
rect -508 1319 -358 1355
rect -306 1319 -294 1355
rect -242 1319 -104 1355
rect -508 1285 -496 1319
rect -462 1285 -409 1319
rect -375 1303 -358 1319
rect -242 1303 -236 1319
rect -375 1285 -322 1303
rect -288 1285 -236 1303
rect -202 1285 -150 1319
rect -116 1285 -104 1319
rect -508 1282 -104 1285
rect -508 1279 -358 1282
tri -413 1266 -400 1279 ne
rect -400 1266 -358 1279
tri -400 1232 -366 1266 ne
rect -366 1232 -358 1266
tri -366 1224 -358 1232 ne
rect -306 1230 -294 1282
rect -242 1279 -104 1282
rect 55 1412 173 1444
rect 55 1378 61 1412
rect 95 1378 133 1412
rect 167 1378 173 1412
rect 55 1339 173 1378
rect 55 1305 61 1339
rect 95 1305 133 1339
rect 167 1305 173 1339
rect -242 1266 -198 1279
tri -198 1266 -185 1279 nw
rect 55 1266 173 1305
rect -242 1232 -232 1266
tri -232 1232 -198 1266 nw
rect 55 1232 61 1266
rect 95 1232 133 1266
rect 167 1232 173 1266
rect -242 1230 -240 1232
rect -358 1224 -240 1230
tri -240 1224 -232 1232 nw
rect 55 1193 173 1232
rect 55 1159 61 1193
rect 95 1159 133 1193
rect 167 1159 173 1193
rect 55 1120 173 1159
rect 55 1086 61 1120
rect 95 1086 133 1120
rect 167 1086 173 1120
rect -509 1048 -104 1054
rect -509 932 -490 1048
rect -118 932 -104 1048
rect -509 657 -104 932
rect -509 623 -497 657
rect -463 623 -410 657
rect -376 623 -323 657
rect -289 623 -236 657
rect -202 623 -150 657
rect -116 623 -104 657
rect -509 579 -104 623
rect -509 545 -497 579
rect -463 545 -410 579
rect -376 545 -323 579
rect -289 545 -236 579
rect -202 545 -150 579
rect -116 545 -104 579
rect -509 501 -104 545
rect -509 467 -497 501
rect -463 467 -410 501
rect -376 467 -323 501
rect -289 467 -236 501
rect -202 467 -150 501
rect -116 467 -104 501
rect -509 461 -104 467
rect 55 1047 173 1086
rect 55 1013 61 1047
rect 95 1013 133 1047
rect 167 1013 173 1047
rect 55 974 173 1013
rect 55 940 61 974
rect 95 940 133 974
rect 167 940 173 974
rect 55 901 173 940
rect 55 867 61 901
rect 95 867 133 901
rect 167 867 173 901
rect 55 828 173 867
rect 55 794 61 828
rect 95 794 133 828
rect 167 794 173 828
rect 55 755 173 794
rect 55 721 61 755
rect 95 721 133 755
rect 167 721 173 755
rect 55 682 173 721
rect 55 648 61 682
rect 95 648 133 682
rect 167 648 173 682
rect 55 609 173 648
rect 55 575 61 609
rect 95 575 133 609
rect 167 575 173 609
rect 55 536 173 575
rect 55 502 61 536
rect 95 502 133 536
rect 167 502 173 536
rect 55 463 173 502
rect 55 429 61 463
rect 95 429 133 463
rect 167 429 173 463
rect 55 390 173 429
rect 55 356 61 390
rect 95 356 133 390
rect 167 356 173 390
rect 55 317 173 356
rect 55 283 61 317
rect 95 283 133 317
rect 167 283 173 317
rect 318 1437 1748 1443
rect 318 1403 402 1437
rect 436 1403 480 1437
rect 514 1403 558 1437
rect 592 1403 636 1437
rect 670 1403 714 1437
rect 748 1403 792 1437
rect 826 1403 870 1437
rect 904 1403 949 1437
rect 983 1403 1059 1437
rect 318 1365 1059 1403
rect 318 1331 324 1365
rect 358 1331 396 1365
rect 430 1331 480 1365
rect 514 1331 558 1365
rect 592 1331 636 1365
rect 670 1331 714 1365
rect 748 1331 792 1365
rect 826 1331 870 1365
rect 904 1331 949 1365
rect 983 1331 1059 1365
rect 1597 1403 1636 1437
rect 1670 1403 1748 1437
rect 1597 1365 1748 1403
rect 1597 1331 1636 1365
rect 1670 1363 1748 1365
rect 1670 1331 1708 1363
rect 318 1329 1708 1331
rect 1742 1329 1748 1363
rect 318 1325 1748 1329
rect 318 1315 473 1325
tri 473 1315 483 1325 nw
tri 1583 1315 1593 1325 ne
rect 1593 1315 1748 1325
rect 318 1305 463 1315
tri 463 1305 473 1315 nw
tri 1593 1305 1603 1315 ne
rect 1603 1305 1748 1315
rect 318 1290 447 1305
rect 318 1256 324 1290
rect 358 1256 396 1290
rect 430 1289 447 1290
tri 447 1289 463 1305 nw
tri 1603 1289 1619 1305 ne
rect 1619 1289 1748 1305
rect 430 1256 436 1289
tri 436 1278 447 1289 nw
tri 1619 1278 1630 1289 ne
rect 318 1215 436 1256
rect 1630 1255 1636 1289
rect 1670 1255 1708 1289
rect 1742 1255 1748 1289
rect 318 1181 324 1215
rect 358 1181 396 1215
rect 430 1181 436 1215
rect 554 1235 1504 1241
rect 554 1201 566 1235
rect 600 1224 641 1235
rect 675 1224 716 1235
rect 750 1224 791 1235
rect 825 1224 866 1235
rect 900 1224 940 1235
rect 600 1201 640 1224
rect 554 1195 640 1201
tri 606 1187 614 1195 ne
rect 614 1187 640 1195
rect 318 1140 436 1181
rect 318 1106 324 1140
rect 358 1106 396 1140
rect 430 1106 436 1140
rect 318 1065 436 1106
rect 318 1049 324 1065
rect 358 1049 396 1065
rect 430 1049 436 1065
rect 318 997 320 1049
rect 372 997 384 1049
rect 318 990 436 997
rect 318 958 324 990
rect 358 958 396 990
rect 430 958 436 990
rect 318 906 320 958
rect 372 906 384 958
rect 318 881 324 906
rect 358 881 396 906
rect 430 881 436 906
rect 318 867 436 881
rect 318 815 320 867
rect 372 815 384 867
rect 318 807 324 815
rect 358 807 396 815
rect 430 807 436 815
rect 318 767 436 807
rect 318 733 324 767
rect 358 733 396 767
rect 430 733 436 767
rect 318 693 436 733
rect 318 659 324 693
rect 358 659 396 693
rect 430 659 436 693
rect 318 619 436 659
rect 318 585 324 619
rect 358 585 396 619
rect 430 585 436 619
rect 318 545 436 585
rect 318 511 324 545
rect 358 511 396 545
rect 430 511 436 545
rect 318 471 436 511
rect 318 437 324 471
rect 358 437 396 471
rect 430 437 436 471
rect 467 1175 519 1187
tri 614 1181 620 1187 ne
rect 620 1181 640 1187
rect 467 1141 476 1175
rect 510 1141 519 1175
tri 620 1167 634 1181 ne
rect 634 1172 640 1181
rect 692 1172 712 1224
rect 764 1172 784 1224
rect 836 1172 855 1224
rect 907 1201 940 1224
rect 974 1201 1014 1235
rect 1048 1201 1088 1235
rect 1122 1201 1162 1235
rect 1196 1201 1236 1235
rect 1270 1201 1310 1235
rect 1344 1201 1384 1235
rect 1418 1201 1458 1235
rect 1492 1201 1504 1235
rect 907 1195 1504 1201
rect 1630 1215 1748 1255
rect 907 1181 927 1195
tri 927 1181 941 1195 nw
rect 1630 1181 1636 1215
rect 1670 1181 1708 1215
rect 1742 1181 1748 1215
rect 907 1172 913 1181
rect 467 1102 519 1141
rect 467 1068 476 1102
rect 510 1068 519 1102
rect 467 1029 519 1068
rect 467 995 476 1029
rect 510 995 519 1029
rect 467 956 519 995
rect 467 922 476 956
rect 510 922 519 956
rect 634 1160 913 1172
tri 913 1167 927 1181 nw
rect 634 1108 640 1160
rect 692 1108 712 1160
rect 764 1108 784 1160
rect 836 1108 855 1160
rect 907 1108 913 1160
rect 1630 1141 1748 1181
tri 624 945 634 955 se
rect 634 945 913 1108
rect 1112 1081 1118 1133
rect 1170 1081 1195 1133
rect 1247 1081 1272 1133
rect 1324 1081 1348 1133
rect 1400 1081 1424 1133
rect 1476 1081 1500 1133
rect 1552 1081 1558 1133
rect 1112 1076 1558 1081
rect 1112 1055 1124 1076
rect 1158 1055 1202 1076
rect 1236 1055 1280 1076
rect 1314 1055 1358 1076
rect 1392 1055 1435 1076
rect 1469 1055 1512 1076
rect 1546 1055 1558 1076
rect 1112 1003 1118 1055
rect 1170 1003 1195 1055
rect 1247 1003 1272 1055
rect 1324 1003 1348 1055
rect 1400 1003 1424 1055
rect 1476 1003 1500 1055
rect 1552 1003 1558 1055
rect 1630 1107 1636 1141
rect 1670 1107 1708 1141
rect 1742 1107 1748 1141
rect 1630 1067 1748 1107
rect 1630 1033 1636 1067
rect 1670 1033 1708 1067
rect 1742 1033 1748 1067
rect 1630 993 1748 1033
rect 1630 959 1636 993
rect 1670 959 1708 993
rect 1742 959 1748 993
tri 913 945 924 956 sw
tri 619 940 624 945 se
rect 624 940 924 945
tri 924 940 929 945 sw
tri 606 927 619 940 se
rect 619 927 929 940
tri 929 927 942 940 sw
rect 1630 931 1748 959
rect 467 883 519 922
rect 467 849 476 883
rect 510 849 519 883
rect 554 921 1504 927
rect 554 887 566 921
rect 600 887 641 921
rect 675 887 716 921
rect 750 887 791 921
rect 825 887 866 921
rect 900 887 940 921
rect 974 887 1014 921
rect 1048 887 1088 921
rect 1122 887 1162 921
rect 1196 887 1236 921
rect 1270 887 1310 921
rect 1344 887 1384 921
rect 1418 887 1458 921
rect 1492 887 1504 921
rect 554 881 1504 887
rect 467 810 519 849
rect 467 776 476 810
rect 510 776 519 810
rect 1630 815 1631 931
rect 1747 815 1748 931
rect 1630 811 1636 815
rect 1670 811 1708 815
rect 1742 811 1748 815
rect 467 738 519 776
rect 554 790 1504 796
rect 554 756 566 790
rect 600 759 641 790
rect 675 759 716 790
rect 750 759 791 790
rect 825 759 866 790
rect 900 759 940 790
rect 600 756 640 759
rect 554 750 640 756
rect 467 704 476 738
rect 510 704 519 738
tri 596 736 610 750 ne
rect 610 736 640 750
tri 610 723 623 736 ne
rect 623 723 640 736
tri 623 722 624 723 ne
rect 624 722 640 723
tri 624 721 625 722 ne
rect 625 721 640 722
tri 625 717 629 721 ne
rect 467 666 519 704
rect 467 632 476 666
rect 510 632 519 666
rect 467 594 519 632
rect 467 560 476 594
rect 510 560 519 594
rect 467 522 519 560
rect 467 496 476 522
rect 510 496 519 522
rect 629 707 640 721
rect 692 707 712 759
rect 764 707 784 759
rect 836 707 855 759
rect 907 756 940 759
rect 974 756 1014 790
rect 1048 756 1088 790
rect 1122 756 1162 790
rect 1196 756 1236 790
rect 1270 756 1310 790
rect 1344 756 1384 790
rect 1418 756 1458 790
rect 1492 756 1504 790
rect 907 750 1504 756
rect 1630 770 1748 811
rect 907 736 928 750
tri 928 736 942 750 nw
rect 1630 736 1636 770
rect 1670 736 1708 770
rect 1742 736 1748 770
rect 907 723 915 736
tri 915 723 928 736 nw
rect 907 707 914 723
tri 914 722 915 723 nw
rect 629 695 914 707
rect 629 643 640 695
rect 692 643 712 695
rect 764 643 784 695
rect 836 643 855 695
rect 907 643 914 695
rect 1630 695 1748 736
rect 629 511 914 643
rect 1111 630 1117 682
rect 1169 630 1194 682
rect 1246 630 1271 682
rect 1323 630 1348 682
rect 1400 630 1424 682
rect 1476 630 1500 682
rect 1552 630 1558 682
rect 1111 604 1123 630
rect 1157 604 1201 630
rect 1235 604 1279 630
rect 1313 604 1357 630
rect 1391 604 1435 630
rect 1469 604 1512 630
rect 1546 604 1558 630
rect 1111 552 1117 604
rect 1169 552 1194 604
rect 1246 552 1271 604
rect 1323 552 1348 604
rect 1400 552 1424 604
rect 1476 552 1500 604
rect 1552 552 1558 604
rect 1630 661 1636 695
rect 1670 661 1708 695
rect 1742 661 1748 695
rect 1630 620 1748 661
rect 1630 586 1636 620
rect 1670 586 1708 620
rect 1742 586 1748 620
rect 1630 545 1748 586
tri 914 511 915 512 sw
rect 1630 511 1636 545
rect 1670 511 1708 545
rect 1742 511 1748 545
rect 629 501 915 511
tri 915 501 925 511 sw
rect 629 496 925 501
tri 925 496 930 501 sw
rect 467 444 473 496
rect 525 444 537 496
rect 589 444 595 496
rect 629 484 930 496
tri 930 484 942 496 sw
rect 629 478 1504 484
rect 629 444 641 478
rect 675 444 716 478
rect 750 444 791 478
rect 825 444 866 478
rect 900 444 940 478
rect 974 444 1014 478
rect 1048 444 1088 478
rect 1122 444 1162 478
rect 1196 444 1236 478
rect 1270 444 1310 478
rect 1344 444 1384 478
rect 1418 444 1458 478
rect 1492 444 1504 478
rect 1630 470 1748 511
rect 629 438 1504 444
tri 1620 438 1630 448 se
rect 1630 438 1636 470
rect 318 428 436 437
tri 1618 436 1620 438 se
rect 1620 436 1636 438
rect 1670 436 1708 470
rect 1742 436 1748 470
tri 1616 434 1618 436 se
rect 1618 434 1748 436
tri 436 428 442 434 sw
tri 1610 428 1616 434 se
rect 1616 428 1748 434
rect 318 401 442 428
tri 442 401 469 428 sw
tri 1583 401 1610 428 se
rect 1610 401 1748 428
rect 318 397 1748 401
rect 318 363 324 397
rect 358 395 1748 397
rect 358 363 396 395
rect 318 361 396 363
rect 430 361 469 395
rect 503 361 542 395
rect 576 361 615 395
rect 649 361 688 395
rect 722 361 761 395
rect 795 361 834 395
rect 868 361 907 395
rect 941 361 980 395
rect 1014 361 1053 395
rect 1087 361 1126 395
rect 1160 361 1199 395
rect 1233 361 1272 395
rect 1306 361 1345 395
rect 1379 361 1418 395
rect 1452 361 1491 395
rect 1525 361 1564 395
rect 318 323 1564 361
rect 318 289 396 323
rect 430 289 469 323
rect 503 289 542 323
rect 576 289 615 323
rect 649 289 688 323
rect 722 289 761 323
rect 795 289 834 323
rect 868 289 907 323
rect 941 289 980 323
rect 1014 289 1053 323
rect 1087 289 1126 323
rect 1160 289 1199 323
rect 1233 289 1272 323
rect 1306 289 1345 323
rect 1379 289 1418 323
rect 1452 289 1491 323
rect 1525 289 1564 323
rect 1670 361 1708 395
rect 1742 361 1748 395
rect 1670 289 1748 361
rect 318 283 1748 289
rect 1898 1438 2016 1455
rect 1898 1423 1931 1438
rect 1983 1423 2016 1438
rect 1898 1389 1904 1423
rect 2010 1389 2016 1423
rect 1898 1386 1931 1389
rect 1983 1386 2016 1389
rect 1898 1365 2016 1386
rect 1898 1349 1931 1365
rect 1983 1349 2016 1365
rect 1898 1315 1904 1349
rect 2010 1315 2016 1349
rect 1898 1313 1931 1315
rect 1983 1313 2016 1315
rect 1898 1291 2016 1313
rect 1898 1275 1931 1291
rect 1983 1275 2016 1291
rect 1898 1241 1904 1275
rect 2010 1241 2016 1275
rect 1898 1239 1931 1241
rect 1983 1239 2016 1241
rect 1898 1201 2016 1239
rect 1898 1167 1904 1201
rect 1938 1167 1976 1201
rect 2010 1167 2016 1201
rect 1898 1127 2016 1167
rect 1898 1093 1904 1127
rect 1938 1093 1976 1127
rect 2010 1093 2016 1127
rect 1898 1053 2016 1093
rect 1898 1019 1904 1053
rect 1938 1019 1976 1053
rect 2010 1019 2016 1053
rect 1898 979 2016 1019
rect 1898 945 1904 979
rect 1938 945 1976 979
rect 2010 945 2016 979
rect 1898 905 2016 945
rect 1898 871 1904 905
rect 1938 871 1976 905
rect 2010 871 2016 905
rect 1898 831 2016 871
rect 1898 797 1904 831
rect 1938 797 1976 831
rect 2010 797 2016 831
rect 1898 757 2016 797
rect 1898 723 1904 757
rect 1938 723 1976 757
rect 2010 723 2016 757
rect 1898 683 2016 723
rect 1898 649 1904 683
rect 1938 649 1976 683
rect 2010 649 2016 683
rect 1898 609 2016 649
rect 1898 575 1904 609
rect 1938 575 1976 609
rect 2010 575 2016 609
rect 1898 535 2016 575
rect 1898 501 1904 535
rect 1938 501 1976 535
rect 2010 501 2016 535
rect 1898 462 2016 501
rect 1898 428 1904 462
rect 1938 428 1976 462
rect 2010 428 2016 462
rect 1898 389 2016 428
rect 1898 355 1904 389
rect 1938 355 1976 389
rect 2010 355 2016 389
rect 1898 316 2016 355
rect 55 244 173 283
rect 55 210 61 244
rect 95 210 133 244
rect 167 210 173 244
rect 1898 282 1904 316
rect 1938 282 1976 316
rect 2010 282 2016 316
rect 1898 243 2016 282
rect 2153 1450 3599 1456
rect 3651 1450 3665 1456
rect 3717 1450 3731 1456
rect 3783 1450 3797 1456
rect 3849 1450 3863 1456
rect 3915 1450 3929 1456
rect 3981 1450 3995 1456
rect 2153 1416 2237 1450
rect 2271 1416 2315 1450
rect 2349 1416 2393 1450
rect 2427 1416 2471 1450
rect 2505 1416 2549 1450
rect 2583 1416 2627 1450
rect 2661 1416 2705 1450
rect 2739 1416 2784 1450
rect 2818 1416 2894 1450
rect 2928 1416 2967 1450
rect 3001 1416 3040 1450
rect 3074 1416 3113 1450
rect 3147 1416 3186 1450
rect 3220 1416 3259 1450
rect 3293 1416 3332 1450
rect 3366 1416 3405 1450
rect 3439 1416 3478 1450
rect 3512 1416 3551 1450
rect 3585 1416 3599 1450
rect 3658 1416 3665 1450
rect 3915 1416 3916 1450
rect 3981 1416 3989 1450
rect 2153 1404 3599 1416
rect 3651 1404 3665 1416
rect 3717 1404 3731 1416
rect 3783 1404 3797 1416
rect 3849 1404 3863 1416
rect 3915 1404 3929 1416
rect 3981 1404 3995 1416
rect 4047 1404 4061 1456
rect 4113 1404 4127 1456
rect 4179 1404 4193 1456
rect 4245 1404 4259 1456
rect 4311 1450 4325 1456
rect 4377 1450 4391 1456
rect 4443 1450 4457 1456
rect 4509 1450 4523 1456
rect 4575 1450 4589 1456
rect 4641 1450 4655 1456
rect 4707 1450 4721 1456
rect 4315 1416 4325 1450
rect 4388 1416 4391 1450
rect 4641 1416 4646 1450
rect 4707 1416 4719 1450
rect 4311 1404 4325 1416
rect 4377 1404 4391 1416
rect 4443 1404 4457 1416
rect 4509 1404 4523 1416
rect 4575 1404 4589 1416
rect 4641 1404 4655 1416
rect 4707 1404 4721 1416
rect 4773 1404 4786 1456
rect 4838 1404 4851 1456
rect 4903 1404 4916 1456
rect 4968 1450 4981 1456
rect 5033 1450 5046 1456
rect 5098 1450 5111 1456
rect 5163 1450 5176 1456
rect 5228 1450 5241 1456
rect 5293 1450 6626 1456
rect 4972 1416 4981 1450
rect 5045 1416 5046 1450
rect 5228 1416 5230 1450
rect 5293 1416 5303 1450
rect 5337 1416 5376 1450
rect 5410 1416 5449 1450
rect 5483 1416 5522 1450
rect 5556 1416 5595 1450
rect 5629 1416 5668 1450
rect 5702 1416 5741 1450
rect 5775 1416 5814 1450
rect 5848 1416 5887 1450
rect 5921 1416 5961 1450
rect 5995 1416 6035 1450
rect 6069 1416 6109 1450
rect 6143 1416 6183 1450
rect 6217 1416 6257 1450
rect 6291 1416 6331 1450
rect 6365 1416 6405 1450
rect 6439 1416 6479 1450
rect 6513 1416 6553 1450
rect 6587 1416 6626 1450
rect 4968 1404 4981 1416
rect 5033 1404 5046 1416
rect 5098 1404 5111 1416
rect 5163 1404 5176 1416
rect 5228 1404 5241 1416
rect 5293 1404 6626 1416
rect 6678 1404 6731 1456
rect 6783 1404 6789 1456
rect 6876 1424 6994 1456
rect 8735 1446 8741 1454
rect 2153 1392 6789 1404
rect 2153 1378 3599 1392
rect 3651 1378 3665 1392
rect 3717 1378 3731 1392
rect 3783 1378 3797 1392
rect 3849 1378 3863 1392
rect 3915 1378 3929 1392
rect 3981 1378 3995 1392
rect 2153 1344 2159 1378
rect 2193 1344 2231 1378
rect 2265 1344 2315 1378
rect 2349 1344 2393 1378
rect 2427 1344 2471 1378
rect 2505 1344 2549 1378
rect 2583 1344 2627 1378
rect 2661 1344 2705 1378
rect 2739 1344 2784 1378
rect 2818 1344 2894 1378
rect 2928 1344 2967 1378
rect 3001 1344 3040 1378
rect 3074 1344 3113 1378
rect 3147 1344 3186 1378
rect 3220 1344 3259 1378
rect 3293 1344 3332 1378
rect 3366 1344 3405 1378
rect 3439 1344 3478 1378
rect 3512 1344 3551 1378
rect 3585 1344 3599 1378
rect 3658 1344 3665 1378
rect 3915 1344 3916 1378
rect 3981 1344 3989 1378
rect 2153 1340 3599 1344
rect 3651 1340 3665 1344
rect 3717 1340 3731 1344
rect 3783 1340 3797 1344
rect 3849 1340 3863 1344
rect 3915 1340 3929 1344
rect 3981 1340 3995 1344
rect 4047 1340 4061 1392
rect 4113 1340 4127 1392
rect 4179 1340 4193 1392
rect 4245 1340 4259 1392
rect 4311 1378 4325 1392
rect 4377 1378 4391 1392
rect 4443 1378 4457 1392
rect 4509 1378 4523 1392
rect 4575 1378 4589 1392
rect 4641 1378 4655 1392
rect 4707 1378 4721 1392
rect 4315 1344 4325 1378
rect 4388 1344 4391 1378
rect 4641 1344 4646 1378
rect 4707 1344 4719 1378
rect 4311 1340 4325 1344
rect 4377 1340 4391 1344
rect 4443 1340 4457 1344
rect 4509 1340 4523 1344
rect 4575 1340 4589 1344
rect 4641 1340 4655 1344
rect 4707 1340 4721 1344
rect 4773 1340 4786 1392
rect 4838 1340 4851 1392
rect 4903 1340 4916 1392
rect 4968 1378 4981 1392
rect 5033 1378 5046 1392
rect 5098 1378 5111 1392
rect 5163 1378 5176 1392
rect 5228 1378 5241 1392
rect 5293 1378 6626 1392
rect 6678 1378 6731 1392
rect 6783 1390 6789 1392
tri 6789 1390 6805 1406 sw
rect 6876 1390 6882 1424
rect 6916 1390 6954 1424
rect 6988 1390 6994 1424
rect 4972 1344 4981 1378
rect 5045 1344 5046 1378
rect 5228 1344 5230 1378
rect 5293 1344 5303 1378
rect 5337 1344 5376 1378
rect 5410 1344 5449 1378
rect 5483 1344 5522 1378
rect 5556 1344 5595 1378
rect 5629 1344 5668 1378
rect 5702 1344 5741 1378
rect 5775 1344 5814 1378
rect 5848 1344 5887 1378
rect 5921 1344 5961 1378
rect 5995 1344 6035 1378
rect 6069 1344 6109 1378
rect 6143 1344 6183 1378
rect 6217 1344 6257 1378
rect 6291 1344 6331 1378
rect 6365 1344 6405 1378
rect 6439 1344 6479 1378
rect 6513 1344 6553 1378
rect 6587 1344 6626 1378
rect 4968 1340 4981 1344
rect 5033 1340 5046 1344
rect 5098 1340 5111 1344
rect 5163 1340 5176 1344
rect 5228 1340 5241 1344
rect 5293 1340 6626 1344
rect 6783 1368 6805 1390
tri 6805 1368 6827 1390 sw
rect 6783 1355 6827 1368
tri 6827 1355 6840 1368 sw
rect 6783 1340 6840 1355
rect 2153 1338 6627 1340
rect 2153 1305 2271 1338
rect 2153 1271 2159 1305
rect 2193 1271 2231 1305
rect 2265 1271 2271 1305
tri 2271 1291 2318 1338 nw
tri 6556 1291 6603 1338 ne
rect 6603 1328 6627 1338
rect 6733 1328 6840 1340
rect 6603 1291 6626 1328
tri 6603 1276 6618 1291 ne
rect 6618 1276 6626 1291
rect 6783 1276 6840 1328
tri 6618 1273 6621 1276 ne
rect 2153 1232 2271 1271
tri 3127 1264 3130 1267 se
rect 3130 1264 3136 1267
rect 2153 1206 2159 1232
rect 2193 1206 2231 1232
rect 2265 1206 2271 1232
rect 2389 1258 3136 1264
rect 2389 1224 2401 1258
rect 2435 1224 2475 1258
rect 2509 1224 2549 1258
rect 2583 1224 2623 1258
rect 2657 1224 2697 1258
rect 2731 1224 2771 1258
rect 2805 1224 2845 1258
rect 2879 1224 2919 1258
rect 2953 1224 2993 1258
rect 3027 1224 3067 1258
rect 3101 1224 3136 1258
rect 2389 1218 3136 1224
tri 3127 1215 3130 1218 ne
rect 3130 1215 3136 1218
rect 3188 1215 3203 1267
rect 3255 1215 3269 1267
rect 3321 1258 3335 1267
rect 3387 1258 3401 1267
rect 3453 1264 3459 1267
tri 3459 1264 3462 1267 sw
tri 5816 1264 5819 1267 se
rect 5819 1264 5870 1267
rect 3453 1258 4359 1264
rect 3323 1224 3335 1258
rect 3397 1224 3401 1258
rect 3471 1224 3510 1258
rect 3544 1224 3583 1258
rect 3617 1224 3656 1258
rect 3690 1224 3729 1258
rect 3763 1224 3802 1258
rect 3836 1224 3875 1258
rect 3909 1224 3948 1258
rect 3982 1224 4021 1258
rect 4055 1224 4094 1258
rect 4128 1224 4167 1258
rect 4201 1224 4240 1258
rect 4274 1224 4313 1258
rect 4347 1224 4359 1258
rect 3321 1215 3335 1224
rect 3387 1215 3401 1224
rect 3453 1218 4359 1224
rect 4533 1258 5870 1264
rect 4533 1224 4545 1258
rect 4579 1224 4618 1258
rect 4652 1224 4691 1258
rect 4725 1224 4764 1258
rect 4798 1224 4837 1258
rect 4871 1224 4910 1258
rect 4944 1224 4983 1258
rect 5017 1224 5056 1258
rect 5090 1224 5129 1258
rect 5163 1224 5202 1258
rect 5236 1224 5275 1258
rect 5309 1224 5348 1258
rect 5382 1224 5421 1258
rect 5455 1224 5495 1258
rect 5529 1224 5569 1258
rect 5603 1224 5643 1258
rect 5677 1224 5717 1258
rect 5751 1224 5791 1258
rect 5825 1224 5865 1258
rect 4533 1218 5870 1224
rect 3453 1215 3459 1218
tri 3459 1215 3462 1218 nw
tri 5816 1215 5819 1218 ne
rect 5819 1215 5870 1218
rect 5922 1215 5935 1267
rect 5987 1215 5999 1267
rect 6051 1215 6063 1267
rect 6115 1258 6127 1267
rect 6179 1258 6191 1267
rect 6243 1258 6255 1267
rect 6307 1258 6319 1267
rect 6121 1224 6127 1258
rect 6307 1224 6309 1258
rect 6115 1215 6127 1224
rect 6179 1215 6191 1224
rect 6243 1215 6255 1224
rect 6307 1215 6319 1224
rect 6371 1215 6383 1267
rect 6435 1215 6447 1267
rect 6499 1215 6505 1267
rect 2153 1154 2154 1206
rect 2206 1154 2218 1206
rect 2270 1154 2271 1206
rect 2153 1140 2159 1154
rect 2193 1140 2231 1154
rect 2265 1140 2271 1154
rect 2153 1088 2154 1140
rect 2206 1088 2218 1140
rect 2270 1088 2271 1140
rect 2153 1086 2271 1088
rect 2153 1074 2159 1086
rect 2193 1074 2231 1086
rect 2265 1074 2271 1086
rect 2153 1022 2154 1074
rect 2206 1022 2218 1074
rect 2270 1022 2271 1074
rect 2153 1013 2271 1022
rect 2153 979 2159 1013
rect 2193 979 2231 1013
rect 2265 979 2271 1013
rect 2153 940 2271 979
rect 2153 906 2159 940
rect 2193 906 2231 940
rect 2265 906 2271 940
rect 2153 867 2271 906
rect 2153 833 2159 867
rect 2193 833 2231 867
rect 2265 833 2271 867
rect 2153 794 2271 833
rect 2153 760 2159 794
rect 2193 760 2231 794
rect 2265 760 2271 794
rect 2153 721 2271 760
rect 2153 687 2159 721
rect 2193 687 2231 721
rect 2265 687 2271 721
rect 2153 648 2271 687
rect 2305 1207 2357 1213
rect 2305 1137 2357 1155
rect 6539 1207 6591 1213
rect 6539 1137 6591 1155
tri 3590 1108 3593 1111 se
rect 3593 1108 3599 1111
rect 2305 1067 2357 1085
rect 2389 1102 3599 1108
rect 3651 1102 3670 1111
rect 3722 1102 3741 1111
rect 3793 1102 3811 1111
rect 3863 1102 3881 1111
rect 3933 1102 3951 1111
rect 2389 1068 2401 1102
rect 2435 1068 2475 1102
rect 2509 1068 2549 1102
rect 2583 1068 2623 1102
rect 2657 1068 2697 1102
rect 2731 1068 2771 1102
rect 2805 1068 2845 1102
rect 2879 1068 2919 1102
rect 2953 1068 2993 1102
rect 3027 1068 3067 1102
rect 3101 1068 3141 1102
rect 3175 1068 3215 1102
rect 3249 1068 3289 1102
rect 3323 1068 3363 1102
rect 3397 1068 3437 1102
rect 3471 1068 3510 1102
rect 3544 1068 3583 1102
rect 3651 1068 3656 1102
rect 3722 1068 3729 1102
rect 3793 1068 3802 1102
rect 3863 1068 3875 1102
rect 3933 1068 3948 1102
rect 2389 1062 3599 1068
tri 3590 1059 3593 1062 ne
rect 3593 1059 3599 1062
rect 3651 1059 3670 1068
rect 3722 1059 3741 1068
rect 3793 1059 3811 1068
rect 3863 1059 3881 1068
rect 3933 1059 3951 1068
rect 4003 1059 4021 1111
rect 4073 1059 4091 1111
rect 4143 1059 4161 1111
rect 4213 1059 4231 1111
rect 4283 1059 4301 1111
rect 4353 1059 4359 1111
rect 4533 1059 4539 1111
rect 4591 1059 4609 1111
rect 4661 1059 4679 1111
rect 4731 1059 4749 1111
rect 4801 1059 4819 1111
rect 4871 1059 4889 1111
rect 4941 1102 4959 1111
rect 5011 1102 5029 1111
rect 5081 1102 5099 1111
rect 5151 1102 5170 1111
rect 5222 1102 5241 1111
rect 5293 1108 5299 1111
tri 5299 1108 5302 1111 sw
rect 5293 1102 6503 1108
rect 4944 1068 4959 1102
rect 5017 1068 5029 1102
rect 5090 1068 5099 1102
rect 5163 1068 5170 1102
rect 5236 1068 5241 1102
rect 5309 1068 5348 1102
rect 5382 1068 5421 1102
rect 5455 1068 5495 1102
rect 5529 1068 5569 1102
rect 5603 1068 5643 1102
rect 5677 1068 5717 1102
rect 5751 1068 5791 1102
rect 5825 1068 5865 1102
rect 5899 1068 5939 1102
rect 5973 1068 6013 1102
rect 6047 1068 6087 1102
rect 6121 1068 6161 1102
rect 6195 1068 6235 1102
rect 6269 1068 6309 1102
rect 6343 1068 6383 1102
rect 6417 1068 6457 1102
rect 6491 1068 6503 1102
rect 4941 1059 4959 1068
rect 5011 1059 5029 1068
rect 5081 1059 5099 1068
rect 5151 1059 5170 1068
rect 5222 1059 5241 1068
rect 5293 1062 6503 1068
rect 6539 1084 6547 1085
rect 6581 1084 6591 1085
rect 6539 1067 6591 1084
rect 5293 1059 5299 1062
tri 5299 1059 5302 1062 nw
rect 2305 1004 2311 1015
rect 2345 1004 2357 1015
rect 2305 998 2357 1004
rect 6539 1001 6547 1015
rect 6581 1001 6591 1015
rect 6539 996 6591 1001
tri 3127 952 3130 955 se
rect 3130 952 3136 955
rect 2305 929 2311 946
rect 2345 929 2357 946
rect 2389 946 3136 952
rect 2389 912 2401 946
rect 2435 912 2475 946
rect 2509 912 2549 946
rect 2583 912 2623 946
rect 2657 912 2697 946
rect 2731 912 2771 946
rect 2805 912 2845 946
rect 2879 912 2919 946
rect 2953 912 2993 946
rect 3027 912 3067 946
rect 3101 912 3136 946
rect 2389 906 3136 912
tri 3127 903 3130 906 ne
rect 3130 903 3136 906
rect 3188 903 3203 955
rect 3255 903 3269 955
rect 3321 946 3335 955
rect 3387 946 3401 955
rect 3453 952 3459 955
tri 3459 952 3462 955 sw
tri 5816 952 5819 955 se
rect 5819 952 5870 955
rect 3453 946 4359 952
rect 3323 912 3335 946
rect 3397 912 3401 946
rect 3471 912 3510 946
rect 3544 912 3583 946
rect 3617 912 3656 946
rect 3690 912 3729 946
rect 3763 912 3802 946
rect 3836 912 3875 946
rect 3909 912 3948 946
rect 3982 912 4021 946
rect 4055 912 4094 946
rect 4128 912 4167 946
rect 4201 912 4240 946
rect 4274 912 4313 946
rect 4347 912 4359 946
rect 3321 903 3335 912
rect 3387 903 3401 912
rect 3453 906 4359 912
rect 4533 946 5870 952
rect 4533 912 4545 946
rect 4579 912 4618 946
rect 4652 912 4691 946
rect 4725 912 4764 946
rect 4798 912 4837 946
rect 4871 912 4910 946
rect 4944 912 4983 946
rect 5017 912 5056 946
rect 5090 912 5129 946
rect 5163 912 5202 946
rect 5236 912 5275 946
rect 5309 912 5348 946
rect 5382 912 5421 946
rect 5455 912 5495 946
rect 5529 912 5569 946
rect 5603 912 5643 946
rect 5677 912 5717 946
rect 5751 912 5791 946
rect 5825 912 5865 946
rect 4533 906 5870 912
rect 3453 903 3459 906
tri 3459 903 3462 906 nw
tri 5816 903 5819 906 ne
rect 5819 903 5870 906
rect 5922 903 5935 955
rect 5987 903 5999 955
rect 6051 903 6063 955
rect 6115 946 6127 955
rect 6179 946 6191 955
rect 6243 946 6255 955
rect 6307 946 6319 955
rect 6121 912 6127 946
rect 6307 912 6309 946
rect 6115 903 6127 912
rect 6179 903 6191 912
rect 6243 903 6255 912
rect 6307 903 6319 912
rect 6371 903 6383 955
rect 6435 903 6447 955
rect 6499 903 6505 955
rect 6539 925 6547 944
rect 6581 925 6591 944
rect 2305 874 2357 877
rect 2305 860 2311 874
rect 2345 860 2357 874
rect 2305 792 2357 808
rect 6539 868 6591 873
rect 6539 854 6547 868
rect 6581 854 6591 868
tri 3590 796 3593 799 se
rect 3593 796 3599 799
rect 2305 791 2311 792
rect 2345 791 2357 792
rect 2389 790 3599 796
rect 3651 790 3670 799
rect 3722 790 3741 799
rect 3793 790 3811 799
rect 3863 790 3881 799
rect 3933 790 3951 799
rect 2389 756 2401 790
rect 2435 756 2475 790
rect 2509 756 2549 790
rect 2583 756 2623 790
rect 2657 756 2697 790
rect 2731 756 2771 790
rect 2805 756 2845 790
rect 2879 756 2919 790
rect 2953 756 2993 790
rect 3027 756 3067 790
rect 3101 756 3141 790
rect 3175 756 3215 790
rect 3249 756 3289 790
rect 3323 756 3363 790
rect 3397 756 3437 790
rect 3471 756 3510 790
rect 3544 756 3583 790
rect 3651 756 3656 790
rect 3722 756 3729 790
rect 3793 756 3802 790
rect 3863 756 3875 790
rect 3933 756 3948 790
rect 2389 750 3599 756
tri 3590 747 3593 750 ne
rect 3593 747 3599 750
rect 3651 747 3670 756
rect 3722 747 3741 756
rect 3793 747 3811 756
rect 3863 747 3881 756
rect 3933 747 3951 756
rect 4003 747 4021 799
rect 4073 747 4091 799
rect 4143 747 4161 799
rect 4213 747 4231 799
rect 4283 747 4301 799
rect 4353 747 4359 799
rect 4533 747 4539 799
rect 4591 747 4609 799
rect 4661 747 4679 799
rect 4731 747 4749 799
rect 4801 747 4819 799
rect 4871 747 4889 799
rect 4941 790 4959 799
rect 5011 790 5029 799
rect 5081 790 5099 799
rect 5151 790 5170 799
rect 5222 790 5241 799
rect 5293 796 5299 799
tri 5299 796 5302 799 sw
rect 5293 790 6503 796
rect 4944 756 4959 790
rect 5017 756 5029 790
rect 5090 756 5099 790
rect 5163 756 5170 790
rect 5236 756 5241 790
rect 5309 756 5348 790
rect 5382 756 5421 790
rect 5455 756 5495 790
rect 5529 756 5569 790
rect 5603 756 5643 790
rect 5677 756 5717 790
rect 5751 756 5791 790
rect 5825 756 5865 790
rect 5899 756 5939 790
rect 5973 756 6013 790
rect 6047 756 6087 790
rect 6121 756 6161 790
rect 6195 756 6235 790
rect 6269 756 6309 790
rect 6343 756 6383 790
rect 6417 756 6457 790
rect 6491 756 6503 790
rect 4941 747 4959 756
rect 5011 747 5029 756
rect 5081 747 5099 756
rect 5151 747 5170 756
rect 5222 747 5241 756
rect 5293 750 6503 756
rect 6539 784 6591 802
rect 6539 783 6547 784
rect 6581 783 6591 784
rect 5293 747 5299 750
tri 5299 747 5302 750 nw
rect 2305 722 2357 739
rect 2305 664 2357 670
rect 6539 712 6591 731
rect 6539 654 6591 660
rect 6621 1200 6627 1276
rect 6733 1200 6840 1276
rect 6621 1161 6840 1200
rect 6621 1127 6627 1161
rect 6661 1127 6699 1161
rect 6733 1127 6840 1161
rect 6621 1088 6840 1127
rect 6621 1054 6627 1088
rect 6661 1054 6699 1088
rect 6733 1054 6840 1088
rect 6621 1015 6840 1054
rect 6621 981 6627 1015
rect 6661 981 6699 1015
rect 6733 981 6840 1015
rect 6621 942 6840 981
rect 6621 908 6627 942
rect 6661 908 6699 942
rect 6733 908 6840 942
rect 6621 869 6840 908
rect 6621 835 6627 869
rect 6661 835 6699 869
rect 6733 835 6840 869
rect 6621 796 6840 835
rect 6621 762 6627 796
rect 6661 762 6699 796
rect 6733 762 6840 796
rect 6621 723 6840 762
rect 6621 689 6627 723
rect 6661 689 6699 723
rect 6733 689 6840 723
rect 2153 614 2159 648
rect 2193 614 2231 648
rect 2265 614 2271 648
rect 6621 650 6840 689
tri 3127 640 3130 643 se
rect 3130 640 3136 643
rect 2389 634 3136 640
rect 2153 600 2271 614
tri 2271 600 2303 632 sw
rect 2389 600 2401 634
rect 2435 600 2475 634
rect 2509 600 2549 634
rect 2583 600 2623 634
rect 2657 600 2697 634
rect 2731 600 2771 634
rect 2805 600 2845 634
rect 2879 600 2919 634
rect 2953 600 2993 634
rect 3027 600 3067 634
rect 3101 600 3136 634
rect 2153 594 2303 600
tri 2303 594 2309 600 sw
rect 2389 594 3136 600
rect 2153 579 2309 594
tri 2309 579 2324 594 sw
tri 3127 591 3130 594 ne
rect 3130 591 3136 594
rect 3188 591 3203 643
rect 3255 591 3269 643
rect 3321 634 3335 643
rect 3387 634 3401 643
rect 3453 640 3459 643
tri 3459 640 3462 643 sw
tri 5816 640 5819 643 se
rect 5819 640 5870 643
rect 3453 634 4359 640
rect 3323 600 3335 634
rect 3397 600 3401 634
rect 3471 600 3510 634
rect 3544 600 3583 634
rect 3617 600 3656 634
rect 3690 600 3729 634
rect 3763 600 3802 634
rect 3836 600 3875 634
rect 3909 600 3948 634
rect 3982 600 4021 634
rect 4055 600 4094 634
rect 4128 600 4167 634
rect 4201 600 4240 634
rect 4274 600 4313 634
rect 4347 600 4359 634
rect 3321 591 3335 600
rect 3387 591 3401 600
rect 3453 594 4359 600
rect 4533 634 5870 640
rect 4533 600 4545 634
rect 4579 600 4618 634
rect 4652 600 4691 634
rect 4725 600 4764 634
rect 4798 600 4837 634
rect 4871 600 4910 634
rect 4944 600 4983 634
rect 5017 600 5056 634
rect 5090 600 5129 634
rect 5163 600 5202 634
rect 5236 600 5275 634
rect 5309 600 5348 634
rect 5382 600 5421 634
rect 5455 600 5495 634
rect 5529 600 5569 634
rect 5603 600 5643 634
rect 5677 600 5717 634
rect 5751 600 5791 634
rect 5825 600 5865 634
rect 4533 594 5870 600
rect 3453 591 3459 594
tri 3459 591 3462 594 nw
tri 5816 591 5819 594 ne
rect 5819 591 5870 594
rect 5922 591 5935 643
rect 5987 591 5999 643
rect 6051 591 6063 643
rect 6115 634 6127 643
rect 6179 634 6191 643
rect 6243 634 6255 643
rect 6307 634 6319 643
rect 6121 600 6127 634
rect 6307 600 6309 634
rect 6115 591 6127 600
rect 6179 591 6191 600
rect 6243 591 6255 600
rect 6307 591 6319 600
rect 6371 591 6383 643
rect 6435 591 6447 643
rect 6499 591 6505 643
tri 6605 616 6621 632 se
rect 6621 616 6627 650
rect 6661 616 6699 650
rect 6733 616 6840 650
tri 6602 613 6605 616 se
rect 6605 613 6840 616
tri 6583 594 6602 613 se
rect 6602 594 6840 613
tri 6580 591 6583 594 se
rect 6583 591 6840 594
tri 6568 579 6580 591 se
rect 6580 579 6840 591
rect 2153 577 2324 579
tri 2324 577 2326 579 sw
tri 6566 577 6568 579 se
rect 6568 577 6840 579
rect 2153 575 2326 577
rect 2153 541 2159 575
rect 2193 541 2231 575
rect 2265 543 2326 575
tri 2326 543 2360 577 sw
tri 6532 543 6566 577 se
rect 6566 543 6627 577
rect 6661 543 6699 577
rect 6733 543 6840 577
rect 2265 541 2360 543
rect 2153 539 2360 541
tri 2360 539 2364 543 sw
tri 6528 539 6532 543 se
rect 6532 539 6840 543
rect 2153 505 2364 539
tri 2364 505 2398 539 sw
tri 6494 505 6528 539 se
rect 6528 505 6840 539
rect 2153 504 2398 505
tri 2398 504 2399 505 sw
tri 6493 504 6494 505 se
rect 6494 504 6840 505
rect 2153 502 2399 504
rect 2153 324 2159 502
rect 2265 484 2399 502
tri 2399 484 2419 504 sw
tri 6476 487 6493 504 se
rect 6493 487 6627 504
rect 6661 493 6699 504
rect 6733 493 6840 504
tri 3587 484 3590 487 se
rect 3590 484 3599 487
rect 2265 478 3599 484
rect 3651 478 3670 487
rect 3722 478 3741 487
rect 3793 478 3811 487
rect 3863 478 3881 487
rect 3933 478 3951 487
rect 2265 444 2401 478
rect 2435 444 2475 478
rect 2509 444 2549 478
rect 2583 444 2623 478
rect 2657 444 2697 478
rect 2731 444 2771 478
rect 2805 444 2845 478
rect 2879 444 2919 478
rect 2953 444 2993 478
rect 3027 444 3067 478
rect 3101 444 3141 478
rect 3175 444 3215 478
rect 3249 444 3289 478
rect 3323 444 3363 478
rect 3397 444 3437 478
rect 3471 444 3510 478
rect 3544 444 3583 478
rect 3651 444 3656 478
rect 3722 444 3729 478
rect 3793 444 3802 478
rect 3863 444 3875 478
rect 3933 444 3948 478
rect 2265 435 3599 444
rect 3651 435 3670 444
rect 3722 435 3741 444
rect 3793 435 3811 444
rect 3863 435 3881 444
rect 3933 435 3951 444
rect 4003 435 4021 487
rect 4073 435 4091 487
rect 4143 435 4161 487
rect 4213 435 4231 487
rect 4283 435 4301 487
rect 4353 435 4539 487
rect 4591 435 4609 487
rect 4661 435 4679 487
rect 4731 435 4749 487
rect 4801 435 4819 487
rect 4871 435 4889 487
rect 4941 478 4959 487
rect 5011 478 5029 487
rect 5081 478 5099 487
rect 5151 478 5170 487
rect 5222 478 5241 487
rect 5293 484 5304 487
tri 5304 484 5307 487 sw
tri 6473 484 6476 487 se
rect 6476 484 6627 487
rect 5293 478 6627 484
rect 4944 444 4959 478
rect 5017 444 5029 478
rect 5090 444 5099 478
rect 5163 444 5170 478
rect 5236 444 5241 478
rect 5309 444 5348 478
rect 5382 444 5421 478
rect 5455 444 5495 478
rect 5529 444 5569 478
rect 5603 444 5643 478
rect 5677 444 5717 478
rect 5751 444 5791 478
rect 5825 444 5865 478
rect 5899 444 5939 478
rect 5973 444 6013 478
rect 6047 444 6087 478
rect 6121 444 6161 478
rect 6195 444 6235 478
rect 6269 444 6309 478
rect 6343 444 6383 478
rect 6417 444 6457 478
rect 6491 470 6627 478
rect 6733 470 6760 493
rect 6491 444 6655 470
rect 4941 435 4959 444
rect 5011 435 5029 444
rect 5081 435 5099 444
rect 5151 435 5170 444
rect 5222 435 5241 444
rect 5293 441 6655 444
rect 6707 441 6760 470
rect 6812 441 6840 493
rect 5293 435 6840 441
rect 2265 431 6840 435
rect 2265 419 6627 431
rect 6661 429 6699 431
rect 6733 429 6840 431
rect 2265 367 3599 419
rect 3651 367 3665 419
rect 3717 367 3731 419
rect 3783 367 3797 419
rect 3849 367 3863 419
rect 3915 367 3929 419
rect 3981 367 3995 419
rect 4047 367 4061 419
rect 4113 367 4127 419
rect 4179 367 4193 419
rect 4245 367 4259 419
rect 4311 367 4325 419
rect 4377 367 4391 419
rect 4443 367 4457 419
rect 4509 367 4523 419
rect 4575 367 4589 419
rect 4641 367 4655 419
rect 4707 367 4721 419
rect 4773 367 4786 419
rect 4838 367 4851 419
rect 4903 367 4916 419
rect 4968 367 4981 419
rect 5033 367 5046 419
rect 5098 367 5111 419
rect 5163 367 5176 419
rect 5228 367 5241 419
rect 5293 397 6627 419
rect 6733 397 6760 429
rect 5293 377 6655 397
rect 6707 377 6760 397
rect 6812 377 6840 429
rect 5293 367 6840 377
rect 2265 365 6840 367
rect 2265 358 6655 365
rect 6707 358 6760 365
rect 2265 324 2304 358
rect 2338 324 2377 358
rect 2411 324 2450 358
rect 2484 324 2523 358
rect 2153 286 2523 324
rect 6733 324 6760 358
rect 6707 313 6760 324
rect 6812 313 6840 365
rect 2153 252 2231 286
rect 2265 252 2304 286
rect 2338 252 2377 286
rect 2411 252 2450 286
rect 2484 252 2523 286
rect 6661 252 6840 313
rect 2153 246 6840 252
rect 6876 1351 6994 1390
rect 6876 1317 6882 1351
rect 6916 1317 6954 1351
rect 6988 1317 6994 1351
rect 6876 1278 6994 1317
rect 6876 1244 6882 1278
rect 6916 1244 6954 1278
rect 6988 1244 6994 1278
rect 6876 1205 6994 1244
rect 6876 1171 6882 1205
rect 6916 1171 6954 1205
rect 6988 1171 6994 1205
rect 6876 1131 6994 1171
rect 6876 1097 6882 1131
rect 6916 1097 6954 1131
rect 6988 1097 6994 1131
rect 6876 1057 6994 1097
rect 6876 1023 6882 1057
rect 6916 1023 6954 1057
rect 6988 1023 6994 1057
rect 6876 983 6994 1023
rect 6876 949 6882 983
rect 6916 949 6954 983
rect 6988 949 6994 983
rect 6876 942 6994 949
rect 6876 909 6909 942
rect 6961 909 6994 942
rect 6876 875 6882 909
rect 6916 876 6954 890
rect 6988 875 6994 909
rect 6876 835 6909 875
rect 6961 835 6994 875
rect 6876 801 6882 835
rect 6916 810 6954 824
rect 6988 801 6994 835
rect 6876 761 6909 801
rect 6961 761 6994 801
rect 6876 727 6882 761
rect 6916 744 6954 758
rect 6988 727 6994 761
rect 6876 692 6909 727
rect 6961 692 6994 727
rect 6876 687 6994 692
rect 6876 653 6882 687
rect 6916 677 6954 687
rect 6988 653 6994 687
rect 6876 625 6909 653
rect 6961 625 6994 653
rect 6876 613 6994 625
rect 6876 579 6882 613
rect 6916 579 6954 613
rect 6988 579 6994 613
rect 6876 539 6994 579
rect 6876 505 6882 539
rect 6916 505 6954 539
rect 6988 505 6994 539
rect 6876 465 6994 505
rect 6876 431 6882 465
rect 6916 431 6954 465
rect 6988 431 6994 465
rect 6876 391 6994 431
rect 6876 357 6882 391
rect 6916 357 6954 391
rect 6988 357 6994 391
rect 6876 317 6994 357
rect 6876 283 6882 317
rect 6916 283 6954 317
rect 6988 283 6994 317
rect 55 209 173 210
tri 173 209 188 224 sw
tri 1883 209 1898 224 se
rect 1898 209 1904 243
rect 1938 209 1976 243
rect 2010 209 2016 243
rect 6876 243 6994 283
rect 55 177 188 209
tri 188 177 220 209 sw
tri 1851 177 1883 209 se
rect 1883 177 2016 209
tri 2016 177 2063 224 sw
tri 6842 177 6876 211 se
rect 6876 177 6882 243
rect 55 171 6882 177
rect 6988 177 6994 243
rect 7157 1440 8741 1446
rect 8793 1440 8808 1454
rect 8860 1440 8874 1454
rect 8926 1440 8940 1454
rect 8992 1440 9006 1454
rect 9058 1440 9072 1454
rect 9124 1440 9138 1454
rect 9190 1440 9204 1454
rect 9256 1440 9270 1454
rect 9322 1440 9336 1454
rect 9388 1440 9402 1454
rect 9454 1440 9468 1454
rect 9520 1440 9534 1454
rect 9586 1440 9600 1454
rect 9652 1440 9666 1454
rect 9718 1440 9732 1454
rect 9784 1440 9798 1454
rect 9850 1440 9864 1454
rect 9916 1440 9930 1454
rect 9982 1440 9996 1454
rect 10048 1440 10062 1454
rect 10114 1440 10128 1454
rect 10180 1440 10194 1454
rect 10246 1440 10260 1454
rect 10312 1446 10318 1454
rect 10312 1440 11757 1446
rect 7157 1406 7241 1440
rect 7275 1406 7319 1440
rect 7353 1406 7397 1440
rect 7431 1406 7475 1440
rect 7509 1406 7553 1440
rect 7587 1406 7631 1440
rect 7665 1406 7709 1440
rect 7743 1406 7788 1440
rect 7822 1406 7898 1440
rect 7157 1368 7898 1406
rect 11460 1406 11499 1440
rect 11533 1406 11572 1440
rect 11606 1406 11645 1440
rect 11679 1406 11757 1440
rect 7157 1334 7163 1368
rect 7197 1334 7235 1368
rect 7269 1334 7319 1368
rect 7353 1334 7397 1368
rect 7431 1334 7475 1368
rect 7509 1334 7553 1368
rect 7587 1334 7631 1368
rect 7665 1334 7709 1368
rect 7743 1334 7788 1368
rect 7822 1334 7898 1368
rect 11460 1368 11757 1406
rect 11460 1334 11499 1368
rect 11533 1334 11572 1368
rect 11606 1334 11645 1368
rect 7157 1328 11645 1334
rect 7157 1295 7275 1328
rect 7157 1261 7163 1295
rect 7197 1261 7235 1295
rect 7269 1261 7275 1295
tri 7275 1294 7309 1328 nw
tri 11605 1294 11639 1328 ne
tri 7415 1264 7418 1267 se
rect 7418 1264 8030 1267
rect 7157 1222 7275 1261
rect 7157 324 7163 1222
rect 7269 397 7275 1222
rect 7408 1258 8030 1264
rect 8082 1258 8095 1267
rect 7408 1224 7420 1258
rect 7454 1224 7494 1258
rect 7528 1224 7568 1258
rect 7602 1224 7642 1258
rect 7676 1224 7716 1258
rect 7750 1224 7790 1258
rect 7824 1224 7864 1258
rect 7898 1224 7938 1258
rect 7972 1224 8012 1258
rect 8082 1224 8086 1258
rect 7408 1218 8030 1224
tri 7415 1215 7418 1218 ne
rect 7418 1215 8030 1218
rect 8082 1215 8095 1224
rect 8147 1215 8159 1267
rect 8211 1215 8223 1267
rect 8275 1215 8287 1267
rect 8339 1258 8351 1267
rect 8403 1258 8415 1267
rect 8467 1258 8479 1267
rect 8531 1258 8543 1267
rect 8595 1258 8607 1267
rect 8659 1264 8665 1267
tri 10449 1264 10452 1267 se
rect 10452 1264 10458 1267
rect 8659 1258 9378 1264
rect 8342 1224 8351 1258
rect 8595 1224 8602 1258
rect 8659 1224 8675 1258
rect 8709 1224 8748 1258
rect 8782 1224 8821 1258
rect 8855 1224 8894 1258
rect 8928 1224 8967 1258
rect 9001 1224 9040 1258
rect 9074 1224 9113 1258
rect 9147 1224 9186 1258
rect 9220 1224 9259 1258
rect 9293 1224 9332 1258
rect 9366 1224 9378 1258
rect 8339 1215 8351 1224
rect 8403 1215 8415 1224
rect 8467 1215 8479 1224
rect 8531 1215 8543 1224
rect 8595 1215 8607 1224
rect 8659 1218 9378 1224
rect 9552 1258 10458 1264
rect 10510 1258 10525 1267
rect 10577 1258 10591 1267
rect 9552 1224 9564 1258
rect 9598 1224 9637 1258
rect 9671 1224 9710 1258
rect 9744 1224 9783 1258
rect 9817 1224 9856 1258
rect 9890 1224 9929 1258
rect 9963 1224 10002 1258
rect 10036 1224 10075 1258
rect 10109 1224 10148 1258
rect 10182 1224 10221 1258
rect 10255 1224 10294 1258
rect 10328 1224 10367 1258
rect 10401 1224 10440 1258
rect 10510 1224 10514 1258
rect 10577 1224 10588 1258
rect 9552 1218 10458 1224
rect 8659 1215 8665 1218
tri 10449 1215 10452 1218 ne
rect 10452 1215 10458 1218
rect 10510 1215 10525 1224
rect 10577 1215 10591 1224
rect 10643 1215 10657 1267
rect 10709 1215 10723 1267
rect 10775 1264 10781 1267
tri 10781 1264 10784 1267 sw
rect 10775 1258 11522 1264
rect 10775 1224 10810 1258
rect 10844 1224 10884 1258
rect 10918 1224 10958 1258
rect 10992 1224 11032 1258
rect 11066 1224 11106 1258
rect 11140 1224 11180 1258
rect 11214 1224 11254 1258
rect 11288 1224 11328 1258
rect 11362 1224 11402 1258
rect 11436 1224 11476 1258
rect 11510 1224 11522 1258
rect 10775 1218 11522 1224
rect 10775 1215 10781 1218
tri 10781 1215 10784 1218 nw
rect 7322 1207 7374 1213
rect 7322 1141 7374 1155
rect 11558 1207 11610 1213
rect 11558 1141 11610 1155
tri 8732 1108 8735 1111 se
rect 8735 1108 8741 1111
rect 7322 1075 7374 1089
rect 7408 1102 8741 1108
rect 7408 1068 7420 1102
rect 7454 1068 7494 1102
rect 7528 1068 7568 1102
rect 7602 1068 7642 1102
rect 7676 1068 7716 1102
rect 7750 1068 7790 1102
rect 7824 1068 7864 1102
rect 7898 1068 7938 1102
rect 7972 1068 8012 1102
rect 8046 1068 8086 1102
rect 8120 1068 8160 1102
rect 8194 1068 8234 1102
rect 8268 1068 8308 1102
rect 8342 1068 8382 1102
rect 8416 1068 8456 1102
rect 8490 1068 8529 1102
rect 8563 1068 8602 1102
rect 8636 1068 8675 1102
rect 8709 1068 8741 1102
rect 7408 1062 8741 1068
tri 8732 1059 8735 1062 ne
rect 8735 1059 8741 1062
rect 8793 1059 8806 1111
rect 8858 1059 8871 1111
rect 8923 1102 8936 1111
rect 8988 1102 9000 1111
rect 9052 1102 9064 1111
rect 9116 1102 9128 1111
rect 9180 1102 9192 1111
rect 8928 1068 8936 1102
rect 9180 1068 9186 1102
rect 8923 1059 8936 1068
rect 8988 1059 9000 1068
rect 9052 1059 9064 1068
rect 9116 1059 9128 1068
rect 9180 1059 9192 1068
rect 9244 1059 9256 1111
rect 9308 1059 9320 1111
rect 9372 1059 9378 1111
rect 9552 1059 9558 1111
rect 9610 1059 9628 1111
rect 9680 1059 9698 1111
rect 9750 1059 9768 1111
rect 9820 1059 9838 1111
rect 9890 1059 9908 1111
rect 9960 1102 9978 1111
rect 10030 1102 10048 1111
rect 10100 1102 10118 1111
rect 10170 1102 10189 1111
rect 10241 1102 10260 1111
rect 10312 1108 10318 1111
tri 10318 1108 10321 1111 sw
rect 10312 1102 11522 1108
rect 9963 1068 9978 1102
rect 10036 1068 10048 1102
rect 10109 1068 10118 1102
rect 10182 1068 10189 1102
rect 10255 1068 10260 1102
rect 10328 1068 10367 1102
rect 10401 1068 10440 1102
rect 10474 1068 10514 1102
rect 10548 1068 10588 1102
rect 10622 1068 10662 1102
rect 10696 1068 10736 1102
rect 10770 1068 10810 1102
rect 10844 1068 10884 1102
rect 10918 1068 10958 1102
rect 10992 1068 11032 1102
rect 11066 1068 11106 1102
rect 11140 1068 11180 1102
rect 11214 1068 11254 1102
rect 11288 1068 11328 1102
rect 11362 1068 11402 1102
rect 11436 1068 11476 1102
rect 11510 1068 11522 1102
rect 9960 1059 9978 1068
rect 10030 1059 10048 1068
rect 10100 1059 10118 1068
rect 10170 1059 10189 1068
rect 10241 1059 10260 1068
rect 10312 1062 11522 1068
rect 11558 1075 11610 1089
rect 10312 1059 10318 1062
tri 10318 1059 10321 1062 nw
rect 7322 1019 7330 1023
rect 7364 1019 7374 1023
rect 7322 1009 7374 1019
rect 7322 945 7330 957
rect 7364 945 7374 957
rect 11558 1019 11566 1023
rect 11600 1019 11610 1023
rect 11558 1009 11610 1019
tri 7415 952 7418 955 se
rect 7418 952 8027 955
rect 7322 943 7374 945
rect 7408 946 8027 952
rect 8079 946 8092 955
rect 7408 912 7420 946
rect 7454 912 7494 946
rect 7528 912 7568 946
rect 7602 912 7642 946
rect 7676 912 7716 946
rect 7750 912 7790 946
rect 7824 912 7864 946
rect 7898 912 7938 946
rect 7972 912 8012 946
rect 8079 912 8086 946
rect 7408 906 8027 912
tri 7415 905 7416 906 ne
rect 7416 905 8027 906
tri 7416 903 7418 905 ne
rect 7418 903 8027 905
rect 8079 903 8092 912
rect 8144 903 8156 955
rect 8208 903 8220 955
rect 8272 903 8284 955
rect 8336 946 8348 955
rect 8400 946 8412 955
rect 8464 946 8476 955
rect 8528 946 8540 955
rect 8592 946 8604 955
rect 8656 952 8662 955
tri 10449 952 10452 955 se
rect 10452 952 10458 955
rect 8656 946 9378 952
rect 8342 912 8348 946
rect 8528 912 8529 946
rect 8592 912 8602 946
rect 8656 912 8675 946
rect 8709 912 8748 946
rect 8782 912 8821 946
rect 8855 912 8894 946
rect 8928 912 8967 946
rect 9001 912 9040 946
rect 9074 912 9113 946
rect 9147 912 9186 946
rect 9220 912 9259 946
rect 9293 912 9332 946
rect 9366 912 9378 946
rect 8336 903 8348 912
rect 8400 903 8412 912
rect 8464 903 8476 912
rect 8528 903 8540 912
rect 8592 903 8604 912
rect 8656 906 9378 912
rect 9552 946 10458 952
rect 10510 946 10525 955
rect 10577 946 10591 955
rect 9552 912 9564 946
rect 9598 912 9637 946
rect 9671 912 9710 946
rect 9744 912 9783 946
rect 9817 912 9856 946
rect 9890 912 9929 946
rect 9963 912 10002 946
rect 10036 912 10075 946
rect 10109 912 10148 946
rect 10182 912 10221 946
rect 10255 912 10294 946
rect 10328 912 10367 946
rect 10401 912 10440 946
rect 10510 912 10514 946
rect 10577 912 10588 946
rect 9552 906 10458 912
rect 8656 903 8662 906
tri 10449 905 10450 906 ne
rect 10450 905 10458 906
tri 10450 903 10452 905 ne
rect 10452 903 10458 905
rect 10510 903 10525 912
rect 10577 903 10591 912
rect 10643 903 10657 955
rect 10709 903 10723 955
rect 10775 952 10781 955
tri 10781 952 10784 955 sw
rect 10775 946 11522 952
rect 10775 912 10810 946
rect 10844 912 10884 946
rect 10918 912 10958 946
rect 10992 912 11032 946
rect 11066 912 11106 946
rect 11140 912 11180 946
rect 11214 912 11254 946
rect 11288 912 11328 946
rect 11362 912 11402 946
rect 11436 912 11476 946
rect 11510 912 11522 946
rect 10775 906 11522 912
rect 11558 945 11566 957
rect 11600 945 11610 957
rect 11558 943 11610 945
rect 10775 905 10783 906
tri 10783 905 10784 906 nw
rect 10775 903 10781 905
tri 10781 903 10783 905 nw
rect 7322 877 7330 891
rect 7364 877 7374 891
rect 7322 811 7330 825
rect 7364 811 7374 825
rect 11558 877 11566 891
rect 11600 877 11610 891
rect 11558 811 11566 825
rect 11600 811 11610 825
tri 8733 797 8735 799 se
rect 8735 797 8741 799
tri 8732 796 8733 797 se
rect 8733 796 8741 797
rect 7322 757 7374 759
rect 7322 745 7330 757
rect 7364 745 7374 757
rect 7408 790 8741 796
rect 7408 756 7420 790
rect 7454 756 7494 790
rect 7528 756 7568 790
rect 7602 756 7642 790
rect 7676 756 7716 790
rect 7750 756 7790 790
rect 7824 756 7864 790
rect 7898 756 7938 790
rect 7972 756 8012 790
rect 8046 756 8086 790
rect 8120 756 8160 790
rect 8194 756 8234 790
rect 8268 756 8308 790
rect 8342 756 8382 790
rect 8416 756 8456 790
rect 8490 756 8529 790
rect 8563 756 8602 790
rect 8636 756 8675 790
rect 8709 756 8741 790
rect 7408 750 8741 756
tri 8732 747 8735 750 ne
rect 8735 747 8741 750
rect 8793 747 8806 799
rect 8858 747 8871 799
rect 8923 790 8936 799
rect 8988 790 9000 799
rect 9052 790 9064 799
rect 9116 790 9128 799
rect 9180 790 9192 799
rect 8928 756 8936 790
rect 9180 756 9186 790
rect 8923 747 8936 756
rect 8988 747 9000 756
rect 9052 747 9064 756
rect 9116 747 9128 756
rect 9180 747 9192 756
rect 9244 747 9256 799
rect 9308 747 9320 799
rect 9372 747 9378 799
rect 9552 747 9558 799
rect 9610 747 9628 799
rect 9680 747 9698 799
rect 9750 747 9768 799
rect 9820 747 9838 799
rect 9890 747 9908 799
rect 9960 790 9978 799
rect 10030 790 10048 799
rect 10100 790 10118 799
rect 10170 790 10189 799
rect 10241 790 10260 799
rect 10312 797 10318 799
tri 10318 797 10320 799 sw
rect 10312 796 10320 797
tri 10320 796 10321 797 sw
rect 10312 790 11522 796
rect 9963 756 9978 790
rect 10036 756 10048 790
rect 10109 756 10118 790
rect 10182 756 10189 790
rect 10255 756 10260 790
rect 10328 756 10367 790
rect 10401 756 10440 790
rect 10474 756 10514 790
rect 10548 756 10588 790
rect 10622 756 10662 790
rect 10696 756 10736 790
rect 10770 756 10810 790
rect 10844 756 10884 790
rect 10918 756 10958 790
rect 10992 756 11032 790
rect 11066 756 11106 790
rect 11140 756 11180 790
rect 11214 756 11254 790
rect 11288 756 11328 790
rect 11362 756 11402 790
rect 11436 756 11476 790
rect 11510 756 11522 790
rect 9960 747 9978 756
rect 10030 747 10048 756
rect 10100 747 10118 756
rect 10170 747 10189 756
rect 10241 747 10260 756
rect 10312 750 11522 756
rect 11558 757 11610 759
rect 10312 747 10318 750
tri 10318 747 10321 750 nw
rect 7322 683 7374 693
rect 7322 679 7330 683
rect 7364 679 7374 683
rect 11558 745 11566 757
rect 11600 745 11610 757
rect 11558 683 11610 693
rect 11558 679 11566 683
rect 11600 679 11610 683
tri 7415 640 7418 643 se
rect 7418 640 8027 643
rect 7322 613 7374 627
rect 7408 634 8027 640
rect 8079 634 8092 643
rect 7408 600 7420 634
rect 7454 600 7494 634
rect 7528 600 7568 634
rect 7602 600 7642 634
rect 7676 600 7716 634
rect 7750 600 7790 634
rect 7824 600 7864 634
rect 7898 600 7938 634
rect 7972 600 8012 634
rect 8079 600 8086 634
rect 7408 594 8027 600
tri 7415 591 7418 594 ne
rect 7418 591 8027 594
rect 8079 591 8092 600
rect 8144 591 8156 643
rect 8208 591 8220 643
rect 8272 591 8284 643
rect 8336 634 8348 643
rect 8400 634 8412 643
rect 8464 634 8476 643
rect 8528 634 8540 643
rect 8592 634 8604 643
rect 8656 640 8662 643
tri 10449 640 10452 643 se
rect 10452 640 10458 643
rect 8656 634 9378 640
rect 8342 600 8348 634
rect 8528 600 8529 634
rect 8592 600 8602 634
rect 8656 600 8675 634
rect 8709 600 8748 634
rect 8782 600 8821 634
rect 8855 600 8894 634
rect 8928 600 8967 634
rect 9001 600 9040 634
rect 9074 600 9113 634
rect 9147 600 9186 634
rect 9220 600 9259 634
rect 9293 600 9332 634
rect 9366 600 9378 634
rect 8336 591 8348 600
rect 8400 591 8412 600
rect 8464 591 8476 600
rect 8528 591 8540 600
rect 8592 591 8604 600
rect 8656 594 9378 600
rect 9552 634 10458 640
rect 10510 634 10525 643
rect 10577 634 10591 643
rect 9552 600 9564 634
rect 9598 600 9637 634
rect 9671 600 9710 634
rect 9744 600 9783 634
rect 9817 600 9856 634
rect 9890 600 9929 634
rect 9963 600 10002 634
rect 10036 600 10075 634
rect 10109 600 10148 634
rect 10182 600 10221 634
rect 10255 600 10294 634
rect 10328 600 10367 634
rect 10401 600 10440 634
rect 10510 600 10514 634
rect 10577 600 10588 634
rect 9552 594 10458 600
rect 8656 591 8662 594
tri 10449 591 10452 594 ne
rect 10452 591 10458 594
rect 10510 591 10525 600
rect 10577 591 10591 600
rect 10643 591 10657 643
rect 10709 591 10723 643
rect 10775 640 10781 643
tri 10781 640 10784 643 sw
rect 10775 634 11522 640
rect 10775 600 10810 634
rect 10844 600 10884 634
rect 10918 600 10958 634
rect 10992 600 11032 634
rect 11066 600 11106 634
rect 11140 600 11180 634
rect 11214 600 11254 634
rect 11288 600 11328 634
rect 11362 600 11402 634
rect 11436 600 11476 634
rect 11510 600 11522 634
rect 10775 594 11522 600
rect 11558 613 11610 627
rect 10775 591 10781 594
tri 10781 591 10784 594 nw
rect 7322 547 7374 561
rect 7322 489 7374 495
rect 11558 547 11610 561
rect 11558 489 11610 495
tri 8732 484 8735 487 se
rect 8735 484 8741 487
rect 7408 478 8741 484
rect 7408 444 7420 478
rect 7454 444 7494 478
rect 7528 444 7568 478
rect 7602 444 7642 478
rect 7676 444 7716 478
rect 7750 444 7790 478
rect 7824 444 7864 478
rect 7898 444 7938 478
rect 7972 444 8012 478
rect 8046 444 8086 478
rect 8120 444 8160 478
rect 8194 444 8234 478
rect 8268 444 8308 478
rect 8342 444 8382 478
rect 8416 444 8456 478
rect 8490 444 8529 478
rect 8563 444 8602 478
rect 8636 444 8675 478
rect 8709 444 8741 478
rect 7408 438 8741 444
tri 8732 435 8735 438 ne
rect 8735 435 8741 438
rect 8793 435 8806 487
rect 8858 435 8871 487
rect 8923 478 8936 487
rect 8988 478 9000 487
rect 9052 478 9064 487
rect 9116 478 9128 487
rect 9180 478 9192 487
rect 8928 444 8936 478
rect 9180 444 9186 478
rect 8923 435 8936 444
rect 8988 435 9000 444
rect 9052 435 9064 444
rect 9116 435 9128 444
rect 9180 435 9192 444
rect 9244 435 9256 487
rect 9308 435 9320 487
rect 9372 435 9378 487
rect 9552 435 9558 487
rect 9610 435 9628 487
rect 9680 435 9698 487
rect 9750 435 9768 487
rect 9820 435 9838 487
rect 9890 435 9908 487
rect 9960 478 9978 487
rect 10030 478 10048 487
rect 10100 478 10118 487
rect 10170 478 10189 487
rect 10241 478 10260 487
rect 10312 484 10318 487
tri 10318 484 10321 487 sw
rect 10312 478 11522 484
rect 9963 444 9978 478
rect 10036 444 10048 478
rect 10109 444 10118 478
rect 10182 444 10189 478
rect 10255 444 10260 478
rect 10328 444 10367 478
rect 10401 444 10440 478
rect 10474 444 10514 478
rect 10548 444 10588 478
rect 10622 444 10662 478
rect 10696 444 10736 478
rect 10770 444 10810 478
rect 10844 444 10884 478
rect 10918 444 10958 478
rect 10992 444 11032 478
rect 11066 444 11106 478
rect 11140 444 11180 478
rect 11214 444 11254 478
rect 11288 444 11328 478
rect 11362 444 11402 478
rect 11436 444 11476 478
rect 11510 444 11522 478
rect 9960 435 9978 444
rect 10030 435 10048 444
rect 10100 435 10118 444
rect 10170 435 10189 444
rect 10241 435 10260 444
rect 10312 438 11522 444
rect 11639 470 11645 1328
rect 11751 470 11757 1368
rect 10312 435 10318 438
tri 10318 435 10321 438 nw
rect 11639 431 11757 470
tri 7275 397 7276 398 sw
tri 11638 397 11639 398 se
rect 11639 397 11645 431
rect 11679 397 11717 431
rect 11751 397 11757 431
rect 7269 383 7276 397
tri 7276 383 7290 397 sw
tri 11624 383 11638 397 se
rect 11638 383 11757 397
rect 7269 364 7290 383
tri 7290 364 7309 383 sw
tri 8716 364 8735 383 se
rect 8735 364 8741 383
rect 7269 358 8741 364
rect 8793 358 8808 383
rect 8860 358 8874 383
rect 8926 358 8940 383
rect 8992 358 9006 383
rect 9058 358 9072 383
rect 9124 358 9138 383
rect 9190 358 9204 383
rect 9256 358 9270 383
rect 9322 358 9336 383
rect 9388 358 9402 383
rect 9454 358 9468 383
rect 9520 358 9534 383
rect 9586 358 9600 383
rect 9652 358 9666 383
rect 9718 358 9732 383
rect 9784 358 9798 383
rect 9850 358 9864 383
rect 9916 358 9930 383
rect 9982 358 9996 383
rect 10048 358 10062 383
rect 10114 358 10128 383
rect 10180 358 10194 383
rect 10246 358 10260 383
rect 10312 364 10318 383
tri 10318 364 10337 383 sw
tri 11605 364 11624 383 se
rect 11624 364 11757 383
rect 10312 358 11757 364
rect 7269 324 7308 358
rect 7342 324 7381 358
rect 7415 324 7454 358
rect 7488 324 7527 358
rect 7561 324 7600 358
rect 7634 324 7673 358
rect 7707 324 7746 358
rect 7780 324 7819 358
rect 7853 324 7892 358
rect 7926 324 7965 358
rect 7999 324 8038 358
rect 8072 324 8111 358
rect 8145 324 8184 358
rect 8218 324 8257 358
rect 8291 324 8330 358
rect 8364 324 8403 358
rect 8437 324 8476 358
rect 8510 324 8549 358
rect 7157 286 8549 324
rect 11679 324 11717 358
rect 11751 324 11757 358
rect 7157 266 7235 286
rect 7269 266 7308 286
rect 7342 266 7381 286
rect 7415 266 7454 286
rect 7488 266 7527 286
rect 7561 266 7600 286
rect 7634 266 7673 286
rect 7707 266 7746 286
rect 7780 266 7819 286
rect 7853 266 7892 286
rect 7926 266 7965 286
rect 7999 266 8038 286
rect 8072 266 8111 286
rect 7157 214 7163 266
rect 7215 214 7229 266
rect 7281 214 7295 266
rect 7347 214 7361 266
rect 7415 252 7426 266
rect 7488 252 7491 266
rect 7738 252 7746 266
rect 7413 214 7426 252
rect 7478 214 7491 252
rect 7543 214 7556 252
rect 7608 214 7621 252
rect 7673 214 7686 252
rect 7738 214 7751 252
rect 7803 214 7816 266
rect 7868 214 7881 266
rect 7933 214 7946 266
rect 7999 252 8011 266
rect 8072 252 8076 266
rect 8145 252 8184 286
rect 8218 252 8257 286
rect 8291 252 8330 286
rect 8364 252 8403 286
rect 8437 252 8476 286
rect 8510 252 8549 286
rect 11679 252 11757 324
rect 7998 214 8011 252
rect 8063 214 8076 252
rect 8128 246 11757 252
rect 8128 224 8144 246
tri 8144 224 8166 246 nw
rect 8128 214 8134 224
tri 8134 214 8144 224 nw
tri 6994 177 7028 211 sw
tri 11860 177 11894 211 se
rect 6988 175 11894 177
rect 6988 171 10880 175
rect 10932 171 10946 175
rect 10998 171 11012 175
rect 11064 171 11078 175
rect 11130 171 11894 175
rect 55 137 61 171
rect 95 137 133 171
rect 167 137 206 171
rect 240 137 279 171
rect 313 137 352 171
rect 386 137 425 171
rect 459 137 498 171
rect 532 137 571 171
rect 605 137 644 171
rect 678 137 717 171
rect 751 137 790 171
rect 824 137 863 171
rect 897 137 936 171
rect 970 137 1009 171
rect 1043 137 1082 171
rect 1116 137 1155 171
rect 1189 137 1228 171
rect 1262 137 1301 171
rect 1335 137 1374 171
rect 1408 137 1447 171
rect 1481 137 1520 171
rect 1554 137 1593 171
rect 1627 137 1666 171
rect 1700 137 1739 171
rect 1773 137 1812 171
rect 1846 137 1885 171
rect 1919 137 1958 171
rect 1992 137 2031 171
rect 2065 137 2104 171
rect 2138 137 2177 171
rect 2211 137 2250 171
rect 2284 137 2323 171
rect 55 99 2323 137
rect 55 65 133 99
rect 167 65 206 99
rect 240 65 279 99
rect 313 65 352 99
rect 386 65 425 99
rect 459 65 498 99
rect 532 65 571 99
rect 605 65 644 99
rect 678 65 717 99
rect 751 65 790 99
rect 824 65 863 99
rect 897 65 936 99
rect 970 65 1009 99
rect 1043 65 1082 99
rect 1116 65 1155 99
rect 1189 65 1228 99
rect 1262 65 1301 99
rect 1335 65 1374 99
rect 1408 65 1447 99
rect 1481 65 1520 99
rect 1554 65 1593 99
rect 1627 65 1666 99
rect 1700 65 1739 99
rect 1773 65 1812 99
rect 1846 65 1885 99
rect 1919 65 1958 99
rect 1992 65 2031 99
rect 2065 65 2104 99
rect 2138 65 2177 99
rect 2211 65 2250 99
rect 2284 65 2323 99
rect 11861 65 11894 171
rect 55 59 11894 65
rect -508 -183 37 -177
rect -508 -217 -496 -183
rect -462 -217 -409 -183
rect -375 -217 -322 -183
rect -288 -217 -236 -183
rect -202 -217 -150 -183
rect -116 -184 37 -183
rect -116 -217 -79 -184
rect -508 -236 -79 -217
rect -27 -236 -15 -184
rect -508 -252 37 -236
rect -508 -293 -79 -252
rect -508 -327 -496 -293
rect -462 -327 -409 -293
rect -375 -327 -322 -293
rect -288 -327 -236 -293
rect -202 -327 -150 -293
rect -116 -304 -79 -293
rect -27 -304 -15 -252
rect -116 -327 37 -304
rect -508 -333 37 -327
rect 6402 -1153 8791 -1138
rect 6402 -1187 6483 -1153
rect 6517 -1187 6558 -1153
rect 6592 -1187 6633 -1153
rect 6667 -1187 6708 -1153
rect 6742 -1187 6783 -1153
rect 6817 -1187 6859 -1153
rect 6893 -1187 6935 -1153
rect 6969 -1187 7011 -1153
rect 7045 -1187 7087 -1153
rect 7121 -1187 7197 -1153
rect 7231 -1187 7271 -1153
rect 7305 -1187 7345 -1153
rect 7379 -1187 7419 -1153
rect 7453 -1187 7493 -1153
rect 7527 -1187 7567 -1153
rect 7601 -1187 7641 -1153
rect 7675 -1187 7715 -1153
rect 7749 -1187 7789 -1153
rect 7823 -1187 7863 -1153
rect 7897 -1187 7937 -1153
rect 7971 -1187 8011 -1153
rect 8045 -1187 8085 -1153
rect 8119 -1187 8159 -1153
rect 8193 -1187 8233 -1153
rect 8267 -1187 8307 -1153
rect 8341 -1187 8381 -1153
rect 8415 -1187 8455 -1153
rect 8489 -1187 8529 -1153
rect 8563 -1187 8604 -1153
rect 8638 -1187 8679 -1153
rect 8713 -1187 8791 -1153
rect 6402 -1202 8791 -1187
rect 6402 -1216 6466 -1202
rect 6402 -1250 6417 -1216
rect 6451 -1250 6466 -1216
rect 6402 -1294 6466 -1250
rect 8727 -1217 8791 -1202
rect 8727 -1251 8742 -1217
rect 8776 -1251 8791 -1217
rect 6402 -1328 6417 -1294
rect 6451 -1328 6466 -1294
rect 6640 -1313 6646 -1261
rect 6698 -1313 6711 -1261
rect 6763 -1313 6776 -1261
rect 6828 -1270 6841 -1261
rect 6893 -1270 6906 -1261
rect 6958 -1270 6971 -1261
rect 7023 -1270 7036 -1261
rect 6836 -1304 6841 -1270
rect 7023 -1304 7027 -1270
rect 6828 -1313 6841 -1304
rect 6893 -1313 6906 -1304
rect 6958 -1313 6971 -1304
rect 7023 -1313 7036 -1304
rect 7088 -1313 7101 -1261
rect 7153 -1313 7165 -1261
rect 7217 -1313 7229 -1261
rect 7281 -1270 7293 -1261
rect 7345 -1270 7357 -1261
rect 7409 -1270 7421 -1261
rect 7473 -1270 7485 -1261
rect 7286 -1304 7293 -1270
rect 7473 -1304 7476 -1270
rect 7281 -1313 7293 -1304
rect 7345 -1313 7357 -1304
rect 7409 -1313 7421 -1304
rect 7473 -1313 7485 -1304
rect 7537 -1313 7549 -1261
rect 7601 -1313 7613 -1261
rect 7665 -1313 7677 -1261
rect 7729 -1270 7741 -1261
rect 7793 -1270 7805 -1261
rect 7857 -1270 7869 -1261
rect 7921 -1270 7933 -1261
rect 7985 -1270 7997 -1261
rect 7732 -1304 7741 -1270
rect 7985 -1304 7994 -1270
rect 7729 -1313 7741 -1304
rect 7793 -1313 7805 -1304
rect 7857 -1313 7869 -1304
rect 7921 -1313 7933 -1304
rect 7985 -1313 7997 -1304
rect 8049 -1313 8061 -1261
rect 8113 -1313 8125 -1261
rect 8177 -1313 8189 -1261
rect 8241 -1270 8253 -1261
rect 8305 -1270 8317 -1261
rect 8369 -1270 8381 -1261
rect 8433 -1270 8445 -1261
rect 8250 -1304 8253 -1270
rect 8433 -1304 8438 -1270
rect 8241 -1313 8253 -1304
rect 8305 -1313 8317 -1304
rect 8369 -1313 8381 -1304
rect 8433 -1313 8445 -1304
rect 8497 -1313 8509 -1261
rect 8561 -1313 8573 -1261
rect 8625 -1264 8631 -1261
rect 8625 -1310 8632 -1264
rect 8727 -1290 8791 -1251
rect 8625 -1313 8631 -1310
rect 6402 -1372 6466 -1328
rect 6402 -1406 6417 -1372
rect 6451 -1406 6466 -1372
rect 6402 -1450 6466 -1406
rect 6522 -1321 6574 -1315
rect 6522 -1385 6574 -1373
rect 8727 -1324 8742 -1290
rect 8776 -1324 8791 -1290
rect 8727 -1363 8791 -1324
rect 8727 -1397 8742 -1363
rect 8776 -1397 8791 -1363
rect 6522 -1443 6574 -1437
rect 6402 -1484 6417 -1450
rect 6451 -1484 6466 -1450
rect 6402 -1528 6466 -1484
rect 6402 -1562 6417 -1528
rect 6451 -1562 6466 -1528
rect 6402 -1606 6466 -1562
rect 6402 -1640 6417 -1606
rect 6451 -1640 6466 -1606
rect 6402 -1684 6466 -1640
rect 6402 -1718 6417 -1684
rect 6451 -1718 6466 -1684
rect 6402 -1762 6466 -1718
rect 6402 -1796 6417 -1762
rect 6451 -1796 6466 -1762
rect 6402 -1840 6466 -1796
rect 6402 -1874 6417 -1840
rect 6451 -1874 6466 -1840
rect 6402 -1918 6466 -1874
rect 6528 -1472 6574 -1443
rect 6640 -1469 6646 -1417
rect 6698 -1469 6711 -1417
rect 6763 -1469 6776 -1417
rect 6828 -1426 6841 -1417
rect 6893 -1426 6906 -1417
rect 6958 -1426 6971 -1417
rect 7023 -1426 7036 -1417
rect 6836 -1460 6841 -1426
rect 7023 -1460 7027 -1426
rect 6828 -1469 6841 -1460
rect 6893 -1469 6906 -1460
rect 6958 -1469 6971 -1460
rect 7023 -1469 7036 -1460
rect 7088 -1469 7101 -1417
rect 7153 -1469 7165 -1417
rect 7217 -1469 7229 -1417
rect 7281 -1426 7293 -1417
rect 7345 -1426 7357 -1417
rect 7409 -1426 7421 -1417
rect 7473 -1426 7485 -1417
rect 7286 -1460 7293 -1426
rect 7473 -1460 7476 -1426
rect 7281 -1469 7293 -1460
rect 7345 -1469 7357 -1460
rect 7409 -1469 7421 -1460
rect 7473 -1469 7485 -1460
rect 7537 -1469 7549 -1417
rect 7601 -1469 7613 -1417
rect 7665 -1469 7677 -1417
rect 7729 -1426 7741 -1417
rect 7793 -1426 7805 -1417
rect 7857 -1426 7869 -1417
rect 7921 -1426 7933 -1417
rect 7985 -1426 7997 -1417
rect 7732 -1460 7741 -1426
rect 7985 -1460 7994 -1426
rect 7729 -1469 7741 -1460
rect 7793 -1469 7805 -1460
rect 7857 -1469 7869 -1460
rect 7921 -1469 7933 -1460
rect 7985 -1469 7997 -1460
rect 8049 -1469 8061 -1417
rect 8113 -1469 8125 -1417
rect 8177 -1469 8189 -1417
rect 8241 -1426 8253 -1417
rect 8305 -1426 8317 -1417
rect 8369 -1426 8381 -1417
rect 8433 -1426 8445 -1417
rect 8250 -1460 8253 -1426
rect 8433 -1460 8438 -1426
rect 8241 -1469 8253 -1460
rect 8305 -1469 8317 -1460
rect 8369 -1469 8381 -1460
rect 8433 -1469 8445 -1460
rect 8497 -1469 8509 -1417
rect 8561 -1469 8573 -1417
rect 8625 -1420 8631 -1417
rect 8625 -1466 8632 -1420
rect 8727 -1436 8791 -1397
rect 8625 -1469 8631 -1466
rect 6528 -1506 6534 -1472
rect 6568 -1506 6574 -1472
rect 6528 -1545 6574 -1506
rect 6528 -1579 6534 -1545
rect 6568 -1579 6574 -1545
rect 8727 -1470 8742 -1436
rect 8776 -1470 8791 -1436
rect 8727 -1509 8791 -1470
rect 8727 -1543 8742 -1509
rect 8776 -1543 8791 -1509
rect 6528 -1618 6574 -1579
rect 6528 -1652 6534 -1618
rect 6568 -1652 6574 -1618
rect 6640 -1625 6646 -1573
rect 6698 -1625 6711 -1573
rect 6763 -1625 6776 -1573
rect 6828 -1582 6841 -1573
rect 6893 -1582 6906 -1573
rect 6958 -1582 6971 -1573
rect 7023 -1582 7036 -1573
rect 6836 -1616 6841 -1582
rect 7023 -1616 7027 -1582
rect 6828 -1625 6841 -1616
rect 6893 -1625 6906 -1616
rect 6958 -1625 6971 -1616
rect 7023 -1625 7036 -1616
rect 7088 -1625 7101 -1573
rect 7153 -1625 7165 -1573
rect 7217 -1625 7229 -1573
rect 7281 -1582 7293 -1573
rect 7345 -1582 7357 -1573
rect 7409 -1582 7421 -1573
rect 7473 -1582 7485 -1573
rect 7286 -1616 7293 -1582
rect 7473 -1616 7476 -1582
rect 7281 -1625 7293 -1616
rect 7345 -1625 7357 -1616
rect 7409 -1625 7421 -1616
rect 7473 -1625 7485 -1616
rect 7537 -1625 7549 -1573
rect 7601 -1625 7613 -1573
rect 7665 -1625 7677 -1573
rect 7729 -1582 7741 -1573
rect 7793 -1582 7805 -1573
rect 7857 -1582 7869 -1573
rect 7921 -1582 7933 -1573
rect 7985 -1582 7997 -1573
rect 7732 -1616 7741 -1582
rect 7985 -1616 7994 -1582
rect 7729 -1625 7741 -1616
rect 7793 -1625 7805 -1616
rect 7857 -1625 7869 -1616
rect 7921 -1625 7933 -1616
rect 7985 -1625 7997 -1616
rect 8049 -1625 8061 -1573
rect 8113 -1625 8125 -1573
rect 8177 -1625 8189 -1573
rect 8241 -1582 8253 -1573
rect 8305 -1582 8317 -1573
rect 8369 -1582 8381 -1573
rect 8433 -1582 8445 -1573
rect 8250 -1616 8253 -1582
rect 8433 -1616 8438 -1582
rect 8241 -1625 8253 -1616
rect 8305 -1625 8317 -1616
rect 8369 -1625 8381 -1616
rect 8433 -1625 8445 -1616
rect 8497 -1625 8509 -1573
rect 8561 -1625 8573 -1573
rect 8625 -1576 8631 -1573
rect 8625 -1622 8632 -1576
rect 8727 -1582 8791 -1543
rect 8727 -1616 8742 -1582
rect 8776 -1616 8791 -1582
rect 8625 -1625 8631 -1622
rect 6528 -1691 6574 -1652
rect 6528 -1725 6534 -1691
rect 6568 -1725 6574 -1691
rect 6528 -1764 6574 -1725
rect 8727 -1655 8791 -1616
rect 8727 -1689 8742 -1655
rect 8776 -1689 8791 -1655
rect 8727 -1728 8791 -1689
rect 6528 -1798 6534 -1764
rect 6568 -1798 6574 -1764
rect 6640 -1781 6646 -1729
rect 6698 -1781 6711 -1729
rect 6763 -1781 6776 -1729
rect 6828 -1738 6841 -1729
rect 6893 -1738 6906 -1729
rect 6958 -1738 6971 -1729
rect 7023 -1738 7036 -1729
rect 6836 -1772 6841 -1738
rect 7023 -1772 7027 -1738
rect 6828 -1781 6841 -1772
rect 6893 -1781 6906 -1772
rect 6958 -1781 6971 -1772
rect 7023 -1781 7036 -1772
rect 7088 -1781 7101 -1729
rect 7153 -1781 7165 -1729
rect 7217 -1781 7229 -1729
rect 7281 -1738 7293 -1729
rect 7345 -1738 7357 -1729
rect 7409 -1738 7421 -1729
rect 7473 -1738 7485 -1729
rect 7286 -1772 7293 -1738
rect 7473 -1772 7476 -1738
rect 7281 -1781 7293 -1772
rect 7345 -1781 7357 -1772
rect 7409 -1781 7421 -1772
rect 7473 -1781 7485 -1772
rect 7537 -1781 7549 -1729
rect 7601 -1781 7613 -1729
rect 7665 -1781 7677 -1729
rect 7729 -1738 7741 -1729
rect 7793 -1738 7805 -1729
rect 7857 -1738 7869 -1729
rect 7921 -1738 7933 -1729
rect 7985 -1738 7997 -1729
rect 7732 -1772 7741 -1738
rect 7985 -1772 7994 -1738
rect 7729 -1781 7741 -1772
rect 7793 -1781 7805 -1772
rect 7857 -1781 7869 -1772
rect 7921 -1781 7933 -1772
rect 7985 -1781 7997 -1772
rect 8049 -1781 8061 -1729
rect 8113 -1781 8125 -1729
rect 8177 -1781 8189 -1729
rect 8241 -1738 8253 -1729
rect 8305 -1738 8317 -1729
rect 8369 -1738 8381 -1729
rect 8433 -1738 8445 -1729
rect 8250 -1772 8253 -1738
rect 8433 -1772 8438 -1738
rect 8241 -1781 8253 -1772
rect 8305 -1781 8317 -1772
rect 8369 -1781 8381 -1772
rect 8433 -1781 8445 -1772
rect 8497 -1781 8509 -1729
rect 8561 -1781 8573 -1729
rect 8625 -1732 8631 -1729
rect 8625 -1778 8632 -1732
rect 8727 -1762 8742 -1728
rect 8776 -1762 8791 -1728
rect 8625 -1781 8631 -1778
rect 6528 -1837 6574 -1798
rect 6528 -1871 6534 -1837
rect 6568 -1871 6574 -1837
rect 6528 -1883 6574 -1871
rect 8727 -1801 8791 -1762
rect 8727 -1835 8742 -1801
rect 8776 -1835 8791 -1801
rect 8727 -1874 8791 -1835
rect 6402 -1952 6417 -1918
rect 6451 -1952 6466 -1918
rect 6640 -1937 6646 -1885
rect 6698 -1937 6711 -1885
rect 6763 -1937 6776 -1885
rect 6828 -1894 6841 -1885
rect 6893 -1894 6906 -1885
rect 6958 -1894 6971 -1885
rect 7023 -1894 7036 -1885
rect 6836 -1928 6841 -1894
rect 7023 -1928 7027 -1894
rect 6828 -1937 6841 -1928
rect 6893 -1937 6906 -1928
rect 6958 -1937 6971 -1928
rect 7023 -1937 7036 -1928
rect 7088 -1937 7101 -1885
rect 7153 -1937 7165 -1885
rect 7217 -1937 7229 -1885
rect 7281 -1894 7293 -1885
rect 7345 -1894 7357 -1885
rect 7409 -1894 7421 -1885
rect 7473 -1894 7485 -1885
rect 7286 -1928 7293 -1894
rect 7473 -1928 7476 -1894
rect 7281 -1937 7293 -1928
rect 7345 -1937 7357 -1928
rect 7409 -1937 7421 -1928
rect 7473 -1937 7485 -1928
rect 7537 -1937 7549 -1885
rect 7601 -1937 7613 -1885
rect 7665 -1937 7677 -1885
rect 7729 -1894 7741 -1885
rect 7793 -1894 7805 -1885
rect 7857 -1894 7869 -1885
rect 7921 -1894 7933 -1885
rect 7985 -1894 7997 -1885
rect 7732 -1928 7741 -1894
rect 7985 -1928 7994 -1894
rect 7729 -1937 7741 -1928
rect 7793 -1937 7805 -1928
rect 7857 -1937 7869 -1928
rect 7921 -1937 7933 -1928
rect 7985 -1937 7997 -1928
rect 8049 -1937 8061 -1885
rect 8113 -1937 8125 -1885
rect 8177 -1937 8189 -1885
rect 8241 -1894 8253 -1885
rect 8305 -1894 8317 -1885
rect 8369 -1894 8381 -1885
rect 8433 -1894 8445 -1885
rect 8250 -1928 8253 -1894
rect 8433 -1928 8438 -1894
rect 8241 -1937 8253 -1928
rect 8305 -1937 8317 -1928
rect 8369 -1937 8381 -1928
rect 8433 -1937 8445 -1928
rect 8497 -1937 8509 -1885
rect 8561 -1937 8573 -1885
rect 8625 -1888 8631 -1885
rect 8625 -1934 8632 -1888
rect 8727 -1908 8742 -1874
rect 8776 -1908 8791 -1874
rect 8625 -1937 8631 -1934
rect 6402 -1971 6466 -1952
rect 8727 -1947 8791 -1908
rect 6402 -1986 6721 -1971
rect 6402 -2020 6480 -1986
rect 6514 -2020 6581 -1986
rect 6615 -1995 6721 -1986
rect 8727 -1981 8742 -1947
rect 8776 -1981 8791 -1947
rect 8727 -1995 8791 -1981
rect 6615 -2010 8791 -1995
rect 6615 -2020 6735 -2010
rect 6402 -2035 6735 -2020
rect 6657 -2044 6735 -2035
rect 6769 -2044 6807 -2010
rect 6841 -2044 6879 -2010
rect 6913 -2044 6951 -2010
rect 6985 -2044 7023 -2010
rect 7057 -2044 7095 -2010
rect 7129 -2044 7167 -2010
rect 7201 -2044 7239 -2010
rect 7273 -2044 7311 -2010
rect 7345 -2044 7383 -2010
rect 7417 -2044 7455 -2010
rect 7489 -2044 7527 -2010
rect 7561 -2044 7599 -2010
rect 7633 -2044 7671 -2010
rect 7705 -2044 7743 -2010
rect 7777 -2044 7815 -2010
rect 7849 -2044 7887 -2010
rect 7921 -2044 7959 -2010
rect 7993 -2044 8031 -2010
rect 8065 -2044 8103 -2010
rect 8137 -2044 8175 -2010
rect 8209 -2044 8247 -2010
rect 8281 -2044 8319 -2010
rect 8353 -2044 8391 -2010
rect 8425 -2044 8463 -2010
rect 8497 -2044 8535 -2010
rect 8569 -2044 8607 -2010
rect 8641 -2044 8679 -2010
rect 8713 -2044 8791 -2010
rect 6657 -2059 8791 -2044
<< via1 >>
rect -358 1395 -322 1428
rect -322 1395 -306 1428
rect -294 1395 -288 1428
rect -288 1395 -242 1428
rect -358 1376 -306 1395
rect -294 1376 -242 1395
rect -358 1319 -306 1355
rect -294 1319 -242 1355
rect -358 1303 -322 1319
rect -322 1303 -306 1319
rect -294 1303 -288 1319
rect -288 1303 -242 1319
rect -358 1230 -306 1282
rect -294 1230 -242 1282
rect -490 932 -118 1048
rect 640 1201 641 1224
rect 641 1201 675 1224
rect 675 1201 692 1224
rect 320 1031 324 1049
rect 324 1031 358 1049
rect 358 1031 372 1049
rect 320 997 372 1031
rect 384 1031 396 1049
rect 396 1031 430 1049
rect 430 1031 436 1049
rect 384 997 436 1031
rect 320 956 324 958
rect 324 956 358 958
rect 358 956 372 958
rect 320 915 372 956
rect 320 906 324 915
rect 324 906 358 915
rect 358 906 372 915
rect 384 956 396 958
rect 396 956 430 958
rect 430 956 436 958
rect 384 915 436 956
rect 384 906 396 915
rect 396 906 430 915
rect 430 906 436 915
rect 320 841 372 867
rect 320 815 324 841
rect 324 815 358 841
rect 358 815 372 841
rect 384 841 436 867
rect 384 815 396 841
rect 396 815 430 841
rect 430 815 436 841
rect 640 1172 692 1201
rect 712 1201 716 1224
rect 716 1201 750 1224
rect 750 1201 764 1224
rect 712 1172 764 1201
rect 784 1201 791 1224
rect 791 1201 825 1224
rect 825 1201 836 1224
rect 784 1172 836 1201
rect 855 1201 866 1224
rect 866 1201 900 1224
rect 900 1201 907 1224
rect 855 1172 907 1201
rect 640 1108 692 1160
rect 712 1108 764 1160
rect 784 1108 836 1160
rect 855 1108 907 1160
rect 1118 1081 1170 1133
rect 1195 1081 1247 1133
rect 1272 1081 1324 1133
rect 1348 1081 1400 1133
rect 1424 1081 1476 1133
rect 1500 1081 1552 1133
rect 1118 1042 1124 1055
rect 1124 1042 1158 1055
rect 1158 1042 1170 1055
rect 1118 1003 1170 1042
rect 1195 1042 1202 1055
rect 1202 1042 1236 1055
rect 1236 1042 1247 1055
rect 1195 1003 1247 1042
rect 1272 1042 1280 1055
rect 1280 1042 1314 1055
rect 1314 1042 1324 1055
rect 1272 1003 1324 1042
rect 1348 1042 1358 1055
rect 1358 1042 1392 1055
rect 1392 1042 1400 1055
rect 1348 1003 1400 1042
rect 1424 1042 1435 1055
rect 1435 1042 1469 1055
rect 1469 1042 1476 1055
rect 1424 1003 1476 1042
rect 1500 1042 1512 1055
rect 1512 1042 1546 1055
rect 1546 1042 1552 1055
rect 1500 1003 1552 1042
rect 1631 919 1747 931
rect 1631 885 1636 919
rect 1636 885 1670 919
rect 1670 885 1708 919
rect 1708 885 1742 919
rect 1742 885 1747 919
rect 1631 845 1747 885
rect 1631 815 1636 845
rect 1636 815 1670 845
rect 1670 815 1708 845
rect 1708 815 1742 845
rect 1742 815 1747 845
rect 640 756 641 759
rect 641 756 675 759
rect 675 756 692 759
rect 640 707 692 756
rect 712 756 716 759
rect 716 756 750 759
rect 750 756 764 759
rect 712 707 764 756
rect 784 756 791 759
rect 791 756 825 759
rect 825 756 836 759
rect 784 707 836 756
rect 855 756 866 759
rect 866 756 900 759
rect 900 756 907 759
rect 855 707 907 756
rect 640 643 692 695
rect 712 643 764 695
rect 784 643 836 695
rect 855 643 907 695
rect 1117 634 1169 682
rect 1117 630 1123 634
rect 1123 630 1157 634
rect 1157 630 1169 634
rect 1194 634 1246 682
rect 1194 630 1201 634
rect 1201 630 1235 634
rect 1235 630 1246 634
rect 1271 634 1323 682
rect 1271 630 1279 634
rect 1279 630 1313 634
rect 1313 630 1323 634
rect 1348 634 1400 682
rect 1348 630 1357 634
rect 1357 630 1391 634
rect 1391 630 1400 634
rect 1424 634 1476 682
rect 1424 630 1435 634
rect 1435 630 1469 634
rect 1469 630 1476 634
rect 1500 634 1552 682
rect 1500 630 1512 634
rect 1512 630 1546 634
rect 1546 630 1552 634
rect 1117 600 1123 604
rect 1123 600 1157 604
rect 1157 600 1169 604
rect 1117 552 1169 600
rect 1194 600 1201 604
rect 1201 600 1235 604
rect 1235 600 1246 604
rect 1194 552 1246 600
rect 1271 600 1279 604
rect 1279 600 1313 604
rect 1313 600 1323 604
rect 1271 552 1323 600
rect 1348 600 1357 604
rect 1357 600 1391 604
rect 1391 600 1400 604
rect 1348 552 1400 600
rect 1424 600 1435 604
rect 1435 600 1469 604
rect 1469 600 1476 604
rect 1424 552 1476 600
rect 1500 600 1512 604
rect 1512 600 1546 604
rect 1546 600 1552 604
rect 1500 552 1552 600
rect 473 488 476 496
rect 476 488 510 496
rect 510 488 525 496
rect 473 444 525 488
rect 537 444 589 496
rect 1931 1423 1983 1438
rect 1931 1389 1938 1423
rect 1938 1389 1976 1423
rect 1976 1389 1983 1423
rect 1931 1386 1983 1389
rect 1931 1349 1983 1365
rect 1931 1315 1938 1349
rect 1938 1315 1976 1349
rect 1976 1315 1983 1349
rect 1931 1313 1983 1315
rect 1931 1275 1983 1291
rect 1931 1241 1938 1275
rect 1938 1241 1976 1275
rect 1976 1241 1983 1275
rect 1931 1239 1983 1241
rect 3599 1450 3651 1456
rect 3665 1450 3717 1456
rect 3731 1450 3783 1456
rect 3797 1450 3849 1456
rect 3863 1450 3915 1456
rect 3929 1450 3981 1456
rect 3995 1450 4047 1456
rect 3599 1416 3624 1450
rect 3624 1416 3651 1450
rect 3665 1416 3697 1450
rect 3697 1416 3717 1450
rect 3731 1416 3770 1450
rect 3770 1416 3783 1450
rect 3797 1416 3804 1450
rect 3804 1416 3843 1450
rect 3843 1416 3849 1450
rect 3863 1416 3877 1450
rect 3877 1416 3915 1450
rect 3929 1416 3950 1450
rect 3950 1416 3981 1450
rect 3995 1416 4023 1450
rect 4023 1416 4047 1450
rect 3599 1404 3651 1416
rect 3665 1404 3717 1416
rect 3731 1404 3783 1416
rect 3797 1404 3849 1416
rect 3863 1404 3915 1416
rect 3929 1404 3981 1416
rect 3995 1404 4047 1416
rect 4061 1450 4113 1456
rect 4061 1416 4062 1450
rect 4062 1416 4096 1450
rect 4096 1416 4113 1450
rect 4061 1404 4113 1416
rect 4127 1450 4179 1456
rect 4127 1416 4135 1450
rect 4135 1416 4169 1450
rect 4169 1416 4179 1450
rect 4127 1404 4179 1416
rect 4193 1450 4245 1456
rect 4193 1416 4208 1450
rect 4208 1416 4242 1450
rect 4242 1416 4245 1450
rect 4193 1404 4245 1416
rect 4259 1450 4311 1456
rect 4325 1450 4377 1456
rect 4391 1450 4443 1456
rect 4457 1450 4509 1456
rect 4523 1450 4575 1456
rect 4589 1450 4641 1456
rect 4655 1450 4707 1456
rect 4721 1450 4773 1456
rect 4259 1416 4281 1450
rect 4281 1416 4311 1450
rect 4325 1416 4354 1450
rect 4354 1416 4377 1450
rect 4391 1416 4427 1450
rect 4427 1416 4443 1450
rect 4457 1416 4461 1450
rect 4461 1416 4500 1450
rect 4500 1416 4509 1450
rect 4523 1416 4534 1450
rect 4534 1416 4573 1450
rect 4573 1416 4575 1450
rect 4589 1416 4607 1450
rect 4607 1416 4641 1450
rect 4655 1416 4680 1450
rect 4680 1416 4707 1450
rect 4721 1416 4753 1450
rect 4753 1416 4773 1450
rect 4259 1404 4311 1416
rect 4325 1404 4377 1416
rect 4391 1404 4443 1416
rect 4457 1404 4509 1416
rect 4523 1404 4575 1416
rect 4589 1404 4641 1416
rect 4655 1404 4707 1416
rect 4721 1404 4773 1416
rect 4786 1450 4838 1456
rect 4786 1416 4792 1450
rect 4792 1416 4826 1450
rect 4826 1416 4838 1450
rect 4786 1404 4838 1416
rect 4851 1450 4903 1456
rect 4851 1416 4865 1450
rect 4865 1416 4899 1450
rect 4899 1416 4903 1450
rect 4851 1404 4903 1416
rect 4916 1450 4968 1456
rect 4981 1450 5033 1456
rect 5046 1450 5098 1456
rect 5111 1450 5163 1456
rect 5176 1450 5228 1456
rect 5241 1450 5293 1456
rect 6626 1450 6678 1456
rect 4916 1416 4938 1450
rect 4938 1416 4968 1450
rect 4981 1416 5011 1450
rect 5011 1416 5033 1450
rect 5046 1416 5084 1450
rect 5084 1416 5098 1450
rect 5111 1416 5118 1450
rect 5118 1416 5157 1450
rect 5157 1416 5163 1450
rect 5176 1416 5191 1450
rect 5191 1416 5228 1450
rect 5241 1416 5264 1450
rect 5264 1416 5293 1450
rect 6626 1416 6627 1450
rect 6627 1416 6661 1450
rect 6661 1416 6678 1450
rect 4916 1404 4968 1416
rect 4981 1404 5033 1416
rect 5046 1404 5098 1416
rect 5111 1404 5163 1416
rect 5176 1404 5228 1416
rect 5241 1404 5293 1416
rect 6626 1404 6678 1416
rect 6731 1404 6783 1456
rect 3599 1378 3651 1392
rect 3665 1378 3717 1392
rect 3731 1378 3783 1392
rect 3797 1378 3849 1392
rect 3863 1378 3915 1392
rect 3929 1378 3981 1392
rect 3995 1378 4047 1392
rect 3599 1344 3624 1378
rect 3624 1344 3651 1378
rect 3665 1344 3697 1378
rect 3697 1344 3717 1378
rect 3731 1344 3770 1378
rect 3770 1344 3783 1378
rect 3797 1344 3804 1378
rect 3804 1344 3843 1378
rect 3843 1344 3849 1378
rect 3863 1344 3877 1378
rect 3877 1344 3915 1378
rect 3929 1344 3950 1378
rect 3950 1344 3981 1378
rect 3995 1344 4023 1378
rect 4023 1344 4047 1378
rect 3599 1340 3651 1344
rect 3665 1340 3717 1344
rect 3731 1340 3783 1344
rect 3797 1340 3849 1344
rect 3863 1340 3915 1344
rect 3929 1340 3981 1344
rect 3995 1340 4047 1344
rect 4061 1378 4113 1392
rect 4061 1344 4062 1378
rect 4062 1344 4096 1378
rect 4096 1344 4113 1378
rect 4061 1340 4113 1344
rect 4127 1378 4179 1392
rect 4127 1344 4135 1378
rect 4135 1344 4169 1378
rect 4169 1344 4179 1378
rect 4127 1340 4179 1344
rect 4193 1378 4245 1392
rect 4193 1344 4208 1378
rect 4208 1344 4242 1378
rect 4242 1344 4245 1378
rect 4193 1340 4245 1344
rect 4259 1378 4311 1392
rect 4325 1378 4377 1392
rect 4391 1378 4443 1392
rect 4457 1378 4509 1392
rect 4523 1378 4575 1392
rect 4589 1378 4641 1392
rect 4655 1378 4707 1392
rect 4721 1378 4773 1392
rect 4259 1344 4281 1378
rect 4281 1344 4311 1378
rect 4325 1344 4354 1378
rect 4354 1344 4377 1378
rect 4391 1344 4427 1378
rect 4427 1344 4443 1378
rect 4457 1344 4461 1378
rect 4461 1344 4500 1378
rect 4500 1344 4509 1378
rect 4523 1344 4534 1378
rect 4534 1344 4573 1378
rect 4573 1344 4575 1378
rect 4589 1344 4607 1378
rect 4607 1344 4641 1378
rect 4655 1344 4680 1378
rect 4680 1344 4707 1378
rect 4721 1344 4753 1378
rect 4753 1344 4773 1378
rect 4259 1340 4311 1344
rect 4325 1340 4377 1344
rect 4391 1340 4443 1344
rect 4457 1340 4509 1344
rect 4523 1340 4575 1344
rect 4589 1340 4641 1344
rect 4655 1340 4707 1344
rect 4721 1340 4773 1344
rect 4786 1378 4838 1392
rect 4786 1344 4792 1378
rect 4792 1344 4826 1378
rect 4826 1344 4838 1378
rect 4786 1340 4838 1344
rect 4851 1378 4903 1392
rect 4851 1344 4865 1378
rect 4865 1344 4899 1378
rect 4899 1344 4903 1378
rect 4851 1340 4903 1344
rect 4916 1378 4968 1392
rect 4981 1378 5033 1392
rect 5046 1378 5098 1392
rect 5111 1378 5163 1392
rect 5176 1378 5228 1392
rect 5241 1378 5293 1392
rect 6626 1378 6678 1392
rect 6731 1378 6783 1392
rect 4916 1344 4938 1378
rect 4938 1344 4968 1378
rect 4981 1344 5011 1378
rect 5011 1344 5033 1378
rect 5046 1344 5084 1378
rect 5084 1344 5098 1378
rect 5111 1344 5118 1378
rect 5118 1344 5157 1378
rect 5157 1344 5163 1378
rect 5176 1344 5191 1378
rect 5191 1344 5228 1378
rect 5241 1344 5264 1378
rect 5264 1344 5293 1378
rect 4916 1340 4968 1344
rect 4981 1340 5033 1344
rect 5046 1340 5098 1344
rect 5111 1340 5163 1344
rect 5176 1340 5228 1344
rect 5241 1340 5293 1344
rect 6626 1340 6627 1378
rect 6627 1340 6678 1378
rect 6731 1340 6733 1378
rect 6733 1340 6783 1378
rect 6626 1276 6627 1328
rect 6627 1276 6678 1328
rect 6731 1276 6733 1328
rect 6733 1276 6783 1328
rect 3136 1258 3188 1267
rect 3136 1224 3141 1258
rect 3141 1224 3175 1258
rect 3175 1224 3188 1258
rect 3136 1215 3188 1224
rect 3203 1258 3255 1267
rect 3203 1224 3215 1258
rect 3215 1224 3249 1258
rect 3249 1224 3255 1258
rect 3203 1215 3255 1224
rect 3269 1258 3321 1267
rect 3335 1258 3387 1267
rect 3401 1258 3453 1267
rect 3269 1224 3289 1258
rect 3289 1224 3321 1258
rect 3335 1224 3363 1258
rect 3363 1224 3387 1258
rect 3401 1224 3437 1258
rect 3437 1224 3453 1258
rect 3269 1215 3321 1224
rect 3335 1215 3387 1224
rect 3401 1215 3453 1224
rect 5870 1258 5922 1267
rect 5870 1224 5899 1258
rect 5899 1224 5922 1258
rect 5870 1215 5922 1224
rect 5935 1258 5987 1267
rect 5935 1224 5939 1258
rect 5939 1224 5973 1258
rect 5973 1224 5987 1258
rect 5935 1215 5987 1224
rect 5999 1258 6051 1267
rect 5999 1224 6013 1258
rect 6013 1224 6047 1258
rect 6047 1224 6051 1258
rect 5999 1215 6051 1224
rect 6063 1258 6115 1267
rect 6127 1258 6179 1267
rect 6191 1258 6243 1267
rect 6255 1258 6307 1267
rect 6319 1258 6371 1267
rect 6063 1224 6087 1258
rect 6087 1224 6115 1258
rect 6127 1224 6161 1258
rect 6161 1224 6179 1258
rect 6191 1224 6195 1258
rect 6195 1224 6235 1258
rect 6235 1224 6243 1258
rect 6255 1224 6269 1258
rect 6269 1224 6307 1258
rect 6319 1224 6343 1258
rect 6343 1224 6371 1258
rect 6063 1215 6115 1224
rect 6127 1215 6179 1224
rect 6191 1215 6243 1224
rect 6255 1215 6307 1224
rect 6319 1215 6371 1224
rect 6383 1258 6435 1267
rect 6383 1224 6417 1258
rect 6417 1224 6435 1258
rect 6383 1215 6435 1224
rect 6447 1258 6499 1267
rect 6447 1224 6457 1258
rect 6457 1224 6491 1258
rect 6491 1224 6499 1258
rect 6447 1215 6499 1224
rect 2154 1198 2159 1206
rect 2159 1198 2193 1206
rect 2193 1198 2206 1206
rect 2154 1159 2206 1198
rect 2154 1154 2159 1159
rect 2159 1154 2193 1159
rect 2193 1154 2206 1159
rect 2218 1198 2231 1206
rect 2231 1198 2265 1206
rect 2265 1198 2270 1206
rect 2218 1159 2270 1198
rect 2218 1154 2231 1159
rect 2231 1154 2265 1159
rect 2265 1154 2270 1159
rect 2154 1125 2159 1140
rect 2159 1125 2193 1140
rect 2193 1125 2206 1140
rect 2154 1088 2206 1125
rect 2218 1125 2231 1140
rect 2231 1125 2265 1140
rect 2265 1125 2270 1140
rect 2218 1088 2270 1125
rect 2154 1052 2159 1074
rect 2159 1052 2193 1074
rect 2193 1052 2206 1074
rect 2154 1022 2206 1052
rect 2218 1052 2231 1074
rect 2231 1052 2265 1074
rect 2265 1052 2270 1074
rect 2218 1022 2270 1052
rect 2305 1201 2357 1207
rect 2305 1167 2311 1201
rect 2311 1167 2345 1201
rect 2345 1167 2357 1201
rect 2305 1155 2357 1167
rect 2305 1120 2357 1137
rect 2305 1086 2311 1120
rect 2311 1086 2345 1120
rect 2345 1086 2357 1120
rect 6539 1201 6591 1207
rect 6539 1167 6547 1201
rect 6547 1167 6581 1201
rect 6581 1167 6591 1201
rect 6539 1155 6591 1167
rect 6539 1118 6591 1137
rect 2305 1085 2357 1086
rect 2305 1038 2357 1067
rect 3599 1102 3651 1111
rect 3670 1102 3722 1111
rect 3741 1102 3793 1111
rect 3811 1102 3863 1111
rect 3881 1102 3933 1111
rect 3951 1102 4003 1111
rect 3599 1068 3617 1102
rect 3617 1068 3651 1102
rect 3670 1068 3690 1102
rect 3690 1068 3722 1102
rect 3741 1068 3763 1102
rect 3763 1068 3793 1102
rect 3811 1068 3836 1102
rect 3836 1068 3863 1102
rect 3881 1068 3909 1102
rect 3909 1068 3933 1102
rect 3951 1068 3982 1102
rect 3982 1068 4003 1102
rect 3599 1059 3651 1068
rect 3670 1059 3722 1068
rect 3741 1059 3793 1068
rect 3811 1059 3863 1068
rect 3881 1059 3933 1068
rect 3951 1059 4003 1068
rect 4021 1102 4073 1111
rect 4021 1068 4055 1102
rect 4055 1068 4073 1102
rect 4021 1059 4073 1068
rect 4091 1102 4143 1111
rect 4091 1068 4094 1102
rect 4094 1068 4128 1102
rect 4128 1068 4143 1102
rect 4091 1059 4143 1068
rect 4161 1102 4213 1111
rect 4161 1068 4167 1102
rect 4167 1068 4201 1102
rect 4201 1068 4213 1102
rect 4161 1059 4213 1068
rect 4231 1102 4283 1111
rect 4231 1068 4240 1102
rect 4240 1068 4274 1102
rect 4274 1068 4283 1102
rect 4231 1059 4283 1068
rect 4301 1102 4353 1111
rect 4301 1068 4313 1102
rect 4313 1068 4347 1102
rect 4347 1068 4353 1102
rect 4301 1059 4353 1068
rect 4539 1102 4591 1111
rect 4539 1068 4545 1102
rect 4545 1068 4579 1102
rect 4579 1068 4591 1102
rect 4539 1059 4591 1068
rect 4609 1102 4661 1111
rect 4609 1068 4618 1102
rect 4618 1068 4652 1102
rect 4652 1068 4661 1102
rect 4609 1059 4661 1068
rect 4679 1102 4731 1111
rect 4679 1068 4691 1102
rect 4691 1068 4725 1102
rect 4725 1068 4731 1102
rect 4679 1059 4731 1068
rect 4749 1102 4801 1111
rect 4749 1068 4764 1102
rect 4764 1068 4798 1102
rect 4798 1068 4801 1102
rect 4749 1059 4801 1068
rect 4819 1102 4871 1111
rect 4819 1068 4837 1102
rect 4837 1068 4871 1102
rect 4819 1059 4871 1068
rect 4889 1102 4941 1111
rect 4959 1102 5011 1111
rect 5029 1102 5081 1111
rect 5099 1102 5151 1111
rect 5170 1102 5222 1111
rect 5241 1102 5293 1111
rect 4889 1068 4910 1102
rect 4910 1068 4941 1102
rect 4959 1068 4983 1102
rect 4983 1068 5011 1102
rect 5029 1068 5056 1102
rect 5056 1068 5081 1102
rect 5099 1068 5129 1102
rect 5129 1068 5151 1102
rect 5170 1068 5202 1102
rect 5202 1068 5222 1102
rect 5241 1068 5275 1102
rect 5275 1068 5293 1102
rect 4889 1059 4941 1068
rect 4959 1059 5011 1068
rect 5029 1059 5081 1068
rect 5099 1059 5151 1068
rect 5170 1059 5222 1068
rect 5241 1059 5293 1068
rect 6539 1085 6547 1118
rect 6547 1085 6581 1118
rect 6581 1085 6591 1118
rect 2305 1015 2311 1038
rect 2311 1015 2345 1038
rect 2345 1015 2357 1038
rect 2305 956 2357 998
rect 2305 946 2311 956
rect 2311 946 2345 956
rect 2345 946 2357 956
rect 6539 1035 6591 1067
rect 6539 1015 6547 1035
rect 6547 1015 6581 1035
rect 6581 1015 6591 1035
rect 2305 922 2311 929
rect 2311 922 2345 929
rect 2345 922 2357 929
rect 2305 877 2357 922
rect 3136 946 3188 955
rect 3136 912 3141 946
rect 3141 912 3175 946
rect 3175 912 3188 946
rect 3136 903 3188 912
rect 3203 946 3255 955
rect 3203 912 3215 946
rect 3215 912 3249 946
rect 3249 912 3255 946
rect 3203 903 3255 912
rect 3269 946 3321 955
rect 3335 946 3387 955
rect 3401 946 3453 955
rect 3269 912 3289 946
rect 3289 912 3321 946
rect 3335 912 3363 946
rect 3363 912 3387 946
rect 3401 912 3437 946
rect 3437 912 3453 946
rect 3269 903 3321 912
rect 3335 903 3387 912
rect 3401 903 3453 912
rect 5870 946 5922 955
rect 5870 912 5899 946
rect 5899 912 5922 946
rect 5870 903 5922 912
rect 5935 946 5987 955
rect 5935 912 5939 946
rect 5939 912 5973 946
rect 5973 912 5987 946
rect 5935 903 5987 912
rect 5999 946 6051 955
rect 5999 912 6013 946
rect 6013 912 6047 946
rect 6047 912 6051 946
rect 5999 903 6051 912
rect 6063 946 6115 955
rect 6127 946 6179 955
rect 6191 946 6243 955
rect 6255 946 6307 955
rect 6319 946 6371 955
rect 6063 912 6087 946
rect 6087 912 6115 946
rect 6127 912 6161 946
rect 6161 912 6179 946
rect 6191 912 6195 946
rect 6195 912 6235 946
rect 6235 912 6243 946
rect 6255 912 6269 946
rect 6269 912 6307 946
rect 6319 912 6343 946
rect 6343 912 6371 946
rect 6063 903 6115 912
rect 6127 903 6179 912
rect 6191 903 6243 912
rect 6255 903 6307 912
rect 6319 903 6371 912
rect 6383 946 6435 955
rect 6383 912 6417 946
rect 6417 912 6435 946
rect 6383 903 6435 912
rect 6447 946 6499 955
rect 6447 912 6457 946
rect 6457 912 6491 946
rect 6491 912 6499 946
rect 6447 903 6499 912
rect 6539 952 6591 996
rect 6539 944 6547 952
rect 6547 944 6581 952
rect 6581 944 6591 952
rect 6539 918 6547 925
rect 6547 918 6581 925
rect 6581 918 6591 925
rect 2305 840 2311 860
rect 2311 840 2345 860
rect 2345 840 2357 860
rect 2305 808 2357 840
rect 6539 873 6591 918
rect 6539 834 6547 854
rect 6547 834 6581 854
rect 6581 834 6591 854
rect 6539 802 6591 834
rect 2305 758 2311 791
rect 2311 758 2345 791
rect 2345 758 2357 791
rect 2305 739 2357 758
rect 3599 790 3651 799
rect 3670 790 3722 799
rect 3741 790 3793 799
rect 3811 790 3863 799
rect 3881 790 3933 799
rect 3951 790 4003 799
rect 3599 756 3617 790
rect 3617 756 3651 790
rect 3670 756 3690 790
rect 3690 756 3722 790
rect 3741 756 3763 790
rect 3763 756 3793 790
rect 3811 756 3836 790
rect 3836 756 3863 790
rect 3881 756 3909 790
rect 3909 756 3933 790
rect 3951 756 3982 790
rect 3982 756 4003 790
rect 3599 747 3651 756
rect 3670 747 3722 756
rect 3741 747 3793 756
rect 3811 747 3863 756
rect 3881 747 3933 756
rect 3951 747 4003 756
rect 4021 790 4073 799
rect 4021 756 4055 790
rect 4055 756 4073 790
rect 4021 747 4073 756
rect 4091 790 4143 799
rect 4091 756 4094 790
rect 4094 756 4128 790
rect 4128 756 4143 790
rect 4091 747 4143 756
rect 4161 790 4213 799
rect 4161 756 4167 790
rect 4167 756 4201 790
rect 4201 756 4213 790
rect 4161 747 4213 756
rect 4231 790 4283 799
rect 4231 756 4240 790
rect 4240 756 4274 790
rect 4274 756 4283 790
rect 4231 747 4283 756
rect 4301 790 4353 799
rect 4301 756 4313 790
rect 4313 756 4347 790
rect 4347 756 4353 790
rect 4301 747 4353 756
rect 4539 790 4591 799
rect 4539 756 4545 790
rect 4545 756 4579 790
rect 4579 756 4591 790
rect 4539 747 4591 756
rect 4609 790 4661 799
rect 4609 756 4618 790
rect 4618 756 4652 790
rect 4652 756 4661 790
rect 4609 747 4661 756
rect 4679 790 4731 799
rect 4679 756 4691 790
rect 4691 756 4725 790
rect 4725 756 4731 790
rect 4679 747 4731 756
rect 4749 790 4801 799
rect 4749 756 4764 790
rect 4764 756 4798 790
rect 4798 756 4801 790
rect 4749 747 4801 756
rect 4819 790 4871 799
rect 4819 756 4837 790
rect 4837 756 4871 790
rect 4819 747 4871 756
rect 4889 790 4941 799
rect 4959 790 5011 799
rect 5029 790 5081 799
rect 5099 790 5151 799
rect 5170 790 5222 799
rect 5241 790 5293 799
rect 4889 756 4910 790
rect 4910 756 4941 790
rect 4959 756 4983 790
rect 4983 756 5011 790
rect 5029 756 5056 790
rect 5056 756 5081 790
rect 5099 756 5129 790
rect 5129 756 5151 790
rect 5170 756 5202 790
rect 5202 756 5222 790
rect 5241 756 5275 790
rect 5275 756 5293 790
rect 4889 747 4941 756
rect 4959 747 5011 756
rect 5029 747 5081 756
rect 5099 747 5151 756
rect 5170 747 5222 756
rect 5241 747 5293 756
rect 6539 750 6547 783
rect 6547 750 6581 783
rect 6581 750 6591 783
rect 2305 710 2357 722
rect 2305 676 2311 710
rect 2311 676 2345 710
rect 2345 676 2357 710
rect 2305 670 2357 676
rect 6539 731 6591 750
rect 6539 700 6591 712
rect 6539 666 6547 700
rect 6547 666 6581 700
rect 6581 666 6591 700
rect 6539 660 6591 666
rect 3136 634 3188 643
rect 3136 600 3141 634
rect 3141 600 3175 634
rect 3175 600 3188 634
rect 3136 591 3188 600
rect 3203 634 3255 643
rect 3203 600 3215 634
rect 3215 600 3249 634
rect 3249 600 3255 634
rect 3203 591 3255 600
rect 3269 634 3321 643
rect 3335 634 3387 643
rect 3401 634 3453 643
rect 3269 600 3289 634
rect 3289 600 3321 634
rect 3335 600 3363 634
rect 3363 600 3387 634
rect 3401 600 3437 634
rect 3437 600 3453 634
rect 3269 591 3321 600
rect 3335 591 3387 600
rect 3401 591 3453 600
rect 5870 634 5922 643
rect 5870 600 5899 634
rect 5899 600 5922 634
rect 5870 591 5922 600
rect 5935 634 5987 643
rect 5935 600 5939 634
rect 5939 600 5973 634
rect 5973 600 5987 634
rect 5935 591 5987 600
rect 5999 634 6051 643
rect 5999 600 6013 634
rect 6013 600 6047 634
rect 6047 600 6051 634
rect 5999 591 6051 600
rect 6063 634 6115 643
rect 6127 634 6179 643
rect 6191 634 6243 643
rect 6255 634 6307 643
rect 6319 634 6371 643
rect 6063 600 6087 634
rect 6087 600 6115 634
rect 6127 600 6161 634
rect 6161 600 6179 634
rect 6191 600 6195 634
rect 6195 600 6235 634
rect 6235 600 6243 634
rect 6255 600 6269 634
rect 6269 600 6307 634
rect 6319 600 6343 634
rect 6343 600 6371 634
rect 6063 591 6115 600
rect 6127 591 6179 600
rect 6191 591 6243 600
rect 6255 591 6307 600
rect 6319 591 6371 600
rect 6383 634 6435 643
rect 6383 600 6417 634
rect 6417 600 6435 634
rect 6383 591 6435 600
rect 6447 634 6499 643
rect 6447 600 6457 634
rect 6457 600 6491 634
rect 6491 600 6499 634
rect 6447 591 6499 600
rect 3599 478 3651 487
rect 3670 478 3722 487
rect 3741 478 3793 487
rect 3811 478 3863 487
rect 3881 478 3933 487
rect 3951 478 4003 487
rect 3599 444 3617 478
rect 3617 444 3651 478
rect 3670 444 3690 478
rect 3690 444 3722 478
rect 3741 444 3763 478
rect 3763 444 3793 478
rect 3811 444 3836 478
rect 3836 444 3863 478
rect 3881 444 3909 478
rect 3909 444 3933 478
rect 3951 444 3982 478
rect 3982 444 4003 478
rect 3599 435 3651 444
rect 3670 435 3722 444
rect 3741 435 3793 444
rect 3811 435 3863 444
rect 3881 435 3933 444
rect 3951 435 4003 444
rect 4021 478 4073 487
rect 4021 444 4055 478
rect 4055 444 4073 478
rect 4021 435 4073 444
rect 4091 478 4143 487
rect 4091 444 4094 478
rect 4094 444 4128 478
rect 4128 444 4143 478
rect 4091 435 4143 444
rect 4161 478 4213 487
rect 4161 444 4167 478
rect 4167 444 4201 478
rect 4201 444 4213 478
rect 4161 435 4213 444
rect 4231 478 4283 487
rect 4231 444 4240 478
rect 4240 444 4274 478
rect 4274 444 4283 478
rect 4231 435 4283 444
rect 4301 478 4353 487
rect 4301 444 4313 478
rect 4313 444 4347 478
rect 4347 444 4353 478
rect 4301 435 4353 444
rect 4539 478 4591 487
rect 4539 444 4545 478
rect 4545 444 4579 478
rect 4579 444 4591 478
rect 4539 435 4591 444
rect 4609 478 4661 487
rect 4609 444 4618 478
rect 4618 444 4652 478
rect 4652 444 4661 478
rect 4609 435 4661 444
rect 4679 478 4731 487
rect 4679 444 4691 478
rect 4691 444 4725 478
rect 4725 444 4731 478
rect 4679 435 4731 444
rect 4749 478 4801 487
rect 4749 444 4764 478
rect 4764 444 4798 478
rect 4798 444 4801 478
rect 4749 435 4801 444
rect 4819 478 4871 487
rect 4819 444 4837 478
rect 4837 444 4871 478
rect 4819 435 4871 444
rect 4889 478 4941 487
rect 4959 478 5011 487
rect 5029 478 5081 487
rect 5099 478 5151 487
rect 5170 478 5222 487
rect 5241 478 5293 487
rect 4889 444 4910 478
rect 4910 444 4941 478
rect 4959 444 4983 478
rect 4983 444 5011 478
rect 5029 444 5056 478
rect 5056 444 5081 478
rect 5099 444 5129 478
rect 5129 444 5151 478
rect 5170 444 5202 478
rect 5202 444 5222 478
rect 5241 444 5275 478
rect 5275 444 5293 478
rect 6655 470 6661 493
rect 6661 470 6699 493
rect 6699 470 6707 493
rect 4889 435 4941 444
rect 4959 435 5011 444
rect 5029 435 5081 444
rect 5099 435 5151 444
rect 5170 435 5222 444
rect 5241 435 5293 444
rect 6655 441 6707 470
rect 6760 441 6812 493
rect 3599 367 3651 419
rect 3665 367 3717 419
rect 3731 367 3783 419
rect 3797 367 3849 419
rect 3863 367 3915 419
rect 3929 367 3981 419
rect 3995 367 4047 419
rect 4061 367 4113 419
rect 4127 367 4179 419
rect 4193 367 4245 419
rect 4259 367 4311 419
rect 4325 367 4377 419
rect 4391 367 4443 419
rect 4457 367 4509 419
rect 4523 367 4575 419
rect 4589 367 4641 419
rect 4655 367 4707 419
rect 4721 367 4773 419
rect 4786 367 4838 419
rect 4851 367 4903 419
rect 4916 367 4968 419
rect 4981 367 5033 419
rect 5046 367 5098 419
rect 5111 367 5163 419
rect 5176 367 5228 419
rect 5241 367 5293 419
rect 6655 397 6661 429
rect 6661 397 6699 429
rect 6699 397 6707 429
rect 6655 377 6707 397
rect 6760 377 6812 429
rect 6655 358 6707 365
rect 6655 313 6661 358
rect 6661 324 6699 358
rect 6699 324 6707 358
rect 6661 313 6707 324
rect 6760 313 6812 365
rect 6909 909 6961 942
rect 6909 890 6916 909
rect 6916 890 6954 909
rect 6954 890 6961 909
rect 6909 875 6916 876
rect 6916 875 6954 876
rect 6954 875 6961 876
rect 6909 835 6961 875
rect 6909 824 6916 835
rect 6916 824 6954 835
rect 6954 824 6961 835
rect 6909 801 6916 810
rect 6916 801 6954 810
rect 6954 801 6961 810
rect 6909 761 6961 801
rect 6909 758 6916 761
rect 6916 758 6954 761
rect 6954 758 6961 761
rect 6909 727 6916 744
rect 6916 727 6954 744
rect 6954 727 6961 744
rect 6909 692 6961 727
rect 6909 653 6916 677
rect 6916 653 6954 677
rect 6954 653 6961 677
rect 6909 625 6961 653
rect 8741 1440 8793 1454
rect 8808 1440 8860 1454
rect 8874 1440 8926 1454
rect 8940 1440 8992 1454
rect 9006 1440 9058 1454
rect 9072 1440 9124 1454
rect 9138 1440 9190 1454
rect 9204 1440 9256 1454
rect 9270 1440 9322 1454
rect 9336 1440 9388 1454
rect 9402 1440 9454 1454
rect 9468 1440 9520 1454
rect 9534 1440 9586 1454
rect 9600 1440 9652 1454
rect 9666 1440 9718 1454
rect 9732 1440 9784 1454
rect 9798 1440 9850 1454
rect 9864 1440 9916 1454
rect 9930 1440 9982 1454
rect 9996 1440 10048 1454
rect 10062 1440 10114 1454
rect 10128 1440 10180 1454
rect 10194 1440 10246 1454
rect 10260 1440 10312 1454
rect 8741 1402 8793 1440
rect 8808 1402 8860 1440
rect 8874 1402 8926 1440
rect 8940 1402 8992 1440
rect 9006 1402 9058 1440
rect 9072 1402 9124 1440
rect 9138 1402 9190 1440
rect 9204 1402 9256 1440
rect 9270 1402 9322 1440
rect 9336 1402 9388 1440
rect 9402 1402 9454 1440
rect 9468 1402 9520 1440
rect 9534 1402 9586 1440
rect 9600 1402 9652 1440
rect 9666 1402 9718 1440
rect 9732 1402 9784 1440
rect 9798 1402 9850 1440
rect 9864 1402 9916 1440
rect 9930 1402 9982 1440
rect 9996 1402 10048 1440
rect 10062 1402 10114 1440
rect 10128 1402 10180 1440
rect 10194 1402 10246 1440
rect 10260 1402 10312 1440
rect 8741 1338 8793 1390
rect 8808 1338 8860 1390
rect 8874 1338 8926 1390
rect 8940 1338 8992 1390
rect 9006 1338 9058 1390
rect 9072 1338 9124 1390
rect 9138 1338 9190 1390
rect 9204 1338 9256 1390
rect 9270 1338 9322 1390
rect 9336 1338 9388 1390
rect 9402 1338 9454 1390
rect 9468 1338 9520 1390
rect 9534 1338 9586 1390
rect 9600 1338 9652 1390
rect 9666 1338 9718 1390
rect 9732 1338 9784 1390
rect 9798 1338 9850 1390
rect 9864 1338 9916 1390
rect 9930 1338 9982 1390
rect 9996 1338 10048 1390
rect 10062 1338 10114 1390
rect 10128 1338 10180 1390
rect 10194 1338 10246 1390
rect 10260 1338 10312 1390
rect 8030 1258 8082 1267
rect 8095 1258 8147 1267
rect 8030 1224 8046 1258
rect 8046 1224 8082 1258
rect 8095 1224 8120 1258
rect 8120 1224 8147 1258
rect 8030 1215 8082 1224
rect 8095 1215 8147 1224
rect 8159 1258 8211 1267
rect 8159 1224 8160 1258
rect 8160 1224 8194 1258
rect 8194 1224 8211 1258
rect 8159 1215 8211 1224
rect 8223 1258 8275 1267
rect 8223 1224 8234 1258
rect 8234 1224 8268 1258
rect 8268 1224 8275 1258
rect 8223 1215 8275 1224
rect 8287 1258 8339 1267
rect 8351 1258 8403 1267
rect 8415 1258 8467 1267
rect 8479 1258 8531 1267
rect 8543 1258 8595 1267
rect 8607 1258 8659 1267
rect 8287 1224 8308 1258
rect 8308 1224 8339 1258
rect 8351 1224 8382 1258
rect 8382 1224 8403 1258
rect 8415 1224 8416 1258
rect 8416 1224 8456 1258
rect 8456 1224 8467 1258
rect 8479 1224 8490 1258
rect 8490 1224 8529 1258
rect 8529 1224 8531 1258
rect 8543 1224 8563 1258
rect 8563 1224 8595 1258
rect 8607 1224 8636 1258
rect 8636 1224 8659 1258
rect 8287 1215 8339 1224
rect 8351 1215 8403 1224
rect 8415 1215 8467 1224
rect 8479 1215 8531 1224
rect 8543 1215 8595 1224
rect 8607 1215 8659 1224
rect 10458 1258 10510 1267
rect 10525 1258 10577 1267
rect 10591 1258 10643 1267
rect 10458 1224 10474 1258
rect 10474 1224 10510 1258
rect 10525 1224 10548 1258
rect 10548 1224 10577 1258
rect 10591 1224 10622 1258
rect 10622 1224 10643 1258
rect 10458 1215 10510 1224
rect 10525 1215 10577 1224
rect 10591 1215 10643 1224
rect 10657 1258 10709 1267
rect 10657 1224 10662 1258
rect 10662 1224 10696 1258
rect 10696 1224 10709 1258
rect 10657 1215 10709 1224
rect 10723 1258 10775 1267
rect 10723 1224 10736 1258
rect 10736 1224 10770 1258
rect 10770 1224 10775 1258
rect 10723 1215 10775 1224
rect 7322 1201 7374 1207
rect 7322 1167 7330 1201
rect 7330 1167 7364 1201
rect 7364 1167 7374 1201
rect 7322 1155 7374 1167
rect 7322 1127 7374 1141
rect 7322 1093 7330 1127
rect 7330 1093 7364 1127
rect 7364 1093 7374 1127
rect 11558 1201 11610 1207
rect 11558 1167 11566 1201
rect 11566 1167 11600 1201
rect 11600 1167 11610 1201
rect 11558 1155 11610 1167
rect 11558 1127 11610 1141
rect 7322 1089 7374 1093
rect 7322 1053 7374 1075
rect 8741 1102 8793 1111
rect 8741 1068 8748 1102
rect 8748 1068 8782 1102
rect 8782 1068 8793 1102
rect 8741 1059 8793 1068
rect 8806 1102 8858 1111
rect 8806 1068 8821 1102
rect 8821 1068 8855 1102
rect 8855 1068 8858 1102
rect 8806 1059 8858 1068
rect 8871 1102 8923 1111
rect 8936 1102 8988 1111
rect 9000 1102 9052 1111
rect 9064 1102 9116 1111
rect 9128 1102 9180 1111
rect 9192 1102 9244 1111
rect 8871 1068 8894 1102
rect 8894 1068 8923 1102
rect 8936 1068 8967 1102
rect 8967 1068 8988 1102
rect 9000 1068 9001 1102
rect 9001 1068 9040 1102
rect 9040 1068 9052 1102
rect 9064 1068 9074 1102
rect 9074 1068 9113 1102
rect 9113 1068 9116 1102
rect 9128 1068 9147 1102
rect 9147 1068 9180 1102
rect 9192 1068 9220 1102
rect 9220 1068 9244 1102
rect 8871 1059 8923 1068
rect 8936 1059 8988 1068
rect 9000 1059 9052 1068
rect 9064 1059 9116 1068
rect 9128 1059 9180 1068
rect 9192 1059 9244 1068
rect 9256 1102 9308 1111
rect 9256 1068 9259 1102
rect 9259 1068 9293 1102
rect 9293 1068 9308 1102
rect 9256 1059 9308 1068
rect 9320 1102 9372 1111
rect 9320 1068 9332 1102
rect 9332 1068 9366 1102
rect 9366 1068 9372 1102
rect 9320 1059 9372 1068
rect 9558 1102 9610 1111
rect 9558 1068 9564 1102
rect 9564 1068 9598 1102
rect 9598 1068 9610 1102
rect 9558 1059 9610 1068
rect 9628 1102 9680 1111
rect 9628 1068 9637 1102
rect 9637 1068 9671 1102
rect 9671 1068 9680 1102
rect 9628 1059 9680 1068
rect 9698 1102 9750 1111
rect 9698 1068 9710 1102
rect 9710 1068 9744 1102
rect 9744 1068 9750 1102
rect 9698 1059 9750 1068
rect 9768 1102 9820 1111
rect 9768 1068 9783 1102
rect 9783 1068 9817 1102
rect 9817 1068 9820 1102
rect 9768 1059 9820 1068
rect 9838 1102 9890 1111
rect 9838 1068 9856 1102
rect 9856 1068 9890 1102
rect 9838 1059 9890 1068
rect 9908 1102 9960 1111
rect 9978 1102 10030 1111
rect 10048 1102 10100 1111
rect 10118 1102 10170 1111
rect 10189 1102 10241 1111
rect 10260 1102 10312 1111
rect 9908 1068 9929 1102
rect 9929 1068 9960 1102
rect 9978 1068 10002 1102
rect 10002 1068 10030 1102
rect 10048 1068 10075 1102
rect 10075 1068 10100 1102
rect 10118 1068 10148 1102
rect 10148 1068 10170 1102
rect 10189 1068 10221 1102
rect 10221 1068 10241 1102
rect 10260 1068 10294 1102
rect 10294 1068 10312 1102
rect 9908 1059 9960 1068
rect 9978 1059 10030 1068
rect 10048 1059 10100 1068
rect 10118 1059 10170 1068
rect 10189 1059 10241 1068
rect 10260 1059 10312 1068
rect 11558 1093 11566 1127
rect 11566 1093 11600 1127
rect 11600 1093 11610 1127
rect 11558 1089 11610 1093
rect 7322 1023 7330 1053
rect 7330 1023 7364 1053
rect 7364 1023 7374 1053
rect 7322 979 7374 1009
rect 7322 957 7330 979
rect 7330 957 7364 979
rect 7364 957 7374 979
rect 11558 1053 11610 1075
rect 11558 1023 11566 1053
rect 11566 1023 11600 1053
rect 11600 1023 11610 1053
rect 11558 979 11610 1009
rect 11558 957 11566 979
rect 11566 957 11600 979
rect 11600 957 11610 979
rect 7322 905 7374 943
rect 8027 946 8079 955
rect 8092 946 8144 955
rect 8027 912 8046 946
rect 8046 912 8079 946
rect 8092 912 8120 946
rect 8120 912 8144 946
rect 7322 891 7330 905
rect 7330 891 7364 905
rect 7364 891 7374 905
rect 8027 903 8079 912
rect 8092 903 8144 912
rect 8156 946 8208 955
rect 8156 912 8160 946
rect 8160 912 8194 946
rect 8194 912 8208 946
rect 8156 903 8208 912
rect 8220 946 8272 955
rect 8220 912 8234 946
rect 8234 912 8268 946
rect 8268 912 8272 946
rect 8220 903 8272 912
rect 8284 946 8336 955
rect 8348 946 8400 955
rect 8412 946 8464 955
rect 8476 946 8528 955
rect 8540 946 8592 955
rect 8604 946 8656 955
rect 8284 912 8308 946
rect 8308 912 8336 946
rect 8348 912 8382 946
rect 8382 912 8400 946
rect 8412 912 8416 946
rect 8416 912 8456 946
rect 8456 912 8464 946
rect 8476 912 8490 946
rect 8490 912 8528 946
rect 8540 912 8563 946
rect 8563 912 8592 946
rect 8604 912 8636 946
rect 8636 912 8656 946
rect 8284 903 8336 912
rect 8348 903 8400 912
rect 8412 903 8464 912
rect 8476 903 8528 912
rect 8540 903 8592 912
rect 8604 903 8656 912
rect 10458 946 10510 955
rect 10525 946 10577 955
rect 10591 946 10643 955
rect 10458 912 10474 946
rect 10474 912 10510 946
rect 10525 912 10548 946
rect 10548 912 10577 946
rect 10591 912 10622 946
rect 10622 912 10643 946
rect 10458 903 10510 912
rect 10525 903 10577 912
rect 10591 903 10643 912
rect 10657 946 10709 955
rect 10657 912 10662 946
rect 10662 912 10696 946
rect 10696 912 10709 946
rect 10657 903 10709 912
rect 10723 946 10775 955
rect 10723 912 10736 946
rect 10736 912 10770 946
rect 10770 912 10775 946
rect 10723 903 10775 912
rect 11558 905 11610 943
rect 7322 871 7330 877
rect 7330 871 7364 877
rect 7364 871 7374 877
rect 7322 831 7374 871
rect 7322 825 7330 831
rect 7330 825 7364 831
rect 7364 825 7374 831
rect 7322 797 7330 811
rect 7330 797 7364 811
rect 7364 797 7374 811
rect 11558 891 11566 905
rect 11566 891 11600 905
rect 11600 891 11610 905
rect 11558 871 11566 877
rect 11566 871 11600 877
rect 11600 871 11610 877
rect 11558 831 11610 871
rect 11558 825 11566 831
rect 11566 825 11600 831
rect 11600 825 11610 831
rect 7322 759 7374 797
rect 8741 790 8793 799
rect 8741 756 8748 790
rect 8748 756 8782 790
rect 8782 756 8793 790
rect 8741 747 8793 756
rect 8806 790 8858 799
rect 8806 756 8821 790
rect 8821 756 8855 790
rect 8855 756 8858 790
rect 8806 747 8858 756
rect 8871 790 8923 799
rect 8936 790 8988 799
rect 9000 790 9052 799
rect 9064 790 9116 799
rect 9128 790 9180 799
rect 9192 790 9244 799
rect 8871 756 8894 790
rect 8894 756 8923 790
rect 8936 756 8967 790
rect 8967 756 8988 790
rect 9000 756 9001 790
rect 9001 756 9040 790
rect 9040 756 9052 790
rect 9064 756 9074 790
rect 9074 756 9113 790
rect 9113 756 9116 790
rect 9128 756 9147 790
rect 9147 756 9180 790
rect 9192 756 9220 790
rect 9220 756 9244 790
rect 8871 747 8923 756
rect 8936 747 8988 756
rect 9000 747 9052 756
rect 9064 747 9116 756
rect 9128 747 9180 756
rect 9192 747 9244 756
rect 9256 790 9308 799
rect 9256 756 9259 790
rect 9259 756 9293 790
rect 9293 756 9308 790
rect 9256 747 9308 756
rect 9320 790 9372 799
rect 9320 756 9332 790
rect 9332 756 9366 790
rect 9366 756 9372 790
rect 9320 747 9372 756
rect 9558 790 9610 799
rect 9558 756 9564 790
rect 9564 756 9598 790
rect 9598 756 9610 790
rect 9558 747 9610 756
rect 9628 790 9680 799
rect 9628 756 9637 790
rect 9637 756 9671 790
rect 9671 756 9680 790
rect 9628 747 9680 756
rect 9698 790 9750 799
rect 9698 756 9710 790
rect 9710 756 9744 790
rect 9744 756 9750 790
rect 9698 747 9750 756
rect 9768 790 9820 799
rect 9768 756 9783 790
rect 9783 756 9817 790
rect 9817 756 9820 790
rect 9768 747 9820 756
rect 9838 790 9890 799
rect 9838 756 9856 790
rect 9856 756 9890 790
rect 9838 747 9890 756
rect 9908 790 9960 799
rect 9978 790 10030 799
rect 10048 790 10100 799
rect 10118 790 10170 799
rect 10189 790 10241 799
rect 10260 790 10312 799
rect 11558 797 11566 811
rect 11566 797 11600 811
rect 11600 797 11610 811
rect 9908 756 9929 790
rect 9929 756 9960 790
rect 9978 756 10002 790
rect 10002 756 10030 790
rect 10048 756 10075 790
rect 10075 756 10100 790
rect 10118 756 10148 790
rect 10148 756 10170 790
rect 10189 756 10221 790
rect 10221 756 10241 790
rect 10260 756 10294 790
rect 10294 756 10312 790
rect 9908 747 9960 756
rect 9978 747 10030 756
rect 10048 747 10100 756
rect 10118 747 10170 756
rect 10189 747 10241 756
rect 10260 747 10312 756
rect 11558 759 11610 797
rect 7322 723 7330 745
rect 7330 723 7364 745
rect 7364 723 7374 745
rect 7322 693 7374 723
rect 7322 649 7330 679
rect 7330 649 7364 679
rect 7364 649 7374 679
rect 7322 627 7374 649
rect 11558 723 11566 745
rect 11566 723 11600 745
rect 11600 723 11610 745
rect 11558 693 11610 723
rect 11558 649 11566 679
rect 11566 649 11600 679
rect 11600 649 11610 679
rect 7322 609 7374 613
rect 7322 575 7330 609
rect 7330 575 7364 609
rect 7364 575 7374 609
rect 8027 634 8079 643
rect 8092 634 8144 643
rect 8027 600 8046 634
rect 8046 600 8079 634
rect 8092 600 8120 634
rect 8120 600 8144 634
rect 8027 591 8079 600
rect 8092 591 8144 600
rect 8156 634 8208 643
rect 8156 600 8160 634
rect 8160 600 8194 634
rect 8194 600 8208 634
rect 8156 591 8208 600
rect 8220 634 8272 643
rect 8220 600 8234 634
rect 8234 600 8268 634
rect 8268 600 8272 634
rect 8220 591 8272 600
rect 8284 634 8336 643
rect 8348 634 8400 643
rect 8412 634 8464 643
rect 8476 634 8528 643
rect 8540 634 8592 643
rect 8604 634 8656 643
rect 8284 600 8308 634
rect 8308 600 8336 634
rect 8348 600 8382 634
rect 8382 600 8400 634
rect 8412 600 8416 634
rect 8416 600 8456 634
rect 8456 600 8464 634
rect 8476 600 8490 634
rect 8490 600 8528 634
rect 8540 600 8563 634
rect 8563 600 8592 634
rect 8604 600 8636 634
rect 8636 600 8656 634
rect 8284 591 8336 600
rect 8348 591 8400 600
rect 8412 591 8464 600
rect 8476 591 8528 600
rect 8540 591 8592 600
rect 8604 591 8656 600
rect 10458 634 10510 643
rect 10525 634 10577 643
rect 10591 634 10643 643
rect 10458 600 10474 634
rect 10474 600 10510 634
rect 10525 600 10548 634
rect 10548 600 10577 634
rect 10591 600 10622 634
rect 10622 600 10643 634
rect 10458 591 10510 600
rect 10525 591 10577 600
rect 10591 591 10643 600
rect 10657 634 10709 643
rect 10657 600 10662 634
rect 10662 600 10696 634
rect 10696 600 10709 634
rect 10657 591 10709 600
rect 10723 634 10775 643
rect 10723 600 10736 634
rect 10736 600 10770 634
rect 10770 600 10775 634
rect 10723 591 10775 600
rect 11558 627 11610 649
rect 11558 609 11610 613
rect 7322 561 7374 575
rect 7322 535 7374 547
rect 7322 501 7330 535
rect 7330 501 7364 535
rect 7364 501 7374 535
rect 7322 495 7374 501
rect 11558 575 11566 609
rect 11566 575 11600 609
rect 11600 575 11610 609
rect 11558 561 11610 575
rect 11558 535 11610 547
rect 11558 501 11566 535
rect 11566 501 11600 535
rect 11600 501 11610 535
rect 11558 495 11610 501
rect 8741 478 8793 487
rect 8741 444 8748 478
rect 8748 444 8782 478
rect 8782 444 8793 478
rect 8741 435 8793 444
rect 8806 478 8858 487
rect 8806 444 8821 478
rect 8821 444 8855 478
rect 8855 444 8858 478
rect 8806 435 8858 444
rect 8871 478 8923 487
rect 8936 478 8988 487
rect 9000 478 9052 487
rect 9064 478 9116 487
rect 9128 478 9180 487
rect 9192 478 9244 487
rect 8871 444 8894 478
rect 8894 444 8923 478
rect 8936 444 8967 478
rect 8967 444 8988 478
rect 9000 444 9001 478
rect 9001 444 9040 478
rect 9040 444 9052 478
rect 9064 444 9074 478
rect 9074 444 9113 478
rect 9113 444 9116 478
rect 9128 444 9147 478
rect 9147 444 9180 478
rect 9192 444 9220 478
rect 9220 444 9244 478
rect 8871 435 8923 444
rect 8936 435 8988 444
rect 9000 435 9052 444
rect 9064 435 9116 444
rect 9128 435 9180 444
rect 9192 435 9244 444
rect 9256 478 9308 487
rect 9256 444 9259 478
rect 9259 444 9293 478
rect 9293 444 9308 478
rect 9256 435 9308 444
rect 9320 478 9372 487
rect 9320 444 9332 478
rect 9332 444 9366 478
rect 9366 444 9372 478
rect 9320 435 9372 444
rect 9558 478 9610 487
rect 9558 444 9564 478
rect 9564 444 9598 478
rect 9598 444 9610 478
rect 9558 435 9610 444
rect 9628 478 9680 487
rect 9628 444 9637 478
rect 9637 444 9671 478
rect 9671 444 9680 478
rect 9628 435 9680 444
rect 9698 478 9750 487
rect 9698 444 9710 478
rect 9710 444 9744 478
rect 9744 444 9750 478
rect 9698 435 9750 444
rect 9768 478 9820 487
rect 9768 444 9783 478
rect 9783 444 9817 478
rect 9817 444 9820 478
rect 9768 435 9820 444
rect 9838 478 9890 487
rect 9838 444 9856 478
rect 9856 444 9890 478
rect 9838 435 9890 444
rect 9908 478 9960 487
rect 9978 478 10030 487
rect 10048 478 10100 487
rect 10118 478 10170 487
rect 10189 478 10241 487
rect 10260 478 10312 487
rect 9908 444 9929 478
rect 9929 444 9960 478
rect 9978 444 10002 478
rect 10002 444 10030 478
rect 10048 444 10075 478
rect 10075 444 10100 478
rect 10118 444 10148 478
rect 10148 444 10170 478
rect 10189 444 10221 478
rect 10221 444 10241 478
rect 10260 444 10294 478
rect 10294 444 10312 478
rect 9908 435 9960 444
rect 9978 435 10030 444
rect 10048 435 10100 444
rect 10118 435 10170 444
rect 10189 435 10241 444
rect 10260 435 10312 444
rect 8741 358 8793 383
rect 8808 358 8860 383
rect 8874 358 8926 383
rect 8940 358 8992 383
rect 9006 358 9058 383
rect 9072 358 9124 383
rect 9138 358 9190 383
rect 9204 358 9256 383
rect 9270 358 9322 383
rect 9336 358 9388 383
rect 9402 358 9454 383
rect 9468 358 9520 383
rect 9534 358 9586 383
rect 9600 358 9652 383
rect 9666 358 9718 383
rect 9732 358 9784 383
rect 9798 358 9850 383
rect 9864 358 9916 383
rect 9930 358 9982 383
rect 9996 358 10048 383
rect 10062 358 10114 383
rect 10128 358 10180 383
rect 10194 358 10246 383
rect 10260 358 10312 383
rect 8741 331 8793 358
rect 8808 331 8860 358
rect 8874 331 8926 358
rect 8940 331 8992 358
rect 9006 331 9058 358
rect 9072 331 9124 358
rect 9138 331 9190 358
rect 9204 331 9256 358
rect 9270 331 9322 358
rect 9336 331 9388 358
rect 9402 331 9454 358
rect 9468 331 9520 358
rect 9534 331 9586 358
rect 9600 331 9652 358
rect 9666 331 9718 358
rect 9732 331 9784 358
rect 9798 331 9850 358
rect 9864 331 9916 358
rect 9930 331 9982 358
rect 9996 331 10048 358
rect 10062 331 10114 358
rect 10128 331 10180 358
rect 10194 331 10246 358
rect 10260 331 10312 358
rect 7163 214 7215 266
rect 7229 252 7235 266
rect 7235 252 7269 266
rect 7269 252 7281 266
rect 7229 214 7281 252
rect 7295 252 7308 266
rect 7308 252 7342 266
rect 7342 252 7347 266
rect 7295 214 7347 252
rect 7361 252 7381 266
rect 7381 252 7413 266
rect 7426 252 7454 266
rect 7454 252 7478 266
rect 7491 252 7527 266
rect 7527 252 7543 266
rect 7556 252 7561 266
rect 7561 252 7600 266
rect 7600 252 7608 266
rect 7621 252 7634 266
rect 7634 252 7673 266
rect 7686 252 7707 266
rect 7707 252 7738 266
rect 7751 252 7780 266
rect 7780 252 7803 266
rect 7361 214 7413 252
rect 7426 214 7478 252
rect 7491 214 7543 252
rect 7556 214 7608 252
rect 7621 214 7673 252
rect 7686 214 7738 252
rect 7751 214 7803 252
rect 7816 252 7819 266
rect 7819 252 7853 266
rect 7853 252 7868 266
rect 7816 214 7868 252
rect 7881 252 7892 266
rect 7892 252 7926 266
rect 7926 252 7933 266
rect 7881 214 7933 252
rect 7946 252 7965 266
rect 7965 252 7998 266
rect 8011 252 8038 266
rect 8038 252 8063 266
rect 8076 252 8111 266
rect 8111 252 8128 266
rect 8741 267 8793 319
rect 8808 267 8860 319
rect 8874 267 8926 319
rect 8940 267 8992 319
rect 9006 267 9058 319
rect 9072 267 9124 319
rect 9138 267 9190 319
rect 9204 267 9256 319
rect 9270 267 9322 319
rect 9336 267 9388 319
rect 9402 267 9454 319
rect 9468 267 9520 319
rect 9534 267 9586 319
rect 9600 267 9652 319
rect 9666 267 9718 319
rect 9732 267 9784 319
rect 9798 267 9850 319
rect 9864 267 9916 319
rect 9930 267 9982 319
rect 9996 267 10048 319
rect 10062 267 10114 319
rect 10128 267 10180 319
rect 10194 267 10246 319
rect 10260 267 10312 319
rect 7946 214 7998 252
rect 8011 214 8063 252
rect 8076 214 8128 252
rect 10880 171 10932 175
rect 10946 171 10998 175
rect 11012 171 11064 175
rect 11078 171 11130 175
rect 10880 123 10932 171
rect 10946 123 10998 171
rect 11012 123 11064 171
rect 11078 123 11130 171
rect -79 -236 -27 -184
rect -15 -236 37 -184
rect -79 -304 -27 -252
rect -15 -304 37 -252
rect 6646 -1270 6698 -1261
rect 6646 -1304 6652 -1270
rect 6652 -1304 6686 -1270
rect 6686 -1304 6698 -1270
rect 6646 -1313 6698 -1304
rect 6711 -1270 6763 -1261
rect 6711 -1304 6727 -1270
rect 6727 -1304 6761 -1270
rect 6761 -1304 6763 -1270
rect 6711 -1313 6763 -1304
rect 6776 -1270 6828 -1261
rect 6841 -1270 6893 -1261
rect 6906 -1270 6958 -1261
rect 6971 -1270 7023 -1261
rect 7036 -1270 7088 -1261
rect 6776 -1304 6802 -1270
rect 6802 -1304 6828 -1270
rect 6841 -1304 6877 -1270
rect 6877 -1304 6893 -1270
rect 6906 -1304 6911 -1270
rect 6911 -1304 6952 -1270
rect 6952 -1304 6958 -1270
rect 6971 -1304 6986 -1270
rect 6986 -1304 7023 -1270
rect 7036 -1304 7061 -1270
rect 7061 -1304 7088 -1270
rect 6776 -1313 6828 -1304
rect 6841 -1313 6893 -1304
rect 6906 -1313 6958 -1304
rect 6971 -1313 7023 -1304
rect 7036 -1313 7088 -1304
rect 7101 -1270 7153 -1261
rect 7101 -1304 7102 -1270
rect 7102 -1304 7136 -1270
rect 7136 -1304 7153 -1270
rect 7101 -1313 7153 -1304
rect 7165 -1270 7217 -1261
rect 7165 -1304 7177 -1270
rect 7177 -1304 7211 -1270
rect 7211 -1304 7217 -1270
rect 7165 -1313 7217 -1304
rect 7229 -1270 7281 -1261
rect 7293 -1270 7345 -1261
rect 7357 -1270 7409 -1261
rect 7421 -1270 7473 -1261
rect 7485 -1270 7537 -1261
rect 7229 -1304 7252 -1270
rect 7252 -1304 7281 -1270
rect 7293 -1304 7327 -1270
rect 7327 -1304 7345 -1270
rect 7357 -1304 7361 -1270
rect 7361 -1304 7402 -1270
rect 7402 -1304 7409 -1270
rect 7421 -1304 7436 -1270
rect 7436 -1304 7473 -1270
rect 7485 -1304 7510 -1270
rect 7510 -1304 7537 -1270
rect 7229 -1313 7281 -1304
rect 7293 -1313 7345 -1304
rect 7357 -1313 7409 -1304
rect 7421 -1313 7473 -1304
rect 7485 -1313 7537 -1304
rect 7549 -1270 7601 -1261
rect 7549 -1304 7550 -1270
rect 7550 -1304 7584 -1270
rect 7584 -1304 7601 -1270
rect 7549 -1313 7601 -1304
rect 7613 -1270 7665 -1261
rect 7613 -1304 7624 -1270
rect 7624 -1304 7658 -1270
rect 7658 -1304 7665 -1270
rect 7613 -1313 7665 -1304
rect 7677 -1270 7729 -1261
rect 7741 -1270 7793 -1261
rect 7805 -1270 7857 -1261
rect 7869 -1270 7921 -1261
rect 7933 -1270 7985 -1261
rect 7997 -1270 8049 -1261
rect 7677 -1304 7698 -1270
rect 7698 -1304 7729 -1270
rect 7741 -1304 7772 -1270
rect 7772 -1304 7793 -1270
rect 7805 -1304 7806 -1270
rect 7806 -1304 7846 -1270
rect 7846 -1304 7857 -1270
rect 7869 -1304 7880 -1270
rect 7880 -1304 7920 -1270
rect 7920 -1304 7921 -1270
rect 7933 -1304 7954 -1270
rect 7954 -1304 7985 -1270
rect 7997 -1304 8028 -1270
rect 8028 -1304 8049 -1270
rect 7677 -1313 7729 -1304
rect 7741 -1313 7793 -1304
rect 7805 -1313 7857 -1304
rect 7869 -1313 7921 -1304
rect 7933 -1313 7985 -1304
rect 7997 -1313 8049 -1304
rect 8061 -1270 8113 -1261
rect 8061 -1304 8068 -1270
rect 8068 -1304 8102 -1270
rect 8102 -1304 8113 -1270
rect 8061 -1313 8113 -1304
rect 8125 -1270 8177 -1261
rect 8125 -1304 8142 -1270
rect 8142 -1304 8176 -1270
rect 8176 -1304 8177 -1270
rect 8125 -1313 8177 -1304
rect 8189 -1270 8241 -1261
rect 8253 -1270 8305 -1261
rect 8317 -1270 8369 -1261
rect 8381 -1270 8433 -1261
rect 8445 -1270 8497 -1261
rect 8189 -1304 8216 -1270
rect 8216 -1304 8241 -1270
rect 8253 -1304 8290 -1270
rect 8290 -1304 8305 -1270
rect 8317 -1304 8324 -1270
rect 8324 -1304 8364 -1270
rect 8364 -1304 8369 -1270
rect 8381 -1304 8398 -1270
rect 8398 -1304 8433 -1270
rect 8445 -1304 8472 -1270
rect 8472 -1304 8497 -1270
rect 8189 -1313 8241 -1304
rect 8253 -1313 8305 -1304
rect 8317 -1313 8369 -1304
rect 8381 -1313 8433 -1304
rect 8445 -1313 8497 -1304
rect 8509 -1270 8561 -1261
rect 8509 -1304 8512 -1270
rect 8512 -1304 8546 -1270
rect 8546 -1304 8561 -1270
rect 8509 -1313 8561 -1304
rect 8573 -1270 8625 -1261
rect 8573 -1304 8586 -1270
rect 8586 -1304 8620 -1270
rect 8620 -1304 8625 -1270
rect 8573 -1313 8625 -1304
rect 6522 -1327 6574 -1321
rect 6522 -1361 6534 -1327
rect 6534 -1361 6568 -1327
rect 6568 -1361 6574 -1327
rect 6522 -1373 6574 -1361
rect 6522 -1399 6574 -1385
rect 6522 -1433 6534 -1399
rect 6534 -1433 6568 -1399
rect 6568 -1433 6574 -1399
rect 6522 -1437 6574 -1433
rect 6646 -1426 6698 -1417
rect 6646 -1460 6652 -1426
rect 6652 -1460 6686 -1426
rect 6686 -1460 6698 -1426
rect 6646 -1469 6698 -1460
rect 6711 -1426 6763 -1417
rect 6711 -1460 6727 -1426
rect 6727 -1460 6761 -1426
rect 6761 -1460 6763 -1426
rect 6711 -1469 6763 -1460
rect 6776 -1426 6828 -1417
rect 6841 -1426 6893 -1417
rect 6906 -1426 6958 -1417
rect 6971 -1426 7023 -1417
rect 7036 -1426 7088 -1417
rect 6776 -1460 6802 -1426
rect 6802 -1460 6828 -1426
rect 6841 -1460 6877 -1426
rect 6877 -1460 6893 -1426
rect 6906 -1460 6911 -1426
rect 6911 -1460 6952 -1426
rect 6952 -1460 6958 -1426
rect 6971 -1460 6986 -1426
rect 6986 -1460 7023 -1426
rect 7036 -1460 7061 -1426
rect 7061 -1460 7088 -1426
rect 6776 -1469 6828 -1460
rect 6841 -1469 6893 -1460
rect 6906 -1469 6958 -1460
rect 6971 -1469 7023 -1460
rect 7036 -1469 7088 -1460
rect 7101 -1426 7153 -1417
rect 7101 -1460 7102 -1426
rect 7102 -1460 7136 -1426
rect 7136 -1460 7153 -1426
rect 7101 -1469 7153 -1460
rect 7165 -1426 7217 -1417
rect 7165 -1460 7177 -1426
rect 7177 -1460 7211 -1426
rect 7211 -1460 7217 -1426
rect 7165 -1469 7217 -1460
rect 7229 -1426 7281 -1417
rect 7293 -1426 7345 -1417
rect 7357 -1426 7409 -1417
rect 7421 -1426 7473 -1417
rect 7485 -1426 7537 -1417
rect 7229 -1460 7252 -1426
rect 7252 -1460 7281 -1426
rect 7293 -1460 7327 -1426
rect 7327 -1460 7345 -1426
rect 7357 -1460 7361 -1426
rect 7361 -1460 7402 -1426
rect 7402 -1460 7409 -1426
rect 7421 -1460 7436 -1426
rect 7436 -1460 7473 -1426
rect 7485 -1460 7510 -1426
rect 7510 -1460 7537 -1426
rect 7229 -1469 7281 -1460
rect 7293 -1469 7345 -1460
rect 7357 -1469 7409 -1460
rect 7421 -1469 7473 -1460
rect 7485 -1469 7537 -1460
rect 7549 -1426 7601 -1417
rect 7549 -1460 7550 -1426
rect 7550 -1460 7584 -1426
rect 7584 -1460 7601 -1426
rect 7549 -1469 7601 -1460
rect 7613 -1426 7665 -1417
rect 7613 -1460 7624 -1426
rect 7624 -1460 7658 -1426
rect 7658 -1460 7665 -1426
rect 7613 -1469 7665 -1460
rect 7677 -1426 7729 -1417
rect 7741 -1426 7793 -1417
rect 7805 -1426 7857 -1417
rect 7869 -1426 7921 -1417
rect 7933 -1426 7985 -1417
rect 7997 -1426 8049 -1417
rect 7677 -1460 7698 -1426
rect 7698 -1460 7729 -1426
rect 7741 -1460 7772 -1426
rect 7772 -1460 7793 -1426
rect 7805 -1460 7806 -1426
rect 7806 -1460 7846 -1426
rect 7846 -1460 7857 -1426
rect 7869 -1460 7880 -1426
rect 7880 -1460 7920 -1426
rect 7920 -1460 7921 -1426
rect 7933 -1460 7954 -1426
rect 7954 -1460 7985 -1426
rect 7997 -1460 8028 -1426
rect 8028 -1460 8049 -1426
rect 7677 -1469 7729 -1460
rect 7741 -1469 7793 -1460
rect 7805 -1469 7857 -1460
rect 7869 -1469 7921 -1460
rect 7933 -1469 7985 -1460
rect 7997 -1469 8049 -1460
rect 8061 -1426 8113 -1417
rect 8061 -1460 8068 -1426
rect 8068 -1460 8102 -1426
rect 8102 -1460 8113 -1426
rect 8061 -1469 8113 -1460
rect 8125 -1426 8177 -1417
rect 8125 -1460 8142 -1426
rect 8142 -1460 8176 -1426
rect 8176 -1460 8177 -1426
rect 8125 -1469 8177 -1460
rect 8189 -1426 8241 -1417
rect 8253 -1426 8305 -1417
rect 8317 -1426 8369 -1417
rect 8381 -1426 8433 -1417
rect 8445 -1426 8497 -1417
rect 8189 -1460 8216 -1426
rect 8216 -1460 8241 -1426
rect 8253 -1460 8290 -1426
rect 8290 -1460 8305 -1426
rect 8317 -1460 8324 -1426
rect 8324 -1460 8364 -1426
rect 8364 -1460 8369 -1426
rect 8381 -1460 8398 -1426
rect 8398 -1460 8433 -1426
rect 8445 -1460 8472 -1426
rect 8472 -1460 8497 -1426
rect 8189 -1469 8241 -1460
rect 8253 -1469 8305 -1460
rect 8317 -1469 8369 -1460
rect 8381 -1469 8433 -1460
rect 8445 -1469 8497 -1460
rect 8509 -1426 8561 -1417
rect 8509 -1460 8512 -1426
rect 8512 -1460 8546 -1426
rect 8546 -1460 8561 -1426
rect 8509 -1469 8561 -1460
rect 8573 -1426 8625 -1417
rect 8573 -1460 8586 -1426
rect 8586 -1460 8620 -1426
rect 8620 -1460 8625 -1426
rect 8573 -1469 8625 -1460
rect 6646 -1582 6698 -1573
rect 6646 -1616 6652 -1582
rect 6652 -1616 6686 -1582
rect 6686 -1616 6698 -1582
rect 6646 -1625 6698 -1616
rect 6711 -1582 6763 -1573
rect 6711 -1616 6727 -1582
rect 6727 -1616 6761 -1582
rect 6761 -1616 6763 -1582
rect 6711 -1625 6763 -1616
rect 6776 -1582 6828 -1573
rect 6841 -1582 6893 -1573
rect 6906 -1582 6958 -1573
rect 6971 -1582 7023 -1573
rect 7036 -1582 7088 -1573
rect 6776 -1616 6802 -1582
rect 6802 -1616 6828 -1582
rect 6841 -1616 6877 -1582
rect 6877 -1616 6893 -1582
rect 6906 -1616 6911 -1582
rect 6911 -1616 6952 -1582
rect 6952 -1616 6958 -1582
rect 6971 -1616 6986 -1582
rect 6986 -1616 7023 -1582
rect 7036 -1616 7061 -1582
rect 7061 -1616 7088 -1582
rect 6776 -1625 6828 -1616
rect 6841 -1625 6893 -1616
rect 6906 -1625 6958 -1616
rect 6971 -1625 7023 -1616
rect 7036 -1625 7088 -1616
rect 7101 -1582 7153 -1573
rect 7101 -1616 7102 -1582
rect 7102 -1616 7136 -1582
rect 7136 -1616 7153 -1582
rect 7101 -1625 7153 -1616
rect 7165 -1582 7217 -1573
rect 7165 -1616 7177 -1582
rect 7177 -1616 7211 -1582
rect 7211 -1616 7217 -1582
rect 7165 -1625 7217 -1616
rect 7229 -1582 7281 -1573
rect 7293 -1582 7345 -1573
rect 7357 -1582 7409 -1573
rect 7421 -1582 7473 -1573
rect 7485 -1582 7537 -1573
rect 7229 -1616 7252 -1582
rect 7252 -1616 7281 -1582
rect 7293 -1616 7327 -1582
rect 7327 -1616 7345 -1582
rect 7357 -1616 7361 -1582
rect 7361 -1616 7402 -1582
rect 7402 -1616 7409 -1582
rect 7421 -1616 7436 -1582
rect 7436 -1616 7473 -1582
rect 7485 -1616 7510 -1582
rect 7510 -1616 7537 -1582
rect 7229 -1625 7281 -1616
rect 7293 -1625 7345 -1616
rect 7357 -1625 7409 -1616
rect 7421 -1625 7473 -1616
rect 7485 -1625 7537 -1616
rect 7549 -1582 7601 -1573
rect 7549 -1616 7550 -1582
rect 7550 -1616 7584 -1582
rect 7584 -1616 7601 -1582
rect 7549 -1625 7601 -1616
rect 7613 -1582 7665 -1573
rect 7613 -1616 7624 -1582
rect 7624 -1616 7658 -1582
rect 7658 -1616 7665 -1582
rect 7613 -1625 7665 -1616
rect 7677 -1582 7729 -1573
rect 7741 -1582 7793 -1573
rect 7805 -1582 7857 -1573
rect 7869 -1582 7921 -1573
rect 7933 -1582 7985 -1573
rect 7997 -1582 8049 -1573
rect 7677 -1616 7698 -1582
rect 7698 -1616 7729 -1582
rect 7741 -1616 7772 -1582
rect 7772 -1616 7793 -1582
rect 7805 -1616 7806 -1582
rect 7806 -1616 7846 -1582
rect 7846 -1616 7857 -1582
rect 7869 -1616 7880 -1582
rect 7880 -1616 7920 -1582
rect 7920 -1616 7921 -1582
rect 7933 -1616 7954 -1582
rect 7954 -1616 7985 -1582
rect 7997 -1616 8028 -1582
rect 8028 -1616 8049 -1582
rect 7677 -1625 7729 -1616
rect 7741 -1625 7793 -1616
rect 7805 -1625 7857 -1616
rect 7869 -1625 7921 -1616
rect 7933 -1625 7985 -1616
rect 7997 -1625 8049 -1616
rect 8061 -1582 8113 -1573
rect 8061 -1616 8068 -1582
rect 8068 -1616 8102 -1582
rect 8102 -1616 8113 -1582
rect 8061 -1625 8113 -1616
rect 8125 -1582 8177 -1573
rect 8125 -1616 8142 -1582
rect 8142 -1616 8176 -1582
rect 8176 -1616 8177 -1582
rect 8125 -1625 8177 -1616
rect 8189 -1582 8241 -1573
rect 8253 -1582 8305 -1573
rect 8317 -1582 8369 -1573
rect 8381 -1582 8433 -1573
rect 8445 -1582 8497 -1573
rect 8189 -1616 8216 -1582
rect 8216 -1616 8241 -1582
rect 8253 -1616 8290 -1582
rect 8290 -1616 8305 -1582
rect 8317 -1616 8324 -1582
rect 8324 -1616 8364 -1582
rect 8364 -1616 8369 -1582
rect 8381 -1616 8398 -1582
rect 8398 -1616 8433 -1582
rect 8445 -1616 8472 -1582
rect 8472 -1616 8497 -1582
rect 8189 -1625 8241 -1616
rect 8253 -1625 8305 -1616
rect 8317 -1625 8369 -1616
rect 8381 -1625 8433 -1616
rect 8445 -1625 8497 -1616
rect 8509 -1582 8561 -1573
rect 8509 -1616 8512 -1582
rect 8512 -1616 8546 -1582
rect 8546 -1616 8561 -1582
rect 8509 -1625 8561 -1616
rect 8573 -1582 8625 -1573
rect 8573 -1616 8586 -1582
rect 8586 -1616 8620 -1582
rect 8620 -1616 8625 -1582
rect 8573 -1625 8625 -1616
rect 6646 -1738 6698 -1729
rect 6646 -1772 6652 -1738
rect 6652 -1772 6686 -1738
rect 6686 -1772 6698 -1738
rect 6646 -1781 6698 -1772
rect 6711 -1738 6763 -1729
rect 6711 -1772 6727 -1738
rect 6727 -1772 6761 -1738
rect 6761 -1772 6763 -1738
rect 6711 -1781 6763 -1772
rect 6776 -1738 6828 -1729
rect 6841 -1738 6893 -1729
rect 6906 -1738 6958 -1729
rect 6971 -1738 7023 -1729
rect 7036 -1738 7088 -1729
rect 6776 -1772 6802 -1738
rect 6802 -1772 6828 -1738
rect 6841 -1772 6877 -1738
rect 6877 -1772 6893 -1738
rect 6906 -1772 6911 -1738
rect 6911 -1772 6952 -1738
rect 6952 -1772 6958 -1738
rect 6971 -1772 6986 -1738
rect 6986 -1772 7023 -1738
rect 7036 -1772 7061 -1738
rect 7061 -1772 7088 -1738
rect 6776 -1781 6828 -1772
rect 6841 -1781 6893 -1772
rect 6906 -1781 6958 -1772
rect 6971 -1781 7023 -1772
rect 7036 -1781 7088 -1772
rect 7101 -1738 7153 -1729
rect 7101 -1772 7102 -1738
rect 7102 -1772 7136 -1738
rect 7136 -1772 7153 -1738
rect 7101 -1781 7153 -1772
rect 7165 -1738 7217 -1729
rect 7165 -1772 7177 -1738
rect 7177 -1772 7211 -1738
rect 7211 -1772 7217 -1738
rect 7165 -1781 7217 -1772
rect 7229 -1738 7281 -1729
rect 7293 -1738 7345 -1729
rect 7357 -1738 7409 -1729
rect 7421 -1738 7473 -1729
rect 7485 -1738 7537 -1729
rect 7229 -1772 7252 -1738
rect 7252 -1772 7281 -1738
rect 7293 -1772 7327 -1738
rect 7327 -1772 7345 -1738
rect 7357 -1772 7361 -1738
rect 7361 -1772 7402 -1738
rect 7402 -1772 7409 -1738
rect 7421 -1772 7436 -1738
rect 7436 -1772 7473 -1738
rect 7485 -1772 7510 -1738
rect 7510 -1772 7537 -1738
rect 7229 -1781 7281 -1772
rect 7293 -1781 7345 -1772
rect 7357 -1781 7409 -1772
rect 7421 -1781 7473 -1772
rect 7485 -1781 7537 -1772
rect 7549 -1738 7601 -1729
rect 7549 -1772 7550 -1738
rect 7550 -1772 7584 -1738
rect 7584 -1772 7601 -1738
rect 7549 -1781 7601 -1772
rect 7613 -1738 7665 -1729
rect 7613 -1772 7624 -1738
rect 7624 -1772 7658 -1738
rect 7658 -1772 7665 -1738
rect 7613 -1781 7665 -1772
rect 7677 -1738 7729 -1729
rect 7741 -1738 7793 -1729
rect 7805 -1738 7857 -1729
rect 7869 -1738 7921 -1729
rect 7933 -1738 7985 -1729
rect 7997 -1738 8049 -1729
rect 7677 -1772 7698 -1738
rect 7698 -1772 7729 -1738
rect 7741 -1772 7772 -1738
rect 7772 -1772 7793 -1738
rect 7805 -1772 7806 -1738
rect 7806 -1772 7846 -1738
rect 7846 -1772 7857 -1738
rect 7869 -1772 7880 -1738
rect 7880 -1772 7920 -1738
rect 7920 -1772 7921 -1738
rect 7933 -1772 7954 -1738
rect 7954 -1772 7985 -1738
rect 7997 -1772 8028 -1738
rect 8028 -1772 8049 -1738
rect 7677 -1781 7729 -1772
rect 7741 -1781 7793 -1772
rect 7805 -1781 7857 -1772
rect 7869 -1781 7921 -1772
rect 7933 -1781 7985 -1772
rect 7997 -1781 8049 -1772
rect 8061 -1738 8113 -1729
rect 8061 -1772 8068 -1738
rect 8068 -1772 8102 -1738
rect 8102 -1772 8113 -1738
rect 8061 -1781 8113 -1772
rect 8125 -1738 8177 -1729
rect 8125 -1772 8142 -1738
rect 8142 -1772 8176 -1738
rect 8176 -1772 8177 -1738
rect 8125 -1781 8177 -1772
rect 8189 -1738 8241 -1729
rect 8253 -1738 8305 -1729
rect 8317 -1738 8369 -1729
rect 8381 -1738 8433 -1729
rect 8445 -1738 8497 -1729
rect 8189 -1772 8216 -1738
rect 8216 -1772 8241 -1738
rect 8253 -1772 8290 -1738
rect 8290 -1772 8305 -1738
rect 8317 -1772 8324 -1738
rect 8324 -1772 8364 -1738
rect 8364 -1772 8369 -1738
rect 8381 -1772 8398 -1738
rect 8398 -1772 8433 -1738
rect 8445 -1772 8472 -1738
rect 8472 -1772 8497 -1738
rect 8189 -1781 8241 -1772
rect 8253 -1781 8305 -1772
rect 8317 -1781 8369 -1772
rect 8381 -1781 8433 -1772
rect 8445 -1781 8497 -1772
rect 8509 -1738 8561 -1729
rect 8509 -1772 8512 -1738
rect 8512 -1772 8546 -1738
rect 8546 -1772 8561 -1738
rect 8509 -1781 8561 -1772
rect 8573 -1738 8625 -1729
rect 8573 -1772 8586 -1738
rect 8586 -1772 8620 -1738
rect 8620 -1772 8625 -1738
rect 8573 -1781 8625 -1772
rect 6646 -1894 6698 -1885
rect 6646 -1928 6652 -1894
rect 6652 -1928 6686 -1894
rect 6686 -1928 6698 -1894
rect 6646 -1937 6698 -1928
rect 6711 -1894 6763 -1885
rect 6711 -1928 6727 -1894
rect 6727 -1928 6761 -1894
rect 6761 -1928 6763 -1894
rect 6711 -1937 6763 -1928
rect 6776 -1894 6828 -1885
rect 6841 -1894 6893 -1885
rect 6906 -1894 6958 -1885
rect 6971 -1894 7023 -1885
rect 7036 -1894 7088 -1885
rect 6776 -1928 6802 -1894
rect 6802 -1928 6828 -1894
rect 6841 -1928 6877 -1894
rect 6877 -1928 6893 -1894
rect 6906 -1928 6911 -1894
rect 6911 -1928 6952 -1894
rect 6952 -1928 6958 -1894
rect 6971 -1928 6986 -1894
rect 6986 -1928 7023 -1894
rect 7036 -1928 7061 -1894
rect 7061 -1928 7088 -1894
rect 6776 -1937 6828 -1928
rect 6841 -1937 6893 -1928
rect 6906 -1937 6958 -1928
rect 6971 -1937 7023 -1928
rect 7036 -1937 7088 -1928
rect 7101 -1894 7153 -1885
rect 7101 -1928 7102 -1894
rect 7102 -1928 7136 -1894
rect 7136 -1928 7153 -1894
rect 7101 -1937 7153 -1928
rect 7165 -1894 7217 -1885
rect 7165 -1928 7177 -1894
rect 7177 -1928 7211 -1894
rect 7211 -1928 7217 -1894
rect 7165 -1937 7217 -1928
rect 7229 -1894 7281 -1885
rect 7293 -1894 7345 -1885
rect 7357 -1894 7409 -1885
rect 7421 -1894 7473 -1885
rect 7485 -1894 7537 -1885
rect 7229 -1928 7252 -1894
rect 7252 -1928 7281 -1894
rect 7293 -1928 7327 -1894
rect 7327 -1928 7345 -1894
rect 7357 -1928 7361 -1894
rect 7361 -1928 7402 -1894
rect 7402 -1928 7409 -1894
rect 7421 -1928 7436 -1894
rect 7436 -1928 7473 -1894
rect 7485 -1928 7510 -1894
rect 7510 -1928 7537 -1894
rect 7229 -1937 7281 -1928
rect 7293 -1937 7345 -1928
rect 7357 -1937 7409 -1928
rect 7421 -1937 7473 -1928
rect 7485 -1937 7537 -1928
rect 7549 -1894 7601 -1885
rect 7549 -1928 7550 -1894
rect 7550 -1928 7584 -1894
rect 7584 -1928 7601 -1894
rect 7549 -1937 7601 -1928
rect 7613 -1894 7665 -1885
rect 7613 -1928 7624 -1894
rect 7624 -1928 7658 -1894
rect 7658 -1928 7665 -1894
rect 7613 -1937 7665 -1928
rect 7677 -1894 7729 -1885
rect 7741 -1894 7793 -1885
rect 7805 -1894 7857 -1885
rect 7869 -1894 7921 -1885
rect 7933 -1894 7985 -1885
rect 7997 -1894 8049 -1885
rect 7677 -1928 7698 -1894
rect 7698 -1928 7729 -1894
rect 7741 -1928 7772 -1894
rect 7772 -1928 7793 -1894
rect 7805 -1928 7806 -1894
rect 7806 -1928 7846 -1894
rect 7846 -1928 7857 -1894
rect 7869 -1928 7880 -1894
rect 7880 -1928 7920 -1894
rect 7920 -1928 7921 -1894
rect 7933 -1928 7954 -1894
rect 7954 -1928 7985 -1894
rect 7997 -1928 8028 -1894
rect 8028 -1928 8049 -1894
rect 7677 -1937 7729 -1928
rect 7741 -1937 7793 -1928
rect 7805 -1937 7857 -1928
rect 7869 -1937 7921 -1928
rect 7933 -1937 7985 -1928
rect 7997 -1937 8049 -1928
rect 8061 -1894 8113 -1885
rect 8061 -1928 8068 -1894
rect 8068 -1928 8102 -1894
rect 8102 -1928 8113 -1894
rect 8061 -1937 8113 -1928
rect 8125 -1894 8177 -1885
rect 8125 -1928 8142 -1894
rect 8142 -1928 8176 -1894
rect 8176 -1928 8177 -1894
rect 8125 -1937 8177 -1928
rect 8189 -1894 8241 -1885
rect 8253 -1894 8305 -1885
rect 8317 -1894 8369 -1885
rect 8381 -1894 8433 -1885
rect 8445 -1894 8497 -1885
rect 8189 -1928 8216 -1894
rect 8216 -1928 8241 -1894
rect 8253 -1928 8290 -1894
rect 8290 -1928 8305 -1894
rect 8317 -1928 8324 -1894
rect 8324 -1928 8364 -1894
rect 8364 -1928 8369 -1894
rect 8381 -1928 8398 -1894
rect 8398 -1928 8433 -1894
rect 8445 -1928 8472 -1894
rect 8472 -1928 8497 -1894
rect 8189 -1937 8241 -1928
rect 8253 -1937 8305 -1928
rect 8317 -1937 8369 -1928
rect 8381 -1937 8433 -1928
rect 8445 -1937 8497 -1928
rect 8509 -1894 8561 -1885
rect 8509 -1928 8512 -1894
rect 8512 -1928 8546 -1894
rect 8546 -1928 8561 -1894
rect 8509 -1937 8561 -1928
rect 8573 -1894 8625 -1885
rect 8573 -1928 8586 -1894
rect 8586 -1928 8620 -1894
rect 8620 -1928 8625 -1894
rect 8573 -1937 8625 -1928
<< metal2 >>
rect 1934 2803 1990 2812
rect 1934 2703 1990 2747
rect 1934 2603 1990 2647
rect 1934 2503 1990 2547
rect 1990 2447 3889 2494
rect 1934 2438 3889 2447
rect 3945 2438 3970 2494
rect 4026 2438 4051 2494
rect 4107 2438 4132 2494
rect 4188 2438 4213 2494
rect 4269 2438 4294 2494
rect 4350 2438 4376 2494
rect 4432 2438 4458 2494
rect 4514 2438 4540 2494
rect 4596 2438 4622 2494
rect 4678 2438 4704 2494
rect 4760 2438 4769 2494
rect -298 1736 11953 1856
rect -298 1580 11953 1700
tri 3103 1553 3130 1580 ne
rect 1900 1438 2014 1444
rect -359 1428 -242 1434
rect -359 1376 -358 1428
rect -306 1376 -294 1428
rect -359 1355 -242 1376
rect -359 1303 -358 1355
rect -306 1303 -294 1355
rect 1900 1432 1931 1438
rect 1983 1432 2014 1438
rect 1900 1376 1929 1432
rect 1985 1376 2014 1432
rect 1900 1365 2014 1376
rect 1900 1313 1931 1365
rect 1983 1313 2014 1365
rect -359 1291 -242 1303
tri -242 1291 -225 1308 sw
rect 1900 1300 2014 1313
rect -359 1282 -225 1291
rect -359 1230 -358 1282
rect -306 1230 -294 1282
rect -242 1239 -225 1282
tri -225 1239 -173 1291 sw
rect 1900 1244 1929 1300
rect 1985 1244 2014 1300
rect 1900 1239 1931 1244
rect 1983 1239 2014 1244
rect -242 1233 -173 1239
tri -173 1233 -167 1239 sw
rect 1900 1233 2014 1239
rect 3130 1267 3459 1580
tri 3459 1553 3486 1580 nw
rect -242 1230 -167 1233
rect -359 1224 -167 1230
tri -167 1224 -158 1233 sw
rect -359 1172 640 1224
rect 692 1172 712 1224
rect 764 1172 784 1224
rect 836 1172 855 1224
rect 907 1172 913 1224
rect 3130 1215 3136 1267
rect 3188 1215 3203 1267
rect 3255 1215 3269 1267
rect 3321 1215 3335 1267
rect 3387 1215 3401 1267
rect 3453 1215 3459 1267
tri 2149 1207 2154 1212 se
rect 2154 1207 2270 1212
tri 2148 1206 2149 1207 se
rect 2149 1206 2270 1207
rect -359 1160 913 1172
tri 2108 1166 2148 1206 se
rect 2148 1166 2154 1206
rect -359 1108 640 1160
rect 692 1108 712 1160
rect 764 1108 784 1160
rect 836 1108 855 1160
rect 907 1108 913 1160
rect 1112 1154 2154 1166
rect 2206 1154 2218 1206
rect 1112 1140 2270 1154
rect 1112 1133 2154 1140
rect 1112 1081 1118 1133
rect 1170 1081 1195 1133
rect 1247 1081 1272 1133
rect 1324 1081 1348 1133
rect 1400 1081 1424 1133
rect 1476 1081 1500 1133
rect 1552 1088 2154 1133
rect 2206 1088 2218 1140
rect 1552 1081 2270 1088
rect 1112 1074 2270 1081
rect 1112 1055 2154 1074
rect -490 1049 436 1055
rect -490 1048 320 1049
rect -118 997 320 1048
rect 372 997 384 1049
rect 1112 1003 1118 1055
rect 1170 1003 1195 1055
rect 1247 1003 1272 1055
rect 1324 1003 1348 1055
rect 1400 1003 1424 1055
rect 1476 1003 1500 1055
rect 1552 1022 2154 1055
rect 2206 1022 2218 1074
rect 1552 1016 2270 1022
rect 2305 1207 2361 1213
rect 2357 1155 2361 1207
rect 2305 1137 2361 1155
rect 2357 1085 2361 1137
rect 2305 1067 2361 1085
rect 1552 1015 1570 1016
tri 1570 1015 1571 1016 nw
rect 2357 1015 2361 1067
rect 1552 1009 1564 1015
tri 1564 1009 1570 1015 nw
rect 1552 1003 1558 1009
tri 1558 1003 1564 1009 nw
rect -118 958 436 997
rect -118 932 320 958
rect -490 926 320 932
tri 203 906 223 926 ne
rect 223 906 320 926
rect 372 906 384 958
rect 2305 998 2361 1015
rect 2357 946 2361 998
tri 223 867 262 906 ne
rect 262 867 436 906
tri 262 815 314 867 ne
rect 314 815 320 867
rect 372 815 384 867
tri 314 809 320 815 ne
rect 320 809 436 815
rect 1631 931 1747 937
rect 1631 809 1747 815
rect 2305 929 2361 946
rect 2357 877 2361 929
rect 2305 860 2361 877
rect 2357 808 2361 860
rect 2305 791 2361 808
rect 3130 955 3459 1215
rect 3130 903 3136 955
rect 3188 903 3203 955
rect 3255 903 3269 955
rect 3321 903 3335 955
rect 3387 903 3401 955
rect 3453 903 3459 955
rect 3130 791 3459 903
rect 3593 1404 3599 1456
rect 3651 1404 3665 1456
rect 3717 1404 3731 1456
rect 3783 1404 3797 1456
rect 3849 1404 3863 1456
rect 3915 1404 3929 1456
rect 3981 1404 3995 1456
rect 4047 1404 4061 1456
rect 4113 1404 4127 1456
rect 4179 1404 4193 1456
rect 4245 1404 4259 1456
rect 4311 1404 4325 1456
rect 4377 1404 4391 1456
rect 4443 1404 4457 1456
rect 4509 1404 4523 1456
rect 4575 1404 4589 1456
rect 4641 1404 4655 1456
rect 4707 1404 4721 1456
rect 4773 1404 4786 1456
rect 4838 1404 4851 1456
rect 4903 1404 4916 1456
rect 4968 1404 4981 1456
rect 5033 1404 5046 1456
rect 5098 1404 5111 1456
rect 5163 1404 5176 1456
rect 5228 1404 5241 1456
rect 5293 1404 5299 1456
rect 3593 1392 5299 1404
rect 3593 1340 3599 1392
rect 3651 1340 3665 1392
rect 3717 1340 3731 1392
rect 3783 1340 3797 1392
rect 3849 1340 3863 1392
rect 3915 1340 3929 1392
rect 3981 1340 3995 1392
rect 4047 1340 4061 1392
rect 4113 1340 4127 1392
rect 4179 1340 4193 1392
rect 4245 1340 4259 1392
rect 4311 1340 4325 1392
rect 4377 1340 4391 1392
rect 4443 1340 4457 1392
rect 4509 1340 4523 1392
rect 4575 1340 4589 1392
rect 4641 1340 4655 1392
rect 4707 1340 4721 1392
rect 4773 1340 4786 1392
rect 4838 1340 4851 1392
rect 4903 1340 4916 1392
rect 4968 1340 4981 1392
rect 5033 1340 5046 1392
rect 5098 1340 5111 1392
rect 5163 1340 5176 1392
rect 5228 1340 5241 1392
rect 5293 1340 5299 1392
rect 3593 1111 5299 1340
rect 6620 1404 6626 1456
rect 6678 1404 6731 1456
rect 6783 1445 7463 1456
rect 6783 1404 7247 1445
rect 6620 1392 7247 1404
rect 6620 1340 6626 1392
rect 6678 1340 6731 1392
rect 6783 1389 7247 1392
rect 7303 1389 7327 1445
rect 7383 1389 7407 1445
rect 6783 1343 7463 1389
rect 6783 1340 7247 1343
rect 6620 1328 7247 1340
rect 6620 1276 6626 1328
rect 6678 1276 6731 1328
rect 6783 1287 7247 1328
rect 7303 1287 7327 1343
rect 7383 1287 7407 1343
rect 6783 1276 7463 1287
rect 8735 1402 8741 1454
rect 8793 1402 8808 1454
rect 8860 1402 8874 1454
rect 8926 1402 8940 1454
rect 8992 1402 9006 1454
rect 9058 1402 9072 1454
rect 9124 1402 9138 1454
rect 9190 1402 9204 1454
rect 9256 1402 9270 1454
rect 9322 1402 9336 1454
rect 9388 1402 9402 1454
rect 9454 1402 9468 1454
rect 9520 1402 9534 1454
rect 9586 1402 9600 1454
rect 9652 1402 9666 1454
rect 9718 1402 9732 1454
rect 9784 1402 9798 1454
rect 9850 1402 9864 1454
rect 9916 1402 9930 1454
rect 9982 1402 9996 1454
rect 10048 1402 10062 1454
rect 10114 1402 10128 1454
rect 10180 1402 10194 1454
rect 10246 1402 10260 1454
rect 10312 1402 10318 1454
rect 8735 1390 10318 1402
rect 8735 1338 8741 1390
rect 8793 1338 8808 1390
rect 8860 1338 8874 1390
rect 8926 1338 8940 1390
rect 8992 1338 9006 1390
rect 9058 1338 9072 1390
rect 9124 1338 9138 1390
rect 9190 1338 9204 1390
rect 9256 1338 9270 1390
rect 9322 1338 9336 1390
rect 9388 1338 9402 1390
rect 9454 1338 9468 1390
rect 9520 1338 9534 1390
rect 9586 1338 9600 1390
rect 9652 1338 9666 1390
rect 9718 1338 9732 1390
rect 9784 1338 9798 1390
rect 9850 1338 9864 1390
rect 9916 1338 9930 1390
rect 9982 1338 9996 1390
rect 10048 1338 10062 1390
rect 10114 1338 10128 1390
rect 10180 1338 10194 1390
rect 10246 1338 10260 1390
rect 10312 1338 10318 1390
rect 5864 1267 5873 1269
rect 5929 1267 5954 1269
rect 6010 1267 6034 1269
rect 6090 1267 6114 1269
rect 6170 1267 6194 1269
rect 6250 1267 6274 1269
rect 6330 1267 6354 1269
rect 6410 1267 6434 1269
rect 6490 1267 6505 1269
rect 5864 1215 5870 1267
rect 5929 1215 5935 1267
rect 6179 1215 6191 1267
rect 6250 1215 6255 1267
rect 6499 1215 6505 1267
rect 5864 1213 5873 1215
rect 5929 1213 5954 1215
rect 6010 1213 6034 1215
rect 6090 1213 6114 1215
rect 6170 1213 6194 1215
rect 6250 1213 6274 1215
rect 6330 1213 6354 1215
rect 6410 1213 6434 1215
rect 6490 1213 6505 1215
rect 8024 1267 8033 1269
rect 8089 1267 8114 1269
rect 8170 1267 8195 1269
rect 8251 1267 8276 1269
rect 8332 1267 8357 1269
rect 8413 1267 8438 1269
rect 8494 1267 8519 1269
rect 8575 1267 8600 1269
rect 8656 1267 8665 1269
rect 8024 1215 8030 1267
rect 8089 1215 8095 1267
rect 8275 1215 8276 1267
rect 8339 1215 8351 1267
rect 8413 1215 8415 1267
rect 8595 1215 8600 1267
rect 8659 1215 8665 1267
rect 8024 1213 8033 1215
rect 8089 1213 8114 1215
rect 8170 1213 8195 1215
rect 8251 1213 8276 1215
rect 8332 1213 8357 1215
rect 8413 1213 8438 1215
rect 8494 1213 8519 1215
rect 8575 1213 8600 1215
rect 8656 1213 8665 1215
rect 3593 1059 3599 1111
rect 3651 1059 3670 1111
rect 3722 1059 3741 1111
rect 3793 1059 3811 1111
rect 3863 1059 3881 1111
rect 3933 1059 3951 1111
rect 4003 1059 4021 1111
rect 4073 1059 4091 1111
rect 4143 1059 4161 1111
rect 4213 1059 4231 1111
rect 4283 1059 4301 1111
rect 4353 1059 4539 1111
rect 4591 1059 4609 1111
rect 4661 1059 4679 1111
rect 4731 1059 4749 1111
rect 4801 1059 4819 1111
rect 4871 1059 4889 1111
rect 4941 1059 4959 1111
rect 5011 1059 5029 1111
rect 5081 1059 5099 1111
rect 5151 1059 5170 1111
rect 5222 1059 5241 1111
rect 5293 1059 5299 1111
rect 3593 799 5299 1059
rect 6535 1207 7374 1213
rect 6535 1155 6539 1207
rect 6591 1165 7322 1207
rect 6591 1155 6732 1165
rect 6535 1137 6732 1155
rect 6535 1085 6539 1137
rect 6591 1109 6732 1137
rect 6788 1155 7322 1165
rect 6788 1141 7374 1155
rect 6788 1109 7322 1141
rect 6591 1089 7322 1109
rect 6591 1085 7374 1089
rect 6535 1067 6732 1085
rect 6535 1015 6539 1067
rect 6591 1029 6732 1067
rect 6788 1075 7374 1085
rect 6788 1029 7322 1075
rect 6591 1023 7322 1029
rect 6591 1020 7374 1023
rect 6535 996 6591 1015
rect 5864 955 5873 957
rect 5929 955 5954 957
rect 6010 955 6034 957
rect 6090 955 6114 957
rect 6170 955 6194 957
rect 6250 955 6274 957
rect 6330 955 6354 957
rect 6410 955 6434 957
rect 6490 955 6505 957
rect 5864 903 5870 955
rect 5929 903 5935 955
rect 6179 903 6191 955
rect 6250 903 6255 955
rect 6499 903 6505 955
rect 5864 901 5873 903
rect 5929 901 5954 903
rect 6010 901 6034 903
rect 6090 901 6114 903
rect 6170 901 6194 903
rect 6250 901 6274 903
rect 6330 901 6354 903
rect 6410 901 6434 903
rect 6490 901 6505 903
rect 6535 944 6539 996
rect 7318 1009 7374 1020
rect 7318 957 7322 1009
rect 8735 1111 10318 1338
rect 10452 1267 10461 1269
rect 10517 1267 10546 1269
rect 10602 1267 10631 1269
rect 10687 1267 10716 1269
rect 10772 1267 10781 1269
rect 10452 1215 10458 1267
rect 10517 1215 10525 1267
rect 10709 1215 10716 1267
rect 10775 1215 10781 1267
rect 10452 1213 10461 1215
rect 10517 1213 10546 1215
rect 10602 1213 10631 1215
rect 10687 1213 10716 1215
rect 10772 1213 10781 1215
rect 8735 1059 8741 1111
rect 8793 1059 8806 1111
rect 8858 1059 8871 1111
rect 8923 1059 8936 1111
rect 8988 1059 9000 1111
rect 9052 1059 9064 1111
rect 9116 1059 9128 1111
rect 9180 1059 9192 1111
rect 9244 1059 9256 1111
rect 9308 1059 9320 1111
rect 9372 1059 9558 1111
rect 9610 1059 9628 1111
rect 9680 1059 9698 1111
rect 9750 1059 9768 1111
rect 9820 1059 9838 1111
rect 9890 1059 9908 1111
rect 9960 1059 9978 1111
rect 10030 1059 10048 1111
rect 10100 1059 10118 1111
rect 10170 1059 10189 1111
rect 10241 1059 10260 1111
rect 10312 1059 10318 1111
rect 6535 925 6591 944
tri -28 707 24 759 se
rect 24 707 640 759
rect 692 707 712 759
rect 764 707 784 759
rect 836 707 855 759
rect 907 707 913 759
tri -40 695 -28 707 se
rect -28 695 913 707
tri -53 682 -40 695 se
rect -40 682 640 695
tri -79 656 -53 682 se
rect -53 656 640 682
rect -79 643 640 656
rect 692 643 712 695
rect 764 643 784 695
rect 836 643 855 695
rect 907 643 913 695
rect 2357 739 2361 791
rect 2305 722 2361 739
rect -79 630 78 643
tri 78 630 91 643 nw
rect 1111 630 1117 682
rect 1169 630 1194 682
rect 1246 630 1271 682
rect 1323 630 1348 682
rect 1400 630 1424 682
rect 1476 630 1500 682
rect 1552 630 1558 682
rect -79 604 52 630
tri 52 604 78 630 nw
rect 1111 604 1558 630
rect -79 -184 37 604
tri 37 589 52 604 nw
rect 1111 552 1117 604
rect 1169 552 1194 604
rect 1246 552 1271 604
rect 1323 552 1348 604
rect 1400 552 1424 604
rect 1476 552 1500 604
rect 1552 552 1558 604
rect 467 444 473 496
rect 525 444 537 496
rect 589 444 595 496
rect 467 212 519 444
rect 1111 367 1558 552
rect 2357 670 2361 722
tri 1558 367 1568 377 sw
rect 1111 365 1568 367
tri 1568 365 1570 367 sw
rect 1111 313 1570 365
tri 1570 313 1622 365 sw
rect 2305 327 2361 670
rect 3130 643 3459 753
rect 3130 591 3136 643
rect 3188 591 3203 643
rect 3255 591 3269 643
rect 3321 591 3335 643
rect 3387 591 3401 643
rect 3453 591 3459 643
rect 3130 438 3459 591
rect 3593 747 3599 799
rect 3651 747 3670 799
rect 3722 747 3741 799
rect 3793 747 3811 799
rect 3863 747 3881 799
rect 3933 747 3951 799
rect 4003 747 4021 799
rect 4073 747 4091 799
rect 4143 747 4161 799
rect 4213 747 4231 799
rect 4283 747 4301 799
rect 4353 747 4539 799
rect 4591 747 4609 799
rect 4661 747 4679 799
rect 4731 747 4749 799
rect 4801 747 4819 799
rect 4871 747 4889 799
rect 4941 747 4959 799
rect 5011 747 5029 799
rect 5081 747 5099 799
rect 5151 747 5170 799
rect 5222 747 5241 799
rect 5293 747 5299 799
rect 3593 487 5299 747
rect 6535 873 6539 925
rect 6535 854 6591 873
rect 6535 802 6539 854
rect 6535 783 6591 802
rect 6535 731 6539 783
rect 6535 712 6591 731
rect 6535 660 6539 712
rect 6535 654 6591 660
rect 6885 942 6985 948
rect 6885 939 6909 942
rect 6961 939 6985 942
rect 6885 883 6907 939
rect 6963 883 6985 939
rect 6885 876 6985 883
rect 6885 824 6909 876
rect 6961 824 6985 876
rect 6885 812 6985 824
rect 6885 756 6907 812
rect 6963 756 6985 812
rect 6885 744 6985 756
rect 6885 692 6909 744
rect 6961 692 6985 744
rect 6885 684 6985 692
rect 5864 643 5873 645
rect 5929 643 5954 645
rect 6010 643 6034 645
rect 6090 643 6114 645
rect 6170 643 6194 645
rect 6250 643 6274 645
rect 6330 643 6354 645
rect 6410 643 6434 645
rect 6490 643 6505 645
rect 5864 591 5870 643
rect 5929 591 5935 643
rect 6179 591 6191 643
rect 6250 591 6255 643
rect 6499 591 6505 643
rect 6885 628 6907 684
rect 6963 628 6985 684
rect 6885 625 6909 628
rect 6961 625 6985 628
rect 6885 619 6985 625
rect 7318 943 7374 957
rect 7318 891 7322 943
rect 8021 955 8030 957
rect 8086 955 8111 957
rect 8167 955 8192 957
rect 8248 955 8273 957
rect 8329 955 8354 957
rect 8410 955 8435 957
rect 8491 955 8516 957
rect 8572 955 8597 957
rect 8653 955 8662 957
rect 8021 903 8027 955
rect 8086 903 8092 955
rect 8272 903 8273 955
rect 8336 903 8348 955
rect 8410 903 8412 955
rect 8592 903 8597 955
rect 8656 903 8662 955
rect 8021 901 8030 903
rect 8086 901 8111 903
rect 8167 901 8192 903
rect 8248 901 8273 903
rect 8329 901 8354 903
rect 8410 901 8435 903
rect 8491 901 8516 903
rect 8572 901 8597 903
rect 8653 901 8662 903
rect 7318 877 7374 891
rect 7318 825 7322 877
rect 7318 811 7374 825
rect 7318 759 7322 811
rect 7318 745 7374 759
rect 7318 693 7322 745
rect 7318 679 7374 693
rect 7318 627 7322 679
rect 8735 799 10318 1059
rect 11554 1207 11610 1213
rect 11554 1155 11558 1207
rect 11554 1141 11610 1155
rect 11554 1089 11558 1141
rect 11554 1075 11610 1089
rect 11554 1023 11558 1075
rect 11554 1009 11610 1023
rect 11554 957 11558 1009
rect 10452 955 10461 957
rect 10517 955 10546 957
rect 10602 955 10631 957
rect 10687 955 10716 957
rect 10772 955 10781 957
rect 10452 903 10458 955
rect 10517 903 10525 955
rect 10709 903 10716 955
rect 10775 903 10781 955
rect 10452 901 10461 903
rect 10517 901 10546 903
rect 10602 901 10631 903
rect 10687 901 10716 903
rect 10772 901 10781 903
rect 11554 943 11610 957
rect 8735 747 8741 799
rect 8793 747 8806 799
rect 8858 747 8871 799
rect 8923 747 8936 799
rect 8988 747 9000 799
rect 9052 747 9064 799
rect 9116 747 9128 799
rect 9180 747 9192 799
rect 9244 747 9256 799
rect 9308 747 9320 799
rect 9372 747 9558 799
rect 9610 747 9628 799
rect 9680 747 9698 799
rect 9750 747 9768 799
rect 9820 747 9838 799
rect 9890 747 9908 799
rect 9960 747 9978 799
rect 10030 747 10048 799
rect 10100 747 10118 799
rect 10170 747 10189 799
rect 10241 747 10260 799
rect 10312 747 10318 799
rect 5864 589 5873 591
rect 5929 589 5954 591
rect 6010 589 6034 591
rect 6090 589 6114 591
rect 6170 589 6194 591
rect 6250 589 6274 591
rect 6330 589 6354 591
rect 6410 589 6434 591
rect 6490 589 6505 591
rect 7318 613 7374 627
rect 7318 561 7322 613
rect 8021 643 8030 645
rect 8086 643 8111 645
rect 8167 643 8192 645
rect 8248 643 8273 645
rect 8329 643 8354 645
rect 8410 643 8435 645
rect 8491 643 8516 645
rect 8572 643 8597 645
rect 8653 643 8662 645
rect 8021 591 8027 643
rect 8086 591 8092 643
rect 8272 591 8273 643
rect 8336 591 8348 643
rect 8410 591 8412 643
rect 8592 591 8597 643
rect 8656 591 8662 643
rect 8021 589 8030 591
rect 8086 589 8111 591
rect 8167 589 8192 591
rect 8248 589 8273 591
rect 8329 589 8354 591
rect 8410 589 8435 591
rect 8491 589 8516 591
rect 8572 589 8597 591
rect 8653 589 8662 591
rect 7318 547 7374 561
rect 7318 495 7322 547
rect 3593 435 3599 487
rect 3651 435 3670 487
rect 3722 435 3741 487
rect 3793 435 3811 487
rect 3863 435 3881 487
rect 3933 435 3951 487
rect 4003 435 4021 487
rect 4073 435 4091 487
rect 4143 435 4161 487
rect 4213 435 4231 487
rect 4283 435 4301 487
rect 4353 435 4539 487
rect 4591 435 4609 487
rect 4661 435 4679 487
rect 4731 435 4749 487
rect 4801 435 4819 487
rect 4871 435 4889 487
rect 4941 435 4959 487
rect 5011 435 5029 487
rect 5081 435 5099 487
rect 5151 435 5170 487
rect 5222 435 5241 487
rect 5293 435 5299 487
rect 3593 419 5299 435
rect 3593 367 3599 419
rect 3651 367 3665 419
rect 3717 367 3731 419
rect 3783 367 3797 419
rect 3849 367 3863 419
rect 3915 367 3929 419
rect 3981 367 3995 419
rect 4047 367 4061 419
rect 4113 367 4127 419
rect 4179 367 4193 419
rect 4245 367 4259 419
rect 4311 367 4325 419
rect 4377 367 4391 419
rect 4443 367 4457 419
rect 4509 367 4523 419
rect 4575 367 4589 419
rect 4641 367 4655 419
rect 4707 367 4721 419
rect 4773 367 4786 419
rect 4838 367 4851 419
rect 4903 367 4916 419
rect 4968 367 4981 419
rect 5033 367 5046 419
rect 5098 367 5111 419
rect 5163 367 5176 419
rect 5228 367 5241 419
rect 5293 367 5299 419
rect 6649 441 6655 493
rect 6707 441 6760 493
rect 6812 441 6818 493
rect 7318 489 7374 495
rect 8735 487 10318 747
rect 11554 891 11558 943
rect 11554 877 11610 891
rect 11554 825 11558 877
rect 11554 811 11610 825
rect 11554 759 11558 811
rect 11554 745 11610 759
rect 11554 693 11558 745
rect 11554 679 11610 693
rect 10452 643 10461 645
rect 10517 643 10546 645
rect 10602 643 10631 645
rect 10687 643 10716 645
rect 10772 643 10781 645
rect 10452 591 10458 643
rect 10517 591 10525 643
rect 10709 591 10716 643
rect 10775 591 10781 643
rect 10452 589 10461 591
rect 10517 589 10546 591
rect 10602 589 10631 591
rect 10687 589 10716 591
rect 10772 589 10781 591
rect 11554 627 11558 679
rect 11554 613 11610 627
rect 6649 435 6818 441
tri 6818 435 6855 472 sw
rect 8735 435 8741 487
rect 8793 435 8806 487
rect 8858 435 8871 487
rect 8923 435 8936 487
rect 8988 435 9000 487
rect 9052 435 9064 487
rect 9116 435 9128 487
rect 9180 435 9192 487
rect 9244 435 9256 487
rect 9308 435 9320 487
rect 9372 435 9558 487
rect 9610 435 9628 487
rect 9680 435 9698 487
rect 9750 435 9768 487
rect 9820 435 9838 487
rect 9890 435 9908 487
rect 9960 435 9978 487
rect 10030 435 10048 487
rect 10100 435 10118 487
rect 10170 435 10189 487
rect 10241 435 10260 487
rect 10312 435 10318 487
rect 6649 434 6855 435
tri 6855 434 6856 435 sw
rect 6649 429 7446 434
rect 6649 377 6655 429
rect 6707 377 6760 429
rect 6812 423 7446 429
rect 6812 377 7246 423
rect 6649 367 7246 377
rect 7302 367 7390 423
rect 6649 365 7446 367
tri 2361 327 2370 336 sw
rect 2305 313 2370 327
tri 2370 313 2384 327 sw
rect 6649 313 6655 365
rect 6707 313 6760 365
rect 6812 358 7446 365
rect 8735 383 10318 435
rect 6812 336 6836 358
tri 6836 336 6858 358 nw
rect 6812 331 6831 336
tri 6831 331 6836 336 nw
rect 8735 331 8741 383
rect 8793 331 8808 383
rect 8860 331 8874 383
rect 8926 331 8940 383
rect 8992 331 9006 383
rect 9058 331 9072 383
rect 9124 331 9138 383
rect 9190 331 9204 383
rect 9256 331 9270 383
rect 9322 331 9336 383
rect 9388 331 9402 383
rect 9454 331 9468 383
rect 9520 331 9534 383
rect 9586 331 9600 383
rect 9652 331 9666 383
rect 9718 331 9732 383
rect 9784 331 9798 383
rect 9850 331 9864 383
rect 9916 331 9930 383
rect 9982 331 9996 383
rect 10048 331 10062 383
rect 10114 331 10128 383
rect 10180 331 10194 383
rect 10246 331 10260 383
rect 10312 331 10318 383
rect 11554 561 11558 613
rect 11554 547 11610 561
rect 11554 495 11558 547
rect 6812 327 6827 331
tri 6827 327 6831 331 nw
rect 6812 319 6819 327
tri 6819 319 6827 327 nw
tri 7042 319 7050 327 se
rect 7050 319 8372 327
tri 8372 319 8380 327 sw
rect 8735 319 10318 331
rect 6812 313 6818 319
tri 6818 318 6819 319 nw
tri 7041 318 7042 319 se
rect 7042 318 8380 319
tri 7036 313 7041 318 se
rect 7041 313 8380 318
rect 1111 267 1622 313
tri 1622 267 1668 313 sw
rect 2305 296 2384 313
tri 2384 296 2401 313 sw
tri 7019 296 7036 313 se
rect 7036 296 8380 313
tri 8380 296 8403 319 sw
rect 2305 292 3494 296
tri 3494 292 3498 296 sw
tri 7015 292 7019 296 se
rect 7019 295 8403 296
rect 7019 292 7075 295
tri 7075 292 7078 295 nw
tri 8323 292 8326 295 ne
rect 8326 292 8403 295
tri 8403 292 8407 296 sw
rect 2305 280 3498 292
tri 3498 280 3510 292 sw
tri 7003 280 7015 292 se
rect 7015 280 7063 292
tri 7063 280 7075 292 nw
tri 8326 280 8338 292 ne
rect 8338 280 8407 292
rect 2305 267 7050 280
tri 7050 267 7063 280 nw
tri 8338 267 8351 280 ne
rect 8351 267 8407 280
tri 8407 267 8432 292 sw
rect 8735 267 8741 319
rect 8793 267 8808 319
rect 8860 267 8874 319
rect 8926 267 8940 319
rect 8992 267 9006 319
rect 9058 267 9072 319
rect 9124 267 9138 319
rect 9190 267 9204 319
rect 9256 267 9270 319
rect 9322 267 9336 319
rect 9388 267 9402 319
rect 9454 267 9468 319
rect 9520 267 9534 319
rect 9586 267 9600 319
rect 9652 267 9666 319
rect 9718 267 9732 319
rect 9784 267 9798 319
rect 9850 267 9864 319
rect 9916 267 9930 319
rect 9982 267 9996 319
rect 10048 267 10062 319
rect 10114 267 10128 319
rect 10180 267 10194 319
rect 10246 267 10260 319
rect 10312 267 10318 319
tri 11512 296 11554 338 se
rect 11554 296 11610 495
tri 10523 267 10552 296 se
rect 10552 267 11610 296
rect 1111 266 1668 267
tri 1668 266 1669 267 sw
rect 2305 266 7049 267
tri 7049 266 7050 267 nw
tri 8351 266 8352 267 ne
rect 8352 266 8432 267
tri 8432 266 8433 267 sw
tri 10522 266 10523 267 se
rect 10523 266 11610 267
rect 1111 220 1669 266
tri 1669 220 1715 266 sw
rect 2305 264 7047 266
tri 7047 264 7049 266 nw
tri 7097 264 7099 266 se
rect 7099 264 7163 266
tri 3445 248 3461 264 ne
rect 3461 248 7031 264
tri 7031 248 7047 264 nw
tri 7081 248 7097 264 se
rect 7097 248 7163 264
tri 7053 220 7081 248 se
rect 7081 220 7163 248
rect 1111 214 7163 220
rect 7215 214 7229 266
rect 7281 214 7295 266
rect 7347 214 7361 266
rect 7413 214 7426 266
rect 7478 214 7491 266
rect 7543 214 7556 266
rect 7608 214 7621 266
rect 7673 214 7686 266
rect 7738 214 7751 266
rect 7803 214 7816 266
rect 7868 214 7881 266
rect 7933 214 7946 266
rect 7998 214 8011 266
rect 8063 214 8076 266
rect 8128 214 8134 266
tri 8352 246 8372 266 ne
rect 8372 246 8433 266
tri 8372 220 8398 246 ne
rect 8398 220 8433 246
tri 8433 220 8479 266 sw
tri 10476 220 10522 266 se
rect 10522 264 11610 266
rect 10522 220 10552 264
rect 1111 143 8134 214
tri 8398 211 8407 220 ne
rect 8407 215 8479 220
tri 8479 215 8484 220 sw
tri 10471 215 10476 220 se
rect 10476 215 10552 220
tri 10552 215 10601 264 nw
rect 8407 211 8484 215
tri 8484 211 8488 215 sw
tri 10467 211 10471 215 se
rect 10471 211 10548 215
tri 10548 211 10552 215 nw
tri 8407 179 8439 211 ne
rect 8439 179 10516 211
tri 10516 179 10548 211 nw
rect 1111 140 6409 143
tri 6409 140 6412 143 nw
tri 7125 140 7128 143 ne
rect 7128 140 8134 143
rect 10874 175 10883 179
rect 10939 175 10977 179
rect 11033 175 11071 179
rect 11127 175 11136 179
rect 10874 123 10880 175
rect 10939 123 10946 175
rect 11064 123 11071 175
rect 11130 123 11136 175
rect -27 -236 -15 -184
rect -79 -252 37 -236
rect -27 -304 -15 -252
rect -79 -310 37 -304
rect 6522 -1321 6574 -813
rect 6640 -1261 6649 -1259
rect 6705 -1261 6742 -1259
rect 6798 -1261 6834 -1259
rect 6890 -1261 6899 -1259
rect 8038 -1261 8047 -1259
rect 8103 -1261 8135 -1259
rect 8191 -1261 8222 -1259
rect 8278 -1261 8309 -1259
rect 8365 -1261 8396 -1259
rect 8452 -1261 8483 -1259
rect 8539 -1261 8570 -1259
rect 6640 -1313 6646 -1261
rect 6705 -1313 6711 -1261
rect 6828 -1313 6834 -1261
rect 6893 -1313 6906 -1261
rect 6958 -1313 6971 -1261
rect 7023 -1313 7036 -1261
rect 7088 -1313 7101 -1261
rect 7153 -1313 7165 -1261
rect 7217 -1313 7229 -1261
rect 7281 -1313 7293 -1261
rect 7345 -1313 7357 -1261
rect 7409 -1313 7421 -1261
rect 7473 -1313 7485 -1261
rect 7537 -1313 7549 -1261
rect 7601 -1313 7613 -1261
rect 7665 -1313 7677 -1261
rect 7729 -1313 7741 -1261
rect 7793 -1313 7805 -1261
rect 7857 -1313 7869 -1261
rect 7921 -1313 7933 -1261
rect 7985 -1313 7997 -1261
rect 8113 -1313 8125 -1261
rect 8305 -1313 8309 -1261
rect 8369 -1313 8381 -1261
rect 8561 -1313 8570 -1261
rect 6640 -1315 6649 -1313
rect 6705 -1315 6742 -1313
rect 6798 -1315 6834 -1313
rect 6890 -1315 6899 -1313
rect 8038 -1315 8047 -1313
rect 8103 -1315 8135 -1313
rect 8191 -1315 8222 -1313
rect 8278 -1315 8309 -1313
rect 8365 -1315 8396 -1313
rect 8452 -1315 8483 -1313
rect 8539 -1315 8570 -1313
rect 8626 -1315 8635 -1259
rect 6522 -1385 6574 -1373
rect 7230 -1417 7239 -1415
rect 7295 -1417 7394 -1415
rect 7450 -1417 7459 -1415
rect 6522 -1443 6574 -1437
rect 6640 -1469 6646 -1417
rect 6698 -1469 6711 -1417
rect 6763 -1469 6776 -1417
rect 6828 -1469 6841 -1417
rect 6893 -1469 6906 -1417
rect 6958 -1469 6971 -1417
rect 7023 -1469 7036 -1417
rect 7088 -1469 7101 -1417
rect 7153 -1469 7165 -1417
rect 7217 -1469 7229 -1417
rect 7345 -1469 7357 -1417
rect 7473 -1469 7485 -1417
rect 7537 -1469 7549 -1417
rect 7601 -1469 7613 -1417
rect 7665 -1469 7677 -1417
rect 7729 -1469 7741 -1417
rect 7793 -1469 7805 -1417
rect 7857 -1469 7869 -1417
rect 7921 -1469 7933 -1417
rect 7985 -1469 7997 -1417
rect 8049 -1469 8061 -1417
rect 8113 -1469 8125 -1417
rect 8177 -1469 8189 -1417
rect 8241 -1469 8253 -1417
rect 8305 -1469 8317 -1417
rect 8369 -1469 8381 -1417
rect 8433 -1469 8445 -1417
rect 8497 -1469 8509 -1417
rect 8561 -1469 8573 -1417
rect 8625 -1469 8631 -1417
rect 7230 -1471 7239 -1469
rect 7295 -1471 7394 -1469
rect 7450 -1471 7459 -1469
rect 6592 -1627 6601 -1571
rect 6657 -1573 6683 -1571
rect 6739 -1573 6764 -1571
rect 6820 -1573 6845 -1571
rect 6901 -1573 6910 -1571
rect 8038 -1573 8047 -1571
rect 8103 -1573 8135 -1571
rect 8191 -1573 8222 -1571
rect 8278 -1573 8309 -1571
rect 8365 -1573 8396 -1571
rect 8452 -1573 8483 -1571
rect 8539 -1573 8570 -1571
rect 6763 -1625 6764 -1573
rect 6828 -1625 6841 -1573
rect 6901 -1625 6906 -1573
rect 6958 -1625 6971 -1573
rect 7023 -1625 7036 -1573
rect 7088 -1625 7101 -1573
rect 7153 -1625 7165 -1573
rect 7217 -1625 7229 -1573
rect 7281 -1625 7293 -1573
rect 7345 -1625 7357 -1573
rect 7409 -1625 7421 -1573
rect 7473 -1625 7485 -1573
rect 7537 -1625 7549 -1573
rect 7601 -1625 7613 -1573
rect 7665 -1625 7677 -1573
rect 7729 -1625 7741 -1573
rect 7793 -1625 7805 -1573
rect 7857 -1625 7869 -1573
rect 7921 -1625 7933 -1573
rect 7985 -1625 7997 -1573
rect 8113 -1625 8125 -1573
rect 8305 -1625 8309 -1573
rect 8369 -1625 8381 -1573
rect 8561 -1625 8570 -1573
rect 6657 -1627 6683 -1625
rect 6739 -1627 6764 -1625
rect 6820 -1627 6845 -1625
rect 6901 -1627 6910 -1625
rect 8038 -1627 8047 -1625
rect 8103 -1627 8135 -1625
rect 8191 -1627 8222 -1625
rect 8278 -1627 8309 -1625
rect 8365 -1627 8396 -1625
rect 8452 -1627 8483 -1625
rect 8539 -1627 8570 -1625
rect 8626 -1627 8635 -1571
rect 7230 -1729 7239 -1727
rect 7295 -1729 7394 -1727
rect 7450 -1729 7459 -1727
rect 6640 -1781 6646 -1729
rect 6698 -1781 6711 -1729
rect 6763 -1781 6776 -1729
rect 6828 -1781 6841 -1729
rect 6893 -1781 6906 -1729
rect 6958 -1781 6971 -1729
rect 7023 -1781 7036 -1729
rect 7088 -1781 7101 -1729
rect 7153 -1781 7165 -1729
rect 7217 -1781 7229 -1729
rect 7345 -1781 7357 -1729
rect 7473 -1781 7485 -1729
rect 7537 -1781 7549 -1729
rect 7601 -1781 7613 -1729
rect 7665 -1781 7677 -1729
rect 7729 -1781 7741 -1729
rect 7793 -1781 7805 -1729
rect 7857 -1781 7869 -1729
rect 7921 -1781 7933 -1729
rect 7985 -1781 7997 -1729
rect 8049 -1781 8061 -1729
rect 8113 -1781 8125 -1729
rect 8177 -1781 8189 -1729
rect 8241 -1781 8253 -1729
rect 8305 -1781 8317 -1729
rect 8369 -1781 8381 -1729
rect 8433 -1781 8445 -1729
rect 8497 -1781 8509 -1729
rect 8561 -1781 8573 -1729
rect 8625 -1781 8631 -1729
rect 7230 -1783 7239 -1781
rect 7295 -1783 7394 -1781
rect 7450 -1783 7459 -1781
rect 6592 -1939 6601 -1883
rect 6657 -1885 6683 -1883
rect 6739 -1885 6764 -1883
rect 6820 -1885 6845 -1883
rect 6901 -1885 6910 -1883
rect 8038 -1885 8047 -1883
rect 8103 -1885 8135 -1883
rect 8191 -1885 8222 -1883
rect 8278 -1885 8309 -1883
rect 8365 -1885 8396 -1883
rect 8452 -1885 8483 -1883
rect 8539 -1885 8570 -1883
rect 6763 -1937 6764 -1885
rect 6828 -1937 6841 -1885
rect 6901 -1937 6906 -1885
rect 6958 -1937 6971 -1885
rect 7023 -1937 7036 -1885
rect 7088 -1937 7101 -1885
rect 7153 -1937 7165 -1885
rect 7217 -1937 7229 -1885
rect 7281 -1937 7293 -1885
rect 7345 -1937 7357 -1885
rect 7409 -1937 7421 -1885
rect 7473 -1937 7485 -1885
rect 7537 -1937 7549 -1885
rect 7601 -1937 7613 -1885
rect 7665 -1937 7677 -1885
rect 7729 -1937 7741 -1885
rect 7793 -1937 7805 -1885
rect 7857 -1937 7869 -1885
rect 7921 -1937 7933 -1885
rect 7985 -1937 7997 -1885
rect 8113 -1937 8125 -1885
rect 8305 -1937 8309 -1885
rect 8369 -1937 8381 -1885
rect 8561 -1937 8570 -1885
rect 6657 -1939 6683 -1937
rect 6739 -1939 6764 -1937
rect 6820 -1939 6845 -1937
rect 6901 -1939 6910 -1937
rect 8038 -1939 8047 -1937
rect 8103 -1939 8135 -1937
rect 8191 -1939 8222 -1937
rect 8278 -1939 8309 -1937
rect 8365 -1939 8396 -1937
rect 8452 -1939 8483 -1937
rect 8539 -1939 8570 -1937
rect 8626 -1939 8635 -1883
<< via2 >>
rect 1934 2747 1990 2803
rect 1934 2647 1990 2703
rect 1934 2547 1990 2603
rect 1934 2447 1990 2503
rect 3889 2438 3945 2494
rect 3970 2438 4026 2494
rect 4051 2438 4107 2494
rect 4132 2438 4188 2494
rect 4213 2438 4269 2494
rect 4294 2438 4350 2494
rect 4376 2438 4432 2494
rect 4458 2438 4514 2494
rect 4540 2438 4596 2494
rect 4622 2438 4678 2494
rect 4704 2438 4760 2494
rect 1929 1386 1931 1432
rect 1931 1386 1983 1432
rect 1983 1386 1985 1432
rect 1929 1376 1985 1386
rect 1929 1291 1985 1300
rect 1929 1244 1931 1291
rect 1931 1244 1983 1291
rect 1983 1244 1985 1291
rect 7247 1389 7303 1445
rect 7327 1389 7383 1445
rect 7407 1389 7463 1445
rect 7247 1287 7303 1343
rect 7327 1287 7383 1343
rect 7407 1287 7463 1343
rect 5873 1267 5929 1269
rect 5954 1267 6010 1269
rect 6034 1267 6090 1269
rect 6114 1267 6170 1269
rect 6194 1267 6250 1269
rect 6274 1267 6330 1269
rect 6354 1267 6410 1269
rect 6434 1267 6490 1269
rect 5873 1215 5922 1267
rect 5922 1215 5929 1267
rect 5954 1215 5987 1267
rect 5987 1215 5999 1267
rect 5999 1215 6010 1267
rect 6034 1215 6051 1267
rect 6051 1215 6063 1267
rect 6063 1215 6090 1267
rect 6114 1215 6115 1267
rect 6115 1215 6127 1267
rect 6127 1215 6170 1267
rect 6194 1215 6243 1267
rect 6243 1215 6250 1267
rect 6274 1215 6307 1267
rect 6307 1215 6319 1267
rect 6319 1215 6330 1267
rect 6354 1215 6371 1267
rect 6371 1215 6383 1267
rect 6383 1215 6410 1267
rect 6434 1215 6435 1267
rect 6435 1215 6447 1267
rect 6447 1215 6490 1267
rect 5873 1213 5929 1215
rect 5954 1213 6010 1215
rect 6034 1213 6090 1215
rect 6114 1213 6170 1215
rect 6194 1213 6250 1215
rect 6274 1213 6330 1215
rect 6354 1213 6410 1215
rect 6434 1213 6490 1215
rect 8033 1267 8089 1269
rect 8114 1267 8170 1269
rect 8195 1267 8251 1269
rect 8276 1267 8332 1269
rect 8357 1267 8413 1269
rect 8438 1267 8494 1269
rect 8519 1267 8575 1269
rect 8600 1267 8656 1269
rect 8033 1215 8082 1267
rect 8082 1215 8089 1267
rect 8114 1215 8147 1267
rect 8147 1215 8159 1267
rect 8159 1215 8170 1267
rect 8195 1215 8211 1267
rect 8211 1215 8223 1267
rect 8223 1215 8251 1267
rect 8276 1215 8287 1267
rect 8287 1215 8332 1267
rect 8357 1215 8403 1267
rect 8403 1215 8413 1267
rect 8438 1215 8467 1267
rect 8467 1215 8479 1267
rect 8479 1215 8494 1267
rect 8519 1215 8531 1267
rect 8531 1215 8543 1267
rect 8543 1215 8575 1267
rect 8600 1215 8607 1267
rect 8607 1215 8656 1267
rect 8033 1213 8089 1215
rect 8114 1213 8170 1215
rect 8195 1213 8251 1215
rect 8276 1213 8332 1215
rect 8357 1213 8413 1215
rect 8438 1213 8494 1215
rect 8519 1213 8575 1215
rect 8600 1213 8656 1215
rect 6732 1109 6788 1165
rect 6732 1029 6788 1085
rect 5873 955 5929 957
rect 5954 955 6010 957
rect 6034 955 6090 957
rect 6114 955 6170 957
rect 6194 955 6250 957
rect 6274 955 6330 957
rect 6354 955 6410 957
rect 6434 955 6490 957
rect 5873 903 5922 955
rect 5922 903 5929 955
rect 5954 903 5987 955
rect 5987 903 5999 955
rect 5999 903 6010 955
rect 6034 903 6051 955
rect 6051 903 6063 955
rect 6063 903 6090 955
rect 6114 903 6115 955
rect 6115 903 6127 955
rect 6127 903 6170 955
rect 6194 903 6243 955
rect 6243 903 6250 955
rect 6274 903 6307 955
rect 6307 903 6319 955
rect 6319 903 6330 955
rect 6354 903 6371 955
rect 6371 903 6383 955
rect 6383 903 6410 955
rect 6434 903 6435 955
rect 6435 903 6447 955
rect 6447 903 6490 955
rect 5873 901 5929 903
rect 5954 901 6010 903
rect 6034 901 6090 903
rect 6114 901 6170 903
rect 6194 901 6250 903
rect 6274 901 6330 903
rect 6354 901 6410 903
rect 6434 901 6490 903
rect 10461 1267 10517 1269
rect 10546 1267 10602 1269
rect 10631 1267 10687 1269
rect 10716 1267 10772 1269
rect 10461 1215 10510 1267
rect 10510 1215 10517 1267
rect 10546 1215 10577 1267
rect 10577 1215 10591 1267
rect 10591 1215 10602 1267
rect 10631 1215 10643 1267
rect 10643 1215 10657 1267
rect 10657 1215 10687 1267
rect 10716 1215 10723 1267
rect 10723 1215 10772 1267
rect 10461 1213 10517 1215
rect 10546 1213 10602 1215
rect 10631 1213 10687 1215
rect 10716 1213 10772 1215
rect 6907 890 6909 939
rect 6909 890 6961 939
rect 6961 890 6963 939
rect 6907 883 6963 890
rect 6907 810 6963 812
rect 6907 758 6909 810
rect 6909 758 6961 810
rect 6961 758 6963 810
rect 6907 756 6963 758
rect 5873 643 5929 645
rect 5954 643 6010 645
rect 6034 643 6090 645
rect 6114 643 6170 645
rect 6194 643 6250 645
rect 6274 643 6330 645
rect 6354 643 6410 645
rect 6434 643 6490 645
rect 5873 591 5922 643
rect 5922 591 5929 643
rect 5954 591 5987 643
rect 5987 591 5999 643
rect 5999 591 6010 643
rect 6034 591 6051 643
rect 6051 591 6063 643
rect 6063 591 6090 643
rect 6114 591 6115 643
rect 6115 591 6127 643
rect 6127 591 6170 643
rect 6194 591 6243 643
rect 6243 591 6250 643
rect 6274 591 6307 643
rect 6307 591 6319 643
rect 6319 591 6330 643
rect 6354 591 6371 643
rect 6371 591 6383 643
rect 6383 591 6410 643
rect 6434 591 6435 643
rect 6435 591 6447 643
rect 6447 591 6490 643
rect 6907 677 6963 684
rect 6907 628 6909 677
rect 6909 628 6961 677
rect 6961 628 6963 677
rect 8030 955 8086 957
rect 8111 955 8167 957
rect 8192 955 8248 957
rect 8273 955 8329 957
rect 8354 955 8410 957
rect 8435 955 8491 957
rect 8516 955 8572 957
rect 8597 955 8653 957
rect 8030 903 8079 955
rect 8079 903 8086 955
rect 8111 903 8144 955
rect 8144 903 8156 955
rect 8156 903 8167 955
rect 8192 903 8208 955
rect 8208 903 8220 955
rect 8220 903 8248 955
rect 8273 903 8284 955
rect 8284 903 8329 955
rect 8354 903 8400 955
rect 8400 903 8410 955
rect 8435 903 8464 955
rect 8464 903 8476 955
rect 8476 903 8491 955
rect 8516 903 8528 955
rect 8528 903 8540 955
rect 8540 903 8572 955
rect 8597 903 8604 955
rect 8604 903 8653 955
rect 8030 901 8086 903
rect 8111 901 8167 903
rect 8192 901 8248 903
rect 8273 901 8329 903
rect 8354 901 8410 903
rect 8435 901 8491 903
rect 8516 901 8572 903
rect 8597 901 8653 903
rect 10461 955 10517 957
rect 10546 955 10602 957
rect 10631 955 10687 957
rect 10716 955 10772 957
rect 10461 903 10510 955
rect 10510 903 10517 955
rect 10546 903 10577 955
rect 10577 903 10591 955
rect 10591 903 10602 955
rect 10631 903 10643 955
rect 10643 903 10657 955
rect 10657 903 10687 955
rect 10716 903 10723 955
rect 10723 903 10772 955
rect 10461 901 10517 903
rect 10546 901 10602 903
rect 10631 901 10687 903
rect 10716 901 10772 903
rect 5873 589 5929 591
rect 5954 589 6010 591
rect 6034 589 6090 591
rect 6114 589 6170 591
rect 6194 589 6250 591
rect 6274 589 6330 591
rect 6354 589 6410 591
rect 6434 589 6490 591
rect 8030 643 8086 645
rect 8111 643 8167 645
rect 8192 643 8248 645
rect 8273 643 8329 645
rect 8354 643 8410 645
rect 8435 643 8491 645
rect 8516 643 8572 645
rect 8597 643 8653 645
rect 8030 591 8079 643
rect 8079 591 8086 643
rect 8111 591 8144 643
rect 8144 591 8156 643
rect 8156 591 8167 643
rect 8192 591 8208 643
rect 8208 591 8220 643
rect 8220 591 8248 643
rect 8273 591 8284 643
rect 8284 591 8329 643
rect 8354 591 8400 643
rect 8400 591 8410 643
rect 8435 591 8464 643
rect 8464 591 8476 643
rect 8476 591 8491 643
rect 8516 591 8528 643
rect 8528 591 8540 643
rect 8540 591 8572 643
rect 8597 591 8604 643
rect 8604 591 8653 643
rect 8030 589 8086 591
rect 8111 589 8167 591
rect 8192 589 8248 591
rect 8273 589 8329 591
rect 8354 589 8410 591
rect 8435 589 8491 591
rect 8516 589 8572 591
rect 8597 589 8653 591
rect 10461 643 10517 645
rect 10546 643 10602 645
rect 10631 643 10687 645
rect 10716 643 10772 645
rect 10461 591 10510 643
rect 10510 591 10517 643
rect 10546 591 10577 643
rect 10577 591 10591 643
rect 10591 591 10602 643
rect 10631 591 10643 643
rect 10643 591 10657 643
rect 10657 591 10687 643
rect 10716 591 10723 643
rect 10723 591 10772 643
rect 10461 589 10517 591
rect 10546 589 10602 591
rect 10631 589 10687 591
rect 10716 589 10772 591
rect 7246 367 7302 423
rect 7390 367 7446 423
rect 10883 175 10939 179
rect 10977 175 11033 179
rect 11071 175 11127 179
rect 10883 123 10932 175
rect 10932 123 10939 175
rect 10977 123 10998 175
rect 10998 123 11012 175
rect 11012 123 11033 175
rect 11071 123 11078 175
rect 11078 123 11127 175
rect 6649 -1261 6705 -1259
rect 6742 -1261 6798 -1259
rect 6834 -1261 6890 -1259
rect 8047 -1261 8103 -1259
rect 8135 -1261 8191 -1259
rect 8222 -1261 8278 -1259
rect 8309 -1261 8365 -1259
rect 8396 -1261 8452 -1259
rect 8483 -1261 8539 -1259
rect 8570 -1261 8626 -1259
rect 6649 -1313 6698 -1261
rect 6698 -1313 6705 -1261
rect 6742 -1313 6763 -1261
rect 6763 -1313 6776 -1261
rect 6776 -1313 6798 -1261
rect 6834 -1313 6841 -1261
rect 6841 -1313 6890 -1261
rect 8047 -1313 8049 -1261
rect 8049 -1313 8061 -1261
rect 8061 -1313 8103 -1261
rect 8135 -1313 8177 -1261
rect 8177 -1313 8189 -1261
rect 8189 -1313 8191 -1261
rect 8222 -1313 8241 -1261
rect 8241 -1313 8253 -1261
rect 8253 -1313 8278 -1261
rect 8309 -1313 8317 -1261
rect 8317 -1313 8365 -1261
rect 8396 -1313 8433 -1261
rect 8433 -1313 8445 -1261
rect 8445 -1313 8452 -1261
rect 8483 -1313 8497 -1261
rect 8497 -1313 8509 -1261
rect 8509 -1313 8539 -1261
rect 8570 -1313 8573 -1261
rect 8573 -1313 8625 -1261
rect 8625 -1313 8626 -1261
rect 6649 -1315 6705 -1313
rect 6742 -1315 6798 -1313
rect 6834 -1315 6890 -1313
rect 8047 -1315 8103 -1313
rect 8135 -1315 8191 -1313
rect 8222 -1315 8278 -1313
rect 8309 -1315 8365 -1313
rect 8396 -1315 8452 -1313
rect 8483 -1315 8539 -1313
rect 8570 -1315 8626 -1313
rect 7239 -1417 7295 -1415
rect 7394 -1417 7450 -1415
rect 7239 -1469 7281 -1417
rect 7281 -1469 7293 -1417
rect 7293 -1469 7295 -1417
rect 7394 -1469 7409 -1417
rect 7409 -1469 7421 -1417
rect 7421 -1469 7450 -1417
rect 7239 -1471 7295 -1469
rect 7394 -1471 7450 -1469
rect 6601 -1573 6657 -1571
rect 6683 -1573 6739 -1571
rect 6764 -1573 6820 -1571
rect 6845 -1573 6901 -1571
rect 8047 -1573 8103 -1571
rect 8135 -1573 8191 -1571
rect 8222 -1573 8278 -1571
rect 8309 -1573 8365 -1571
rect 8396 -1573 8452 -1571
rect 8483 -1573 8539 -1571
rect 8570 -1573 8626 -1571
rect 6601 -1625 6646 -1573
rect 6646 -1625 6657 -1573
rect 6683 -1625 6698 -1573
rect 6698 -1625 6711 -1573
rect 6711 -1625 6739 -1573
rect 6764 -1625 6776 -1573
rect 6776 -1625 6820 -1573
rect 6845 -1625 6893 -1573
rect 6893 -1625 6901 -1573
rect 8047 -1625 8049 -1573
rect 8049 -1625 8061 -1573
rect 8061 -1625 8103 -1573
rect 8135 -1625 8177 -1573
rect 8177 -1625 8189 -1573
rect 8189 -1625 8191 -1573
rect 8222 -1625 8241 -1573
rect 8241 -1625 8253 -1573
rect 8253 -1625 8278 -1573
rect 8309 -1625 8317 -1573
rect 8317 -1625 8365 -1573
rect 8396 -1625 8433 -1573
rect 8433 -1625 8445 -1573
rect 8445 -1625 8452 -1573
rect 8483 -1625 8497 -1573
rect 8497 -1625 8509 -1573
rect 8509 -1625 8539 -1573
rect 8570 -1625 8573 -1573
rect 8573 -1625 8625 -1573
rect 8625 -1625 8626 -1573
rect 6601 -1627 6657 -1625
rect 6683 -1627 6739 -1625
rect 6764 -1627 6820 -1625
rect 6845 -1627 6901 -1625
rect 8047 -1627 8103 -1625
rect 8135 -1627 8191 -1625
rect 8222 -1627 8278 -1625
rect 8309 -1627 8365 -1625
rect 8396 -1627 8452 -1625
rect 8483 -1627 8539 -1625
rect 8570 -1627 8626 -1625
rect 7239 -1729 7295 -1727
rect 7394 -1729 7450 -1727
rect 7239 -1781 7281 -1729
rect 7281 -1781 7293 -1729
rect 7293 -1781 7295 -1729
rect 7394 -1781 7409 -1729
rect 7409 -1781 7421 -1729
rect 7421 -1781 7450 -1729
rect 7239 -1783 7295 -1781
rect 7394 -1783 7450 -1781
rect 6601 -1885 6657 -1883
rect 6683 -1885 6739 -1883
rect 6764 -1885 6820 -1883
rect 6845 -1885 6901 -1883
rect 8047 -1885 8103 -1883
rect 8135 -1885 8191 -1883
rect 8222 -1885 8278 -1883
rect 8309 -1885 8365 -1883
rect 8396 -1885 8452 -1883
rect 8483 -1885 8539 -1883
rect 8570 -1885 8626 -1883
rect 6601 -1937 6646 -1885
rect 6646 -1937 6657 -1885
rect 6683 -1937 6698 -1885
rect 6698 -1937 6711 -1885
rect 6711 -1937 6739 -1885
rect 6764 -1937 6776 -1885
rect 6776 -1937 6820 -1885
rect 6845 -1937 6893 -1885
rect 6893 -1937 6901 -1885
rect 8047 -1937 8049 -1885
rect 8049 -1937 8061 -1885
rect 8061 -1937 8103 -1885
rect 8135 -1937 8177 -1885
rect 8177 -1937 8189 -1885
rect 8189 -1937 8191 -1885
rect 8222 -1937 8241 -1885
rect 8241 -1937 8253 -1885
rect 8253 -1937 8278 -1885
rect 8309 -1937 8317 -1885
rect 8317 -1937 8365 -1885
rect 8396 -1937 8433 -1885
rect 8433 -1937 8445 -1885
rect 8445 -1937 8452 -1885
rect 8483 -1937 8497 -1885
rect 8497 -1937 8509 -1885
rect 8509 -1937 8539 -1885
rect 8570 -1937 8573 -1885
rect 8573 -1937 8625 -1885
rect 8625 -1937 8626 -1885
rect 6601 -1939 6657 -1937
rect 6683 -1939 6739 -1937
rect 6764 -1939 6820 -1937
rect 6845 -1939 6901 -1937
rect 8047 -1939 8103 -1937
rect 8135 -1939 8191 -1937
rect 8222 -1939 8278 -1937
rect 8309 -1939 8365 -1937
rect 8396 -1939 8452 -1937
rect 8483 -1939 8539 -1937
rect 8570 -1939 8626 -1937
<< metal3 >>
rect 1898 2803 2016 2808
rect 1898 2747 1934 2803
rect 1990 2747 2016 2803
rect 1898 2703 2016 2747
rect 1898 2647 1934 2703
rect 1990 2647 2016 2703
rect 1898 2603 2016 2647
rect 1898 2547 1934 2603
rect 1990 2547 2016 2603
rect 1898 2503 2016 2547
rect 1898 2447 1934 2503
rect 1990 2447 2016 2503
rect 1898 1432 2016 2447
rect 3884 2494 4765 2499
rect 3884 2438 3889 2494
rect 3945 2438 3970 2494
rect 4026 2438 4051 2494
rect 4107 2438 4132 2494
rect 4188 2438 4213 2494
rect 4269 2438 4294 2494
rect 4350 2438 4376 2494
rect 4432 2438 4458 2494
rect 4514 2438 4540 2494
rect 4596 2438 4622 2494
rect 4678 2438 4704 2494
rect 4760 2438 4765 2494
rect 3884 2433 4765 2438
tri 10804 1878 10878 1952 ne
rect 10878 1878 11179 1952
tri 11179 1878 11253 1952 nw
tri 6610 1720 6667 1777 sw
rect 6610 1661 6931 1720
tri 6931 1661 6990 1720 sw
rect 6610 1624 6990 1661
tri 6843 1587 6880 1624 ne
rect 1898 1376 1929 1432
rect 1985 1376 2016 1432
rect 1898 1300 2016 1376
rect 1898 1244 1929 1300
rect 1985 1244 2016 1300
rect 1898 1239 2016 1244
rect 5865 1269 6496 1278
rect 5865 1213 5873 1269
rect 5929 1213 5954 1269
rect 6010 1213 6034 1269
rect 6090 1213 6114 1269
rect 6170 1213 6194 1269
rect 6250 1213 6274 1269
rect 6330 1213 6354 1269
rect 6410 1213 6434 1269
rect 6490 1213 6496 1269
rect 5865 957 6496 1213
rect 5865 901 5873 957
rect 5929 901 5954 957
rect 6010 901 6034 957
rect 6090 901 6114 957
rect 6170 901 6194 957
rect 6250 901 6274 957
rect 6330 901 6354 957
rect 6410 901 6434 957
rect 6490 901 6496 957
rect 5865 645 6496 901
rect 5865 589 5873 645
rect 5929 589 5954 645
rect 6010 589 6034 645
rect 6090 589 6114 645
rect 6170 589 6194 645
rect 6250 589 6274 645
rect 6330 589 6354 645
rect 6410 589 6434 645
rect 6490 589 6496 645
rect 5865 -1252 6496 589
rect 6727 1165 6793 1170
rect 6727 1109 6732 1165
rect 6788 1109 6793 1165
rect 6727 1085 6793 1109
rect 6727 1029 6732 1085
rect 6788 1029 6793 1085
rect 6727 -61 6793 1029
rect 6880 939 6990 1624
rect 7242 1445 7468 1450
rect 7242 1443 7247 1445
rect 6880 883 6907 939
rect 6963 883 6990 939
rect 6880 812 6990 883
rect 6880 756 6907 812
rect 6963 756 6990 812
rect 6880 684 6990 756
rect 6880 628 6907 684
rect 6963 628 6990 684
rect 6880 623 6990 628
rect 7234 1389 7247 1443
rect 7303 1389 7327 1445
rect 7383 1389 7407 1445
rect 7463 1389 7468 1445
rect 7234 1343 7468 1389
rect 7234 1287 7247 1343
rect 7303 1287 7327 1343
rect 7383 1287 7407 1343
rect 7463 1287 7468 1343
rect 7234 1282 7468 1287
rect 7234 423 7455 1282
rect 7234 367 7246 423
rect 7302 367 7390 423
rect 7446 367 7455 423
tri 6496 -1252 6683 -1065 sw
rect 5865 -1259 6906 -1252
rect 5865 -1315 6649 -1259
rect 6705 -1315 6742 -1259
rect 6798 -1315 6834 -1259
rect 6890 -1315 6906 -1259
rect 5865 -1571 6906 -1315
rect 5865 -1627 6601 -1571
rect 6657 -1627 6683 -1571
rect 6739 -1627 6764 -1571
rect 6820 -1627 6845 -1571
rect 6901 -1627 6906 -1571
rect 5865 -1883 6906 -1627
rect 7234 -1415 7455 367
rect 7234 -1471 7239 -1415
rect 7295 -1471 7394 -1415
rect 7450 -1471 7455 -1415
rect 7234 -1727 7455 -1471
rect 7234 -1783 7239 -1727
rect 7295 -1783 7394 -1727
rect 7450 -1783 7455 -1727
rect 7234 -1788 7455 -1783
rect 8025 1269 8665 1274
rect 8025 1213 8033 1269
rect 8089 1213 8114 1269
rect 8170 1213 8195 1269
rect 8251 1213 8276 1269
rect 8332 1213 8357 1269
rect 8413 1213 8438 1269
rect 8494 1213 8519 1269
rect 8575 1213 8600 1269
rect 8656 1213 8665 1269
rect 8025 957 8665 1213
rect 8025 901 8030 957
rect 8086 901 8111 957
rect 8167 901 8192 957
rect 8248 901 8273 957
rect 8329 901 8354 957
rect 8410 901 8435 957
rect 8491 901 8516 957
rect 8572 901 8597 957
rect 8653 901 8665 957
rect 8025 645 8665 901
rect 10452 1269 10781 1859
rect 10452 1213 10461 1269
rect 10517 1213 10546 1269
rect 10602 1213 10631 1269
rect 10687 1213 10716 1269
rect 10772 1213 10781 1269
rect 10452 957 10781 1213
rect 10452 901 10461 957
rect 10517 901 10546 957
rect 10602 901 10631 957
rect 10687 901 10716 957
rect 10772 901 10781 957
rect 10452 882 10781 901
rect 8025 589 8030 645
rect 8086 589 8111 645
rect 8167 589 8192 645
rect 8248 589 8273 645
rect 8329 589 8354 645
rect 8410 589 8435 645
rect 8491 589 8516 645
rect 8572 589 8597 645
rect 8653 589 8665 645
rect 8025 -1259 8665 589
rect 10452 645 10781 803
rect 10452 589 10461 645
rect 10517 589 10546 645
rect 10602 589 10631 645
rect 10687 589 10716 645
rect 10772 589 10781 645
rect 10452 438 10781 589
rect 10878 179 11132 1878
tri 11132 1831 11179 1878 nw
rect 10878 123 10883 179
rect 10939 123 10977 179
rect 11033 123 11071 179
rect 11127 123 11132 179
rect 10878 118 11132 123
rect 8025 -1315 8047 -1259
rect 8103 -1315 8135 -1259
rect 8191 -1315 8222 -1259
rect 8278 -1315 8309 -1259
rect 8365 -1315 8396 -1259
rect 8452 -1315 8483 -1259
rect 8539 -1315 8570 -1259
rect 8626 -1315 8665 -1259
rect 8025 -1571 8665 -1315
rect 8025 -1627 8047 -1571
rect 8103 -1627 8135 -1571
rect 8191 -1627 8222 -1571
rect 8278 -1627 8309 -1571
rect 8365 -1627 8396 -1571
rect 8452 -1627 8483 -1571
rect 8539 -1627 8570 -1571
rect 8626 -1627 8665 -1571
rect 5865 -1939 6601 -1883
rect 6657 -1939 6683 -1883
rect 6739 -1939 6764 -1883
rect 6820 -1939 6845 -1883
rect 6901 -1939 6906 -1883
rect 5865 -2139 6906 -1939
rect 8025 -1883 8665 -1627
rect 8025 -1939 8047 -1883
rect 8103 -1939 8135 -1883
rect 8191 -1939 8222 -1883
rect 8278 -1939 8309 -1883
rect 8365 -1939 8396 -1883
rect 8452 -1939 8483 -1883
rect 8539 -1939 8570 -1883
rect 8626 -1939 8665 -1883
rect 8025 -1944 8665 -1939
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_0
timestamp 1644511149
transform 0 -1 -104 -1 0 701
box 0 0 882 404
use sky130_fd_io__res75only_small  sky130_fd_io__res75only_small_1
timestamp 1644511149
transform 0 -1 -104 1 0 551
box 0 0 882 404
use sky130_fd_pr__nfet_01v8__example_55959141808516  sky130_fd_pr__nfet_01v8__example_55959141808516_0
timestamp 1644511149
transform 0 1 558 -1 0 745
box -28 0 284 471
use sky130_fd_pr__nfet_01v8__example_55959141808516  sky130_fd_pr__nfet_01v8__example_55959141808516_1
timestamp 1644511149
transform 0 1 558 -1 0 1187
box -28 0 284 471
use sky130_fd_pr__nfet_01v8__example_55959141808519  sky130_fd_pr__nfet_01v8__example_55959141808519_0
timestamp 1644511149
transform 0 1 2393 1 0 489
box -28 0 284 981
use sky130_fd_pr__nfet_01v8__example_55959141808519  sky130_fd_pr__nfet_01v8__example_55959141808519_1
timestamp 1644511149
transform 0 -1 11518 1 0 489
box -28 0 284 981
use sky130_fd_pr__nfet_01v8__example_55959141808522  sky130_fd_pr__nfet_01v8__example_55959141808522_0
timestamp 1644511149
transform 0 -1 11518 1 0 801
box -28 0 440 981
use sky130_fd_pr__nfet_01v8__example_55959141808522  sky130_fd_pr__nfet_01v8__example_55959141808522_1
timestamp 1644511149
transform 0 1 2393 1 0 801
box -28 0 440 981
use sky130_fd_pr__nfet_01v8__example_55959141808523  sky130_fd_pr__nfet_01v8__example_55959141808523_0
timestamp 1644511149
transform 0 -1 9412 -1 0 1213
box -28 0 752 981
use sky130_fd_pr__nfet_01v8__example_55959141808523  sky130_fd_pr__nfet_01v8__example_55959141808523_1
timestamp 1644511149
transform 0 -1 6499 1 0 489
box -28 0 752 981
use sky130_fd_pr__pfet_01v8__example_55959141808514  sky130_fd_pr__pfet_01v8__example_55959141808514_0
timestamp 1644511149
transform 0 -1 8616 1 0 -1883
box -28 0 596 981
<< labels >>
flabel metal3 s 6727 680 6793 732 3 FreeSans 520 0 0 0 NG_AG_VPMP
port 1 nsew
flabel metal3 s 5870 -611 6492 -234 3 FreeSans 520 0 0 0 AG_HV
port 2 nsew
flabel metal3 s 10455 1022 10772 1149 3 FreeSans 520 0 0 0 PAD_HV_N2
port 3 nsew
flabel metal3 s 10458 533 10775 681 3 FreeSans 520 0 0 0 PAD_HV_N3
port 4 nsew
flabel metal1 s -474 635 -185 762 3 FreeSans 520 0 0 0 VSSA
port 5 nsew
flabel metal2 s 3130 1035 3459 1165 3 FreeSans 520 0 0 0 PAD_HV_N0
port 6 nsew
flabel metal2 s 3131 650 3458 704 3 FreeSans 520 0 0 0 PAD_HV_N1
port 7 nsew
flabel metal2 s 467 448 519 484 3 FreeSans 520 0 0 0 NMID_VDDA
port 8 nsew
flabel metal2 s 2364 264 2472 296 3 FreeSans 520 0 0 0 NG_PAD_VPMP
port 9 nsew
flabel metal2 s 6522 -1427 6571 -1319 3 FreeSans 520 0 0 0 PG_AG_VDDA
port 10 nsew
flabel comment s 7133 547 7133 547 0 FreeSans 440 90 0 0 CONDIODE
flabel comment s 488 404 488 404 0 FreeSans 400 90 0 0 NMID_VDDA
flabel comment s 2136 547 2136 547 0 FreeSans 440 90 0 0 CONDIODE
flabel comment s 292 547 292 547 0 FreeSans 440 90 0 0 CONDIODE
<< properties >>
string GDS_END 48027794
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 47734134
<< end >>
