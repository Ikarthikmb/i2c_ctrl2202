/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/special_nfet_pass_lvt/sky130_fd_pr__special_nfet_pass_lvt__ss.corner.spice