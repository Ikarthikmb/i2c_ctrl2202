magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect 1632 0 3140 490
<< pwell >>
rect 811 328 913 462
<< psubdiff >>
rect 837 412 887 436
rect 837 378 845 412
rect 879 378 887 412
rect 837 354 887 378
<< nsubdiff >>
rect 2361 412 2411 436
rect 2361 378 2369 412
rect 2403 378 2411 412
rect 2361 354 2411 378
<< psubdiffcont >>
rect 845 378 879 412
<< nsubdiffcont >>
rect 2369 378 2403 412
<< poly >>
rect 44 214 110 230
rect 44 180 60 214
rect 94 212 110 214
rect 94 182 136 212
rect 1588 182 1660 212
rect 94 180 110 182
rect 44 164 110 180
<< polycont >>
rect 60 180 94 214
<< locali >>
rect 845 412 879 428
rect 845 362 879 378
rect 2369 412 2403 428
rect 2369 362 2403 378
rect 845 264 879 280
rect 60 214 94 230
rect 845 214 879 230
rect 2369 264 2403 280
rect 2369 214 2403 230
rect 60 164 94 180
rect 829 130 3122 164
<< viali >>
rect 845 378 879 412
rect 2369 378 2403 412
rect 845 230 879 264
rect 2369 230 2403 264
<< metal1 >>
rect 833 412 891 418
rect 833 378 845 412
rect 879 378 891 412
rect 833 372 891 378
rect 2357 412 2415 418
rect 2357 378 2369 412
rect 2403 378 2415 412
rect 2357 372 2415 378
rect 848 270 876 372
rect 2372 270 2400 372
rect 833 264 891 270
rect 833 230 845 264
rect 879 230 891 264
rect 833 224 891 230
rect 2357 264 2415 270
rect 2357 230 2369 264
rect 2403 230 2415 264
rect 2357 224 2415 230
rect 848 0 876 224
rect 2372 0 2400 224
use contact_7  contact_7_0
timestamp 1644511149
transform 1 0 2357 0 1 214
box 0 0 1 1
use contact_7  contact_7_1
timestamp 1644511149
transform 1 0 833 0 1 214
box 0 0 1 1
use contact_7  contact_7_2
timestamp 1644511149
transform 1 0 833 0 1 362
box 0 0 1 1
use contact_7  contact_7_3
timestamp 1644511149
transform 1 0 2357 0 1 362
box 0 0 1 1
use contact_12  contact_12_0
timestamp 1644511149
transform 1 0 44 0 1 164
box 0 0 1 1
use contact_13  contact_13_0
timestamp 1644511149
transform 1 0 2361 0 1 354
box 0 0 1 1
use contact_18  contact_18_0
timestamp 1644511149
transform 1 0 837 0 1 354
box 0 0 1 1
use nmos_m10_w7_000_sli_dli_da_p  nmos_m10_w7_000_sli_dli_da_p_0
timestamp 1644511149
transform 0 1 162 -1 0 272
box -26 -26 176 1426
use pmos_m10_w7_000_sli_dli_da_p  pmos_m10_w7_000_sli_dli_da_p_0
timestamp 1644511149
transform 0 1 1686 -1 0 272
box -59 -54 209 1454
<< labels >>
rlabel locali s 1975 147 1975 147 4 Z
port 2 nsew
rlabel locali s 77 197 77 197 4 A
port 1 nsew
rlabel metal1 s 2386 197 2386 197 4 vdd
port 3 nsew
rlabel metal1 s 862 197 862 197 4 gnd
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 3122 395
string GDS_END 28274
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 26832
<< end >>
