magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< labels >>
flabel comment s 125 150 125 150 0 FreeSans 300 0 0 0 D
flabel comment s -25 150 -25 150 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7186522
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7185882
<< end >>
