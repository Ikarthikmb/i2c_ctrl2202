magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< obsm1 >>
rect 74152 88980 74210 89026
rect 74342 88980 74400 89026
rect 74603 88980 74661 89026
rect 74953 88980 75011 89026
rect 75214 88980 75272 89026
rect 74164 88638 74198 88980
rect 74226 88737 74292 88789
rect 74354 88786 74388 88980
rect 74342 88740 74400 88786
rect 67462 88560 67520 88606
rect 67723 88560 67781 88606
rect 68073 88560 68131 88606
rect 68334 88560 68392 88606
rect 68524 88560 68582 88606
rect 74148 88586 74214 88638
rect 67474 88366 67508 88560
rect 67462 88320 67520 88366
rect 67474 88046 67508 88320
rect 67575 88237 67641 88289
rect 67539 88200 67597 88206
rect 67735 88200 67769 88560
rect 67807 88446 67861 88455
rect 67805 88400 67863 88446
rect 67807 88391 67861 88400
rect 67539 88166 67769 88200
rect 67539 88160 67597 88166
rect 67735 88046 67769 88166
rect 67817 88135 67851 88391
rect 67807 88126 67861 88135
rect 67805 88080 67863 88126
rect 67807 88071 67861 88080
rect 68085 88046 68119 88560
rect 68346 88366 68380 88560
rect 68334 88320 68392 88366
rect 68346 88046 68380 88320
rect 68442 88317 68508 88369
rect 68536 88218 68570 88560
rect 74164 88466 74198 88586
rect 74354 88466 74388 88740
rect 74615 88466 74649 88980
rect 74873 88866 74927 88875
rect 74871 88820 74929 88866
rect 74873 88811 74927 88820
rect 74883 88555 74917 88811
rect 74965 88620 74999 88980
rect 75226 88786 75260 88980
rect 75214 88740 75272 88786
rect 75093 88657 75159 88709
rect 75137 88620 75195 88626
rect 74965 88586 75195 88620
rect 74873 88546 74927 88555
rect 74871 88500 74929 88546
rect 74873 88491 74927 88500
rect 74965 88466 74999 88586
rect 75137 88580 75195 88586
rect 75226 88466 75260 88740
rect 74152 88420 74210 88466
rect 74342 88420 74400 88466
rect 74603 88420 74661 88466
rect 74953 88420 75011 88466
rect 75214 88420 75272 88466
rect 68520 88166 68586 88218
rect 68536 88046 68570 88166
rect 67462 88000 67520 88046
rect 67723 88000 67781 88046
rect 68073 88000 68131 88046
rect 68334 88000 68392 88046
rect 68524 88000 68582 88046
rect 17812 86099 17858 86353
rect 3350 85804 3408 85850
rect 3611 85804 3669 85850
rect 3961 85804 4019 85850
rect 4222 85804 4280 85850
rect 4412 85804 4470 85850
rect 3362 85530 3396 85804
rect 3427 85684 3485 85690
rect 3623 85684 3657 85804
rect 3695 85770 3749 85779
rect 3693 85724 3751 85770
rect 3695 85715 3749 85724
rect 3427 85650 3657 85684
rect 3427 85644 3485 85650
rect 3463 85561 3529 85613
rect 3350 85484 3408 85530
rect 3362 85290 3396 85484
rect 3623 85290 3657 85650
rect 3705 85459 3739 85715
rect 3695 85450 3749 85459
rect 3693 85404 3751 85450
rect 3695 85395 3749 85404
rect 3973 85290 4007 85804
rect 4234 85530 4268 85804
rect 4424 85684 4458 85804
rect 4408 85632 4474 85684
rect 4222 85484 4280 85530
rect 4234 85290 4268 85484
rect 4330 85481 4396 85533
rect 4424 85290 4458 85632
rect 3350 85244 3408 85290
rect 3611 85244 3669 85290
rect 3961 85244 4019 85290
rect 4222 85244 4280 85290
rect 4412 85244 4470 85290
rect 17904 85269 17938 86353
rect 17980 85269 18008 86353
rect 18066 86208 18112 86282
rect 19060 86099 19106 86353
rect 18066 85885 18112 85961
rect 19152 85269 19186 86353
rect 19228 85269 19256 86353
rect 19314 86208 19360 86282
rect 20308 86099 20354 86353
rect 19314 85885 19360 85961
rect 20400 85269 20434 86353
rect 20476 85269 20504 86353
rect 20562 86208 20608 86282
rect 21556 86099 21602 86353
rect 20562 85885 20608 85961
rect 21648 85269 21682 86353
rect 21724 85269 21752 86353
rect 21810 86208 21856 86282
rect 22804 86099 22850 86353
rect 21810 85885 21856 85961
rect 22896 85269 22930 86353
rect 22972 85269 23000 86353
rect 23058 86208 23104 86282
rect 24052 86099 24098 86353
rect 23058 85885 23104 85961
rect 24144 85269 24178 86353
rect 24220 85269 24248 86353
rect 24306 86208 24352 86282
rect 25300 86099 25346 86353
rect 24306 85885 24352 85961
rect 25392 85269 25426 86353
rect 25468 85269 25496 86353
rect 25554 86208 25600 86282
rect 26548 86099 26594 86353
rect 25554 85885 25600 85961
rect 26640 85269 26674 86353
rect 26716 85269 26744 86353
rect 26802 86208 26848 86282
rect 27796 86099 27842 86353
rect 26802 85885 26848 85961
rect 27888 85269 27922 86353
rect 27964 85269 27992 86353
rect 28050 86208 28096 86282
rect 29044 86099 29090 86353
rect 28050 85885 28096 85961
rect 29136 85269 29170 86353
rect 29212 85269 29240 86353
rect 29298 86208 29344 86282
rect 30292 86099 30338 86353
rect 29298 85885 29344 85961
rect 30384 85269 30418 86353
rect 30460 85269 30488 86353
rect 30546 86208 30592 86282
rect 31540 86099 31586 86353
rect 30546 85885 30592 85961
rect 31632 85269 31666 86353
rect 31708 85269 31736 86353
rect 31794 86208 31840 86282
rect 32788 86099 32834 86353
rect 31794 85885 31840 85961
rect 32880 85269 32914 86353
rect 32956 85269 32984 86353
rect 33042 86208 33088 86282
rect 34036 86099 34082 86353
rect 33042 85885 33088 85961
rect 34128 85269 34162 86353
rect 34204 85269 34232 86353
rect 34290 86208 34336 86282
rect 35284 86099 35330 86353
rect 34290 85885 34336 85961
rect 35376 85269 35410 86353
rect 35452 85269 35480 86353
rect 35538 86208 35584 86282
rect 36532 86099 36578 86353
rect 35538 85885 35584 85961
rect 36624 85269 36658 86353
rect 36700 85269 36728 86353
rect 36786 86208 36832 86282
rect 37780 86099 37826 86353
rect 36786 85885 36832 85961
rect 37872 85269 37906 86353
rect 37948 85269 37976 86353
rect 38034 86208 38080 86282
rect 39028 86099 39074 86353
rect 38034 85885 38080 85961
rect 39120 85269 39154 86353
rect 39196 85269 39224 86353
rect 39282 86208 39328 86282
rect 40276 86099 40322 86353
rect 39282 85885 39328 85961
rect 40368 85269 40402 86353
rect 40444 85269 40472 86353
rect 40530 86208 40576 86282
rect 41524 86099 41570 86353
rect 40530 85885 40576 85961
rect 41616 85269 41650 86353
rect 41692 85269 41720 86353
rect 41778 86208 41824 86282
rect 42772 86099 42818 86353
rect 41778 85885 41824 85961
rect 42864 85269 42898 86353
rect 42940 85269 42968 86353
rect 43026 86208 43072 86282
rect 44020 86099 44066 86353
rect 43026 85885 43072 85961
rect 44112 85269 44146 86353
rect 44188 85269 44216 86353
rect 44274 86208 44320 86282
rect 45268 86099 45314 86353
rect 44274 85885 44320 85961
rect 45360 85269 45394 86353
rect 45436 85269 45464 86353
rect 45522 86208 45568 86282
rect 46516 86099 46562 86353
rect 45522 85885 45568 85961
rect 46608 85269 46642 86353
rect 46684 85269 46712 86353
rect 46770 86208 46816 86282
rect 47764 86099 47810 86353
rect 46770 85885 46816 85961
rect 47856 85269 47890 86353
rect 47932 85269 47960 86353
rect 48018 86208 48064 86282
rect 49012 86099 49058 86353
rect 48018 85885 48064 85961
rect 49104 85269 49138 86353
rect 49180 85269 49208 86353
rect 49266 86208 49312 86282
rect 50260 86099 50306 86353
rect 49266 85885 49312 85961
rect 50352 85269 50386 86353
rect 50428 85269 50456 86353
rect 50514 86208 50560 86282
rect 51508 86099 51554 86353
rect 50514 85885 50560 85961
rect 51600 85269 51634 86353
rect 51676 85269 51704 86353
rect 51762 86208 51808 86282
rect 52756 86099 52802 86353
rect 51762 85885 51808 85961
rect 52848 85269 52882 86353
rect 52924 85269 52952 86353
rect 53010 86208 53056 86282
rect 54004 86099 54050 86353
rect 53010 85885 53056 85961
rect 54096 85269 54130 86353
rect 54172 85269 54200 86353
rect 54258 86208 54304 86282
rect 55252 86099 55298 86353
rect 54258 85885 54304 85961
rect 55344 85269 55378 86353
rect 55420 85269 55448 86353
rect 55506 86208 55552 86282
rect 56500 86099 56546 86353
rect 55506 85885 55552 85961
rect 56592 85269 56626 86353
rect 56668 85269 56696 86353
rect 56754 86208 56800 86282
rect 56754 85885 56800 85961
rect 17892 85223 17950 85269
rect 3350 84756 3408 84802
rect 3611 84756 3669 84802
rect 3961 84756 4019 84802
rect 4222 84756 4280 84802
rect 4412 84756 4470 84802
rect 3362 84562 3396 84756
rect 3350 84516 3408 84562
rect 3362 84242 3396 84516
rect 3463 84433 3529 84485
rect 3427 84396 3485 84402
rect 3623 84396 3657 84756
rect 3695 84642 3749 84651
rect 3693 84596 3751 84642
rect 3695 84587 3749 84596
rect 3427 84362 3657 84396
rect 3427 84356 3485 84362
rect 3623 84242 3657 84362
rect 3705 84331 3739 84587
rect 3695 84322 3749 84331
rect 3693 84276 3751 84322
rect 3695 84267 3749 84276
rect 3973 84242 4007 84756
rect 4234 84562 4268 84756
rect 4222 84516 4280 84562
rect 4234 84242 4268 84516
rect 4330 84513 4396 84565
rect 4424 84414 4458 84756
rect 4408 84362 4474 84414
rect 4424 84242 4458 84362
rect 3350 84196 3408 84242
rect 3611 84196 3669 84242
rect 3961 84196 4019 84242
rect 4222 84196 4280 84242
rect 4412 84196 4470 84242
rect 17802 84129 17860 84189
rect 17904 84097 17938 85223
rect 17980 85211 18048 85269
rect 19140 85223 19198 85269
rect 17980 84097 18008 85211
rect 18046 85051 18108 85119
rect 18136 84274 18182 84348
rect 19050 84129 19108 84189
rect 19152 84097 19186 85223
rect 19228 85211 19296 85269
rect 20388 85223 20446 85269
rect 19228 84097 19256 85211
rect 19294 85051 19356 85119
rect 19384 84274 19430 84348
rect 20298 84129 20356 84189
rect 20400 84097 20434 85223
rect 20476 85211 20544 85269
rect 21636 85223 21694 85269
rect 20476 84097 20504 85211
rect 20542 85051 20604 85119
rect 20632 84274 20678 84348
rect 21546 84129 21604 84189
rect 21648 84097 21682 85223
rect 21724 85211 21792 85269
rect 22884 85223 22942 85269
rect 21724 84097 21752 85211
rect 21790 85051 21852 85119
rect 21880 84274 21926 84348
rect 22794 84129 22852 84189
rect 22896 84097 22930 85223
rect 22972 85211 23040 85269
rect 24132 85223 24190 85269
rect 22972 84097 23000 85211
rect 23038 85051 23100 85119
rect 23128 84274 23174 84348
rect 24042 84129 24100 84189
rect 24144 84097 24178 85223
rect 24220 85211 24288 85269
rect 25380 85223 25438 85269
rect 24220 84097 24248 85211
rect 24286 85051 24348 85119
rect 24376 84274 24422 84348
rect 25290 84129 25348 84189
rect 25392 84097 25426 85223
rect 25468 85211 25536 85269
rect 26628 85223 26686 85269
rect 25468 84097 25496 85211
rect 25534 85051 25596 85119
rect 25624 84274 25670 84348
rect 26538 84129 26596 84189
rect 26640 84097 26674 85223
rect 26716 85211 26784 85269
rect 27876 85223 27934 85269
rect 26716 84097 26744 85211
rect 26782 85051 26844 85119
rect 26872 84274 26918 84348
rect 27786 84129 27844 84189
rect 27888 84097 27922 85223
rect 27964 85211 28032 85269
rect 29124 85223 29182 85269
rect 27964 84097 27992 85211
rect 28030 85051 28092 85119
rect 28120 84274 28166 84348
rect 29034 84129 29092 84189
rect 29136 84097 29170 85223
rect 29212 85211 29280 85269
rect 30372 85223 30430 85269
rect 29212 84097 29240 85211
rect 29278 85051 29340 85119
rect 29368 84274 29414 84348
rect 30282 84129 30340 84189
rect 30384 84097 30418 85223
rect 30460 85211 30528 85269
rect 31620 85223 31678 85269
rect 30460 84097 30488 85211
rect 30526 85051 30588 85119
rect 30616 84274 30662 84348
rect 31530 84129 31588 84189
rect 31632 84097 31666 85223
rect 31708 85211 31776 85269
rect 32868 85223 32926 85269
rect 31708 84097 31736 85211
rect 31774 85051 31836 85119
rect 31864 84274 31910 84348
rect 32778 84129 32836 84189
rect 32880 84097 32914 85223
rect 32956 85211 33024 85269
rect 34116 85223 34174 85269
rect 32956 84097 32984 85211
rect 33022 85051 33084 85119
rect 33112 84274 33158 84348
rect 34026 84129 34084 84189
rect 34128 84097 34162 85223
rect 34204 85211 34272 85269
rect 35364 85223 35422 85269
rect 34204 84097 34232 85211
rect 34270 85051 34332 85119
rect 34360 84274 34406 84348
rect 35274 84129 35332 84189
rect 35376 84097 35410 85223
rect 35452 85211 35520 85269
rect 36612 85223 36670 85269
rect 35452 84097 35480 85211
rect 35518 85051 35580 85119
rect 35608 84274 35654 84348
rect 36522 84129 36580 84189
rect 36624 84097 36658 85223
rect 36700 85211 36768 85269
rect 37860 85223 37918 85269
rect 36700 84097 36728 85211
rect 36766 85051 36828 85119
rect 36856 84274 36902 84348
rect 37770 84129 37828 84189
rect 37872 84097 37906 85223
rect 37948 85211 38016 85269
rect 39108 85223 39166 85269
rect 37948 84097 37976 85211
rect 38014 85051 38076 85119
rect 38104 84274 38150 84348
rect 39018 84129 39076 84189
rect 39120 84097 39154 85223
rect 39196 85211 39264 85269
rect 40356 85223 40414 85269
rect 39196 84097 39224 85211
rect 39262 85051 39324 85119
rect 39352 84274 39398 84348
rect 40266 84129 40324 84189
rect 40368 84097 40402 85223
rect 40444 85211 40512 85269
rect 41604 85223 41662 85269
rect 40444 84097 40472 85211
rect 40510 85051 40572 85119
rect 40600 84274 40646 84348
rect 41514 84129 41572 84189
rect 41616 84097 41650 85223
rect 41692 85211 41760 85269
rect 42852 85223 42910 85269
rect 41692 84097 41720 85211
rect 41758 85051 41820 85119
rect 41848 84274 41894 84348
rect 42762 84129 42820 84189
rect 42864 84097 42898 85223
rect 42940 85211 43008 85269
rect 44100 85223 44158 85269
rect 42940 84097 42968 85211
rect 43006 85051 43068 85119
rect 43096 84274 43142 84348
rect 44010 84129 44068 84189
rect 44112 84097 44146 85223
rect 44188 85211 44256 85269
rect 45348 85223 45406 85269
rect 44188 84097 44216 85211
rect 44254 85051 44316 85119
rect 44344 84274 44390 84348
rect 45258 84129 45316 84189
rect 45360 84097 45394 85223
rect 45436 85211 45504 85269
rect 46596 85223 46654 85269
rect 45436 84097 45464 85211
rect 45502 85051 45564 85119
rect 45592 84274 45638 84348
rect 46506 84129 46564 84189
rect 46608 84097 46642 85223
rect 46684 85211 46752 85269
rect 47844 85223 47902 85269
rect 46684 84097 46712 85211
rect 46750 85051 46812 85119
rect 46840 84274 46886 84348
rect 47754 84129 47812 84189
rect 47856 84097 47890 85223
rect 47932 85211 48000 85269
rect 49092 85223 49150 85269
rect 47932 84097 47960 85211
rect 47998 85051 48060 85119
rect 48088 84274 48134 84348
rect 49002 84129 49060 84189
rect 49104 84097 49138 85223
rect 49180 85211 49248 85269
rect 50340 85223 50398 85269
rect 49180 84097 49208 85211
rect 49246 85051 49308 85119
rect 49336 84274 49382 84348
rect 50250 84129 50308 84189
rect 50352 84097 50386 85223
rect 50428 85211 50496 85269
rect 51588 85223 51646 85269
rect 50428 84097 50456 85211
rect 50494 85051 50556 85119
rect 50584 84274 50630 84348
rect 51498 84129 51556 84189
rect 51600 84097 51634 85223
rect 51676 85211 51744 85269
rect 52836 85223 52894 85269
rect 51676 84097 51704 85211
rect 51742 85051 51804 85119
rect 51832 84274 51878 84348
rect 52746 84129 52804 84189
rect 52848 84097 52882 85223
rect 52924 85211 52992 85269
rect 54084 85223 54142 85269
rect 52924 84097 52952 85211
rect 52990 85051 53052 85119
rect 53080 84274 53126 84348
rect 53994 84129 54052 84189
rect 54096 84097 54130 85223
rect 54172 85211 54240 85269
rect 55332 85223 55390 85269
rect 54172 84097 54200 85211
rect 54238 85051 54300 85119
rect 54328 84274 54374 84348
rect 55242 84129 55300 84189
rect 55344 84097 55378 85223
rect 55420 85211 55488 85269
rect 56580 85223 56638 85269
rect 55420 84097 55448 85211
rect 55486 85051 55548 85119
rect 55576 84274 55622 84348
rect 56490 84129 56548 84189
rect 56592 84097 56626 85223
rect 56668 85211 56736 85269
rect 56668 84097 56696 85211
rect 56734 85051 56796 85119
rect 56824 84274 56870 84348
rect 17788 83169 17816 83597
rect 18252 83169 18280 83721
rect 18384 83169 18412 83225
rect 18848 83169 18876 83225
rect 19036 83169 19064 83597
rect 19500 83169 19528 83721
rect 19632 83169 19660 83225
rect 20096 83169 20124 83225
rect 20284 83169 20312 83597
rect 20748 83169 20776 83721
rect 20880 83169 20908 83225
rect 21344 83169 21372 83225
rect 21532 83169 21560 83597
rect 21996 83169 22024 83721
rect 22128 83169 22156 83225
rect 22592 83169 22620 83225
rect 22780 83169 22808 83597
rect 23244 83169 23272 83721
rect 23376 83169 23404 83225
rect 23840 83169 23868 83225
rect 24028 83169 24056 83597
rect 24492 83169 24520 83721
rect 24624 83169 24652 83225
rect 25088 83169 25116 83225
rect 25276 83169 25304 83597
rect 25740 83169 25768 83721
rect 25872 83169 25900 83225
rect 26336 83169 26364 83225
rect 26524 83169 26552 83597
rect 26988 83169 27016 83721
rect 27120 83169 27148 83225
rect 27584 83169 27612 83225
rect 27772 83169 27800 83597
rect 28236 83169 28264 83721
rect 28368 83169 28396 83225
rect 28832 83169 28860 83225
rect 29020 83169 29048 83597
rect 29484 83169 29512 83721
rect 29616 83169 29644 83225
rect 30080 83169 30108 83225
rect 30268 83169 30296 83597
rect 30732 83169 30760 83721
rect 30864 83169 30892 83225
rect 31328 83169 31356 83225
rect 31516 83169 31544 83597
rect 31980 83169 32008 83721
rect 32112 83169 32140 83225
rect 32576 83169 32604 83225
rect 32764 83169 32792 83597
rect 33228 83169 33256 83721
rect 33360 83169 33388 83225
rect 33824 83169 33852 83225
rect 34012 83169 34040 83597
rect 34476 83169 34504 83721
rect 34608 83169 34636 83225
rect 35072 83169 35100 83225
rect 35260 83169 35288 83597
rect 35724 83169 35752 83721
rect 35856 83169 35884 83225
rect 36320 83169 36348 83225
rect 36508 83169 36536 83597
rect 36972 83169 37000 83721
rect 37104 83169 37132 83225
rect 37568 83169 37596 83225
rect 37756 83169 37784 83597
rect 38220 83169 38248 83721
rect 38352 83169 38380 83225
rect 38816 83169 38844 83225
rect 39004 83169 39032 83597
rect 39468 83169 39496 83721
rect 39600 83169 39628 83225
rect 40064 83169 40092 83225
rect 40252 83169 40280 83597
rect 40716 83169 40744 83721
rect 40848 83169 40876 83225
rect 41312 83169 41340 83225
rect 41500 83169 41528 83597
rect 41964 83169 41992 83721
rect 42096 83169 42124 83225
rect 42560 83169 42588 83225
rect 42748 83169 42776 83597
rect 43212 83169 43240 83721
rect 43344 83169 43372 83225
rect 43808 83169 43836 83225
rect 43996 83169 44024 83597
rect 44460 83169 44488 83721
rect 44592 83169 44620 83225
rect 45056 83169 45084 83225
rect 45244 83169 45272 83597
rect 45708 83169 45736 83721
rect 45840 83169 45868 83225
rect 46304 83169 46332 83225
rect 46492 83169 46520 83597
rect 46956 83169 46984 83721
rect 47088 83169 47116 83225
rect 47552 83169 47580 83225
rect 47740 83169 47768 83597
rect 48204 83169 48232 83721
rect 48336 83169 48364 83225
rect 48800 83169 48828 83225
rect 48988 83169 49016 83597
rect 49452 83169 49480 83721
rect 49584 83169 49612 83225
rect 50048 83169 50076 83225
rect 50236 83169 50264 83597
rect 50700 83169 50728 83721
rect 50832 83169 50860 83225
rect 51296 83169 51324 83225
rect 51484 83169 51512 83597
rect 51948 83169 51976 83721
rect 52080 83169 52108 83225
rect 52544 83169 52572 83225
rect 52732 83169 52760 83597
rect 53196 83169 53224 83721
rect 53328 83169 53356 83225
rect 53792 83169 53820 83225
rect 53980 83169 54008 83597
rect 54444 83169 54472 83721
rect 54576 83169 54604 83225
rect 55040 83169 55068 83225
rect 55228 83169 55256 83597
rect 55692 83169 55720 83721
rect 55824 83169 55852 83225
rect 56288 83169 56316 83225
rect 56476 83169 56504 83597
rect 56940 83169 56968 83721
rect 57072 83169 57100 83225
rect 57536 83169 57564 83225
rect 3350 82976 3408 83022
rect 3611 82976 3669 83022
rect 3961 82976 4019 83022
rect 4222 82976 4280 83022
rect 4412 82976 4470 83022
rect 3362 82702 3396 82976
rect 3427 82856 3485 82862
rect 3623 82856 3657 82976
rect 3695 82942 3749 82951
rect 3693 82896 3751 82942
rect 3695 82887 3749 82896
rect 3427 82822 3657 82856
rect 3427 82816 3485 82822
rect 3463 82733 3529 82785
rect 3350 82656 3408 82702
rect 3362 82462 3396 82656
rect 3623 82462 3657 82822
rect 3705 82631 3739 82887
rect 3695 82622 3749 82631
rect 3693 82576 3751 82622
rect 3695 82567 3749 82576
rect 3973 82462 4007 82976
rect 4234 82702 4268 82976
rect 4424 82856 4458 82976
rect 4408 82804 4474 82856
rect 4222 82656 4280 82702
rect 4234 82462 4268 82656
rect 4330 82653 4396 82705
rect 4424 82462 4458 82804
rect 3350 82416 3408 82462
rect 3611 82416 3669 82462
rect 3961 82416 4019 82462
rect 4222 82416 4280 82462
rect 4412 82416 4470 82462
rect 3350 81928 3408 81974
rect 3611 81928 3669 81974
rect 3961 81928 4019 81974
rect 4222 81928 4280 81974
rect 4412 81928 4470 81974
rect 3362 81734 3396 81928
rect 3350 81688 3408 81734
rect 3362 81414 3396 81688
rect 3463 81605 3529 81657
rect 3427 81568 3485 81574
rect 3623 81568 3657 81928
rect 3695 81814 3749 81823
rect 3693 81768 3751 81814
rect 3695 81759 3749 81768
rect 3427 81534 3657 81568
rect 3427 81528 3485 81534
rect 3623 81414 3657 81534
rect 3705 81503 3739 81759
rect 3695 81494 3749 81503
rect 3693 81448 3751 81494
rect 3695 81439 3749 81448
rect 3973 81414 4007 81928
rect 4234 81734 4268 81928
rect 4222 81688 4280 81734
rect 4234 81414 4268 81688
rect 4330 81685 4396 81737
rect 4424 81586 4458 81928
rect 17788 81861 17816 81917
rect 18252 81861 18280 81917
rect 18384 81861 18412 81917
rect 18848 81861 18876 81917
rect 19036 81861 19064 81917
rect 19500 81861 19528 81917
rect 19632 81861 19660 81917
rect 20096 81861 20124 81917
rect 20284 81861 20312 81917
rect 20748 81861 20776 81917
rect 20880 81861 20908 81917
rect 21344 81861 21372 81917
rect 21532 81861 21560 81917
rect 21996 81861 22024 81917
rect 22128 81861 22156 81917
rect 22592 81861 22620 81917
rect 22780 81861 22808 81917
rect 23244 81861 23272 81917
rect 23376 81861 23404 81917
rect 23840 81861 23868 81917
rect 24028 81861 24056 81917
rect 24492 81861 24520 81917
rect 24624 81861 24652 81917
rect 25088 81861 25116 81917
rect 25276 81861 25304 81917
rect 25740 81861 25768 81917
rect 25872 81861 25900 81917
rect 26336 81861 26364 81917
rect 26524 81861 26552 81917
rect 26988 81861 27016 81917
rect 27120 81861 27148 81917
rect 27584 81861 27612 81917
rect 27772 81861 27800 81917
rect 28236 81861 28264 81917
rect 28368 81861 28396 81917
rect 28832 81861 28860 81917
rect 29020 81861 29048 81917
rect 29484 81861 29512 81917
rect 29616 81861 29644 81917
rect 30080 81861 30108 81917
rect 30268 81861 30296 81917
rect 30732 81861 30760 81917
rect 30864 81861 30892 81917
rect 31328 81861 31356 81917
rect 31516 81861 31544 81917
rect 31980 81861 32008 81917
rect 32112 81861 32140 81917
rect 32576 81861 32604 81917
rect 32764 81861 32792 81917
rect 33228 81861 33256 81917
rect 33360 81861 33388 81917
rect 33824 81861 33852 81917
rect 34012 81861 34040 81917
rect 34476 81861 34504 81917
rect 34608 81861 34636 81917
rect 35072 81861 35100 81917
rect 35260 81861 35288 81917
rect 35724 81861 35752 81917
rect 35856 81861 35884 81917
rect 36320 81861 36348 81917
rect 36508 81861 36536 81917
rect 36972 81861 37000 81917
rect 37104 81861 37132 81917
rect 37568 81861 37596 81917
rect 37756 81861 37784 81917
rect 38220 81861 38248 81917
rect 38352 81861 38380 81917
rect 38816 81861 38844 81917
rect 39004 81861 39032 81917
rect 39468 81861 39496 81917
rect 39600 81861 39628 81917
rect 40064 81861 40092 81917
rect 40252 81861 40280 81917
rect 40716 81861 40744 81917
rect 40848 81861 40876 81917
rect 41312 81861 41340 81917
rect 41500 81861 41528 81917
rect 41964 81861 41992 81917
rect 42096 81861 42124 81917
rect 42560 81861 42588 81917
rect 42748 81861 42776 81917
rect 43212 81861 43240 81917
rect 43344 81861 43372 81917
rect 43808 81861 43836 81917
rect 43996 81861 44024 81917
rect 44460 81861 44488 81917
rect 44592 81861 44620 81917
rect 45056 81861 45084 81917
rect 45244 81861 45272 81917
rect 45708 81861 45736 81917
rect 45840 81861 45868 81917
rect 46304 81861 46332 81917
rect 46492 81861 46520 81917
rect 46956 81861 46984 81917
rect 47088 81861 47116 81917
rect 47552 81861 47580 81917
rect 47740 81861 47768 81917
rect 48204 81861 48232 81917
rect 48336 81861 48364 81917
rect 48800 81861 48828 81917
rect 48988 81861 49016 81917
rect 49452 81861 49480 81917
rect 49584 81861 49612 81917
rect 50048 81861 50076 81917
rect 50236 81861 50264 81917
rect 50700 81861 50728 81917
rect 50832 81861 50860 81917
rect 51296 81861 51324 81917
rect 51484 81861 51512 81917
rect 51948 81861 51976 81917
rect 52080 81861 52108 81917
rect 52544 81861 52572 81917
rect 52732 81861 52760 81917
rect 53196 81861 53224 81917
rect 53328 81861 53356 81917
rect 53792 81861 53820 81917
rect 53980 81861 54008 81917
rect 54444 81861 54472 81917
rect 54576 81861 54604 81917
rect 55040 81861 55068 81917
rect 55228 81861 55256 81917
rect 55692 81861 55720 81917
rect 55824 81861 55852 81917
rect 56288 81861 56316 81917
rect 56476 81861 56504 81917
rect 56940 81861 56968 81917
rect 57072 81861 57100 81917
rect 57536 81861 57564 81917
rect 4408 81534 4474 81586
rect 4424 81414 4458 81534
rect 3350 81368 3408 81414
rect 3611 81368 3669 81414
rect 3961 81368 4019 81414
rect 4222 81368 4280 81414
rect 4412 81368 4470 81414
rect 17774 80855 17802 81609
rect 18238 80855 18266 81609
rect 18398 80855 18426 81609
rect 18862 80855 18890 81609
rect 19022 80855 19050 81609
rect 19486 80855 19514 81609
rect 19646 80855 19674 81609
rect 20110 80855 20138 81609
rect 20270 80855 20298 81609
rect 20734 80855 20762 81609
rect 20894 80855 20922 81609
rect 21358 80855 21386 81609
rect 21518 80855 21546 81609
rect 21982 80855 22010 81609
rect 22142 80855 22170 81609
rect 22606 80855 22634 81609
rect 22766 80855 22794 81609
rect 23230 80855 23258 81609
rect 23390 80855 23418 81609
rect 23854 80855 23882 81609
rect 24014 80855 24042 81609
rect 24478 80855 24506 81609
rect 24638 80855 24666 81609
rect 25102 80855 25130 81609
rect 25262 80855 25290 81609
rect 25726 80855 25754 81609
rect 25886 80855 25914 81609
rect 26350 80855 26378 81609
rect 26510 80855 26538 81609
rect 26974 80855 27002 81609
rect 27134 80855 27162 81609
rect 27598 80855 27626 81609
rect 27758 80855 27786 81609
rect 28222 80855 28250 81609
rect 28382 80855 28410 81609
rect 28846 80855 28874 81609
rect 29006 80855 29034 81609
rect 29470 80855 29498 81609
rect 29630 80855 29658 81609
rect 30094 80855 30122 81609
rect 30254 80855 30282 81609
rect 30718 80855 30746 81609
rect 30878 80855 30906 81609
rect 31342 80855 31370 81609
rect 31502 80855 31530 81609
rect 31966 80855 31994 81609
rect 32126 80855 32154 81609
rect 32590 80855 32618 81609
rect 32750 80855 32778 81609
rect 33214 80855 33242 81609
rect 33374 80855 33402 81609
rect 33838 80855 33866 81609
rect 33998 80855 34026 81609
rect 34462 80855 34490 81609
rect 34622 80855 34650 81609
rect 35086 80855 35114 81609
rect 35246 80855 35274 81609
rect 35710 80855 35738 81609
rect 35870 80855 35898 81609
rect 36334 80855 36362 81609
rect 36494 80855 36522 81609
rect 36958 80855 36986 81609
rect 37118 80855 37146 81609
rect 37582 80855 37610 81609
rect 37742 80855 37770 81609
rect 38206 80855 38234 81609
rect 38366 80855 38394 81609
rect 38830 80855 38858 81609
rect 38990 80855 39018 81609
rect 39454 80855 39482 81609
rect 39614 80855 39642 81609
rect 40078 80855 40106 81609
rect 40238 80855 40266 81609
rect 40702 80855 40730 81609
rect 40862 80855 40890 81609
rect 41326 80855 41354 81609
rect 41486 80855 41514 81609
rect 41950 80855 41978 81609
rect 42110 80855 42138 81609
rect 42574 80855 42602 81609
rect 42734 80855 42762 81609
rect 43198 80855 43226 81609
rect 43358 80855 43386 81609
rect 43822 80855 43850 81609
rect 43982 80855 44010 81609
rect 44446 80855 44474 81609
rect 44606 80855 44634 81609
rect 45070 80855 45098 81609
rect 45230 80855 45258 81609
rect 45694 80855 45722 81609
rect 45854 80855 45882 81609
rect 46318 80855 46346 81609
rect 46478 80855 46506 81609
rect 46942 80855 46970 81609
rect 47102 80855 47130 81609
rect 47566 80855 47594 81609
rect 47726 80855 47754 81609
rect 48190 80855 48218 81609
rect 48350 80855 48378 81609
rect 48814 80855 48842 81609
rect 48974 80855 49002 81609
rect 49438 80855 49466 81609
rect 49598 80855 49626 81609
rect 50062 80855 50090 81609
rect 50222 80855 50250 81609
rect 50686 80855 50714 81609
rect 50846 80855 50874 81609
rect 51310 80855 51338 81609
rect 51470 80855 51498 81609
rect 51934 80855 51962 81609
rect 52094 80855 52122 81609
rect 52558 80855 52586 81609
rect 52718 80855 52746 81609
rect 53182 80855 53210 81609
rect 53342 80855 53370 81609
rect 53806 80855 53834 81609
rect 53966 80855 53994 81609
rect 54430 80855 54458 81609
rect 54590 80855 54618 81609
rect 55054 80855 55082 81609
rect 55214 80855 55242 81609
rect 55678 80855 55706 81609
rect 55838 80855 55866 81609
rect 56302 80855 56330 81609
rect 56462 80855 56490 81609
rect 56926 80855 56954 81609
rect 57086 80855 57114 81609
rect 57550 80855 57578 81609
rect 57710 80855 57738 81609
rect 58174 80855 58202 81609
rect 3350 80148 3408 80194
rect 3611 80148 3669 80194
rect 3961 80148 4019 80194
rect 4222 80148 4280 80194
rect 4412 80148 4470 80194
rect 3362 79874 3396 80148
rect 3427 80028 3485 80034
rect 3623 80028 3657 80148
rect 3695 80114 3749 80123
rect 3693 80068 3751 80114
rect 3695 80059 3749 80068
rect 3427 79994 3657 80028
rect 3427 79988 3485 79994
rect 3463 79905 3529 79957
rect 3350 79828 3408 79874
rect 3362 79634 3396 79828
rect 3623 79634 3657 79994
rect 3705 79803 3739 80059
rect 3695 79794 3749 79803
rect 3693 79748 3751 79794
rect 3695 79739 3749 79748
rect 3973 79634 4007 80148
rect 4234 79874 4268 80148
rect 4424 80028 4458 80148
rect 17084 80091 17141 80233
rect 17177 80124 17270 80190
tri 17177 80108 17193 80124 ne
rect 17193 80108 17270 80124
rect 4408 79976 4474 80028
rect 17084 80009 17158 80091
rect 4222 79828 4280 79874
rect 4234 79634 4268 79828
rect 4330 79825 4396 79877
rect 4424 79634 4458 79976
rect 3350 79588 3408 79634
rect 3611 79588 3669 79634
rect 3961 79588 4019 79634
rect 4222 79588 4280 79634
rect 4412 79588 4470 79634
rect 3350 79100 3408 79146
rect 3611 79100 3669 79146
rect 3961 79100 4019 79146
rect 4222 79100 4280 79146
rect 4412 79100 4470 79146
rect 3362 78906 3396 79100
rect 3350 78860 3408 78906
rect 3362 78586 3396 78860
rect 3463 78777 3529 78829
rect 3427 78740 3485 78746
rect 3623 78740 3657 79100
rect 3695 78986 3749 78995
rect 3693 78940 3751 78986
rect 3695 78931 3749 78940
rect 3427 78706 3657 78740
rect 3427 78700 3485 78706
rect 3623 78586 3657 78706
rect 3705 78675 3739 78931
rect 3695 78666 3749 78675
rect 3693 78620 3751 78666
rect 3695 78611 3749 78620
rect 3973 78586 4007 79100
rect 4234 78906 4268 79100
rect 4222 78860 4280 78906
rect 4234 78586 4268 78860
rect 4330 78857 4396 78909
rect 4424 78758 4458 79100
rect 4408 78706 4474 78758
rect 4424 78586 4458 78706
rect 3350 78540 3408 78586
rect 3611 78540 3669 78586
rect 3961 78540 4019 78586
rect 4222 78540 4280 78586
rect 4412 78540 4470 78586
rect 3350 77320 3408 77366
rect 3611 77320 3669 77366
rect 3961 77320 4019 77366
rect 4222 77320 4280 77366
rect 4412 77320 4470 77366
rect 3362 77046 3396 77320
rect 3427 77200 3485 77206
rect 3623 77200 3657 77320
rect 3695 77286 3749 77295
rect 3693 77240 3751 77286
rect 3695 77231 3749 77240
rect 3427 77166 3657 77200
rect 3427 77160 3485 77166
rect 3463 77077 3529 77129
rect 3350 77000 3408 77046
rect 3362 76806 3396 77000
rect 3623 76806 3657 77166
rect 3705 76975 3739 77231
rect 3695 76966 3749 76975
rect 3693 76920 3751 76966
rect 3695 76911 3749 76920
rect 3973 76806 4007 77320
rect 4234 77046 4268 77320
rect 4424 77200 4458 77320
rect 4408 77148 4474 77200
rect 4222 77000 4280 77046
rect 4234 76806 4268 77000
rect 4330 76997 4396 77049
rect 4424 76806 4458 77148
rect 3350 76760 3408 76806
rect 3611 76760 3669 76806
rect 3961 76760 4019 76806
rect 4222 76760 4280 76806
rect 4412 76760 4470 76806
rect 4680 29282 4708 37182
rect 4760 29282 4788 37182
rect 4840 29282 4868 37182
rect 4920 29282 4948 37182
rect 5000 29282 5028 37182
rect 5080 29282 5108 37182
rect 5160 29282 5188 37182
rect 5496 34977 5548 35041
rect 5416 34583 5468 34647
rect 5336 34187 5388 34251
rect 5852 34022 5880 35207
rect 6124 34022 6152 35207
rect 7174 33978 7220 37226
rect 7598 36406 7646 37168
rect 8030 36406 8078 37168
rect 7598 35616 7646 36378
rect 8030 35616 8078 36378
rect 7598 34826 7646 35588
rect 8030 34826 8078 35588
rect 7598 34036 7646 34798
rect 8030 34036 8078 34798
rect 8422 34022 8450 37182
rect 8694 34022 8722 37182
rect 6092 32213 6144 32277
rect 6012 31817 6064 31881
rect 6448 31652 6476 32442
rect 6720 31652 6748 32442
rect 7608 31622 7656 33262
rect 8032 31620 8082 33264
rect 8422 31652 8450 33232
rect 8694 31652 8722 33232
rect 6092 29843 6144 29907
rect 6012 29447 6064 29511
rect 6448 29282 6476 30072
rect 6720 29282 6748 30072
rect 7608 29252 7656 30892
rect 8032 29250 8082 30894
rect 8422 29282 8450 30862
rect 8694 29282 8722 30862
rect 10464 29238 10510 79886
rect 17084 79851 17141 80009
tri 17177 79976 17193 79992 se
rect 17193 79976 17270 79992
rect 17177 79910 17270 79976
rect 10888 79066 10936 79828
rect 11320 79066 11368 79828
rect 10888 78276 10936 79038
rect 11320 78276 11368 79038
rect 10888 77486 10936 78248
rect 11320 77486 11368 78248
rect 10888 76696 10936 77458
rect 11320 76696 11368 77458
rect 10888 75906 10936 76668
rect 11320 75906 11368 76668
rect 10888 75116 10936 75878
rect 11320 75116 11368 75878
rect 10888 74326 10936 75088
rect 11320 74326 11368 75088
rect 10888 73536 10936 74298
rect 11320 73536 11368 74298
rect 10888 72746 10936 73508
rect 11320 72746 11368 73508
rect 10888 71956 10936 72718
rect 11320 71956 11368 72718
rect 10888 71166 10936 71928
rect 11320 71166 11368 71928
rect 10888 70376 10936 71138
rect 11320 70376 11368 71138
rect 10888 69586 10936 70348
rect 11320 69586 11368 70348
rect 10888 68796 10936 69558
rect 11320 68796 11368 69558
rect 10888 68006 10936 68768
rect 11320 68006 11368 68768
rect 10888 67216 10936 67978
rect 11320 67216 11368 67978
rect 10888 66426 10936 67188
rect 11320 66426 11368 67188
rect 10888 65636 10936 66398
rect 11320 65636 11368 66398
rect 10888 64846 10936 65608
rect 11320 64846 11368 65608
rect 10888 64056 10936 64818
rect 11320 64056 11368 64818
rect 10888 63266 10936 64028
rect 11320 63266 11368 64028
rect 10888 62476 10936 63238
rect 11320 62476 11368 63238
rect 10888 61686 10936 62448
rect 11320 61686 11368 62448
rect 10888 60896 10936 61658
rect 11320 60896 11368 61658
rect 10888 60106 10936 60868
rect 11320 60106 11368 60868
rect 10888 59316 10936 60078
rect 11320 59316 11368 60078
rect 10888 58526 10936 59288
rect 11320 58526 11368 59288
rect 10888 57736 10936 58498
rect 11320 57736 11368 58498
rect 10888 56946 10936 57708
rect 11320 56946 11368 57708
rect 10888 56156 10936 56918
rect 11320 56156 11368 56918
rect 10888 55366 10936 56128
rect 11320 55366 11368 56128
rect 10888 54576 10936 55338
rect 11320 54576 11368 55338
rect 10888 53786 10936 54548
rect 11320 53786 11368 54548
rect 10888 52996 10936 53758
rect 11320 52996 11368 53758
rect 10888 52206 10936 52968
rect 11320 52206 11368 52968
rect 10888 51416 10936 52178
rect 11320 51416 11368 52178
rect 10888 50626 10936 51388
rect 11320 50626 11368 51388
rect 10888 49836 10936 50598
rect 11320 49836 11368 50598
rect 10888 49046 10936 49808
rect 11320 49046 11368 49808
rect 10888 48256 10936 49018
rect 11320 48256 11368 49018
rect 10888 47466 10936 48228
rect 11320 47466 11368 48228
rect 10888 46676 10936 47438
rect 11320 46676 11368 47438
rect 10888 45886 10936 46648
rect 11320 45886 11368 46648
rect 10888 45096 10936 45858
rect 11320 45096 11368 45858
rect 10888 44306 10936 45068
rect 11320 44306 11368 45068
rect 10888 43516 10936 44278
rect 11320 43516 11368 44278
rect 10888 42726 10936 43488
rect 11320 42726 11368 43488
rect 10888 41936 10936 42698
rect 11320 41936 11368 42698
rect 10888 41146 10936 41908
rect 11320 41146 11368 41908
rect 10888 40356 10936 41118
rect 11320 40356 11368 41118
rect 10888 39566 10936 40328
rect 11320 39566 11368 40328
rect 10888 38776 10936 39538
rect 11320 38776 11368 39538
rect 10888 37986 10936 38748
rect 11320 37986 11368 38748
rect 10888 37196 10936 37958
rect 11320 37196 11368 37958
rect 10888 36406 10936 37168
rect 11320 36406 11368 37168
rect 10888 35616 10936 36378
rect 11320 35616 11368 36378
rect 10888 34826 10936 35588
rect 11320 34826 11368 35588
rect 10888 34036 10936 34798
rect 11320 34036 11368 34798
rect 10888 33246 10936 34008
rect 11320 33246 11368 34008
rect 10888 32456 10936 33218
rect 11320 32456 11368 33218
rect 10888 31666 10936 32428
rect 11320 31666 11368 32428
rect 10888 30876 10936 31638
rect 11320 30876 11368 31638
rect 10888 30086 10936 30848
rect 11320 30086 11368 30848
rect 10888 29296 10936 30058
rect 11320 29296 11368 30058
rect 11712 29282 11740 79842
rect 11984 29282 12012 79842
rect 12420 29223 12468 79843
rect 12844 29221 12894 79845
rect 13898 29253 13926 79813
rect 15422 29253 15450 79813
rect 17084 79775 17270 79851
rect 17084 79617 17141 79775
rect 17177 79650 17270 79716
tri 17177 79634 17193 79650 ne
rect 17193 79634 17270 79650
rect 17084 79535 17158 79617
rect 17084 79301 17141 79535
tri 17177 79502 17193 79518 se
rect 17193 79502 17270 79518
rect 17177 79436 17270 79502
rect 17177 79334 17270 79400
tri 17177 79318 17193 79334 ne
rect 17193 79318 17270 79334
rect 17084 79219 17158 79301
rect 17084 79061 17141 79219
tri 17177 79186 17193 79202 se
rect 17193 79186 17270 79202
rect 17177 79120 17270 79186
rect 17084 78985 17270 79061
rect 17084 78827 17141 78985
rect 17177 78860 17270 78926
tri 17177 78844 17193 78860 ne
rect 17193 78844 17270 78860
rect 17084 78745 17158 78827
rect 17084 78511 17141 78745
tri 17177 78712 17193 78728 se
rect 17193 78712 17270 78728
rect 17177 78646 17270 78712
rect 17177 78544 17270 78610
tri 17177 78528 17193 78544 ne
rect 17193 78528 17270 78544
rect 17084 78429 17158 78511
rect 17084 78271 17141 78429
tri 17177 78396 17193 78412 se
rect 17193 78396 17270 78412
rect 17177 78330 17270 78396
rect 17084 78195 17270 78271
rect 17084 78037 17141 78195
rect 17177 78070 17270 78136
tri 17177 78054 17193 78070 ne
rect 17193 78054 17270 78070
rect 17084 77955 17158 78037
rect 17084 77721 17141 77955
tri 17177 77922 17193 77938 se
rect 17193 77922 17270 77938
rect 17177 77856 17270 77922
rect 17177 77754 17270 77820
tri 17177 77738 17193 77754 ne
rect 17193 77738 17270 77754
rect 17084 77639 17158 77721
rect 17084 77481 17141 77639
tri 17177 77606 17193 77622 se
rect 17193 77606 17270 77622
rect 17177 77540 17270 77606
rect 17084 77405 17270 77481
rect 17084 77247 17141 77405
rect 17177 77280 17270 77346
tri 17177 77264 17193 77280 ne
rect 17193 77264 17270 77280
rect 17084 77165 17158 77247
rect 17084 76931 17141 77165
tri 17177 77132 17193 77148 se
rect 17193 77132 17270 77148
rect 17177 77066 17270 77132
rect 17177 76964 17270 77030
tri 17177 76948 17193 76964 ne
rect 17193 76948 17270 76964
rect 17084 76849 17158 76931
rect 17084 76691 17141 76849
tri 17177 76816 17193 76832 se
rect 17193 76816 17270 76832
rect 17177 76750 17270 76816
rect 17084 76615 17270 76691
rect 17084 76457 17141 76615
rect 17177 76490 17270 76556
tri 17177 76474 17193 76490 ne
rect 17193 76474 17270 76490
rect 17084 76375 17158 76457
rect 17084 76141 17141 76375
tri 17177 76342 17193 76358 se
rect 17193 76342 17270 76358
rect 17177 76276 17270 76342
rect 17177 76174 17270 76240
tri 17177 76158 17193 76174 ne
rect 17193 76158 17270 76174
rect 17084 76059 17158 76141
rect 17084 75901 17141 76059
tri 17177 76026 17193 76042 se
rect 17193 76026 17270 76042
rect 17177 75960 17270 76026
rect 17084 75825 17270 75901
rect 17084 75667 17141 75825
rect 17177 75700 17270 75766
tri 17177 75684 17193 75700 ne
rect 17193 75684 17270 75700
rect 17084 75585 17158 75667
rect 17084 75351 17141 75585
tri 17177 75552 17193 75568 se
rect 17193 75552 17270 75568
rect 17177 75486 17270 75552
rect 17177 75384 17270 75450
tri 17177 75368 17193 75384 ne
rect 17193 75368 17270 75384
rect 17084 75269 17158 75351
rect 17084 75111 17141 75269
tri 17177 75236 17193 75252 se
rect 17193 75236 17270 75252
rect 17177 75170 17270 75236
rect 17084 75035 17270 75111
rect 17084 74877 17141 75035
rect 17177 74910 17270 74976
tri 17177 74894 17193 74910 ne
rect 17193 74894 17270 74910
rect 17084 74795 17158 74877
rect 17084 74561 17141 74795
tri 17177 74762 17193 74778 se
rect 17193 74762 17270 74778
rect 17177 74696 17270 74762
rect 17177 74594 17270 74660
tri 17177 74578 17193 74594 ne
rect 17193 74578 17270 74594
rect 17084 74479 17158 74561
rect 17084 74321 17141 74479
tri 17177 74446 17193 74462 se
rect 17193 74446 17270 74462
rect 17177 74380 17270 74446
rect 17084 74245 17270 74321
rect 17084 74087 17141 74245
rect 17177 74120 17270 74186
tri 17177 74104 17193 74120 ne
rect 17193 74104 17270 74120
rect 17084 74005 17158 74087
rect 17084 73771 17141 74005
tri 17177 73972 17193 73988 se
rect 17193 73972 17270 73988
rect 17177 73906 17270 73972
rect 17177 73804 17270 73870
tri 17177 73788 17193 73804 ne
rect 17193 73788 17270 73804
rect 17084 73689 17158 73771
rect 17084 73531 17141 73689
tri 17177 73656 17193 73672 se
rect 17193 73656 17270 73672
rect 17177 73590 17270 73656
rect 17084 73455 17270 73531
rect 17084 73297 17141 73455
rect 17177 73330 17270 73396
tri 17177 73314 17193 73330 ne
rect 17193 73314 17270 73330
rect 17084 73215 17158 73297
rect 17084 72981 17141 73215
tri 17177 73182 17193 73198 se
rect 17193 73182 17270 73198
rect 17177 73116 17270 73182
rect 17177 73014 17270 73080
tri 17177 72998 17193 73014 ne
rect 17193 72998 17270 73014
rect 17084 72899 17158 72981
rect 17084 72741 17141 72899
tri 17177 72866 17193 72882 se
rect 17193 72866 17270 72882
rect 17177 72800 17270 72866
rect 17084 72665 17270 72741
rect 17084 72507 17141 72665
rect 17177 72540 17270 72606
tri 17177 72524 17193 72540 ne
rect 17193 72524 17270 72540
rect 17084 72425 17158 72507
rect 17084 72191 17141 72425
tri 17177 72392 17193 72408 se
rect 17193 72392 17270 72408
rect 17177 72326 17270 72392
rect 17177 72224 17270 72290
tri 17177 72208 17193 72224 ne
rect 17193 72208 17270 72224
rect 17084 72109 17158 72191
rect 17084 71951 17141 72109
tri 17177 72076 17193 72092 se
rect 17193 72076 17270 72092
rect 17177 72010 17270 72076
rect 17084 71875 17270 71951
rect 17084 71717 17141 71875
rect 17177 71750 17270 71816
tri 17177 71734 17193 71750 ne
rect 17193 71734 17270 71750
rect 17084 71635 17158 71717
rect 17084 71401 17141 71635
tri 17177 71602 17193 71618 se
rect 17193 71602 17270 71618
rect 17177 71536 17270 71602
rect 17177 71434 17270 71500
tri 17177 71418 17193 71434 ne
rect 17193 71418 17270 71434
rect 17084 71319 17158 71401
rect 17084 71161 17141 71319
tri 17177 71286 17193 71302 se
rect 17193 71286 17270 71302
rect 17177 71220 17270 71286
rect 17084 71085 17270 71161
rect 17084 70927 17141 71085
rect 17177 70960 17270 71026
tri 17177 70944 17193 70960 ne
rect 17193 70944 17270 70960
rect 17084 70845 17158 70927
rect 17084 70611 17141 70845
tri 17177 70812 17193 70828 se
rect 17193 70812 17270 70828
rect 17177 70746 17270 70812
rect 17177 70644 17270 70710
tri 17177 70628 17193 70644 ne
rect 17193 70628 17270 70644
rect 17084 70529 17158 70611
rect 17084 70371 17141 70529
tri 17177 70496 17193 70512 se
rect 17193 70496 17270 70512
rect 17177 70430 17270 70496
rect 17084 70295 17270 70371
rect 17084 70137 17141 70295
rect 17177 70170 17270 70236
tri 17177 70154 17193 70170 ne
rect 17193 70154 17270 70170
rect 17084 70055 17158 70137
rect 17084 69821 17141 70055
tri 17177 70022 17193 70038 se
rect 17193 70022 17270 70038
rect 17177 69956 17270 70022
rect 17177 69854 17270 69920
tri 17177 69838 17193 69854 ne
rect 17193 69838 17270 69854
rect 17084 69739 17158 69821
rect 17084 69581 17141 69739
tri 17177 69706 17193 69722 se
rect 17193 69706 17270 69722
rect 17177 69640 17270 69706
rect 17084 69505 17270 69581
rect 17084 69347 17141 69505
rect 17177 69380 17270 69446
tri 17177 69364 17193 69380 ne
rect 17193 69364 17270 69380
rect 17084 69265 17158 69347
rect 17084 69031 17141 69265
tri 17177 69232 17193 69248 se
rect 17193 69232 17270 69248
rect 17177 69166 17270 69232
rect 17177 69064 17270 69130
tri 17177 69048 17193 69064 ne
rect 17193 69048 17270 69064
rect 17084 68949 17158 69031
rect 17084 68791 17141 68949
tri 17177 68916 17193 68932 se
rect 17193 68916 17270 68932
rect 17177 68850 17270 68916
rect 17084 68715 17270 68791
rect 17084 68557 17141 68715
rect 17177 68590 17270 68656
tri 17177 68574 17193 68590 ne
rect 17193 68574 17270 68590
rect 17084 68475 17158 68557
rect 17084 68241 17141 68475
tri 17177 68442 17193 68458 se
rect 17193 68442 17270 68458
rect 17177 68376 17270 68442
rect 17177 68274 17270 68340
tri 17177 68258 17193 68274 ne
rect 17193 68258 17270 68274
rect 17084 68159 17158 68241
rect 17084 68001 17141 68159
tri 17177 68126 17193 68142 se
rect 17193 68126 17270 68142
rect 17177 68060 17270 68126
rect 17084 67925 17270 68001
rect 17084 67767 17141 67925
rect 17177 67800 17270 67866
tri 17177 67784 17193 67800 ne
rect 17193 67784 17270 67800
rect 17084 67685 17158 67767
rect 17084 67451 17141 67685
tri 17177 67652 17193 67668 se
rect 17193 67652 17270 67668
rect 17177 67586 17270 67652
rect 17177 67484 17270 67550
tri 17177 67468 17193 67484 ne
rect 17193 67468 17270 67484
rect 17084 67369 17158 67451
rect 17084 67211 17141 67369
tri 17177 67336 17193 67352 se
rect 17193 67336 17270 67352
rect 17177 67270 17270 67336
rect 17084 67135 17270 67211
rect 17084 66977 17141 67135
rect 17177 67010 17270 67076
tri 17177 66994 17193 67010 ne
rect 17193 66994 17270 67010
rect 17084 66895 17158 66977
rect 17084 66661 17141 66895
tri 17177 66862 17193 66878 se
rect 17193 66862 17270 66878
rect 17177 66796 17270 66862
rect 17177 66694 17270 66760
tri 17177 66678 17193 66694 ne
rect 17193 66678 17270 66694
rect 17084 66579 17158 66661
rect 17084 66421 17141 66579
tri 17177 66546 17193 66562 se
rect 17193 66546 17270 66562
rect 17177 66480 17270 66546
rect 17084 66345 17270 66421
rect 17084 66187 17141 66345
rect 17177 66220 17270 66286
tri 17177 66204 17193 66220 ne
rect 17193 66204 17270 66220
rect 17084 66105 17158 66187
rect 17084 65871 17141 66105
tri 17177 66072 17193 66088 se
rect 17193 66072 17270 66088
rect 17177 66006 17270 66072
rect 17177 65904 17270 65970
tri 17177 65888 17193 65904 ne
rect 17193 65888 17270 65904
rect 17084 65789 17158 65871
rect 17084 65631 17141 65789
tri 17177 65756 17193 65772 se
rect 17193 65756 17270 65772
rect 17177 65690 17270 65756
rect 17084 65555 17270 65631
rect 17084 65397 17141 65555
rect 17177 65430 17270 65496
tri 17177 65414 17193 65430 ne
rect 17193 65414 17270 65430
rect 17084 65315 17158 65397
rect 17084 65081 17141 65315
tri 17177 65282 17193 65298 se
rect 17193 65282 17270 65298
rect 17177 65216 17270 65282
rect 17177 65114 17270 65180
tri 17177 65098 17193 65114 ne
rect 17193 65098 17270 65114
rect 17084 64999 17158 65081
rect 17084 64841 17141 64999
tri 17177 64966 17193 64982 se
rect 17193 64966 17270 64982
rect 17177 64900 17270 64966
rect 17084 64765 17270 64841
rect 17084 64607 17141 64765
rect 17177 64640 17270 64706
tri 17177 64624 17193 64640 ne
rect 17193 64624 17270 64640
rect 17084 64525 17158 64607
rect 17084 64291 17141 64525
tri 17177 64492 17193 64508 se
rect 17193 64492 17270 64508
rect 17177 64426 17270 64492
rect 17177 64324 17270 64390
tri 17177 64308 17193 64324 ne
rect 17193 64308 17270 64324
rect 17084 64209 17158 64291
rect 17084 64051 17141 64209
tri 17177 64176 17193 64192 se
rect 17193 64176 17270 64192
rect 17177 64110 17270 64176
rect 17084 63975 17270 64051
rect 17084 63817 17141 63975
rect 17177 63850 17270 63916
tri 17177 63834 17193 63850 ne
rect 17193 63834 17270 63850
rect 17084 63735 17158 63817
rect 17084 63501 17141 63735
tri 17177 63702 17193 63718 se
rect 17193 63702 17270 63718
rect 17177 63636 17270 63702
rect 17177 63534 17270 63600
tri 17177 63518 17193 63534 ne
rect 17193 63518 17270 63534
rect 17084 63419 17158 63501
rect 17084 63261 17141 63419
tri 17177 63386 17193 63402 se
rect 17193 63386 17270 63402
rect 17177 63320 17270 63386
rect 17084 63185 17270 63261
rect 17084 63027 17141 63185
rect 17177 63060 17270 63126
tri 17177 63044 17193 63060 ne
rect 17193 63044 17270 63060
rect 17084 62945 17158 63027
rect 17084 62711 17141 62945
tri 17177 62912 17193 62928 se
rect 17193 62912 17270 62928
rect 17177 62846 17270 62912
rect 17177 62744 17270 62810
tri 17177 62728 17193 62744 ne
rect 17193 62728 17270 62744
rect 17084 62629 17158 62711
rect 17084 62471 17141 62629
tri 17177 62596 17193 62612 se
rect 17193 62596 17270 62612
rect 17177 62530 17270 62596
rect 17084 62395 17270 62471
rect 17084 62237 17141 62395
rect 17177 62270 17270 62336
tri 17177 62254 17193 62270 ne
rect 17193 62254 17270 62270
rect 17084 62155 17158 62237
rect 17084 61921 17141 62155
tri 17177 62122 17193 62138 se
rect 17193 62122 17270 62138
rect 17177 62056 17270 62122
rect 17177 61954 17270 62020
tri 17177 61938 17193 61954 ne
rect 17193 61938 17270 61954
rect 17084 61839 17158 61921
rect 17084 61681 17141 61839
tri 17177 61806 17193 61822 se
rect 17193 61806 17270 61822
rect 17177 61740 17270 61806
rect 17084 61605 17270 61681
rect 17084 61447 17141 61605
rect 17177 61480 17270 61546
tri 17177 61464 17193 61480 ne
rect 17193 61464 17270 61480
rect 17084 61365 17158 61447
rect 17084 61131 17141 61365
tri 17177 61332 17193 61348 se
rect 17193 61332 17270 61348
rect 17177 61266 17270 61332
rect 17177 61164 17270 61230
tri 17177 61148 17193 61164 ne
rect 17193 61148 17270 61164
rect 17084 61049 17158 61131
rect 17084 60891 17141 61049
tri 17177 61016 17193 61032 se
rect 17193 61016 17270 61032
rect 17177 60950 17270 61016
rect 17084 60815 17270 60891
rect 17084 60657 17141 60815
rect 17177 60690 17270 60756
tri 17177 60674 17193 60690 ne
rect 17193 60674 17270 60690
rect 17084 60575 17158 60657
rect 17084 60341 17141 60575
tri 17177 60542 17193 60558 se
rect 17193 60542 17270 60558
rect 17177 60476 17270 60542
rect 17177 60374 17270 60440
tri 17177 60358 17193 60374 ne
rect 17193 60358 17270 60374
rect 17084 60259 17158 60341
rect 17084 60101 17141 60259
tri 17177 60226 17193 60242 se
rect 17193 60226 17270 60242
rect 17177 60160 17270 60226
rect 17084 60025 17270 60101
rect 17084 59867 17141 60025
rect 17177 59900 17270 59966
tri 17177 59884 17193 59900 ne
rect 17193 59884 17270 59900
rect 17084 59785 17158 59867
rect 17084 59551 17141 59785
tri 17177 59752 17193 59768 se
rect 17193 59752 17270 59768
rect 17177 59686 17270 59752
rect 17177 59584 17270 59650
tri 17177 59568 17193 59584 ne
rect 17193 59568 17270 59584
rect 17084 59469 17158 59551
rect 17084 59311 17141 59469
tri 17177 59436 17193 59452 se
rect 17193 59436 17270 59452
rect 17177 59370 17270 59436
rect 17084 59235 17270 59311
rect 17084 59077 17141 59235
rect 17177 59110 17270 59176
tri 17177 59094 17193 59110 ne
rect 17193 59094 17270 59110
rect 17084 58995 17158 59077
rect 17084 58761 17141 58995
tri 17177 58962 17193 58978 se
rect 17193 58962 17270 58978
rect 17177 58896 17270 58962
rect 17177 58794 17270 58860
tri 17177 58778 17193 58794 ne
rect 17193 58778 17270 58794
rect 17084 58679 17158 58761
rect 17084 58521 17141 58679
tri 17177 58646 17193 58662 se
rect 17193 58646 17270 58662
rect 17177 58580 17270 58646
rect 17084 58445 17270 58521
rect 17084 58287 17141 58445
rect 17177 58320 17270 58386
tri 17177 58304 17193 58320 ne
rect 17193 58304 17270 58320
rect 17084 58205 17158 58287
rect 17084 57971 17141 58205
tri 17177 58172 17193 58188 se
rect 17193 58172 17270 58188
rect 17177 58106 17270 58172
rect 17177 58004 17270 58070
tri 17177 57988 17193 58004 ne
rect 17193 57988 17270 58004
rect 17084 57889 17158 57971
rect 17084 57731 17141 57889
tri 17177 57856 17193 57872 se
rect 17193 57856 17270 57872
rect 17177 57790 17270 57856
rect 17084 57655 17270 57731
rect 17084 57497 17141 57655
rect 17177 57530 17270 57596
tri 17177 57514 17193 57530 ne
rect 17193 57514 17270 57530
rect 17084 57415 17158 57497
rect 17084 57181 17141 57415
tri 17177 57382 17193 57398 se
rect 17193 57382 17270 57398
rect 17177 57316 17270 57382
rect 17177 57214 17270 57280
tri 17177 57198 17193 57214 ne
rect 17193 57198 17270 57214
rect 17084 57099 17158 57181
rect 17084 56941 17141 57099
tri 17177 57066 17193 57082 se
rect 17193 57066 17270 57082
rect 17177 57000 17270 57066
rect 17084 56865 17270 56941
rect 17084 56707 17141 56865
rect 17177 56740 17270 56806
tri 17177 56724 17193 56740 ne
rect 17193 56724 17270 56740
rect 17084 56625 17158 56707
rect 17084 56391 17141 56625
tri 17177 56592 17193 56608 se
rect 17193 56592 17270 56608
rect 17177 56526 17270 56592
rect 17177 56424 17270 56490
tri 17177 56408 17193 56424 ne
rect 17193 56408 17270 56424
rect 17084 56309 17158 56391
rect 17084 56151 17141 56309
tri 17177 56276 17193 56292 se
rect 17193 56276 17270 56292
rect 17177 56210 17270 56276
rect 17084 56075 17270 56151
rect 17084 55917 17141 56075
rect 17177 55950 17270 56016
tri 17177 55934 17193 55950 ne
rect 17193 55934 17270 55950
rect 17084 55835 17158 55917
rect 17084 55601 17141 55835
tri 17177 55802 17193 55818 se
rect 17193 55802 17270 55818
rect 17177 55736 17270 55802
rect 17177 55634 17270 55700
tri 17177 55618 17193 55634 ne
rect 17193 55618 17270 55634
rect 17084 55519 17158 55601
rect 17084 55361 17141 55519
tri 17177 55486 17193 55502 se
rect 17193 55486 17270 55502
rect 17177 55420 17270 55486
rect 17084 55285 17270 55361
rect 17084 55127 17141 55285
rect 17177 55160 17270 55226
tri 17177 55144 17193 55160 ne
rect 17193 55144 17270 55160
rect 17084 55045 17158 55127
rect 17084 54811 17141 55045
tri 17177 55012 17193 55028 se
rect 17193 55012 17270 55028
rect 17177 54946 17270 55012
rect 17177 54844 17270 54910
tri 17177 54828 17193 54844 ne
rect 17193 54828 17270 54844
rect 17084 54729 17158 54811
rect 17084 54571 17141 54729
tri 17177 54696 17193 54712 se
rect 17193 54696 17270 54712
rect 17177 54630 17270 54696
rect 17084 54495 17270 54571
rect 17084 54337 17141 54495
rect 17177 54370 17270 54436
tri 17177 54354 17193 54370 ne
rect 17193 54354 17270 54370
rect 17084 54255 17158 54337
rect 17084 54021 17141 54255
tri 17177 54222 17193 54238 se
rect 17193 54222 17270 54238
rect 17177 54156 17270 54222
rect 17177 54054 17270 54120
tri 17177 54038 17193 54054 ne
rect 17193 54038 17270 54054
rect 17084 53939 17158 54021
rect 17084 53781 17141 53939
tri 17177 53906 17193 53922 se
rect 17193 53906 17270 53922
rect 17177 53840 17270 53906
rect 17084 53705 17270 53781
rect 17084 53547 17141 53705
rect 17177 53580 17270 53646
tri 17177 53564 17193 53580 ne
rect 17193 53564 17270 53580
rect 17084 53465 17158 53547
rect 17084 53231 17141 53465
tri 17177 53432 17193 53448 se
rect 17193 53432 17270 53448
rect 17177 53366 17270 53432
rect 17177 53264 17270 53330
tri 17177 53248 17193 53264 ne
rect 17193 53248 17270 53264
rect 17084 53149 17158 53231
rect 17084 52991 17141 53149
tri 17177 53116 17193 53132 se
rect 17193 53116 17270 53132
rect 17177 53050 17270 53116
rect 17084 52915 17270 52991
rect 17084 52757 17141 52915
rect 17177 52790 17270 52856
tri 17177 52774 17193 52790 ne
rect 17193 52774 17270 52790
rect 17084 52675 17158 52757
rect 17084 52441 17141 52675
tri 17177 52642 17193 52658 se
rect 17193 52642 17270 52658
rect 17177 52576 17270 52642
rect 17177 52474 17270 52540
tri 17177 52458 17193 52474 ne
rect 17193 52458 17270 52474
rect 17084 52359 17158 52441
rect 17084 52201 17141 52359
tri 17177 52326 17193 52342 se
rect 17193 52326 17270 52342
rect 17177 52260 17270 52326
rect 17084 52125 17270 52201
rect 17084 51967 17141 52125
rect 17177 52000 17270 52066
tri 17177 51984 17193 52000 ne
rect 17193 51984 17270 52000
rect 17084 51885 17158 51967
rect 17084 51651 17141 51885
tri 17177 51852 17193 51868 se
rect 17193 51852 17270 51868
rect 17177 51786 17270 51852
rect 17177 51684 17270 51750
tri 17177 51668 17193 51684 ne
rect 17193 51668 17270 51684
rect 17084 51569 17158 51651
rect 17084 51411 17141 51569
tri 17177 51536 17193 51552 se
rect 17193 51536 17270 51552
rect 17177 51470 17270 51536
rect 17084 51335 17270 51411
rect 17084 51177 17141 51335
rect 17177 51210 17270 51276
tri 17177 51194 17193 51210 ne
rect 17193 51194 17270 51210
rect 17084 51095 17158 51177
rect 17084 50861 17141 51095
tri 17177 51062 17193 51078 se
rect 17193 51062 17270 51078
rect 17177 50996 17270 51062
rect 17177 50894 17270 50960
tri 17177 50878 17193 50894 ne
rect 17193 50878 17270 50894
rect 17084 50779 17158 50861
rect 17084 50621 17141 50779
tri 17177 50746 17193 50762 se
rect 17193 50746 17270 50762
rect 17177 50680 17270 50746
rect 17084 50545 17270 50621
rect 17084 50387 17141 50545
rect 17177 50420 17270 50486
tri 17177 50404 17193 50420 ne
rect 17193 50404 17270 50420
rect 17084 50305 17158 50387
rect 17084 50071 17141 50305
tri 17177 50272 17193 50288 se
rect 17193 50272 17270 50288
rect 17177 50206 17270 50272
rect 17177 50104 17270 50170
tri 17177 50088 17193 50104 ne
rect 17193 50088 17270 50104
rect 17084 49989 17158 50071
rect 17084 49831 17141 49989
tri 17177 49956 17193 49972 se
rect 17193 49956 17270 49972
rect 17177 49890 17270 49956
rect 17084 49755 17270 49831
rect 17084 49597 17141 49755
rect 17177 49630 17270 49696
tri 17177 49614 17193 49630 ne
rect 17193 49614 17270 49630
rect 17084 49515 17158 49597
rect 17084 49281 17141 49515
tri 17177 49482 17193 49498 se
rect 17193 49482 17270 49498
rect 17177 49416 17270 49482
rect 17177 49314 17270 49380
tri 17177 49298 17193 49314 ne
rect 17193 49298 17270 49314
rect 17084 49199 17158 49281
rect 17084 49041 17141 49199
tri 17177 49166 17193 49182 se
rect 17193 49166 17270 49182
rect 17177 49100 17270 49166
rect 17084 48965 17270 49041
rect 17084 48807 17141 48965
rect 17177 48840 17270 48906
tri 17177 48824 17193 48840 ne
rect 17193 48824 17270 48840
rect 17084 48725 17158 48807
rect 17084 48491 17141 48725
tri 17177 48692 17193 48708 se
rect 17193 48692 17270 48708
rect 17177 48626 17270 48692
rect 17177 48524 17270 48590
tri 17177 48508 17193 48524 ne
rect 17193 48508 17270 48524
rect 17084 48409 17158 48491
rect 17084 48251 17141 48409
tri 17177 48376 17193 48392 se
rect 17193 48376 17270 48392
rect 17177 48310 17270 48376
rect 17084 48175 17270 48251
rect 17084 48017 17141 48175
rect 17177 48050 17270 48116
tri 17177 48034 17193 48050 ne
rect 17193 48034 17270 48050
rect 17084 47935 17158 48017
rect 17084 47701 17141 47935
tri 17177 47902 17193 47918 se
rect 17193 47902 17270 47918
rect 17177 47836 17270 47902
rect 17177 47734 17270 47800
tri 17177 47718 17193 47734 ne
rect 17193 47718 17270 47734
rect 17084 47619 17158 47701
rect 17084 47461 17141 47619
tri 17177 47586 17193 47602 se
rect 17193 47586 17270 47602
rect 17177 47520 17270 47586
rect 17084 47385 17270 47461
rect 17084 47227 17141 47385
rect 17177 47260 17270 47326
tri 17177 47244 17193 47260 ne
rect 17193 47244 17270 47260
rect 17084 47145 17158 47227
rect 17084 46911 17141 47145
tri 17177 47112 17193 47128 se
rect 17193 47112 17270 47128
rect 17177 47046 17270 47112
rect 17177 46944 17270 47010
tri 17177 46928 17193 46944 ne
rect 17193 46928 17270 46944
rect 17084 46829 17158 46911
rect 17084 46671 17141 46829
tri 17177 46796 17193 46812 se
rect 17193 46796 17270 46812
rect 17177 46730 17270 46796
rect 17084 46595 17270 46671
rect 17084 46437 17141 46595
rect 17177 46470 17270 46536
tri 17177 46454 17193 46470 ne
rect 17193 46454 17270 46470
rect 17084 46355 17158 46437
rect 17084 46121 17141 46355
tri 17177 46322 17193 46338 se
rect 17193 46322 17270 46338
rect 17177 46256 17270 46322
rect 17177 46154 17270 46220
tri 17177 46138 17193 46154 ne
rect 17193 46138 17270 46154
rect 17084 46039 17158 46121
rect 17084 45881 17141 46039
tri 17177 46006 17193 46022 se
rect 17193 46006 17270 46022
rect 17177 45940 17270 46006
rect 17084 45805 17270 45881
rect 17084 45647 17141 45805
rect 17177 45680 17270 45746
tri 17177 45664 17193 45680 ne
rect 17193 45664 17270 45680
rect 17084 45565 17158 45647
rect 17084 45331 17141 45565
tri 17177 45532 17193 45548 se
rect 17193 45532 17270 45548
rect 17177 45466 17270 45532
rect 17177 45364 17270 45430
tri 17177 45348 17193 45364 ne
rect 17193 45348 17270 45364
rect 17084 45249 17158 45331
rect 17084 45091 17141 45249
tri 17177 45216 17193 45232 se
rect 17193 45216 17270 45232
rect 17177 45150 17270 45216
rect 17084 45015 17270 45091
rect 17084 44857 17141 45015
rect 17177 44890 17270 44956
tri 17177 44874 17193 44890 ne
rect 17193 44874 17270 44890
rect 17084 44775 17158 44857
rect 17084 44541 17141 44775
tri 17177 44742 17193 44758 se
rect 17193 44742 17270 44758
rect 17177 44676 17270 44742
rect 17177 44574 17270 44640
tri 17177 44558 17193 44574 ne
rect 17193 44558 17270 44574
rect 17084 44459 17158 44541
rect 17084 44301 17141 44459
tri 17177 44426 17193 44442 se
rect 17193 44426 17270 44442
rect 17177 44360 17270 44426
rect 17084 44225 17270 44301
rect 17084 44067 17141 44225
rect 17177 44100 17270 44166
tri 17177 44084 17193 44100 ne
rect 17193 44084 17270 44100
rect 17084 43985 17158 44067
rect 17084 43751 17141 43985
tri 17177 43952 17193 43968 se
rect 17193 43952 17270 43968
rect 17177 43886 17270 43952
rect 17177 43784 17270 43850
tri 17177 43768 17193 43784 ne
rect 17193 43768 17270 43784
rect 17084 43669 17158 43751
rect 17084 43511 17141 43669
tri 17177 43636 17193 43652 se
rect 17193 43636 17270 43652
rect 17177 43570 17270 43636
rect 17084 43435 17270 43511
rect 17084 43277 17141 43435
rect 17177 43310 17270 43376
tri 17177 43294 17193 43310 ne
rect 17193 43294 17270 43310
rect 17084 43195 17158 43277
rect 17084 42961 17141 43195
tri 17177 43162 17193 43178 se
rect 17193 43162 17270 43178
rect 17177 43096 17270 43162
rect 17177 42994 17270 43060
tri 17177 42978 17193 42994 ne
rect 17193 42978 17270 42994
rect 17084 42879 17158 42961
rect 17084 42721 17141 42879
tri 17177 42846 17193 42862 se
rect 17193 42846 17270 42862
rect 17177 42780 17270 42846
rect 17084 42645 17270 42721
rect 17084 42487 17141 42645
rect 17177 42520 17270 42586
tri 17177 42504 17193 42520 ne
rect 17193 42504 17270 42520
rect 17084 42405 17158 42487
rect 17084 42171 17141 42405
tri 17177 42372 17193 42388 se
rect 17193 42372 17270 42388
rect 17177 42306 17270 42372
rect 17177 42204 17270 42270
tri 17177 42188 17193 42204 ne
rect 17193 42188 17270 42204
rect 17084 42089 17158 42171
rect 17084 41931 17141 42089
tri 17177 42056 17193 42072 se
rect 17193 42056 17270 42072
rect 17177 41990 17270 42056
rect 17084 41855 17270 41931
rect 17084 41697 17141 41855
rect 17177 41730 17270 41796
tri 17177 41714 17193 41730 ne
rect 17193 41714 17270 41730
rect 17084 41615 17158 41697
rect 17084 41381 17141 41615
tri 17177 41582 17193 41598 se
rect 17193 41582 17270 41598
rect 17177 41516 17270 41582
rect 17177 41414 17270 41480
tri 17177 41398 17193 41414 ne
rect 17193 41398 17270 41414
rect 17084 41299 17158 41381
rect 17084 41141 17141 41299
tri 17177 41266 17193 41282 se
rect 17193 41266 17270 41282
rect 17177 41200 17270 41266
rect 17084 41065 17270 41141
rect 17084 40907 17141 41065
rect 17177 40940 17270 41006
tri 17177 40924 17193 40940 ne
rect 17193 40924 17270 40940
rect 17084 40825 17158 40907
rect 17084 40591 17141 40825
tri 17177 40792 17193 40808 se
rect 17193 40792 17270 40808
rect 17177 40726 17270 40792
rect 17177 40624 17270 40690
tri 17177 40608 17193 40624 ne
rect 17193 40608 17270 40624
rect 17084 40509 17158 40591
rect 17084 40351 17141 40509
tri 17177 40476 17193 40492 se
rect 17193 40476 17270 40492
rect 17177 40410 17270 40476
rect 17084 40275 17270 40351
rect 17084 40117 17141 40275
rect 17177 40150 17270 40216
tri 17177 40134 17193 40150 ne
rect 17193 40134 17270 40150
rect 17084 40035 17158 40117
rect 17084 39801 17141 40035
tri 17177 40002 17193 40018 se
rect 17193 40002 17270 40018
rect 17177 39936 17270 40002
rect 17177 39834 17270 39900
tri 17177 39818 17193 39834 ne
rect 17193 39818 17270 39834
rect 17084 39719 17158 39801
rect 17084 39561 17141 39719
tri 17177 39686 17193 39702 se
rect 17193 39686 17270 39702
rect 17177 39620 17270 39686
rect 17084 39485 17270 39561
rect 17084 39327 17141 39485
rect 17177 39360 17270 39426
tri 17177 39344 17193 39360 ne
rect 17193 39344 17270 39360
rect 17084 39245 17158 39327
rect 17084 39011 17141 39245
tri 17177 39212 17193 39228 se
rect 17193 39212 17270 39228
rect 17177 39146 17270 39212
rect 17177 39044 17270 39110
tri 17177 39028 17193 39044 ne
rect 17193 39028 17270 39044
rect 17084 38929 17158 39011
rect 17084 38771 17141 38929
tri 17177 38896 17193 38912 se
rect 17193 38896 17270 38912
rect 17177 38830 17270 38896
rect 17084 38695 17270 38771
rect 17084 38537 17141 38695
rect 17177 38570 17270 38636
tri 17177 38554 17193 38570 ne
rect 17193 38554 17270 38570
rect 17084 38455 17158 38537
rect 17084 38221 17141 38455
tri 17177 38422 17193 38438 se
rect 17193 38422 17270 38438
rect 17177 38356 17270 38422
rect 17177 38254 17270 38320
tri 17177 38238 17193 38254 ne
rect 17193 38238 17270 38254
rect 17084 38139 17158 38221
rect 17084 37981 17141 38139
tri 17177 38106 17193 38122 se
rect 17193 38106 17270 38122
rect 17177 38040 17270 38106
rect 17084 37905 17270 37981
rect 17084 37747 17141 37905
rect 17177 37780 17270 37846
tri 17177 37764 17193 37780 ne
rect 17193 37764 17270 37780
rect 17084 37665 17158 37747
rect 17084 37431 17141 37665
tri 17177 37632 17193 37648 se
rect 17193 37632 17270 37648
rect 17177 37566 17270 37632
rect 17177 37464 17270 37530
tri 17177 37448 17193 37464 ne
rect 17193 37448 17270 37464
rect 17084 37349 17158 37431
rect 17084 37191 17141 37349
tri 17177 37316 17193 37332 se
rect 17193 37316 17270 37332
rect 17177 37250 17270 37316
rect 17084 37115 17270 37191
rect 17084 36957 17141 37115
rect 17177 36990 17270 37056
tri 17177 36974 17193 36990 ne
rect 17193 36974 17270 36990
rect 17084 36875 17158 36957
rect 17084 36641 17141 36875
tri 17177 36842 17193 36858 se
rect 17193 36842 17270 36858
rect 17177 36776 17270 36842
rect 17177 36674 17270 36740
tri 17177 36658 17193 36674 ne
rect 17193 36658 17270 36674
rect 17084 36559 17158 36641
rect 17084 36401 17141 36559
tri 17177 36526 17193 36542 se
rect 17193 36526 17270 36542
rect 17177 36460 17270 36526
rect 17084 36325 17270 36401
rect 17084 36167 17141 36325
rect 17177 36200 17270 36266
tri 17177 36184 17193 36200 ne
rect 17193 36184 17270 36200
rect 17084 36085 17158 36167
rect 17084 35851 17141 36085
tri 17177 36052 17193 36068 se
rect 17193 36052 17270 36068
rect 17177 35986 17270 36052
rect 17177 35884 17270 35950
tri 17177 35868 17193 35884 ne
rect 17193 35868 17270 35884
rect 17084 35769 17158 35851
rect 17084 35611 17141 35769
tri 17177 35736 17193 35752 se
rect 17193 35736 17270 35752
rect 17177 35670 17270 35736
rect 17084 35535 17270 35611
rect 17084 35377 17141 35535
rect 17177 35410 17270 35476
tri 17177 35394 17193 35410 ne
rect 17193 35394 17270 35410
rect 17084 35295 17158 35377
rect 17084 35061 17141 35295
tri 17177 35262 17193 35278 se
rect 17193 35262 17270 35278
rect 17177 35196 17270 35262
rect 17177 35094 17270 35160
tri 17177 35078 17193 35094 ne
rect 17193 35078 17270 35094
rect 17084 34979 17158 35061
rect 17084 34821 17141 34979
tri 17177 34946 17193 34962 se
rect 17193 34946 17270 34962
rect 17177 34880 17270 34946
rect 17084 34745 17270 34821
rect 17084 34587 17141 34745
rect 17177 34620 17270 34686
tri 17177 34604 17193 34620 ne
rect 17193 34604 17270 34620
rect 17084 34505 17158 34587
rect 17084 34271 17141 34505
tri 17177 34472 17193 34488 se
rect 17193 34472 17270 34488
rect 17177 34406 17270 34472
rect 17177 34304 17270 34370
tri 17177 34288 17193 34304 ne
rect 17193 34288 17270 34304
rect 17084 34189 17158 34271
rect 17084 34031 17141 34189
tri 17177 34156 17193 34172 se
rect 17193 34156 17270 34172
rect 17177 34090 17270 34156
rect 17084 33955 17270 34031
rect 17084 33797 17141 33955
rect 17177 33830 17270 33896
tri 17177 33814 17193 33830 ne
rect 17193 33814 17270 33830
rect 17084 33715 17158 33797
rect 17084 33481 17141 33715
tri 17177 33682 17193 33698 se
rect 17193 33682 17270 33698
rect 17177 33616 17270 33682
rect 17177 33514 17270 33580
tri 17177 33498 17193 33514 ne
rect 17193 33498 17270 33514
rect 17084 33399 17158 33481
rect 17084 33241 17141 33399
tri 17177 33366 17193 33382 se
rect 17193 33366 17270 33382
rect 17177 33300 17270 33366
rect 17084 33165 17270 33241
rect 17084 33007 17141 33165
rect 17177 33040 17270 33106
tri 17177 33024 17193 33040 ne
rect 17193 33024 17270 33040
rect 17084 32925 17158 33007
rect 17084 32691 17141 32925
tri 17177 32892 17193 32908 se
rect 17193 32892 17270 32908
rect 17177 32826 17270 32892
rect 17177 32724 17270 32790
tri 17177 32708 17193 32724 ne
rect 17193 32708 17270 32724
rect 17084 32609 17158 32691
rect 17084 32451 17141 32609
tri 17177 32576 17193 32592 se
rect 17193 32576 17270 32592
rect 17177 32510 17270 32576
rect 17084 32375 17270 32451
rect 17084 32217 17141 32375
rect 17177 32250 17270 32316
tri 17177 32234 17193 32250 ne
rect 17193 32234 17270 32250
rect 17084 32135 17158 32217
rect 17084 31901 17141 32135
tri 17177 32102 17193 32118 se
rect 17193 32102 17270 32118
rect 17177 32036 17270 32102
rect 17177 31934 17270 32000
tri 17177 31918 17193 31934 ne
rect 17193 31918 17270 31934
rect 17084 31819 17158 31901
rect 17084 31661 17141 31819
tri 17177 31786 17193 31802 se
rect 17193 31786 17270 31802
rect 17177 31720 17270 31786
rect 17084 31585 17270 31661
rect 17084 31427 17141 31585
rect 17177 31460 17270 31526
tri 17177 31444 17193 31460 ne
rect 17193 31444 17270 31460
rect 17084 31345 17158 31427
rect 17084 31111 17141 31345
tri 17177 31312 17193 31328 se
rect 17193 31312 17270 31328
rect 17177 31246 17270 31312
rect 17177 31144 17270 31210
tri 17177 31128 17193 31144 ne
rect 17193 31128 17270 31144
rect 17084 31029 17158 31111
rect 17084 30871 17141 31029
tri 17177 30996 17193 31012 se
rect 17193 30996 17270 31012
rect 17177 30930 17270 30996
rect 17084 30795 17270 30871
rect 17084 30637 17141 30795
rect 17177 30670 17270 30736
tri 17177 30654 17193 30670 ne
rect 17193 30654 17270 30670
rect 17084 30555 17158 30637
rect 17084 30321 17141 30555
tri 17177 30522 17193 30538 se
rect 17193 30522 17270 30538
rect 17177 30456 17270 30522
rect 17177 30354 17270 30420
tri 17177 30338 17193 30354 ne
rect 17193 30338 17270 30354
rect 17084 30239 17158 30321
rect 17084 30081 17141 30239
tri 17177 30206 17193 30222 se
rect 17193 30206 17270 30222
rect 17177 30140 17270 30206
rect 17084 30005 17270 30081
rect 17084 29847 17141 30005
rect 17177 29880 17270 29946
tri 17177 29864 17193 29880 ne
rect 17193 29864 17270 29880
rect 17084 29765 17158 29847
rect 17084 29531 17141 29765
tri 17177 29732 17193 29748 se
rect 17193 29732 17270 29748
rect 17177 29666 17270 29732
rect 17177 29564 17270 29630
tri 17177 29548 17193 29564 ne
rect 17193 29548 17270 29564
rect 17084 29449 17158 29531
rect 17084 29291 17141 29449
tri 17177 29416 17193 29432 se
rect 17193 29416 17270 29432
rect 17177 29350 17270 29416
rect 17084 29215 17270 29291
rect 17084 29057 17141 29215
rect 17177 29090 17270 29156
tri 17177 29074 17193 29090 ne
rect 17193 29074 17270 29090
rect 17084 28975 17158 29057
rect 17084 28833 17141 28975
tri 17177 28942 17193 28958 se
rect 17193 28942 17270 28958
rect 17177 28876 17270 28942
rect 17306 28463 17342 80603
rect 17378 28463 17414 80603
rect 17450 80445 17486 80603
rect 17442 80303 17494 80445
rect 17450 28763 17486 80303
rect 17442 28621 17494 28763
rect 17450 28463 17486 28621
rect 17522 28463 17558 80603
rect 17594 28463 17630 80603
rect 17666 28833 17750 80233
rect 17786 28463 17822 80603
rect 17858 28463 17894 80603
rect 17930 80445 17966 80603
rect 17922 80303 17974 80445
rect 17930 28763 17966 80303
rect 17922 28621 17974 28763
rect 17930 28463 17966 28621
rect 18002 28463 18038 80603
rect 18074 28463 18110 80603
rect 18146 80124 18239 80190
rect 18146 80108 18223 80124
tri 18223 80108 18239 80124 nw
rect 18275 80091 18389 80233
rect 18425 80124 18518 80190
tri 18425 80108 18441 80124 ne
rect 18441 80108 18518 80124
rect 18258 80009 18406 80091
rect 18146 79976 18223 79992
tri 18223 79976 18239 79992 sw
rect 18146 79910 18239 79976
rect 18275 79851 18389 80009
tri 18425 79976 18441 79992 se
rect 18441 79976 18518 79992
rect 18425 79910 18518 79976
rect 18146 79775 18518 79851
rect 18146 79650 18239 79716
rect 18146 79634 18223 79650
tri 18223 79634 18239 79650 nw
rect 18275 79617 18389 79775
rect 18425 79650 18518 79716
tri 18425 79634 18441 79650 ne
rect 18441 79634 18518 79650
rect 18258 79535 18406 79617
rect 18146 79502 18223 79518
tri 18223 79502 18239 79518 sw
rect 18146 79436 18239 79502
rect 18146 79334 18239 79400
rect 18146 79318 18223 79334
tri 18223 79318 18239 79334 nw
rect 18275 79301 18389 79535
tri 18425 79502 18441 79518 se
rect 18441 79502 18518 79518
rect 18425 79436 18518 79502
rect 18425 79334 18518 79400
tri 18425 79318 18441 79334 ne
rect 18441 79318 18518 79334
rect 18258 79219 18406 79301
rect 18146 79186 18223 79202
tri 18223 79186 18239 79202 sw
rect 18146 79120 18239 79186
rect 18275 79061 18389 79219
tri 18425 79186 18441 79202 se
rect 18441 79186 18518 79202
rect 18425 79120 18518 79186
rect 18146 78985 18518 79061
rect 18146 78860 18239 78926
rect 18146 78844 18223 78860
tri 18223 78844 18239 78860 nw
rect 18275 78827 18389 78985
rect 18425 78860 18518 78926
tri 18425 78844 18441 78860 ne
rect 18441 78844 18518 78860
rect 18258 78745 18406 78827
rect 18146 78712 18223 78728
tri 18223 78712 18239 78728 sw
rect 18146 78646 18239 78712
rect 18146 78544 18239 78610
rect 18146 78528 18223 78544
tri 18223 78528 18239 78544 nw
rect 18275 78511 18389 78745
tri 18425 78712 18441 78728 se
rect 18441 78712 18518 78728
rect 18425 78646 18518 78712
rect 18425 78544 18518 78610
tri 18425 78528 18441 78544 ne
rect 18441 78528 18518 78544
rect 18258 78429 18406 78511
rect 18146 78396 18223 78412
tri 18223 78396 18239 78412 sw
rect 18146 78330 18239 78396
rect 18275 78271 18389 78429
tri 18425 78396 18441 78412 se
rect 18441 78396 18518 78412
rect 18425 78330 18518 78396
rect 18146 78195 18518 78271
rect 18146 78070 18239 78136
rect 18146 78054 18223 78070
tri 18223 78054 18239 78070 nw
rect 18275 78037 18389 78195
rect 18425 78070 18518 78136
tri 18425 78054 18441 78070 ne
rect 18441 78054 18518 78070
rect 18258 77955 18406 78037
rect 18146 77922 18223 77938
tri 18223 77922 18239 77938 sw
rect 18146 77856 18239 77922
rect 18146 77754 18239 77820
rect 18146 77738 18223 77754
tri 18223 77738 18239 77754 nw
rect 18275 77721 18389 77955
tri 18425 77922 18441 77938 se
rect 18441 77922 18518 77938
rect 18425 77856 18518 77922
rect 18425 77754 18518 77820
tri 18425 77738 18441 77754 ne
rect 18441 77738 18518 77754
rect 18258 77639 18406 77721
rect 18146 77606 18223 77622
tri 18223 77606 18239 77622 sw
rect 18146 77540 18239 77606
rect 18275 77481 18389 77639
tri 18425 77606 18441 77622 se
rect 18441 77606 18518 77622
rect 18425 77540 18518 77606
rect 18146 77405 18518 77481
rect 18146 77280 18239 77346
rect 18146 77264 18223 77280
tri 18223 77264 18239 77280 nw
rect 18275 77247 18389 77405
rect 18425 77280 18518 77346
tri 18425 77264 18441 77280 ne
rect 18441 77264 18518 77280
rect 18258 77165 18406 77247
rect 18146 77132 18223 77148
tri 18223 77132 18239 77148 sw
rect 18146 77066 18239 77132
rect 18146 76964 18239 77030
rect 18146 76948 18223 76964
tri 18223 76948 18239 76964 nw
rect 18275 76931 18389 77165
tri 18425 77132 18441 77148 se
rect 18441 77132 18518 77148
rect 18425 77066 18518 77132
rect 18425 76964 18518 77030
tri 18425 76948 18441 76964 ne
rect 18441 76948 18518 76964
rect 18258 76849 18406 76931
rect 18146 76816 18223 76832
tri 18223 76816 18239 76832 sw
rect 18146 76750 18239 76816
rect 18275 76691 18389 76849
tri 18425 76816 18441 76832 se
rect 18441 76816 18518 76832
rect 18425 76750 18518 76816
rect 18146 76615 18518 76691
rect 18146 76490 18239 76556
rect 18146 76474 18223 76490
tri 18223 76474 18239 76490 nw
rect 18275 76457 18389 76615
rect 18425 76490 18518 76556
tri 18425 76474 18441 76490 ne
rect 18441 76474 18518 76490
rect 18258 76375 18406 76457
rect 18146 76342 18223 76358
tri 18223 76342 18239 76358 sw
rect 18146 76276 18239 76342
rect 18146 76174 18239 76240
rect 18146 76158 18223 76174
tri 18223 76158 18239 76174 nw
rect 18275 76141 18389 76375
tri 18425 76342 18441 76358 se
rect 18441 76342 18518 76358
rect 18425 76276 18518 76342
rect 18425 76174 18518 76240
tri 18425 76158 18441 76174 ne
rect 18441 76158 18518 76174
rect 18258 76059 18406 76141
rect 18146 76026 18223 76042
tri 18223 76026 18239 76042 sw
rect 18146 75960 18239 76026
rect 18275 75901 18389 76059
tri 18425 76026 18441 76042 se
rect 18441 76026 18518 76042
rect 18425 75960 18518 76026
rect 18146 75825 18518 75901
rect 18146 75700 18239 75766
rect 18146 75684 18223 75700
tri 18223 75684 18239 75700 nw
rect 18275 75667 18389 75825
rect 18425 75700 18518 75766
tri 18425 75684 18441 75700 ne
rect 18441 75684 18518 75700
rect 18258 75585 18406 75667
rect 18146 75552 18223 75568
tri 18223 75552 18239 75568 sw
rect 18146 75486 18239 75552
rect 18146 75384 18239 75450
rect 18146 75368 18223 75384
tri 18223 75368 18239 75384 nw
rect 18275 75351 18389 75585
tri 18425 75552 18441 75568 se
rect 18441 75552 18518 75568
rect 18425 75486 18518 75552
rect 18425 75384 18518 75450
tri 18425 75368 18441 75384 ne
rect 18441 75368 18518 75384
rect 18258 75269 18406 75351
rect 18146 75236 18223 75252
tri 18223 75236 18239 75252 sw
rect 18146 75170 18239 75236
rect 18275 75111 18389 75269
tri 18425 75236 18441 75252 se
rect 18441 75236 18518 75252
rect 18425 75170 18518 75236
rect 18146 75035 18518 75111
rect 18146 74910 18239 74976
rect 18146 74894 18223 74910
tri 18223 74894 18239 74910 nw
rect 18275 74877 18389 75035
rect 18425 74910 18518 74976
tri 18425 74894 18441 74910 ne
rect 18441 74894 18518 74910
rect 18258 74795 18406 74877
rect 18146 74762 18223 74778
tri 18223 74762 18239 74778 sw
rect 18146 74696 18239 74762
rect 18146 74594 18239 74660
rect 18146 74578 18223 74594
tri 18223 74578 18239 74594 nw
rect 18275 74561 18389 74795
tri 18425 74762 18441 74778 se
rect 18441 74762 18518 74778
rect 18425 74696 18518 74762
rect 18425 74594 18518 74660
tri 18425 74578 18441 74594 ne
rect 18441 74578 18518 74594
rect 18258 74479 18406 74561
rect 18146 74446 18223 74462
tri 18223 74446 18239 74462 sw
rect 18146 74380 18239 74446
rect 18275 74321 18389 74479
tri 18425 74446 18441 74462 se
rect 18441 74446 18518 74462
rect 18425 74380 18518 74446
rect 18146 74245 18518 74321
rect 18146 74120 18239 74186
rect 18146 74104 18223 74120
tri 18223 74104 18239 74120 nw
rect 18275 74087 18389 74245
rect 18425 74120 18518 74186
tri 18425 74104 18441 74120 ne
rect 18441 74104 18518 74120
rect 18258 74005 18406 74087
rect 18146 73972 18223 73988
tri 18223 73972 18239 73988 sw
rect 18146 73906 18239 73972
rect 18146 73804 18239 73870
rect 18146 73788 18223 73804
tri 18223 73788 18239 73804 nw
rect 18275 73771 18389 74005
tri 18425 73972 18441 73988 se
rect 18441 73972 18518 73988
rect 18425 73906 18518 73972
rect 18425 73804 18518 73870
tri 18425 73788 18441 73804 ne
rect 18441 73788 18518 73804
rect 18258 73689 18406 73771
rect 18146 73656 18223 73672
tri 18223 73656 18239 73672 sw
rect 18146 73590 18239 73656
rect 18275 73531 18389 73689
tri 18425 73656 18441 73672 se
rect 18441 73656 18518 73672
rect 18425 73590 18518 73656
rect 18146 73455 18518 73531
rect 18146 73330 18239 73396
rect 18146 73314 18223 73330
tri 18223 73314 18239 73330 nw
rect 18275 73297 18389 73455
rect 18425 73330 18518 73396
tri 18425 73314 18441 73330 ne
rect 18441 73314 18518 73330
rect 18258 73215 18406 73297
rect 18146 73182 18223 73198
tri 18223 73182 18239 73198 sw
rect 18146 73116 18239 73182
rect 18146 73014 18239 73080
rect 18146 72998 18223 73014
tri 18223 72998 18239 73014 nw
rect 18275 72981 18389 73215
tri 18425 73182 18441 73198 se
rect 18441 73182 18518 73198
rect 18425 73116 18518 73182
rect 18425 73014 18518 73080
tri 18425 72998 18441 73014 ne
rect 18441 72998 18518 73014
rect 18258 72899 18406 72981
rect 18146 72866 18223 72882
tri 18223 72866 18239 72882 sw
rect 18146 72800 18239 72866
rect 18275 72741 18389 72899
tri 18425 72866 18441 72882 se
rect 18441 72866 18518 72882
rect 18425 72800 18518 72866
rect 18146 72665 18518 72741
rect 18146 72540 18239 72606
rect 18146 72524 18223 72540
tri 18223 72524 18239 72540 nw
rect 18275 72507 18389 72665
rect 18425 72540 18518 72606
tri 18425 72524 18441 72540 ne
rect 18441 72524 18518 72540
rect 18258 72425 18406 72507
rect 18146 72392 18223 72408
tri 18223 72392 18239 72408 sw
rect 18146 72326 18239 72392
rect 18146 72224 18239 72290
rect 18146 72208 18223 72224
tri 18223 72208 18239 72224 nw
rect 18275 72191 18389 72425
tri 18425 72392 18441 72408 se
rect 18441 72392 18518 72408
rect 18425 72326 18518 72392
rect 18425 72224 18518 72290
tri 18425 72208 18441 72224 ne
rect 18441 72208 18518 72224
rect 18258 72109 18406 72191
rect 18146 72076 18223 72092
tri 18223 72076 18239 72092 sw
rect 18146 72010 18239 72076
rect 18275 71951 18389 72109
tri 18425 72076 18441 72092 se
rect 18441 72076 18518 72092
rect 18425 72010 18518 72076
rect 18146 71875 18518 71951
rect 18146 71750 18239 71816
rect 18146 71734 18223 71750
tri 18223 71734 18239 71750 nw
rect 18275 71717 18389 71875
rect 18425 71750 18518 71816
tri 18425 71734 18441 71750 ne
rect 18441 71734 18518 71750
rect 18258 71635 18406 71717
rect 18146 71602 18223 71618
tri 18223 71602 18239 71618 sw
rect 18146 71536 18239 71602
rect 18146 71434 18239 71500
rect 18146 71418 18223 71434
tri 18223 71418 18239 71434 nw
rect 18275 71401 18389 71635
tri 18425 71602 18441 71618 se
rect 18441 71602 18518 71618
rect 18425 71536 18518 71602
rect 18425 71434 18518 71500
tri 18425 71418 18441 71434 ne
rect 18441 71418 18518 71434
rect 18258 71319 18406 71401
rect 18146 71286 18223 71302
tri 18223 71286 18239 71302 sw
rect 18146 71220 18239 71286
rect 18275 71161 18389 71319
tri 18425 71286 18441 71302 se
rect 18441 71286 18518 71302
rect 18425 71220 18518 71286
rect 18146 71085 18518 71161
rect 18146 70960 18239 71026
rect 18146 70944 18223 70960
tri 18223 70944 18239 70960 nw
rect 18275 70927 18389 71085
rect 18425 70960 18518 71026
tri 18425 70944 18441 70960 ne
rect 18441 70944 18518 70960
rect 18258 70845 18406 70927
rect 18146 70812 18223 70828
tri 18223 70812 18239 70828 sw
rect 18146 70746 18239 70812
rect 18146 70644 18239 70710
rect 18146 70628 18223 70644
tri 18223 70628 18239 70644 nw
rect 18275 70611 18389 70845
tri 18425 70812 18441 70828 se
rect 18441 70812 18518 70828
rect 18425 70746 18518 70812
rect 18425 70644 18518 70710
tri 18425 70628 18441 70644 ne
rect 18441 70628 18518 70644
rect 18258 70529 18406 70611
rect 18146 70496 18223 70512
tri 18223 70496 18239 70512 sw
rect 18146 70430 18239 70496
rect 18275 70371 18389 70529
tri 18425 70496 18441 70512 se
rect 18441 70496 18518 70512
rect 18425 70430 18518 70496
rect 18146 70295 18518 70371
rect 18146 70170 18239 70236
rect 18146 70154 18223 70170
tri 18223 70154 18239 70170 nw
rect 18275 70137 18389 70295
rect 18425 70170 18518 70236
tri 18425 70154 18441 70170 ne
rect 18441 70154 18518 70170
rect 18258 70055 18406 70137
rect 18146 70022 18223 70038
tri 18223 70022 18239 70038 sw
rect 18146 69956 18239 70022
rect 18146 69854 18239 69920
rect 18146 69838 18223 69854
tri 18223 69838 18239 69854 nw
rect 18275 69821 18389 70055
tri 18425 70022 18441 70038 se
rect 18441 70022 18518 70038
rect 18425 69956 18518 70022
rect 18425 69854 18518 69920
tri 18425 69838 18441 69854 ne
rect 18441 69838 18518 69854
rect 18258 69739 18406 69821
rect 18146 69706 18223 69722
tri 18223 69706 18239 69722 sw
rect 18146 69640 18239 69706
rect 18275 69581 18389 69739
tri 18425 69706 18441 69722 se
rect 18441 69706 18518 69722
rect 18425 69640 18518 69706
rect 18146 69505 18518 69581
rect 18146 69380 18239 69446
rect 18146 69364 18223 69380
tri 18223 69364 18239 69380 nw
rect 18275 69347 18389 69505
rect 18425 69380 18518 69446
tri 18425 69364 18441 69380 ne
rect 18441 69364 18518 69380
rect 18258 69265 18406 69347
rect 18146 69232 18223 69248
tri 18223 69232 18239 69248 sw
rect 18146 69166 18239 69232
rect 18146 69064 18239 69130
rect 18146 69048 18223 69064
tri 18223 69048 18239 69064 nw
rect 18275 69031 18389 69265
tri 18425 69232 18441 69248 se
rect 18441 69232 18518 69248
rect 18425 69166 18518 69232
rect 18425 69064 18518 69130
tri 18425 69048 18441 69064 ne
rect 18441 69048 18518 69064
rect 18258 68949 18406 69031
rect 18146 68916 18223 68932
tri 18223 68916 18239 68932 sw
rect 18146 68850 18239 68916
rect 18275 68791 18389 68949
tri 18425 68916 18441 68932 se
rect 18441 68916 18518 68932
rect 18425 68850 18518 68916
rect 18146 68715 18518 68791
rect 18146 68590 18239 68656
rect 18146 68574 18223 68590
tri 18223 68574 18239 68590 nw
rect 18275 68557 18389 68715
rect 18425 68590 18518 68656
tri 18425 68574 18441 68590 ne
rect 18441 68574 18518 68590
rect 18258 68475 18406 68557
rect 18146 68442 18223 68458
tri 18223 68442 18239 68458 sw
rect 18146 68376 18239 68442
rect 18146 68274 18239 68340
rect 18146 68258 18223 68274
tri 18223 68258 18239 68274 nw
rect 18275 68241 18389 68475
tri 18425 68442 18441 68458 se
rect 18441 68442 18518 68458
rect 18425 68376 18518 68442
rect 18425 68274 18518 68340
tri 18425 68258 18441 68274 ne
rect 18441 68258 18518 68274
rect 18258 68159 18406 68241
rect 18146 68126 18223 68142
tri 18223 68126 18239 68142 sw
rect 18146 68060 18239 68126
rect 18275 68001 18389 68159
tri 18425 68126 18441 68142 se
rect 18441 68126 18518 68142
rect 18425 68060 18518 68126
rect 18146 67925 18518 68001
rect 18146 67800 18239 67866
rect 18146 67784 18223 67800
tri 18223 67784 18239 67800 nw
rect 18275 67767 18389 67925
rect 18425 67800 18518 67866
tri 18425 67784 18441 67800 ne
rect 18441 67784 18518 67800
rect 18258 67685 18406 67767
rect 18146 67652 18223 67668
tri 18223 67652 18239 67668 sw
rect 18146 67586 18239 67652
rect 18146 67484 18239 67550
rect 18146 67468 18223 67484
tri 18223 67468 18239 67484 nw
rect 18275 67451 18389 67685
tri 18425 67652 18441 67668 se
rect 18441 67652 18518 67668
rect 18425 67586 18518 67652
rect 18425 67484 18518 67550
tri 18425 67468 18441 67484 ne
rect 18441 67468 18518 67484
rect 18258 67369 18406 67451
rect 18146 67336 18223 67352
tri 18223 67336 18239 67352 sw
rect 18146 67270 18239 67336
rect 18275 67211 18389 67369
tri 18425 67336 18441 67352 se
rect 18441 67336 18518 67352
rect 18425 67270 18518 67336
rect 18146 67135 18518 67211
rect 18146 67010 18239 67076
rect 18146 66994 18223 67010
tri 18223 66994 18239 67010 nw
rect 18275 66977 18389 67135
rect 18425 67010 18518 67076
tri 18425 66994 18441 67010 ne
rect 18441 66994 18518 67010
rect 18258 66895 18406 66977
rect 18146 66862 18223 66878
tri 18223 66862 18239 66878 sw
rect 18146 66796 18239 66862
rect 18146 66694 18239 66760
rect 18146 66678 18223 66694
tri 18223 66678 18239 66694 nw
rect 18275 66661 18389 66895
tri 18425 66862 18441 66878 se
rect 18441 66862 18518 66878
rect 18425 66796 18518 66862
rect 18425 66694 18518 66760
tri 18425 66678 18441 66694 ne
rect 18441 66678 18518 66694
rect 18258 66579 18406 66661
rect 18146 66546 18223 66562
tri 18223 66546 18239 66562 sw
rect 18146 66480 18239 66546
rect 18275 66421 18389 66579
tri 18425 66546 18441 66562 se
rect 18441 66546 18518 66562
rect 18425 66480 18518 66546
rect 18146 66345 18518 66421
rect 18146 66220 18239 66286
rect 18146 66204 18223 66220
tri 18223 66204 18239 66220 nw
rect 18275 66187 18389 66345
rect 18425 66220 18518 66286
tri 18425 66204 18441 66220 ne
rect 18441 66204 18518 66220
rect 18258 66105 18406 66187
rect 18146 66072 18223 66088
tri 18223 66072 18239 66088 sw
rect 18146 66006 18239 66072
rect 18146 65904 18239 65970
rect 18146 65888 18223 65904
tri 18223 65888 18239 65904 nw
rect 18275 65871 18389 66105
tri 18425 66072 18441 66088 se
rect 18441 66072 18518 66088
rect 18425 66006 18518 66072
rect 18425 65904 18518 65970
tri 18425 65888 18441 65904 ne
rect 18441 65888 18518 65904
rect 18258 65789 18406 65871
rect 18146 65756 18223 65772
tri 18223 65756 18239 65772 sw
rect 18146 65690 18239 65756
rect 18275 65631 18389 65789
tri 18425 65756 18441 65772 se
rect 18441 65756 18518 65772
rect 18425 65690 18518 65756
rect 18146 65555 18518 65631
rect 18146 65430 18239 65496
rect 18146 65414 18223 65430
tri 18223 65414 18239 65430 nw
rect 18275 65397 18389 65555
rect 18425 65430 18518 65496
tri 18425 65414 18441 65430 ne
rect 18441 65414 18518 65430
rect 18258 65315 18406 65397
rect 18146 65282 18223 65298
tri 18223 65282 18239 65298 sw
rect 18146 65216 18239 65282
rect 18146 65114 18239 65180
rect 18146 65098 18223 65114
tri 18223 65098 18239 65114 nw
rect 18275 65081 18389 65315
tri 18425 65282 18441 65298 se
rect 18441 65282 18518 65298
rect 18425 65216 18518 65282
rect 18425 65114 18518 65180
tri 18425 65098 18441 65114 ne
rect 18441 65098 18518 65114
rect 18258 64999 18406 65081
rect 18146 64966 18223 64982
tri 18223 64966 18239 64982 sw
rect 18146 64900 18239 64966
rect 18275 64841 18389 64999
tri 18425 64966 18441 64982 se
rect 18441 64966 18518 64982
rect 18425 64900 18518 64966
rect 18146 64765 18518 64841
rect 18146 64640 18239 64706
rect 18146 64624 18223 64640
tri 18223 64624 18239 64640 nw
rect 18275 64607 18389 64765
rect 18425 64640 18518 64706
tri 18425 64624 18441 64640 ne
rect 18441 64624 18518 64640
rect 18258 64525 18406 64607
rect 18146 64492 18223 64508
tri 18223 64492 18239 64508 sw
rect 18146 64426 18239 64492
rect 18146 64324 18239 64390
rect 18146 64308 18223 64324
tri 18223 64308 18239 64324 nw
rect 18275 64291 18389 64525
tri 18425 64492 18441 64508 se
rect 18441 64492 18518 64508
rect 18425 64426 18518 64492
rect 18425 64324 18518 64390
tri 18425 64308 18441 64324 ne
rect 18441 64308 18518 64324
rect 18258 64209 18406 64291
rect 18146 64176 18223 64192
tri 18223 64176 18239 64192 sw
rect 18146 64110 18239 64176
rect 18275 64051 18389 64209
tri 18425 64176 18441 64192 se
rect 18441 64176 18518 64192
rect 18425 64110 18518 64176
rect 18146 63975 18518 64051
rect 18146 63850 18239 63916
rect 18146 63834 18223 63850
tri 18223 63834 18239 63850 nw
rect 18275 63817 18389 63975
rect 18425 63850 18518 63916
tri 18425 63834 18441 63850 ne
rect 18441 63834 18518 63850
rect 18258 63735 18406 63817
rect 18146 63702 18223 63718
tri 18223 63702 18239 63718 sw
rect 18146 63636 18239 63702
rect 18146 63534 18239 63600
rect 18146 63518 18223 63534
tri 18223 63518 18239 63534 nw
rect 18275 63501 18389 63735
tri 18425 63702 18441 63718 se
rect 18441 63702 18518 63718
rect 18425 63636 18518 63702
rect 18425 63534 18518 63600
tri 18425 63518 18441 63534 ne
rect 18441 63518 18518 63534
rect 18258 63419 18406 63501
rect 18146 63386 18223 63402
tri 18223 63386 18239 63402 sw
rect 18146 63320 18239 63386
rect 18275 63261 18389 63419
tri 18425 63386 18441 63402 se
rect 18441 63386 18518 63402
rect 18425 63320 18518 63386
rect 18146 63185 18518 63261
rect 18146 63060 18239 63126
rect 18146 63044 18223 63060
tri 18223 63044 18239 63060 nw
rect 18275 63027 18389 63185
rect 18425 63060 18518 63126
tri 18425 63044 18441 63060 ne
rect 18441 63044 18518 63060
rect 18258 62945 18406 63027
rect 18146 62912 18223 62928
tri 18223 62912 18239 62928 sw
rect 18146 62846 18239 62912
rect 18146 62744 18239 62810
rect 18146 62728 18223 62744
tri 18223 62728 18239 62744 nw
rect 18275 62711 18389 62945
tri 18425 62912 18441 62928 se
rect 18441 62912 18518 62928
rect 18425 62846 18518 62912
rect 18425 62744 18518 62810
tri 18425 62728 18441 62744 ne
rect 18441 62728 18518 62744
rect 18258 62629 18406 62711
rect 18146 62596 18223 62612
tri 18223 62596 18239 62612 sw
rect 18146 62530 18239 62596
rect 18275 62471 18389 62629
tri 18425 62596 18441 62612 se
rect 18441 62596 18518 62612
rect 18425 62530 18518 62596
rect 18146 62395 18518 62471
rect 18146 62270 18239 62336
rect 18146 62254 18223 62270
tri 18223 62254 18239 62270 nw
rect 18275 62237 18389 62395
rect 18425 62270 18518 62336
tri 18425 62254 18441 62270 ne
rect 18441 62254 18518 62270
rect 18258 62155 18406 62237
rect 18146 62122 18223 62138
tri 18223 62122 18239 62138 sw
rect 18146 62056 18239 62122
rect 18146 61954 18239 62020
rect 18146 61938 18223 61954
tri 18223 61938 18239 61954 nw
rect 18275 61921 18389 62155
tri 18425 62122 18441 62138 se
rect 18441 62122 18518 62138
rect 18425 62056 18518 62122
rect 18425 61954 18518 62020
tri 18425 61938 18441 61954 ne
rect 18441 61938 18518 61954
rect 18258 61839 18406 61921
rect 18146 61806 18223 61822
tri 18223 61806 18239 61822 sw
rect 18146 61740 18239 61806
rect 18275 61681 18389 61839
tri 18425 61806 18441 61822 se
rect 18441 61806 18518 61822
rect 18425 61740 18518 61806
rect 18146 61605 18518 61681
rect 18146 61480 18239 61546
rect 18146 61464 18223 61480
tri 18223 61464 18239 61480 nw
rect 18275 61447 18389 61605
rect 18425 61480 18518 61546
tri 18425 61464 18441 61480 ne
rect 18441 61464 18518 61480
rect 18258 61365 18406 61447
rect 18146 61332 18223 61348
tri 18223 61332 18239 61348 sw
rect 18146 61266 18239 61332
rect 18146 61164 18239 61230
rect 18146 61148 18223 61164
tri 18223 61148 18239 61164 nw
rect 18275 61131 18389 61365
tri 18425 61332 18441 61348 se
rect 18441 61332 18518 61348
rect 18425 61266 18518 61332
rect 18425 61164 18518 61230
tri 18425 61148 18441 61164 ne
rect 18441 61148 18518 61164
rect 18258 61049 18406 61131
rect 18146 61016 18223 61032
tri 18223 61016 18239 61032 sw
rect 18146 60950 18239 61016
rect 18275 60891 18389 61049
tri 18425 61016 18441 61032 se
rect 18441 61016 18518 61032
rect 18425 60950 18518 61016
rect 18146 60815 18518 60891
rect 18146 60690 18239 60756
rect 18146 60674 18223 60690
tri 18223 60674 18239 60690 nw
rect 18275 60657 18389 60815
rect 18425 60690 18518 60756
tri 18425 60674 18441 60690 ne
rect 18441 60674 18518 60690
rect 18258 60575 18406 60657
rect 18146 60542 18223 60558
tri 18223 60542 18239 60558 sw
rect 18146 60476 18239 60542
rect 18146 60374 18239 60440
rect 18146 60358 18223 60374
tri 18223 60358 18239 60374 nw
rect 18275 60341 18389 60575
tri 18425 60542 18441 60558 se
rect 18441 60542 18518 60558
rect 18425 60476 18518 60542
rect 18425 60374 18518 60440
tri 18425 60358 18441 60374 ne
rect 18441 60358 18518 60374
rect 18258 60259 18406 60341
rect 18146 60226 18223 60242
tri 18223 60226 18239 60242 sw
rect 18146 60160 18239 60226
rect 18275 60101 18389 60259
tri 18425 60226 18441 60242 se
rect 18441 60226 18518 60242
rect 18425 60160 18518 60226
rect 18146 60025 18518 60101
rect 18146 59900 18239 59966
rect 18146 59884 18223 59900
tri 18223 59884 18239 59900 nw
rect 18275 59867 18389 60025
rect 18425 59900 18518 59966
tri 18425 59884 18441 59900 ne
rect 18441 59884 18518 59900
rect 18258 59785 18406 59867
rect 18146 59752 18223 59768
tri 18223 59752 18239 59768 sw
rect 18146 59686 18239 59752
rect 18146 59584 18239 59650
rect 18146 59568 18223 59584
tri 18223 59568 18239 59584 nw
rect 18275 59551 18389 59785
tri 18425 59752 18441 59768 se
rect 18441 59752 18518 59768
rect 18425 59686 18518 59752
rect 18425 59584 18518 59650
tri 18425 59568 18441 59584 ne
rect 18441 59568 18518 59584
rect 18258 59469 18406 59551
rect 18146 59436 18223 59452
tri 18223 59436 18239 59452 sw
rect 18146 59370 18239 59436
rect 18275 59311 18389 59469
tri 18425 59436 18441 59452 se
rect 18441 59436 18518 59452
rect 18425 59370 18518 59436
rect 18146 59235 18518 59311
rect 18146 59110 18239 59176
rect 18146 59094 18223 59110
tri 18223 59094 18239 59110 nw
rect 18275 59077 18389 59235
rect 18425 59110 18518 59176
tri 18425 59094 18441 59110 ne
rect 18441 59094 18518 59110
rect 18258 58995 18406 59077
rect 18146 58962 18223 58978
tri 18223 58962 18239 58978 sw
rect 18146 58896 18239 58962
rect 18146 58794 18239 58860
rect 18146 58778 18223 58794
tri 18223 58778 18239 58794 nw
rect 18275 58761 18389 58995
tri 18425 58962 18441 58978 se
rect 18441 58962 18518 58978
rect 18425 58896 18518 58962
rect 18425 58794 18518 58860
tri 18425 58778 18441 58794 ne
rect 18441 58778 18518 58794
rect 18258 58679 18406 58761
rect 18146 58646 18223 58662
tri 18223 58646 18239 58662 sw
rect 18146 58580 18239 58646
rect 18275 58521 18389 58679
tri 18425 58646 18441 58662 se
rect 18441 58646 18518 58662
rect 18425 58580 18518 58646
rect 18146 58445 18518 58521
rect 18146 58320 18239 58386
rect 18146 58304 18223 58320
tri 18223 58304 18239 58320 nw
rect 18275 58287 18389 58445
rect 18425 58320 18518 58386
tri 18425 58304 18441 58320 ne
rect 18441 58304 18518 58320
rect 18258 58205 18406 58287
rect 18146 58172 18223 58188
tri 18223 58172 18239 58188 sw
rect 18146 58106 18239 58172
rect 18146 58004 18239 58070
rect 18146 57988 18223 58004
tri 18223 57988 18239 58004 nw
rect 18275 57971 18389 58205
tri 18425 58172 18441 58188 se
rect 18441 58172 18518 58188
rect 18425 58106 18518 58172
rect 18425 58004 18518 58070
tri 18425 57988 18441 58004 ne
rect 18441 57988 18518 58004
rect 18258 57889 18406 57971
rect 18146 57856 18223 57872
tri 18223 57856 18239 57872 sw
rect 18146 57790 18239 57856
rect 18275 57731 18389 57889
tri 18425 57856 18441 57872 se
rect 18441 57856 18518 57872
rect 18425 57790 18518 57856
rect 18146 57655 18518 57731
rect 18146 57530 18239 57596
rect 18146 57514 18223 57530
tri 18223 57514 18239 57530 nw
rect 18275 57497 18389 57655
rect 18425 57530 18518 57596
tri 18425 57514 18441 57530 ne
rect 18441 57514 18518 57530
rect 18258 57415 18406 57497
rect 18146 57382 18223 57398
tri 18223 57382 18239 57398 sw
rect 18146 57316 18239 57382
rect 18146 57214 18239 57280
rect 18146 57198 18223 57214
tri 18223 57198 18239 57214 nw
rect 18275 57181 18389 57415
tri 18425 57382 18441 57398 se
rect 18441 57382 18518 57398
rect 18425 57316 18518 57382
rect 18425 57214 18518 57280
tri 18425 57198 18441 57214 ne
rect 18441 57198 18518 57214
rect 18258 57099 18406 57181
rect 18146 57066 18223 57082
tri 18223 57066 18239 57082 sw
rect 18146 57000 18239 57066
rect 18275 56941 18389 57099
tri 18425 57066 18441 57082 se
rect 18441 57066 18518 57082
rect 18425 57000 18518 57066
rect 18146 56865 18518 56941
rect 18146 56740 18239 56806
rect 18146 56724 18223 56740
tri 18223 56724 18239 56740 nw
rect 18275 56707 18389 56865
rect 18425 56740 18518 56806
tri 18425 56724 18441 56740 ne
rect 18441 56724 18518 56740
rect 18258 56625 18406 56707
rect 18146 56592 18223 56608
tri 18223 56592 18239 56608 sw
rect 18146 56526 18239 56592
rect 18146 56424 18239 56490
rect 18146 56408 18223 56424
tri 18223 56408 18239 56424 nw
rect 18275 56391 18389 56625
tri 18425 56592 18441 56608 se
rect 18441 56592 18518 56608
rect 18425 56526 18518 56592
rect 18425 56424 18518 56490
tri 18425 56408 18441 56424 ne
rect 18441 56408 18518 56424
rect 18258 56309 18406 56391
rect 18146 56276 18223 56292
tri 18223 56276 18239 56292 sw
rect 18146 56210 18239 56276
rect 18275 56151 18389 56309
tri 18425 56276 18441 56292 se
rect 18441 56276 18518 56292
rect 18425 56210 18518 56276
rect 18146 56075 18518 56151
rect 18146 55950 18239 56016
rect 18146 55934 18223 55950
tri 18223 55934 18239 55950 nw
rect 18275 55917 18389 56075
rect 18425 55950 18518 56016
tri 18425 55934 18441 55950 ne
rect 18441 55934 18518 55950
rect 18258 55835 18406 55917
rect 18146 55802 18223 55818
tri 18223 55802 18239 55818 sw
rect 18146 55736 18239 55802
rect 18146 55634 18239 55700
rect 18146 55618 18223 55634
tri 18223 55618 18239 55634 nw
rect 18275 55601 18389 55835
tri 18425 55802 18441 55818 se
rect 18441 55802 18518 55818
rect 18425 55736 18518 55802
rect 18425 55634 18518 55700
tri 18425 55618 18441 55634 ne
rect 18441 55618 18518 55634
rect 18258 55519 18406 55601
rect 18146 55486 18223 55502
tri 18223 55486 18239 55502 sw
rect 18146 55420 18239 55486
rect 18275 55361 18389 55519
tri 18425 55486 18441 55502 se
rect 18441 55486 18518 55502
rect 18425 55420 18518 55486
rect 18146 55285 18518 55361
rect 18146 55160 18239 55226
rect 18146 55144 18223 55160
tri 18223 55144 18239 55160 nw
rect 18275 55127 18389 55285
rect 18425 55160 18518 55226
tri 18425 55144 18441 55160 ne
rect 18441 55144 18518 55160
rect 18258 55045 18406 55127
rect 18146 55012 18223 55028
tri 18223 55012 18239 55028 sw
rect 18146 54946 18239 55012
rect 18146 54844 18239 54910
rect 18146 54828 18223 54844
tri 18223 54828 18239 54844 nw
rect 18275 54811 18389 55045
tri 18425 55012 18441 55028 se
rect 18441 55012 18518 55028
rect 18425 54946 18518 55012
rect 18425 54844 18518 54910
tri 18425 54828 18441 54844 ne
rect 18441 54828 18518 54844
rect 18258 54729 18406 54811
rect 18146 54696 18223 54712
tri 18223 54696 18239 54712 sw
rect 18146 54630 18239 54696
rect 18275 54571 18389 54729
tri 18425 54696 18441 54712 se
rect 18441 54696 18518 54712
rect 18425 54630 18518 54696
rect 18146 54495 18518 54571
rect 18146 54370 18239 54436
rect 18146 54354 18223 54370
tri 18223 54354 18239 54370 nw
rect 18275 54337 18389 54495
rect 18425 54370 18518 54436
tri 18425 54354 18441 54370 ne
rect 18441 54354 18518 54370
rect 18258 54255 18406 54337
rect 18146 54222 18223 54238
tri 18223 54222 18239 54238 sw
rect 18146 54156 18239 54222
rect 18146 54054 18239 54120
rect 18146 54038 18223 54054
tri 18223 54038 18239 54054 nw
rect 18275 54021 18389 54255
tri 18425 54222 18441 54238 se
rect 18441 54222 18518 54238
rect 18425 54156 18518 54222
rect 18425 54054 18518 54120
tri 18425 54038 18441 54054 ne
rect 18441 54038 18518 54054
rect 18258 53939 18406 54021
rect 18146 53906 18223 53922
tri 18223 53906 18239 53922 sw
rect 18146 53840 18239 53906
rect 18275 53781 18389 53939
tri 18425 53906 18441 53922 se
rect 18441 53906 18518 53922
rect 18425 53840 18518 53906
rect 18146 53705 18518 53781
rect 18146 53580 18239 53646
rect 18146 53564 18223 53580
tri 18223 53564 18239 53580 nw
rect 18275 53547 18389 53705
rect 18425 53580 18518 53646
tri 18425 53564 18441 53580 ne
rect 18441 53564 18518 53580
rect 18258 53465 18406 53547
rect 18146 53432 18223 53448
tri 18223 53432 18239 53448 sw
rect 18146 53366 18239 53432
rect 18146 53264 18239 53330
rect 18146 53248 18223 53264
tri 18223 53248 18239 53264 nw
rect 18275 53231 18389 53465
tri 18425 53432 18441 53448 se
rect 18441 53432 18518 53448
rect 18425 53366 18518 53432
rect 18425 53264 18518 53330
tri 18425 53248 18441 53264 ne
rect 18441 53248 18518 53264
rect 18258 53149 18406 53231
rect 18146 53116 18223 53132
tri 18223 53116 18239 53132 sw
rect 18146 53050 18239 53116
rect 18275 52991 18389 53149
tri 18425 53116 18441 53132 se
rect 18441 53116 18518 53132
rect 18425 53050 18518 53116
rect 18146 52915 18518 52991
rect 18146 52790 18239 52856
rect 18146 52774 18223 52790
tri 18223 52774 18239 52790 nw
rect 18275 52757 18389 52915
rect 18425 52790 18518 52856
tri 18425 52774 18441 52790 ne
rect 18441 52774 18518 52790
rect 18258 52675 18406 52757
rect 18146 52642 18223 52658
tri 18223 52642 18239 52658 sw
rect 18146 52576 18239 52642
rect 18146 52474 18239 52540
rect 18146 52458 18223 52474
tri 18223 52458 18239 52474 nw
rect 18275 52441 18389 52675
tri 18425 52642 18441 52658 se
rect 18441 52642 18518 52658
rect 18425 52576 18518 52642
rect 18425 52474 18518 52540
tri 18425 52458 18441 52474 ne
rect 18441 52458 18518 52474
rect 18258 52359 18406 52441
rect 18146 52326 18223 52342
tri 18223 52326 18239 52342 sw
rect 18146 52260 18239 52326
rect 18275 52201 18389 52359
tri 18425 52326 18441 52342 se
rect 18441 52326 18518 52342
rect 18425 52260 18518 52326
rect 18146 52125 18518 52201
rect 18146 52000 18239 52066
rect 18146 51984 18223 52000
tri 18223 51984 18239 52000 nw
rect 18275 51967 18389 52125
rect 18425 52000 18518 52066
tri 18425 51984 18441 52000 ne
rect 18441 51984 18518 52000
rect 18258 51885 18406 51967
rect 18146 51852 18223 51868
tri 18223 51852 18239 51868 sw
rect 18146 51786 18239 51852
rect 18146 51684 18239 51750
rect 18146 51668 18223 51684
tri 18223 51668 18239 51684 nw
rect 18275 51651 18389 51885
tri 18425 51852 18441 51868 se
rect 18441 51852 18518 51868
rect 18425 51786 18518 51852
rect 18425 51684 18518 51750
tri 18425 51668 18441 51684 ne
rect 18441 51668 18518 51684
rect 18258 51569 18406 51651
rect 18146 51536 18223 51552
tri 18223 51536 18239 51552 sw
rect 18146 51470 18239 51536
rect 18275 51411 18389 51569
tri 18425 51536 18441 51552 se
rect 18441 51536 18518 51552
rect 18425 51470 18518 51536
rect 18146 51335 18518 51411
rect 18146 51210 18239 51276
rect 18146 51194 18223 51210
tri 18223 51194 18239 51210 nw
rect 18275 51177 18389 51335
rect 18425 51210 18518 51276
tri 18425 51194 18441 51210 ne
rect 18441 51194 18518 51210
rect 18258 51095 18406 51177
rect 18146 51062 18223 51078
tri 18223 51062 18239 51078 sw
rect 18146 50996 18239 51062
rect 18146 50894 18239 50960
rect 18146 50878 18223 50894
tri 18223 50878 18239 50894 nw
rect 18275 50861 18389 51095
tri 18425 51062 18441 51078 se
rect 18441 51062 18518 51078
rect 18425 50996 18518 51062
rect 18425 50894 18518 50960
tri 18425 50878 18441 50894 ne
rect 18441 50878 18518 50894
rect 18258 50779 18406 50861
rect 18146 50746 18223 50762
tri 18223 50746 18239 50762 sw
rect 18146 50680 18239 50746
rect 18275 50621 18389 50779
tri 18425 50746 18441 50762 se
rect 18441 50746 18518 50762
rect 18425 50680 18518 50746
rect 18146 50545 18518 50621
rect 18146 50420 18239 50486
rect 18146 50404 18223 50420
tri 18223 50404 18239 50420 nw
rect 18275 50387 18389 50545
rect 18425 50420 18518 50486
tri 18425 50404 18441 50420 ne
rect 18441 50404 18518 50420
rect 18258 50305 18406 50387
rect 18146 50272 18223 50288
tri 18223 50272 18239 50288 sw
rect 18146 50206 18239 50272
rect 18146 50104 18239 50170
rect 18146 50088 18223 50104
tri 18223 50088 18239 50104 nw
rect 18275 50071 18389 50305
tri 18425 50272 18441 50288 se
rect 18441 50272 18518 50288
rect 18425 50206 18518 50272
rect 18425 50104 18518 50170
tri 18425 50088 18441 50104 ne
rect 18441 50088 18518 50104
rect 18258 49989 18406 50071
rect 18146 49956 18223 49972
tri 18223 49956 18239 49972 sw
rect 18146 49890 18239 49956
rect 18275 49831 18389 49989
tri 18425 49956 18441 49972 se
rect 18441 49956 18518 49972
rect 18425 49890 18518 49956
rect 18146 49755 18518 49831
rect 18146 49630 18239 49696
rect 18146 49614 18223 49630
tri 18223 49614 18239 49630 nw
rect 18275 49597 18389 49755
rect 18425 49630 18518 49696
tri 18425 49614 18441 49630 ne
rect 18441 49614 18518 49630
rect 18258 49515 18406 49597
rect 18146 49482 18223 49498
tri 18223 49482 18239 49498 sw
rect 18146 49416 18239 49482
rect 18146 49314 18239 49380
rect 18146 49298 18223 49314
tri 18223 49298 18239 49314 nw
rect 18275 49281 18389 49515
tri 18425 49482 18441 49498 se
rect 18441 49482 18518 49498
rect 18425 49416 18518 49482
rect 18425 49314 18518 49380
tri 18425 49298 18441 49314 ne
rect 18441 49298 18518 49314
rect 18258 49199 18406 49281
rect 18146 49166 18223 49182
tri 18223 49166 18239 49182 sw
rect 18146 49100 18239 49166
rect 18275 49041 18389 49199
tri 18425 49166 18441 49182 se
rect 18441 49166 18518 49182
rect 18425 49100 18518 49166
rect 18146 48965 18518 49041
rect 18146 48840 18239 48906
rect 18146 48824 18223 48840
tri 18223 48824 18239 48840 nw
rect 18275 48807 18389 48965
rect 18425 48840 18518 48906
tri 18425 48824 18441 48840 ne
rect 18441 48824 18518 48840
rect 18258 48725 18406 48807
rect 18146 48692 18223 48708
tri 18223 48692 18239 48708 sw
rect 18146 48626 18239 48692
rect 18146 48524 18239 48590
rect 18146 48508 18223 48524
tri 18223 48508 18239 48524 nw
rect 18275 48491 18389 48725
tri 18425 48692 18441 48708 se
rect 18441 48692 18518 48708
rect 18425 48626 18518 48692
rect 18425 48524 18518 48590
tri 18425 48508 18441 48524 ne
rect 18441 48508 18518 48524
rect 18258 48409 18406 48491
rect 18146 48376 18223 48392
tri 18223 48376 18239 48392 sw
rect 18146 48310 18239 48376
rect 18275 48251 18389 48409
tri 18425 48376 18441 48392 se
rect 18441 48376 18518 48392
rect 18425 48310 18518 48376
rect 18146 48175 18518 48251
rect 18146 48050 18239 48116
rect 18146 48034 18223 48050
tri 18223 48034 18239 48050 nw
rect 18275 48017 18389 48175
rect 18425 48050 18518 48116
tri 18425 48034 18441 48050 ne
rect 18441 48034 18518 48050
rect 18258 47935 18406 48017
rect 18146 47902 18223 47918
tri 18223 47902 18239 47918 sw
rect 18146 47836 18239 47902
rect 18146 47734 18239 47800
rect 18146 47718 18223 47734
tri 18223 47718 18239 47734 nw
rect 18275 47701 18389 47935
tri 18425 47902 18441 47918 se
rect 18441 47902 18518 47918
rect 18425 47836 18518 47902
rect 18425 47734 18518 47800
tri 18425 47718 18441 47734 ne
rect 18441 47718 18518 47734
rect 18258 47619 18406 47701
rect 18146 47586 18223 47602
tri 18223 47586 18239 47602 sw
rect 18146 47520 18239 47586
rect 18275 47461 18389 47619
tri 18425 47586 18441 47602 se
rect 18441 47586 18518 47602
rect 18425 47520 18518 47586
rect 18146 47385 18518 47461
rect 18146 47260 18239 47326
rect 18146 47244 18223 47260
tri 18223 47244 18239 47260 nw
rect 18275 47227 18389 47385
rect 18425 47260 18518 47326
tri 18425 47244 18441 47260 ne
rect 18441 47244 18518 47260
rect 18258 47145 18406 47227
rect 18146 47112 18223 47128
tri 18223 47112 18239 47128 sw
rect 18146 47046 18239 47112
rect 18146 46944 18239 47010
rect 18146 46928 18223 46944
tri 18223 46928 18239 46944 nw
rect 18275 46911 18389 47145
tri 18425 47112 18441 47128 se
rect 18441 47112 18518 47128
rect 18425 47046 18518 47112
rect 18425 46944 18518 47010
tri 18425 46928 18441 46944 ne
rect 18441 46928 18518 46944
rect 18258 46829 18406 46911
rect 18146 46796 18223 46812
tri 18223 46796 18239 46812 sw
rect 18146 46730 18239 46796
rect 18275 46671 18389 46829
tri 18425 46796 18441 46812 se
rect 18441 46796 18518 46812
rect 18425 46730 18518 46796
rect 18146 46595 18518 46671
rect 18146 46470 18239 46536
rect 18146 46454 18223 46470
tri 18223 46454 18239 46470 nw
rect 18275 46437 18389 46595
rect 18425 46470 18518 46536
tri 18425 46454 18441 46470 ne
rect 18441 46454 18518 46470
rect 18258 46355 18406 46437
rect 18146 46322 18223 46338
tri 18223 46322 18239 46338 sw
rect 18146 46256 18239 46322
rect 18146 46154 18239 46220
rect 18146 46138 18223 46154
tri 18223 46138 18239 46154 nw
rect 18275 46121 18389 46355
tri 18425 46322 18441 46338 se
rect 18441 46322 18518 46338
rect 18425 46256 18518 46322
rect 18425 46154 18518 46220
tri 18425 46138 18441 46154 ne
rect 18441 46138 18518 46154
rect 18258 46039 18406 46121
rect 18146 46006 18223 46022
tri 18223 46006 18239 46022 sw
rect 18146 45940 18239 46006
rect 18275 45881 18389 46039
tri 18425 46006 18441 46022 se
rect 18441 46006 18518 46022
rect 18425 45940 18518 46006
rect 18146 45805 18518 45881
rect 18146 45680 18239 45746
rect 18146 45664 18223 45680
tri 18223 45664 18239 45680 nw
rect 18275 45647 18389 45805
rect 18425 45680 18518 45746
tri 18425 45664 18441 45680 ne
rect 18441 45664 18518 45680
rect 18258 45565 18406 45647
rect 18146 45532 18223 45548
tri 18223 45532 18239 45548 sw
rect 18146 45466 18239 45532
rect 18146 45364 18239 45430
rect 18146 45348 18223 45364
tri 18223 45348 18239 45364 nw
rect 18275 45331 18389 45565
tri 18425 45532 18441 45548 se
rect 18441 45532 18518 45548
rect 18425 45466 18518 45532
rect 18425 45364 18518 45430
tri 18425 45348 18441 45364 ne
rect 18441 45348 18518 45364
rect 18258 45249 18406 45331
rect 18146 45216 18223 45232
tri 18223 45216 18239 45232 sw
rect 18146 45150 18239 45216
rect 18275 45091 18389 45249
tri 18425 45216 18441 45232 se
rect 18441 45216 18518 45232
rect 18425 45150 18518 45216
rect 18146 45015 18518 45091
rect 18146 44890 18239 44956
rect 18146 44874 18223 44890
tri 18223 44874 18239 44890 nw
rect 18275 44857 18389 45015
rect 18425 44890 18518 44956
tri 18425 44874 18441 44890 ne
rect 18441 44874 18518 44890
rect 18258 44775 18406 44857
rect 18146 44742 18223 44758
tri 18223 44742 18239 44758 sw
rect 18146 44676 18239 44742
rect 18146 44574 18239 44640
rect 18146 44558 18223 44574
tri 18223 44558 18239 44574 nw
rect 18275 44541 18389 44775
tri 18425 44742 18441 44758 se
rect 18441 44742 18518 44758
rect 18425 44676 18518 44742
rect 18425 44574 18518 44640
tri 18425 44558 18441 44574 ne
rect 18441 44558 18518 44574
rect 18258 44459 18406 44541
rect 18146 44426 18223 44442
tri 18223 44426 18239 44442 sw
rect 18146 44360 18239 44426
rect 18275 44301 18389 44459
tri 18425 44426 18441 44442 se
rect 18441 44426 18518 44442
rect 18425 44360 18518 44426
rect 18146 44225 18518 44301
rect 18146 44100 18239 44166
rect 18146 44084 18223 44100
tri 18223 44084 18239 44100 nw
rect 18275 44067 18389 44225
rect 18425 44100 18518 44166
tri 18425 44084 18441 44100 ne
rect 18441 44084 18518 44100
rect 18258 43985 18406 44067
rect 18146 43952 18223 43968
tri 18223 43952 18239 43968 sw
rect 18146 43886 18239 43952
rect 18146 43784 18239 43850
rect 18146 43768 18223 43784
tri 18223 43768 18239 43784 nw
rect 18275 43751 18389 43985
tri 18425 43952 18441 43968 se
rect 18441 43952 18518 43968
rect 18425 43886 18518 43952
rect 18425 43784 18518 43850
tri 18425 43768 18441 43784 ne
rect 18441 43768 18518 43784
rect 18258 43669 18406 43751
rect 18146 43636 18223 43652
tri 18223 43636 18239 43652 sw
rect 18146 43570 18239 43636
rect 18275 43511 18389 43669
tri 18425 43636 18441 43652 se
rect 18441 43636 18518 43652
rect 18425 43570 18518 43636
rect 18146 43435 18518 43511
rect 18146 43310 18239 43376
rect 18146 43294 18223 43310
tri 18223 43294 18239 43310 nw
rect 18275 43277 18389 43435
rect 18425 43310 18518 43376
tri 18425 43294 18441 43310 ne
rect 18441 43294 18518 43310
rect 18258 43195 18406 43277
rect 18146 43162 18223 43178
tri 18223 43162 18239 43178 sw
rect 18146 43096 18239 43162
rect 18146 42994 18239 43060
rect 18146 42978 18223 42994
tri 18223 42978 18239 42994 nw
rect 18275 42961 18389 43195
tri 18425 43162 18441 43178 se
rect 18441 43162 18518 43178
rect 18425 43096 18518 43162
rect 18425 42994 18518 43060
tri 18425 42978 18441 42994 ne
rect 18441 42978 18518 42994
rect 18258 42879 18406 42961
rect 18146 42846 18223 42862
tri 18223 42846 18239 42862 sw
rect 18146 42780 18239 42846
rect 18275 42721 18389 42879
tri 18425 42846 18441 42862 se
rect 18441 42846 18518 42862
rect 18425 42780 18518 42846
rect 18146 42645 18518 42721
rect 18146 42520 18239 42586
rect 18146 42504 18223 42520
tri 18223 42504 18239 42520 nw
rect 18275 42487 18389 42645
rect 18425 42520 18518 42586
tri 18425 42504 18441 42520 ne
rect 18441 42504 18518 42520
rect 18258 42405 18406 42487
rect 18146 42372 18223 42388
tri 18223 42372 18239 42388 sw
rect 18146 42306 18239 42372
rect 18146 42204 18239 42270
rect 18146 42188 18223 42204
tri 18223 42188 18239 42204 nw
rect 18275 42171 18389 42405
tri 18425 42372 18441 42388 se
rect 18441 42372 18518 42388
rect 18425 42306 18518 42372
rect 18425 42204 18518 42270
tri 18425 42188 18441 42204 ne
rect 18441 42188 18518 42204
rect 18258 42089 18406 42171
rect 18146 42056 18223 42072
tri 18223 42056 18239 42072 sw
rect 18146 41990 18239 42056
rect 18275 41931 18389 42089
tri 18425 42056 18441 42072 se
rect 18441 42056 18518 42072
rect 18425 41990 18518 42056
rect 18146 41855 18518 41931
rect 18146 41730 18239 41796
rect 18146 41714 18223 41730
tri 18223 41714 18239 41730 nw
rect 18275 41697 18389 41855
rect 18425 41730 18518 41796
tri 18425 41714 18441 41730 ne
rect 18441 41714 18518 41730
rect 18258 41615 18406 41697
rect 18146 41582 18223 41598
tri 18223 41582 18239 41598 sw
rect 18146 41516 18239 41582
rect 18146 41414 18239 41480
rect 18146 41398 18223 41414
tri 18223 41398 18239 41414 nw
rect 18275 41381 18389 41615
tri 18425 41582 18441 41598 se
rect 18441 41582 18518 41598
rect 18425 41516 18518 41582
rect 18425 41414 18518 41480
tri 18425 41398 18441 41414 ne
rect 18441 41398 18518 41414
rect 18258 41299 18406 41381
rect 18146 41266 18223 41282
tri 18223 41266 18239 41282 sw
rect 18146 41200 18239 41266
rect 18275 41141 18389 41299
tri 18425 41266 18441 41282 se
rect 18441 41266 18518 41282
rect 18425 41200 18518 41266
rect 18146 41065 18518 41141
rect 18146 40940 18239 41006
rect 18146 40924 18223 40940
tri 18223 40924 18239 40940 nw
rect 18275 40907 18389 41065
rect 18425 40940 18518 41006
tri 18425 40924 18441 40940 ne
rect 18441 40924 18518 40940
rect 18258 40825 18406 40907
rect 18146 40792 18223 40808
tri 18223 40792 18239 40808 sw
rect 18146 40726 18239 40792
rect 18146 40624 18239 40690
rect 18146 40608 18223 40624
tri 18223 40608 18239 40624 nw
rect 18275 40591 18389 40825
tri 18425 40792 18441 40808 se
rect 18441 40792 18518 40808
rect 18425 40726 18518 40792
rect 18425 40624 18518 40690
tri 18425 40608 18441 40624 ne
rect 18441 40608 18518 40624
rect 18258 40509 18406 40591
rect 18146 40476 18223 40492
tri 18223 40476 18239 40492 sw
rect 18146 40410 18239 40476
rect 18275 40351 18389 40509
tri 18425 40476 18441 40492 se
rect 18441 40476 18518 40492
rect 18425 40410 18518 40476
rect 18146 40275 18518 40351
rect 18146 40150 18239 40216
rect 18146 40134 18223 40150
tri 18223 40134 18239 40150 nw
rect 18275 40117 18389 40275
rect 18425 40150 18518 40216
tri 18425 40134 18441 40150 ne
rect 18441 40134 18518 40150
rect 18258 40035 18406 40117
rect 18146 40002 18223 40018
tri 18223 40002 18239 40018 sw
rect 18146 39936 18239 40002
rect 18146 39834 18239 39900
rect 18146 39818 18223 39834
tri 18223 39818 18239 39834 nw
rect 18275 39801 18389 40035
tri 18425 40002 18441 40018 se
rect 18441 40002 18518 40018
rect 18425 39936 18518 40002
rect 18425 39834 18518 39900
tri 18425 39818 18441 39834 ne
rect 18441 39818 18518 39834
rect 18258 39719 18406 39801
rect 18146 39686 18223 39702
tri 18223 39686 18239 39702 sw
rect 18146 39620 18239 39686
rect 18275 39561 18389 39719
tri 18425 39686 18441 39702 se
rect 18441 39686 18518 39702
rect 18425 39620 18518 39686
rect 18146 39485 18518 39561
rect 18146 39360 18239 39426
rect 18146 39344 18223 39360
tri 18223 39344 18239 39360 nw
rect 18275 39327 18389 39485
rect 18425 39360 18518 39426
tri 18425 39344 18441 39360 ne
rect 18441 39344 18518 39360
rect 18258 39245 18406 39327
rect 18146 39212 18223 39228
tri 18223 39212 18239 39228 sw
rect 18146 39146 18239 39212
rect 18146 39044 18239 39110
rect 18146 39028 18223 39044
tri 18223 39028 18239 39044 nw
rect 18275 39011 18389 39245
tri 18425 39212 18441 39228 se
rect 18441 39212 18518 39228
rect 18425 39146 18518 39212
rect 18425 39044 18518 39110
tri 18425 39028 18441 39044 ne
rect 18441 39028 18518 39044
rect 18258 38929 18406 39011
rect 18146 38896 18223 38912
tri 18223 38896 18239 38912 sw
rect 18146 38830 18239 38896
rect 18275 38771 18389 38929
tri 18425 38896 18441 38912 se
rect 18441 38896 18518 38912
rect 18425 38830 18518 38896
rect 18146 38695 18518 38771
rect 18146 38570 18239 38636
rect 18146 38554 18223 38570
tri 18223 38554 18239 38570 nw
rect 18275 38537 18389 38695
rect 18425 38570 18518 38636
tri 18425 38554 18441 38570 ne
rect 18441 38554 18518 38570
rect 18258 38455 18406 38537
rect 18146 38422 18223 38438
tri 18223 38422 18239 38438 sw
rect 18146 38356 18239 38422
rect 18146 38254 18239 38320
rect 18146 38238 18223 38254
tri 18223 38238 18239 38254 nw
rect 18275 38221 18389 38455
tri 18425 38422 18441 38438 se
rect 18441 38422 18518 38438
rect 18425 38356 18518 38422
rect 18425 38254 18518 38320
tri 18425 38238 18441 38254 ne
rect 18441 38238 18518 38254
rect 18258 38139 18406 38221
rect 18146 38106 18223 38122
tri 18223 38106 18239 38122 sw
rect 18146 38040 18239 38106
rect 18275 37981 18389 38139
tri 18425 38106 18441 38122 se
rect 18441 38106 18518 38122
rect 18425 38040 18518 38106
rect 18146 37905 18518 37981
rect 18146 37780 18239 37846
rect 18146 37764 18223 37780
tri 18223 37764 18239 37780 nw
rect 18275 37747 18389 37905
rect 18425 37780 18518 37846
tri 18425 37764 18441 37780 ne
rect 18441 37764 18518 37780
rect 18258 37665 18406 37747
rect 18146 37632 18223 37648
tri 18223 37632 18239 37648 sw
rect 18146 37566 18239 37632
rect 18146 37464 18239 37530
rect 18146 37448 18223 37464
tri 18223 37448 18239 37464 nw
rect 18275 37431 18389 37665
tri 18425 37632 18441 37648 se
rect 18441 37632 18518 37648
rect 18425 37566 18518 37632
rect 18425 37464 18518 37530
tri 18425 37448 18441 37464 ne
rect 18441 37448 18518 37464
rect 18258 37349 18406 37431
rect 18146 37316 18223 37332
tri 18223 37316 18239 37332 sw
rect 18146 37250 18239 37316
rect 18275 37191 18389 37349
tri 18425 37316 18441 37332 se
rect 18441 37316 18518 37332
rect 18425 37250 18518 37316
rect 18146 37115 18518 37191
rect 18146 36990 18239 37056
rect 18146 36974 18223 36990
tri 18223 36974 18239 36990 nw
rect 18275 36957 18389 37115
rect 18425 36990 18518 37056
tri 18425 36974 18441 36990 ne
rect 18441 36974 18518 36990
rect 18258 36875 18406 36957
rect 18146 36842 18223 36858
tri 18223 36842 18239 36858 sw
rect 18146 36776 18239 36842
rect 18146 36674 18239 36740
rect 18146 36658 18223 36674
tri 18223 36658 18239 36674 nw
rect 18275 36641 18389 36875
tri 18425 36842 18441 36858 se
rect 18441 36842 18518 36858
rect 18425 36776 18518 36842
rect 18425 36674 18518 36740
tri 18425 36658 18441 36674 ne
rect 18441 36658 18518 36674
rect 18258 36559 18406 36641
rect 18146 36526 18223 36542
tri 18223 36526 18239 36542 sw
rect 18146 36460 18239 36526
rect 18275 36401 18389 36559
tri 18425 36526 18441 36542 se
rect 18441 36526 18518 36542
rect 18425 36460 18518 36526
rect 18146 36325 18518 36401
rect 18146 36200 18239 36266
rect 18146 36184 18223 36200
tri 18223 36184 18239 36200 nw
rect 18275 36167 18389 36325
rect 18425 36200 18518 36266
tri 18425 36184 18441 36200 ne
rect 18441 36184 18518 36200
rect 18258 36085 18406 36167
rect 18146 36052 18223 36068
tri 18223 36052 18239 36068 sw
rect 18146 35986 18239 36052
rect 18146 35884 18239 35950
rect 18146 35868 18223 35884
tri 18223 35868 18239 35884 nw
rect 18275 35851 18389 36085
tri 18425 36052 18441 36068 se
rect 18441 36052 18518 36068
rect 18425 35986 18518 36052
rect 18425 35884 18518 35950
tri 18425 35868 18441 35884 ne
rect 18441 35868 18518 35884
rect 18258 35769 18406 35851
rect 18146 35736 18223 35752
tri 18223 35736 18239 35752 sw
rect 18146 35670 18239 35736
rect 18275 35611 18389 35769
tri 18425 35736 18441 35752 se
rect 18441 35736 18518 35752
rect 18425 35670 18518 35736
rect 18146 35535 18518 35611
rect 18146 35410 18239 35476
rect 18146 35394 18223 35410
tri 18223 35394 18239 35410 nw
rect 18275 35377 18389 35535
rect 18425 35410 18518 35476
tri 18425 35394 18441 35410 ne
rect 18441 35394 18518 35410
rect 18258 35295 18406 35377
rect 18146 35262 18223 35278
tri 18223 35262 18239 35278 sw
rect 18146 35196 18239 35262
rect 18146 35094 18239 35160
rect 18146 35078 18223 35094
tri 18223 35078 18239 35094 nw
rect 18275 35061 18389 35295
tri 18425 35262 18441 35278 se
rect 18441 35262 18518 35278
rect 18425 35196 18518 35262
rect 18425 35094 18518 35160
tri 18425 35078 18441 35094 ne
rect 18441 35078 18518 35094
rect 18258 34979 18406 35061
rect 18146 34946 18223 34962
tri 18223 34946 18239 34962 sw
rect 18146 34880 18239 34946
rect 18275 34821 18389 34979
tri 18425 34946 18441 34962 se
rect 18441 34946 18518 34962
rect 18425 34880 18518 34946
rect 18146 34745 18518 34821
rect 18146 34620 18239 34686
rect 18146 34604 18223 34620
tri 18223 34604 18239 34620 nw
rect 18275 34587 18389 34745
rect 18425 34620 18518 34686
tri 18425 34604 18441 34620 ne
rect 18441 34604 18518 34620
rect 18258 34505 18406 34587
rect 18146 34472 18223 34488
tri 18223 34472 18239 34488 sw
rect 18146 34406 18239 34472
rect 18146 34304 18239 34370
rect 18146 34288 18223 34304
tri 18223 34288 18239 34304 nw
rect 18275 34271 18389 34505
tri 18425 34472 18441 34488 se
rect 18441 34472 18518 34488
rect 18425 34406 18518 34472
rect 18425 34304 18518 34370
tri 18425 34288 18441 34304 ne
rect 18441 34288 18518 34304
rect 18258 34189 18406 34271
rect 18146 34156 18223 34172
tri 18223 34156 18239 34172 sw
rect 18146 34090 18239 34156
rect 18275 34031 18389 34189
tri 18425 34156 18441 34172 se
rect 18441 34156 18518 34172
rect 18425 34090 18518 34156
rect 18146 33955 18518 34031
rect 18146 33830 18239 33896
rect 18146 33814 18223 33830
tri 18223 33814 18239 33830 nw
rect 18275 33797 18389 33955
rect 18425 33830 18518 33896
tri 18425 33814 18441 33830 ne
rect 18441 33814 18518 33830
rect 18258 33715 18406 33797
rect 18146 33682 18223 33698
tri 18223 33682 18239 33698 sw
rect 18146 33616 18239 33682
rect 18146 33514 18239 33580
rect 18146 33498 18223 33514
tri 18223 33498 18239 33514 nw
rect 18275 33481 18389 33715
tri 18425 33682 18441 33698 se
rect 18441 33682 18518 33698
rect 18425 33616 18518 33682
rect 18425 33514 18518 33580
tri 18425 33498 18441 33514 ne
rect 18441 33498 18518 33514
rect 18258 33399 18406 33481
rect 18146 33366 18223 33382
tri 18223 33366 18239 33382 sw
rect 18146 33300 18239 33366
rect 18275 33241 18389 33399
tri 18425 33366 18441 33382 se
rect 18441 33366 18518 33382
rect 18425 33300 18518 33366
rect 18146 33165 18518 33241
rect 18146 33040 18239 33106
rect 18146 33024 18223 33040
tri 18223 33024 18239 33040 nw
rect 18275 33007 18389 33165
rect 18425 33040 18518 33106
tri 18425 33024 18441 33040 ne
rect 18441 33024 18518 33040
rect 18258 32925 18406 33007
rect 18146 32892 18223 32908
tri 18223 32892 18239 32908 sw
rect 18146 32826 18239 32892
rect 18146 32724 18239 32790
rect 18146 32708 18223 32724
tri 18223 32708 18239 32724 nw
rect 18275 32691 18389 32925
tri 18425 32892 18441 32908 se
rect 18441 32892 18518 32908
rect 18425 32826 18518 32892
rect 18425 32724 18518 32790
tri 18425 32708 18441 32724 ne
rect 18441 32708 18518 32724
rect 18258 32609 18406 32691
rect 18146 32576 18223 32592
tri 18223 32576 18239 32592 sw
rect 18146 32510 18239 32576
rect 18275 32451 18389 32609
tri 18425 32576 18441 32592 se
rect 18441 32576 18518 32592
rect 18425 32510 18518 32576
rect 18146 32375 18518 32451
rect 18146 32250 18239 32316
rect 18146 32234 18223 32250
tri 18223 32234 18239 32250 nw
rect 18275 32217 18389 32375
rect 18425 32250 18518 32316
tri 18425 32234 18441 32250 ne
rect 18441 32234 18518 32250
rect 18258 32135 18406 32217
rect 18146 32102 18223 32118
tri 18223 32102 18239 32118 sw
rect 18146 32036 18239 32102
rect 18146 31934 18239 32000
rect 18146 31918 18223 31934
tri 18223 31918 18239 31934 nw
rect 18275 31901 18389 32135
tri 18425 32102 18441 32118 se
rect 18441 32102 18518 32118
rect 18425 32036 18518 32102
rect 18425 31934 18518 32000
tri 18425 31918 18441 31934 ne
rect 18441 31918 18518 31934
rect 18258 31819 18406 31901
rect 18146 31786 18223 31802
tri 18223 31786 18239 31802 sw
rect 18146 31720 18239 31786
rect 18275 31661 18389 31819
tri 18425 31786 18441 31802 se
rect 18441 31786 18518 31802
rect 18425 31720 18518 31786
rect 18146 31585 18518 31661
rect 18146 31460 18239 31526
rect 18146 31444 18223 31460
tri 18223 31444 18239 31460 nw
rect 18275 31427 18389 31585
rect 18425 31460 18518 31526
tri 18425 31444 18441 31460 ne
rect 18441 31444 18518 31460
rect 18258 31345 18406 31427
rect 18146 31312 18223 31328
tri 18223 31312 18239 31328 sw
rect 18146 31246 18239 31312
rect 18146 31144 18239 31210
rect 18146 31128 18223 31144
tri 18223 31128 18239 31144 nw
rect 18275 31111 18389 31345
tri 18425 31312 18441 31328 se
rect 18441 31312 18518 31328
rect 18425 31246 18518 31312
rect 18425 31144 18518 31210
tri 18425 31128 18441 31144 ne
rect 18441 31128 18518 31144
rect 18258 31029 18406 31111
rect 18146 30996 18223 31012
tri 18223 30996 18239 31012 sw
rect 18146 30930 18239 30996
rect 18275 30871 18389 31029
tri 18425 30996 18441 31012 se
rect 18441 30996 18518 31012
rect 18425 30930 18518 30996
rect 18146 30795 18518 30871
rect 18146 30670 18239 30736
rect 18146 30654 18223 30670
tri 18223 30654 18239 30670 nw
rect 18275 30637 18389 30795
rect 18425 30670 18518 30736
tri 18425 30654 18441 30670 ne
rect 18441 30654 18518 30670
rect 18258 30555 18406 30637
rect 18146 30522 18223 30538
tri 18223 30522 18239 30538 sw
rect 18146 30456 18239 30522
rect 18146 30354 18239 30420
rect 18146 30338 18223 30354
tri 18223 30338 18239 30354 nw
rect 18275 30321 18389 30555
tri 18425 30522 18441 30538 se
rect 18441 30522 18518 30538
rect 18425 30456 18518 30522
rect 18425 30354 18518 30420
tri 18425 30338 18441 30354 ne
rect 18441 30338 18518 30354
rect 18258 30239 18406 30321
rect 18146 30206 18223 30222
tri 18223 30206 18239 30222 sw
rect 18146 30140 18239 30206
rect 18275 30081 18389 30239
tri 18425 30206 18441 30222 se
rect 18441 30206 18518 30222
rect 18425 30140 18518 30206
rect 18146 30005 18518 30081
rect 18146 29880 18239 29946
rect 18146 29864 18223 29880
tri 18223 29864 18239 29880 nw
rect 18275 29847 18389 30005
rect 18425 29880 18518 29946
tri 18425 29864 18441 29880 ne
rect 18441 29864 18518 29880
rect 18258 29765 18406 29847
rect 18146 29732 18223 29748
tri 18223 29732 18239 29748 sw
rect 18146 29666 18239 29732
rect 18146 29564 18239 29630
rect 18146 29548 18223 29564
tri 18223 29548 18239 29564 nw
rect 18275 29531 18389 29765
tri 18425 29732 18441 29748 se
rect 18441 29732 18518 29748
rect 18425 29666 18518 29732
rect 18425 29564 18518 29630
tri 18425 29548 18441 29564 ne
rect 18441 29548 18518 29564
rect 18258 29449 18406 29531
rect 18146 29416 18223 29432
tri 18223 29416 18239 29432 sw
rect 18146 29350 18239 29416
rect 18275 29291 18389 29449
tri 18425 29416 18441 29432 se
rect 18441 29416 18518 29432
rect 18425 29350 18518 29416
rect 18146 29215 18518 29291
rect 18146 29090 18239 29156
rect 18146 29074 18223 29090
tri 18223 29074 18239 29090 nw
rect 18275 29057 18389 29215
rect 18425 29090 18518 29156
tri 18425 29074 18441 29090 ne
rect 18441 29074 18518 29090
rect 18258 28975 18406 29057
rect 18146 28942 18223 28958
tri 18223 28942 18239 28958 sw
rect 18146 28876 18239 28942
rect 18275 28833 18389 28975
tri 18425 28942 18441 28958 se
rect 18441 28942 18518 28958
rect 18425 28876 18518 28942
rect 18554 28463 18590 80603
rect 18626 28463 18662 80603
rect 18698 80445 18734 80603
rect 18690 80303 18742 80445
rect 18698 28763 18734 80303
rect 18690 28621 18742 28763
rect 18698 28463 18734 28621
rect 18770 28463 18806 80603
rect 18842 28463 18878 80603
rect 18914 28833 18998 80233
rect 19034 28463 19070 80603
rect 19106 28463 19142 80603
rect 19178 80445 19214 80603
rect 19170 80303 19222 80445
rect 19178 28763 19214 80303
rect 19170 28621 19222 28763
rect 19178 28463 19214 28621
rect 19250 28463 19286 80603
rect 19322 28463 19358 80603
rect 19394 80124 19487 80190
rect 19394 80108 19471 80124
tri 19471 80108 19487 80124 nw
rect 19523 80091 19637 80233
rect 19673 80124 19766 80190
tri 19673 80108 19689 80124 ne
rect 19689 80108 19766 80124
rect 19506 80009 19654 80091
rect 19394 79976 19471 79992
tri 19471 79976 19487 79992 sw
rect 19394 79910 19487 79976
rect 19523 79851 19637 80009
tri 19673 79976 19689 79992 se
rect 19689 79976 19766 79992
rect 19673 79910 19766 79976
rect 19394 79775 19766 79851
rect 19394 79650 19487 79716
rect 19394 79634 19471 79650
tri 19471 79634 19487 79650 nw
rect 19523 79617 19637 79775
rect 19673 79650 19766 79716
tri 19673 79634 19689 79650 ne
rect 19689 79634 19766 79650
rect 19506 79535 19654 79617
rect 19394 79502 19471 79518
tri 19471 79502 19487 79518 sw
rect 19394 79436 19487 79502
rect 19394 79334 19487 79400
rect 19394 79318 19471 79334
tri 19471 79318 19487 79334 nw
rect 19523 79301 19637 79535
tri 19673 79502 19689 79518 se
rect 19689 79502 19766 79518
rect 19673 79436 19766 79502
rect 19673 79334 19766 79400
tri 19673 79318 19689 79334 ne
rect 19689 79318 19766 79334
rect 19506 79219 19654 79301
rect 19394 79186 19471 79202
tri 19471 79186 19487 79202 sw
rect 19394 79120 19487 79186
rect 19523 79061 19637 79219
tri 19673 79186 19689 79202 se
rect 19689 79186 19766 79202
rect 19673 79120 19766 79186
rect 19394 78985 19766 79061
rect 19394 78860 19487 78926
rect 19394 78844 19471 78860
tri 19471 78844 19487 78860 nw
rect 19523 78827 19637 78985
rect 19673 78860 19766 78926
tri 19673 78844 19689 78860 ne
rect 19689 78844 19766 78860
rect 19506 78745 19654 78827
rect 19394 78712 19471 78728
tri 19471 78712 19487 78728 sw
rect 19394 78646 19487 78712
rect 19394 78544 19487 78610
rect 19394 78528 19471 78544
tri 19471 78528 19487 78544 nw
rect 19523 78511 19637 78745
tri 19673 78712 19689 78728 se
rect 19689 78712 19766 78728
rect 19673 78646 19766 78712
rect 19673 78544 19766 78610
tri 19673 78528 19689 78544 ne
rect 19689 78528 19766 78544
rect 19506 78429 19654 78511
rect 19394 78396 19471 78412
tri 19471 78396 19487 78412 sw
rect 19394 78330 19487 78396
rect 19523 78271 19637 78429
tri 19673 78396 19689 78412 se
rect 19689 78396 19766 78412
rect 19673 78330 19766 78396
rect 19394 78195 19766 78271
rect 19394 78070 19487 78136
rect 19394 78054 19471 78070
tri 19471 78054 19487 78070 nw
rect 19523 78037 19637 78195
rect 19673 78070 19766 78136
tri 19673 78054 19689 78070 ne
rect 19689 78054 19766 78070
rect 19506 77955 19654 78037
rect 19394 77922 19471 77938
tri 19471 77922 19487 77938 sw
rect 19394 77856 19487 77922
rect 19394 77754 19487 77820
rect 19394 77738 19471 77754
tri 19471 77738 19487 77754 nw
rect 19523 77721 19637 77955
tri 19673 77922 19689 77938 se
rect 19689 77922 19766 77938
rect 19673 77856 19766 77922
rect 19673 77754 19766 77820
tri 19673 77738 19689 77754 ne
rect 19689 77738 19766 77754
rect 19506 77639 19654 77721
rect 19394 77606 19471 77622
tri 19471 77606 19487 77622 sw
rect 19394 77540 19487 77606
rect 19523 77481 19637 77639
tri 19673 77606 19689 77622 se
rect 19689 77606 19766 77622
rect 19673 77540 19766 77606
rect 19394 77405 19766 77481
rect 19394 77280 19487 77346
rect 19394 77264 19471 77280
tri 19471 77264 19487 77280 nw
rect 19523 77247 19637 77405
rect 19673 77280 19766 77346
tri 19673 77264 19689 77280 ne
rect 19689 77264 19766 77280
rect 19506 77165 19654 77247
rect 19394 77132 19471 77148
tri 19471 77132 19487 77148 sw
rect 19394 77066 19487 77132
rect 19394 76964 19487 77030
rect 19394 76948 19471 76964
tri 19471 76948 19487 76964 nw
rect 19523 76931 19637 77165
tri 19673 77132 19689 77148 se
rect 19689 77132 19766 77148
rect 19673 77066 19766 77132
rect 19673 76964 19766 77030
tri 19673 76948 19689 76964 ne
rect 19689 76948 19766 76964
rect 19506 76849 19654 76931
rect 19394 76816 19471 76832
tri 19471 76816 19487 76832 sw
rect 19394 76750 19487 76816
rect 19523 76691 19637 76849
tri 19673 76816 19689 76832 se
rect 19689 76816 19766 76832
rect 19673 76750 19766 76816
rect 19394 76615 19766 76691
rect 19394 76490 19487 76556
rect 19394 76474 19471 76490
tri 19471 76474 19487 76490 nw
rect 19523 76457 19637 76615
rect 19673 76490 19766 76556
tri 19673 76474 19689 76490 ne
rect 19689 76474 19766 76490
rect 19506 76375 19654 76457
rect 19394 76342 19471 76358
tri 19471 76342 19487 76358 sw
rect 19394 76276 19487 76342
rect 19394 76174 19487 76240
rect 19394 76158 19471 76174
tri 19471 76158 19487 76174 nw
rect 19523 76141 19637 76375
tri 19673 76342 19689 76358 se
rect 19689 76342 19766 76358
rect 19673 76276 19766 76342
rect 19673 76174 19766 76240
tri 19673 76158 19689 76174 ne
rect 19689 76158 19766 76174
rect 19506 76059 19654 76141
rect 19394 76026 19471 76042
tri 19471 76026 19487 76042 sw
rect 19394 75960 19487 76026
rect 19523 75901 19637 76059
tri 19673 76026 19689 76042 se
rect 19689 76026 19766 76042
rect 19673 75960 19766 76026
rect 19394 75825 19766 75901
rect 19394 75700 19487 75766
rect 19394 75684 19471 75700
tri 19471 75684 19487 75700 nw
rect 19523 75667 19637 75825
rect 19673 75700 19766 75766
tri 19673 75684 19689 75700 ne
rect 19689 75684 19766 75700
rect 19506 75585 19654 75667
rect 19394 75552 19471 75568
tri 19471 75552 19487 75568 sw
rect 19394 75486 19487 75552
rect 19394 75384 19487 75450
rect 19394 75368 19471 75384
tri 19471 75368 19487 75384 nw
rect 19523 75351 19637 75585
tri 19673 75552 19689 75568 se
rect 19689 75552 19766 75568
rect 19673 75486 19766 75552
rect 19673 75384 19766 75450
tri 19673 75368 19689 75384 ne
rect 19689 75368 19766 75384
rect 19506 75269 19654 75351
rect 19394 75236 19471 75252
tri 19471 75236 19487 75252 sw
rect 19394 75170 19487 75236
rect 19523 75111 19637 75269
tri 19673 75236 19689 75252 se
rect 19689 75236 19766 75252
rect 19673 75170 19766 75236
rect 19394 75035 19766 75111
rect 19394 74910 19487 74976
rect 19394 74894 19471 74910
tri 19471 74894 19487 74910 nw
rect 19523 74877 19637 75035
rect 19673 74910 19766 74976
tri 19673 74894 19689 74910 ne
rect 19689 74894 19766 74910
rect 19506 74795 19654 74877
rect 19394 74762 19471 74778
tri 19471 74762 19487 74778 sw
rect 19394 74696 19487 74762
rect 19394 74594 19487 74660
rect 19394 74578 19471 74594
tri 19471 74578 19487 74594 nw
rect 19523 74561 19637 74795
tri 19673 74762 19689 74778 se
rect 19689 74762 19766 74778
rect 19673 74696 19766 74762
rect 19673 74594 19766 74660
tri 19673 74578 19689 74594 ne
rect 19689 74578 19766 74594
rect 19506 74479 19654 74561
rect 19394 74446 19471 74462
tri 19471 74446 19487 74462 sw
rect 19394 74380 19487 74446
rect 19523 74321 19637 74479
tri 19673 74446 19689 74462 se
rect 19689 74446 19766 74462
rect 19673 74380 19766 74446
rect 19394 74245 19766 74321
rect 19394 74120 19487 74186
rect 19394 74104 19471 74120
tri 19471 74104 19487 74120 nw
rect 19523 74087 19637 74245
rect 19673 74120 19766 74186
tri 19673 74104 19689 74120 ne
rect 19689 74104 19766 74120
rect 19506 74005 19654 74087
rect 19394 73972 19471 73988
tri 19471 73972 19487 73988 sw
rect 19394 73906 19487 73972
rect 19394 73804 19487 73870
rect 19394 73788 19471 73804
tri 19471 73788 19487 73804 nw
rect 19523 73771 19637 74005
tri 19673 73972 19689 73988 se
rect 19689 73972 19766 73988
rect 19673 73906 19766 73972
rect 19673 73804 19766 73870
tri 19673 73788 19689 73804 ne
rect 19689 73788 19766 73804
rect 19506 73689 19654 73771
rect 19394 73656 19471 73672
tri 19471 73656 19487 73672 sw
rect 19394 73590 19487 73656
rect 19523 73531 19637 73689
tri 19673 73656 19689 73672 se
rect 19689 73656 19766 73672
rect 19673 73590 19766 73656
rect 19394 73455 19766 73531
rect 19394 73330 19487 73396
rect 19394 73314 19471 73330
tri 19471 73314 19487 73330 nw
rect 19523 73297 19637 73455
rect 19673 73330 19766 73396
tri 19673 73314 19689 73330 ne
rect 19689 73314 19766 73330
rect 19506 73215 19654 73297
rect 19394 73182 19471 73198
tri 19471 73182 19487 73198 sw
rect 19394 73116 19487 73182
rect 19394 73014 19487 73080
rect 19394 72998 19471 73014
tri 19471 72998 19487 73014 nw
rect 19523 72981 19637 73215
tri 19673 73182 19689 73198 se
rect 19689 73182 19766 73198
rect 19673 73116 19766 73182
rect 19673 73014 19766 73080
tri 19673 72998 19689 73014 ne
rect 19689 72998 19766 73014
rect 19506 72899 19654 72981
rect 19394 72866 19471 72882
tri 19471 72866 19487 72882 sw
rect 19394 72800 19487 72866
rect 19523 72741 19637 72899
tri 19673 72866 19689 72882 se
rect 19689 72866 19766 72882
rect 19673 72800 19766 72866
rect 19394 72665 19766 72741
rect 19394 72540 19487 72606
rect 19394 72524 19471 72540
tri 19471 72524 19487 72540 nw
rect 19523 72507 19637 72665
rect 19673 72540 19766 72606
tri 19673 72524 19689 72540 ne
rect 19689 72524 19766 72540
rect 19506 72425 19654 72507
rect 19394 72392 19471 72408
tri 19471 72392 19487 72408 sw
rect 19394 72326 19487 72392
rect 19394 72224 19487 72290
rect 19394 72208 19471 72224
tri 19471 72208 19487 72224 nw
rect 19523 72191 19637 72425
tri 19673 72392 19689 72408 se
rect 19689 72392 19766 72408
rect 19673 72326 19766 72392
rect 19673 72224 19766 72290
tri 19673 72208 19689 72224 ne
rect 19689 72208 19766 72224
rect 19506 72109 19654 72191
rect 19394 72076 19471 72092
tri 19471 72076 19487 72092 sw
rect 19394 72010 19487 72076
rect 19523 71951 19637 72109
tri 19673 72076 19689 72092 se
rect 19689 72076 19766 72092
rect 19673 72010 19766 72076
rect 19394 71875 19766 71951
rect 19394 71750 19487 71816
rect 19394 71734 19471 71750
tri 19471 71734 19487 71750 nw
rect 19523 71717 19637 71875
rect 19673 71750 19766 71816
tri 19673 71734 19689 71750 ne
rect 19689 71734 19766 71750
rect 19506 71635 19654 71717
rect 19394 71602 19471 71618
tri 19471 71602 19487 71618 sw
rect 19394 71536 19487 71602
rect 19394 71434 19487 71500
rect 19394 71418 19471 71434
tri 19471 71418 19487 71434 nw
rect 19523 71401 19637 71635
tri 19673 71602 19689 71618 se
rect 19689 71602 19766 71618
rect 19673 71536 19766 71602
rect 19673 71434 19766 71500
tri 19673 71418 19689 71434 ne
rect 19689 71418 19766 71434
rect 19506 71319 19654 71401
rect 19394 71286 19471 71302
tri 19471 71286 19487 71302 sw
rect 19394 71220 19487 71286
rect 19523 71161 19637 71319
tri 19673 71286 19689 71302 se
rect 19689 71286 19766 71302
rect 19673 71220 19766 71286
rect 19394 71085 19766 71161
rect 19394 70960 19487 71026
rect 19394 70944 19471 70960
tri 19471 70944 19487 70960 nw
rect 19523 70927 19637 71085
rect 19673 70960 19766 71026
tri 19673 70944 19689 70960 ne
rect 19689 70944 19766 70960
rect 19506 70845 19654 70927
rect 19394 70812 19471 70828
tri 19471 70812 19487 70828 sw
rect 19394 70746 19487 70812
rect 19394 70644 19487 70710
rect 19394 70628 19471 70644
tri 19471 70628 19487 70644 nw
rect 19523 70611 19637 70845
tri 19673 70812 19689 70828 se
rect 19689 70812 19766 70828
rect 19673 70746 19766 70812
rect 19673 70644 19766 70710
tri 19673 70628 19689 70644 ne
rect 19689 70628 19766 70644
rect 19506 70529 19654 70611
rect 19394 70496 19471 70512
tri 19471 70496 19487 70512 sw
rect 19394 70430 19487 70496
rect 19523 70371 19637 70529
tri 19673 70496 19689 70512 se
rect 19689 70496 19766 70512
rect 19673 70430 19766 70496
rect 19394 70295 19766 70371
rect 19394 70170 19487 70236
rect 19394 70154 19471 70170
tri 19471 70154 19487 70170 nw
rect 19523 70137 19637 70295
rect 19673 70170 19766 70236
tri 19673 70154 19689 70170 ne
rect 19689 70154 19766 70170
rect 19506 70055 19654 70137
rect 19394 70022 19471 70038
tri 19471 70022 19487 70038 sw
rect 19394 69956 19487 70022
rect 19394 69854 19487 69920
rect 19394 69838 19471 69854
tri 19471 69838 19487 69854 nw
rect 19523 69821 19637 70055
tri 19673 70022 19689 70038 se
rect 19689 70022 19766 70038
rect 19673 69956 19766 70022
rect 19673 69854 19766 69920
tri 19673 69838 19689 69854 ne
rect 19689 69838 19766 69854
rect 19506 69739 19654 69821
rect 19394 69706 19471 69722
tri 19471 69706 19487 69722 sw
rect 19394 69640 19487 69706
rect 19523 69581 19637 69739
tri 19673 69706 19689 69722 se
rect 19689 69706 19766 69722
rect 19673 69640 19766 69706
rect 19394 69505 19766 69581
rect 19394 69380 19487 69446
rect 19394 69364 19471 69380
tri 19471 69364 19487 69380 nw
rect 19523 69347 19637 69505
rect 19673 69380 19766 69446
tri 19673 69364 19689 69380 ne
rect 19689 69364 19766 69380
rect 19506 69265 19654 69347
rect 19394 69232 19471 69248
tri 19471 69232 19487 69248 sw
rect 19394 69166 19487 69232
rect 19394 69064 19487 69130
rect 19394 69048 19471 69064
tri 19471 69048 19487 69064 nw
rect 19523 69031 19637 69265
tri 19673 69232 19689 69248 se
rect 19689 69232 19766 69248
rect 19673 69166 19766 69232
rect 19673 69064 19766 69130
tri 19673 69048 19689 69064 ne
rect 19689 69048 19766 69064
rect 19506 68949 19654 69031
rect 19394 68916 19471 68932
tri 19471 68916 19487 68932 sw
rect 19394 68850 19487 68916
rect 19523 68791 19637 68949
tri 19673 68916 19689 68932 se
rect 19689 68916 19766 68932
rect 19673 68850 19766 68916
rect 19394 68715 19766 68791
rect 19394 68590 19487 68656
rect 19394 68574 19471 68590
tri 19471 68574 19487 68590 nw
rect 19523 68557 19637 68715
rect 19673 68590 19766 68656
tri 19673 68574 19689 68590 ne
rect 19689 68574 19766 68590
rect 19506 68475 19654 68557
rect 19394 68442 19471 68458
tri 19471 68442 19487 68458 sw
rect 19394 68376 19487 68442
rect 19394 68274 19487 68340
rect 19394 68258 19471 68274
tri 19471 68258 19487 68274 nw
rect 19523 68241 19637 68475
tri 19673 68442 19689 68458 se
rect 19689 68442 19766 68458
rect 19673 68376 19766 68442
rect 19673 68274 19766 68340
tri 19673 68258 19689 68274 ne
rect 19689 68258 19766 68274
rect 19506 68159 19654 68241
rect 19394 68126 19471 68142
tri 19471 68126 19487 68142 sw
rect 19394 68060 19487 68126
rect 19523 68001 19637 68159
tri 19673 68126 19689 68142 se
rect 19689 68126 19766 68142
rect 19673 68060 19766 68126
rect 19394 67925 19766 68001
rect 19394 67800 19487 67866
rect 19394 67784 19471 67800
tri 19471 67784 19487 67800 nw
rect 19523 67767 19637 67925
rect 19673 67800 19766 67866
tri 19673 67784 19689 67800 ne
rect 19689 67784 19766 67800
rect 19506 67685 19654 67767
rect 19394 67652 19471 67668
tri 19471 67652 19487 67668 sw
rect 19394 67586 19487 67652
rect 19394 67484 19487 67550
rect 19394 67468 19471 67484
tri 19471 67468 19487 67484 nw
rect 19523 67451 19637 67685
tri 19673 67652 19689 67668 se
rect 19689 67652 19766 67668
rect 19673 67586 19766 67652
rect 19673 67484 19766 67550
tri 19673 67468 19689 67484 ne
rect 19689 67468 19766 67484
rect 19506 67369 19654 67451
rect 19394 67336 19471 67352
tri 19471 67336 19487 67352 sw
rect 19394 67270 19487 67336
rect 19523 67211 19637 67369
tri 19673 67336 19689 67352 se
rect 19689 67336 19766 67352
rect 19673 67270 19766 67336
rect 19394 67135 19766 67211
rect 19394 67010 19487 67076
rect 19394 66994 19471 67010
tri 19471 66994 19487 67010 nw
rect 19523 66977 19637 67135
rect 19673 67010 19766 67076
tri 19673 66994 19689 67010 ne
rect 19689 66994 19766 67010
rect 19506 66895 19654 66977
rect 19394 66862 19471 66878
tri 19471 66862 19487 66878 sw
rect 19394 66796 19487 66862
rect 19394 66694 19487 66760
rect 19394 66678 19471 66694
tri 19471 66678 19487 66694 nw
rect 19523 66661 19637 66895
tri 19673 66862 19689 66878 se
rect 19689 66862 19766 66878
rect 19673 66796 19766 66862
rect 19673 66694 19766 66760
tri 19673 66678 19689 66694 ne
rect 19689 66678 19766 66694
rect 19506 66579 19654 66661
rect 19394 66546 19471 66562
tri 19471 66546 19487 66562 sw
rect 19394 66480 19487 66546
rect 19523 66421 19637 66579
tri 19673 66546 19689 66562 se
rect 19689 66546 19766 66562
rect 19673 66480 19766 66546
rect 19394 66345 19766 66421
rect 19394 66220 19487 66286
rect 19394 66204 19471 66220
tri 19471 66204 19487 66220 nw
rect 19523 66187 19637 66345
rect 19673 66220 19766 66286
tri 19673 66204 19689 66220 ne
rect 19689 66204 19766 66220
rect 19506 66105 19654 66187
rect 19394 66072 19471 66088
tri 19471 66072 19487 66088 sw
rect 19394 66006 19487 66072
rect 19394 65904 19487 65970
rect 19394 65888 19471 65904
tri 19471 65888 19487 65904 nw
rect 19523 65871 19637 66105
tri 19673 66072 19689 66088 se
rect 19689 66072 19766 66088
rect 19673 66006 19766 66072
rect 19673 65904 19766 65970
tri 19673 65888 19689 65904 ne
rect 19689 65888 19766 65904
rect 19506 65789 19654 65871
rect 19394 65756 19471 65772
tri 19471 65756 19487 65772 sw
rect 19394 65690 19487 65756
rect 19523 65631 19637 65789
tri 19673 65756 19689 65772 se
rect 19689 65756 19766 65772
rect 19673 65690 19766 65756
rect 19394 65555 19766 65631
rect 19394 65430 19487 65496
rect 19394 65414 19471 65430
tri 19471 65414 19487 65430 nw
rect 19523 65397 19637 65555
rect 19673 65430 19766 65496
tri 19673 65414 19689 65430 ne
rect 19689 65414 19766 65430
rect 19506 65315 19654 65397
rect 19394 65282 19471 65298
tri 19471 65282 19487 65298 sw
rect 19394 65216 19487 65282
rect 19394 65114 19487 65180
rect 19394 65098 19471 65114
tri 19471 65098 19487 65114 nw
rect 19523 65081 19637 65315
tri 19673 65282 19689 65298 se
rect 19689 65282 19766 65298
rect 19673 65216 19766 65282
rect 19673 65114 19766 65180
tri 19673 65098 19689 65114 ne
rect 19689 65098 19766 65114
rect 19506 64999 19654 65081
rect 19394 64966 19471 64982
tri 19471 64966 19487 64982 sw
rect 19394 64900 19487 64966
rect 19523 64841 19637 64999
tri 19673 64966 19689 64982 se
rect 19689 64966 19766 64982
rect 19673 64900 19766 64966
rect 19394 64765 19766 64841
rect 19394 64640 19487 64706
rect 19394 64624 19471 64640
tri 19471 64624 19487 64640 nw
rect 19523 64607 19637 64765
rect 19673 64640 19766 64706
tri 19673 64624 19689 64640 ne
rect 19689 64624 19766 64640
rect 19506 64525 19654 64607
rect 19394 64492 19471 64508
tri 19471 64492 19487 64508 sw
rect 19394 64426 19487 64492
rect 19394 64324 19487 64390
rect 19394 64308 19471 64324
tri 19471 64308 19487 64324 nw
rect 19523 64291 19637 64525
tri 19673 64492 19689 64508 se
rect 19689 64492 19766 64508
rect 19673 64426 19766 64492
rect 19673 64324 19766 64390
tri 19673 64308 19689 64324 ne
rect 19689 64308 19766 64324
rect 19506 64209 19654 64291
rect 19394 64176 19471 64192
tri 19471 64176 19487 64192 sw
rect 19394 64110 19487 64176
rect 19523 64051 19637 64209
tri 19673 64176 19689 64192 se
rect 19689 64176 19766 64192
rect 19673 64110 19766 64176
rect 19394 63975 19766 64051
rect 19394 63850 19487 63916
rect 19394 63834 19471 63850
tri 19471 63834 19487 63850 nw
rect 19523 63817 19637 63975
rect 19673 63850 19766 63916
tri 19673 63834 19689 63850 ne
rect 19689 63834 19766 63850
rect 19506 63735 19654 63817
rect 19394 63702 19471 63718
tri 19471 63702 19487 63718 sw
rect 19394 63636 19487 63702
rect 19394 63534 19487 63600
rect 19394 63518 19471 63534
tri 19471 63518 19487 63534 nw
rect 19523 63501 19637 63735
tri 19673 63702 19689 63718 se
rect 19689 63702 19766 63718
rect 19673 63636 19766 63702
rect 19673 63534 19766 63600
tri 19673 63518 19689 63534 ne
rect 19689 63518 19766 63534
rect 19506 63419 19654 63501
rect 19394 63386 19471 63402
tri 19471 63386 19487 63402 sw
rect 19394 63320 19487 63386
rect 19523 63261 19637 63419
tri 19673 63386 19689 63402 se
rect 19689 63386 19766 63402
rect 19673 63320 19766 63386
rect 19394 63185 19766 63261
rect 19394 63060 19487 63126
rect 19394 63044 19471 63060
tri 19471 63044 19487 63060 nw
rect 19523 63027 19637 63185
rect 19673 63060 19766 63126
tri 19673 63044 19689 63060 ne
rect 19689 63044 19766 63060
rect 19506 62945 19654 63027
rect 19394 62912 19471 62928
tri 19471 62912 19487 62928 sw
rect 19394 62846 19487 62912
rect 19394 62744 19487 62810
rect 19394 62728 19471 62744
tri 19471 62728 19487 62744 nw
rect 19523 62711 19637 62945
tri 19673 62912 19689 62928 se
rect 19689 62912 19766 62928
rect 19673 62846 19766 62912
rect 19673 62744 19766 62810
tri 19673 62728 19689 62744 ne
rect 19689 62728 19766 62744
rect 19506 62629 19654 62711
rect 19394 62596 19471 62612
tri 19471 62596 19487 62612 sw
rect 19394 62530 19487 62596
rect 19523 62471 19637 62629
tri 19673 62596 19689 62612 se
rect 19689 62596 19766 62612
rect 19673 62530 19766 62596
rect 19394 62395 19766 62471
rect 19394 62270 19487 62336
rect 19394 62254 19471 62270
tri 19471 62254 19487 62270 nw
rect 19523 62237 19637 62395
rect 19673 62270 19766 62336
tri 19673 62254 19689 62270 ne
rect 19689 62254 19766 62270
rect 19506 62155 19654 62237
rect 19394 62122 19471 62138
tri 19471 62122 19487 62138 sw
rect 19394 62056 19487 62122
rect 19394 61954 19487 62020
rect 19394 61938 19471 61954
tri 19471 61938 19487 61954 nw
rect 19523 61921 19637 62155
tri 19673 62122 19689 62138 se
rect 19689 62122 19766 62138
rect 19673 62056 19766 62122
rect 19673 61954 19766 62020
tri 19673 61938 19689 61954 ne
rect 19689 61938 19766 61954
rect 19506 61839 19654 61921
rect 19394 61806 19471 61822
tri 19471 61806 19487 61822 sw
rect 19394 61740 19487 61806
rect 19523 61681 19637 61839
tri 19673 61806 19689 61822 se
rect 19689 61806 19766 61822
rect 19673 61740 19766 61806
rect 19394 61605 19766 61681
rect 19394 61480 19487 61546
rect 19394 61464 19471 61480
tri 19471 61464 19487 61480 nw
rect 19523 61447 19637 61605
rect 19673 61480 19766 61546
tri 19673 61464 19689 61480 ne
rect 19689 61464 19766 61480
rect 19506 61365 19654 61447
rect 19394 61332 19471 61348
tri 19471 61332 19487 61348 sw
rect 19394 61266 19487 61332
rect 19394 61164 19487 61230
rect 19394 61148 19471 61164
tri 19471 61148 19487 61164 nw
rect 19523 61131 19637 61365
tri 19673 61332 19689 61348 se
rect 19689 61332 19766 61348
rect 19673 61266 19766 61332
rect 19673 61164 19766 61230
tri 19673 61148 19689 61164 ne
rect 19689 61148 19766 61164
rect 19506 61049 19654 61131
rect 19394 61016 19471 61032
tri 19471 61016 19487 61032 sw
rect 19394 60950 19487 61016
rect 19523 60891 19637 61049
tri 19673 61016 19689 61032 se
rect 19689 61016 19766 61032
rect 19673 60950 19766 61016
rect 19394 60815 19766 60891
rect 19394 60690 19487 60756
rect 19394 60674 19471 60690
tri 19471 60674 19487 60690 nw
rect 19523 60657 19637 60815
rect 19673 60690 19766 60756
tri 19673 60674 19689 60690 ne
rect 19689 60674 19766 60690
rect 19506 60575 19654 60657
rect 19394 60542 19471 60558
tri 19471 60542 19487 60558 sw
rect 19394 60476 19487 60542
rect 19394 60374 19487 60440
rect 19394 60358 19471 60374
tri 19471 60358 19487 60374 nw
rect 19523 60341 19637 60575
tri 19673 60542 19689 60558 se
rect 19689 60542 19766 60558
rect 19673 60476 19766 60542
rect 19673 60374 19766 60440
tri 19673 60358 19689 60374 ne
rect 19689 60358 19766 60374
rect 19506 60259 19654 60341
rect 19394 60226 19471 60242
tri 19471 60226 19487 60242 sw
rect 19394 60160 19487 60226
rect 19523 60101 19637 60259
tri 19673 60226 19689 60242 se
rect 19689 60226 19766 60242
rect 19673 60160 19766 60226
rect 19394 60025 19766 60101
rect 19394 59900 19487 59966
rect 19394 59884 19471 59900
tri 19471 59884 19487 59900 nw
rect 19523 59867 19637 60025
rect 19673 59900 19766 59966
tri 19673 59884 19689 59900 ne
rect 19689 59884 19766 59900
rect 19506 59785 19654 59867
rect 19394 59752 19471 59768
tri 19471 59752 19487 59768 sw
rect 19394 59686 19487 59752
rect 19394 59584 19487 59650
rect 19394 59568 19471 59584
tri 19471 59568 19487 59584 nw
rect 19523 59551 19637 59785
tri 19673 59752 19689 59768 se
rect 19689 59752 19766 59768
rect 19673 59686 19766 59752
rect 19673 59584 19766 59650
tri 19673 59568 19689 59584 ne
rect 19689 59568 19766 59584
rect 19506 59469 19654 59551
rect 19394 59436 19471 59452
tri 19471 59436 19487 59452 sw
rect 19394 59370 19487 59436
rect 19523 59311 19637 59469
tri 19673 59436 19689 59452 se
rect 19689 59436 19766 59452
rect 19673 59370 19766 59436
rect 19394 59235 19766 59311
rect 19394 59110 19487 59176
rect 19394 59094 19471 59110
tri 19471 59094 19487 59110 nw
rect 19523 59077 19637 59235
rect 19673 59110 19766 59176
tri 19673 59094 19689 59110 ne
rect 19689 59094 19766 59110
rect 19506 58995 19654 59077
rect 19394 58962 19471 58978
tri 19471 58962 19487 58978 sw
rect 19394 58896 19487 58962
rect 19394 58794 19487 58860
rect 19394 58778 19471 58794
tri 19471 58778 19487 58794 nw
rect 19523 58761 19637 58995
tri 19673 58962 19689 58978 se
rect 19689 58962 19766 58978
rect 19673 58896 19766 58962
rect 19673 58794 19766 58860
tri 19673 58778 19689 58794 ne
rect 19689 58778 19766 58794
rect 19506 58679 19654 58761
rect 19394 58646 19471 58662
tri 19471 58646 19487 58662 sw
rect 19394 58580 19487 58646
rect 19523 58521 19637 58679
tri 19673 58646 19689 58662 se
rect 19689 58646 19766 58662
rect 19673 58580 19766 58646
rect 19394 58445 19766 58521
rect 19394 58320 19487 58386
rect 19394 58304 19471 58320
tri 19471 58304 19487 58320 nw
rect 19523 58287 19637 58445
rect 19673 58320 19766 58386
tri 19673 58304 19689 58320 ne
rect 19689 58304 19766 58320
rect 19506 58205 19654 58287
rect 19394 58172 19471 58188
tri 19471 58172 19487 58188 sw
rect 19394 58106 19487 58172
rect 19394 58004 19487 58070
rect 19394 57988 19471 58004
tri 19471 57988 19487 58004 nw
rect 19523 57971 19637 58205
tri 19673 58172 19689 58188 se
rect 19689 58172 19766 58188
rect 19673 58106 19766 58172
rect 19673 58004 19766 58070
tri 19673 57988 19689 58004 ne
rect 19689 57988 19766 58004
rect 19506 57889 19654 57971
rect 19394 57856 19471 57872
tri 19471 57856 19487 57872 sw
rect 19394 57790 19487 57856
rect 19523 57731 19637 57889
tri 19673 57856 19689 57872 se
rect 19689 57856 19766 57872
rect 19673 57790 19766 57856
rect 19394 57655 19766 57731
rect 19394 57530 19487 57596
rect 19394 57514 19471 57530
tri 19471 57514 19487 57530 nw
rect 19523 57497 19637 57655
rect 19673 57530 19766 57596
tri 19673 57514 19689 57530 ne
rect 19689 57514 19766 57530
rect 19506 57415 19654 57497
rect 19394 57382 19471 57398
tri 19471 57382 19487 57398 sw
rect 19394 57316 19487 57382
rect 19394 57214 19487 57280
rect 19394 57198 19471 57214
tri 19471 57198 19487 57214 nw
rect 19523 57181 19637 57415
tri 19673 57382 19689 57398 se
rect 19689 57382 19766 57398
rect 19673 57316 19766 57382
rect 19673 57214 19766 57280
tri 19673 57198 19689 57214 ne
rect 19689 57198 19766 57214
rect 19506 57099 19654 57181
rect 19394 57066 19471 57082
tri 19471 57066 19487 57082 sw
rect 19394 57000 19487 57066
rect 19523 56941 19637 57099
tri 19673 57066 19689 57082 se
rect 19689 57066 19766 57082
rect 19673 57000 19766 57066
rect 19394 56865 19766 56941
rect 19394 56740 19487 56806
rect 19394 56724 19471 56740
tri 19471 56724 19487 56740 nw
rect 19523 56707 19637 56865
rect 19673 56740 19766 56806
tri 19673 56724 19689 56740 ne
rect 19689 56724 19766 56740
rect 19506 56625 19654 56707
rect 19394 56592 19471 56608
tri 19471 56592 19487 56608 sw
rect 19394 56526 19487 56592
rect 19394 56424 19487 56490
rect 19394 56408 19471 56424
tri 19471 56408 19487 56424 nw
rect 19523 56391 19637 56625
tri 19673 56592 19689 56608 se
rect 19689 56592 19766 56608
rect 19673 56526 19766 56592
rect 19673 56424 19766 56490
tri 19673 56408 19689 56424 ne
rect 19689 56408 19766 56424
rect 19506 56309 19654 56391
rect 19394 56276 19471 56292
tri 19471 56276 19487 56292 sw
rect 19394 56210 19487 56276
rect 19523 56151 19637 56309
tri 19673 56276 19689 56292 se
rect 19689 56276 19766 56292
rect 19673 56210 19766 56276
rect 19394 56075 19766 56151
rect 19394 55950 19487 56016
rect 19394 55934 19471 55950
tri 19471 55934 19487 55950 nw
rect 19523 55917 19637 56075
rect 19673 55950 19766 56016
tri 19673 55934 19689 55950 ne
rect 19689 55934 19766 55950
rect 19506 55835 19654 55917
rect 19394 55802 19471 55818
tri 19471 55802 19487 55818 sw
rect 19394 55736 19487 55802
rect 19394 55634 19487 55700
rect 19394 55618 19471 55634
tri 19471 55618 19487 55634 nw
rect 19523 55601 19637 55835
tri 19673 55802 19689 55818 se
rect 19689 55802 19766 55818
rect 19673 55736 19766 55802
rect 19673 55634 19766 55700
tri 19673 55618 19689 55634 ne
rect 19689 55618 19766 55634
rect 19506 55519 19654 55601
rect 19394 55486 19471 55502
tri 19471 55486 19487 55502 sw
rect 19394 55420 19487 55486
rect 19523 55361 19637 55519
tri 19673 55486 19689 55502 se
rect 19689 55486 19766 55502
rect 19673 55420 19766 55486
rect 19394 55285 19766 55361
rect 19394 55160 19487 55226
rect 19394 55144 19471 55160
tri 19471 55144 19487 55160 nw
rect 19523 55127 19637 55285
rect 19673 55160 19766 55226
tri 19673 55144 19689 55160 ne
rect 19689 55144 19766 55160
rect 19506 55045 19654 55127
rect 19394 55012 19471 55028
tri 19471 55012 19487 55028 sw
rect 19394 54946 19487 55012
rect 19394 54844 19487 54910
rect 19394 54828 19471 54844
tri 19471 54828 19487 54844 nw
rect 19523 54811 19637 55045
tri 19673 55012 19689 55028 se
rect 19689 55012 19766 55028
rect 19673 54946 19766 55012
rect 19673 54844 19766 54910
tri 19673 54828 19689 54844 ne
rect 19689 54828 19766 54844
rect 19506 54729 19654 54811
rect 19394 54696 19471 54712
tri 19471 54696 19487 54712 sw
rect 19394 54630 19487 54696
rect 19523 54571 19637 54729
tri 19673 54696 19689 54712 se
rect 19689 54696 19766 54712
rect 19673 54630 19766 54696
rect 19394 54495 19766 54571
rect 19394 54370 19487 54436
rect 19394 54354 19471 54370
tri 19471 54354 19487 54370 nw
rect 19523 54337 19637 54495
rect 19673 54370 19766 54436
tri 19673 54354 19689 54370 ne
rect 19689 54354 19766 54370
rect 19506 54255 19654 54337
rect 19394 54222 19471 54238
tri 19471 54222 19487 54238 sw
rect 19394 54156 19487 54222
rect 19394 54054 19487 54120
rect 19394 54038 19471 54054
tri 19471 54038 19487 54054 nw
rect 19523 54021 19637 54255
tri 19673 54222 19689 54238 se
rect 19689 54222 19766 54238
rect 19673 54156 19766 54222
rect 19673 54054 19766 54120
tri 19673 54038 19689 54054 ne
rect 19689 54038 19766 54054
rect 19506 53939 19654 54021
rect 19394 53906 19471 53922
tri 19471 53906 19487 53922 sw
rect 19394 53840 19487 53906
rect 19523 53781 19637 53939
tri 19673 53906 19689 53922 se
rect 19689 53906 19766 53922
rect 19673 53840 19766 53906
rect 19394 53705 19766 53781
rect 19394 53580 19487 53646
rect 19394 53564 19471 53580
tri 19471 53564 19487 53580 nw
rect 19523 53547 19637 53705
rect 19673 53580 19766 53646
tri 19673 53564 19689 53580 ne
rect 19689 53564 19766 53580
rect 19506 53465 19654 53547
rect 19394 53432 19471 53448
tri 19471 53432 19487 53448 sw
rect 19394 53366 19487 53432
rect 19394 53264 19487 53330
rect 19394 53248 19471 53264
tri 19471 53248 19487 53264 nw
rect 19523 53231 19637 53465
tri 19673 53432 19689 53448 se
rect 19689 53432 19766 53448
rect 19673 53366 19766 53432
rect 19673 53264 19766 53330
tri 19673 53248 19689 53264 ne
rect 19689 53248 19766 53264
rect 19506 53149 19654 53231
rect 19394 53116 19471 53132
tri 19471 53116 19487 53132 sw
rect 19394 53050 19487 53116
rect 19523 52991 19637 53149
tri 19673 53116 19689 53132 se
rect 19689 53116 19766 53132
rect 19673 53050 19766 53116
rect 19394 52915 19766 52991
rect 19394 52790 19487 52856
rect 19394 52774 19471 52790
tri 19471 52774 19487 52790 nw
rect 19523 52757 19637 52915
rect 19673 52790 19766 52856
tri 19673 52774 19689 52790 ne
rect 19689 52774 19766 52790
rect 19506 52675 19654 52757
rect 19394 52642 19471 52658
tri 19471 52642 19487 52658 sw
rect 19394 52576 19487 52642
rect 19394 52474 19487 52540
rect 19394 52458 19471 52474
tri 19471 52458 19487 52474 nw
rect 19523 52441 19637 52675
tri 19673 52642 19689 52658 se
rect 19689 52642 19766 52658
rect 19673 52576 19766 52642
rect 19673 52474 19766 52540
tri 19673 52458 19689 52474 ne
rect 19689 52458 19766 52474
rect 19506 52359 19654 52441
rect 19394 52326 19471 52342
tri 19471 52326 19487 52342 sw
rect 19394 52260 19487 52326
rect 19523 52201 19637 52359
tri 19673 52326 19689 52342 se
rect 19689 52326 19766 52342
rect 19673 52260 19766 52326
rect 19394 52125 19766 52201
rect 19394 52000 19487 52066
rect 19394 51984 19471 52000
tri 19471 51984 19487 52000 nw
rect 19523 51967 19637 52125
rect 19673 52000 19766 52066
tri 19673 51984 19689 52000 ne
rect 19689 51984 19766 52000
rect 19506 51885 19654 51967
rect 19394 51852 19471 51868
tri 19471 51852 19487 51868 sw
rect 19394 51786 19487 51852
rect 19394 51684 19487 51750
rect 19394 51668 19471 51684
tri 19471 51668 19487 51684 nw
rect 19523 51651 19637 51885
tri 19673 51852 19689 51868 se
rect 19689 51852 19766 51868
rect 19673 51786 19766 51852
rect 19673 51684 19766 51750
tri 19673 51668 19689 51684 ne
rect 19689 51668 19766 51684
rect 19506 51569 19654 51651
rect 19394 51536 19471 51552
tri 19471 51536 19487 51552 sw
rect 19394 51470 19487 51536
rect 19523 51411 19637 51569
tri 19673 51536 19689 51552 se
rect 19689 51536 19766 51552
rect 19673 51470 19766 51536
rect 19394 51335 19766 51411
rect 19394 51210 19487 51276
rect 19394 51194 19471 51210
tri 19471 51194 19487 51210 nw
rect 19523 51177 19637 51335
rect 19673 51210 19766 51276
tri 19673 51194 19689 51210 ne
rect 19689 51194 19766 51210
rect 19506 51095 19654 51177
rect 19394 51062 19471 51078
tri 19471 51062 19487 51078 sw
rect 19394 50996 19487 51062
rect 19394 50894 19487 50960
rect 19394 50878 19471 50894
tri 19471 50878 19487 50894 nw
rect 19523 50861 19637 51095
tri 19673 51062 19689 51078 se
rect 19689 51062 19766 51078
rect 19673 50996 19766 51062
rect 19673 50894 19766 50960
tri 19673 50878 19689 50894 ne
rect 19689 50878 19766 50894
rect 19506 50779 19654 50861
rect 19394 50746 19471 50762
tri 19471 50746 19487 50762 sw
rect 19394 50680 19487 50746
rect 19523 50621 19637 50779
tri 19673 50746 19689 50762 se
rect 19689 50746 19766 50762
rect 19673 50680 19766 50746
rect 19394 50545 19766 50621
rect 19394 50420 19487 50486
rect 19394 50404 19471 50420
tri 19471 50404 19487 50420 nw
rect 19523 50387 19637 50545
rect 19673 50420 19766 50486
tri 19673 50404 19689 50420 ne
rect 19689 50404 19766 50420
rect 19506 50305 19654 50387
rect 19394 50272 19471 50288
tri 19471 50272 19487 50288 sw
rect 19394 50206 19487 50272
rect 19394 50104 19487 50170
rect 19394 50088 19471 50104
tri 19471 50088 19487 50104 nw
rect 19523 50071 19637 50305
tri 19673 50272 19689 50288 se
rect 19689 50272 19766 50288
rect 19673 50206 19766 50272
rect 19673 50104 19766 50170
tri 19673 50088 19689 50104 ne
rect 19689 50088 19766 50104
rect 19506 49989 19654 50071
rect 19394 49956 19471 49972
tri 19471 49956 19487 49972 sw
rect 19394 49890 19487 49956
rect 19523 49831 19637 49989
tri 19673 49956 19689 49972 se
rect 19689 49956 19766 49972
rect 19673 49890 19766 49956
rect 19394 49755 19766 49831
rect 19394 49630 19487 49696
rect 19394 49614 19471 49630
tri 19471 49614 19487 49630 nw
rect 19523 49597 19637 49755
rect 19673 49630 19766 49696
tri 19673 49614 19689 49630 ne
rect 19689 49614 19766 49630
rect 19506 49515 19654 49597
rect 19394 49482 19471 49498
tri 19471 49482 19487 49498 sw
rect 19394 49416 19487 49482
rect 19394 49314 19487 49380
rect 19394 49298 19471 49314
tri 19471 49298 19487 49314 nw
rect 19523 49281 19637 49515
tri 19673 49482 19689 49498 se
rect 19689 49482 19766 49498
rect 19673 49416 19766 49482
rect 19673 49314 19766 49380
tri 19673 49298 19689 49314 ne
rect 19689 49298 19766 49314
rect 19506 49199 19654 49281
rect 19394 49166 19471 49182
tri 19471 49166 19487 49182 sw
rect 19394 49100 19487 49166
rect 19523 49041 19637 49199
tri 19673 49166 19689 49182 se
rect 19689 49166 19766 49182
rect 19673 49100 19766 49166
rect 19394 48965 19766 49041
rect 19394 48840 19487 48906
rect 19394 48824 19471 48840
tri 19471 48824 19487 48840 nw
rect 19523 48807 19637 48965
rect 19673 48840 19766 48906
tri 19673 48824 19689 48840 ne
rect 19689 48824 19766 48840
rect 19506 48725 19654 48807
rect 19394 48692 19471 48708
tri 19471 48692 19487 48708 sw
rect 19394 48626 19487 48692
rect 19394 48524 19487 48590
rect 19394 48508 19471 48524
tri 19471 48508 19487 48524 nw
rect 19523 48491 19637 48725
tri 19673 48692 19689 48708 se
rect 19689 48692 19766 48708
rect 19673 48626 19766 48692
rect 19673 48524 19766 48590
tri 19673 48508 19689 48524 ne
rect 19689 48508 19766 48524
rect 19506 48409 19654 48491
rect 19394 48376 19471 48392
tri 19471 48376 19487 48392 sw
rect 19394 48310 19487 48376
rect 19523 48251 19637 48409
tri 19673 48376 19689 48392 se
rect 19689 48376 19766 48392
rect 19673 48310 19766 48376
rect 19394 48175 19766 48251
rect 19394 48050 19487 48116
rect 19394 48034 19471 48050
tri 19471 48034 19487 48050 nw
rect 19523 48017 19637 48175
rect 19673 48050 19766 48116
tri 19673 48034 19689 48050 ne
rect 19689 48034 19766 48050
rect 19506 47935 19654 48017
rect 19394 47902 19471 47918
tri 19471 47902 19487 47918 sw
rect 19394 47836 19487 47902
rect 19394 47734 19487 47800
rect 19394 47718 19471 47734
tri 19471 47718 19487 47734 nw
rect 19523 47701 19637 47935
tri 19673 47902 19689 47918 se
rect 19689 47902 19766 47918
rect 19673 47836 19766 47902
rect 19673 47734 19766 47800
tri 19673 47718 19689 47734 ne
rect 19689 47718 19766 47734
rect 19506 47619 19654 47701
rect 19394 47586 19471 47602
tri 19471 47586 19487 47602 sw
rect 19394 47520 19487 47586
rect 19523 47461 19637 47619
tri 19673 47586 19689 47602 se
rect 19689 47586 19766 47602
rect 19673 47520 19766 47586
rect 19394 47385 19766 47461
rect 19394 47260 19487 47326
rect 19394 47244 19471 47260
tri 19471 47244 19487 47260 nw
rect 19523 47227 19637 47385
rect 19673 47260 19766 47326
tri 19673 47244 19689 47260 ne
rect 19689 47244 19766 47260
rect 19506 47145 19654 47227
rect 19394 47112 19471 47128
tri 19471 47112 19487 47128 sw
rect 19394 47046 19487 47112
rect 19394 46944 19487 47010
rect 19394 46928 19471 46944
tri 19471 46928 19487 46944 nw
rect 19523 46911 19637 47145
tri 19673 47112 19689 47128 se
rect 19689 47112 19766 47128
rect 19673 47046 19766 47112
rect 19673 46944 19766 47010
tri 19673 46928 19689 46944 ne
rect 19689 46928 19766 46944
rect 19506 46829 19654 46911
rect 19394 46796 19471 46812
tri 19471 46796 19487 46812 sw
rect 19394 46730 19487 46796
rect 19523 46671 19637 46829
tri 19673 46796 19689 46812 se
rect 19689 46796 19766 46812
rect 19673 46730 19766 46796
rect 19394 46595 19766 46671
rect 19394 46470 19487 46536
rect 19394 46454 19471 46470
tri 19471 46454 19487 46470 nw
rect 19523 46437 19637 46595
rect 19673 46470 19766 46536
tri 19673 46454 19689 46470 ne
rect 19689 46454 19766 46470
rect 19506 46355 19654 46437
rect 19394 46322 19471 46338
tri 19471 46322 19487 46338 sw
rect 19394 46256 19487 46322
rect 19394 46154 19487 46220
rect 19394 46138 19471 46154
tri 19471 46138 19487 46154 nw
rect 19523 46121 19637 46355
tri 19673 46322 19689 46338 se
rect 19689 46322 19766 46338
rect 19673 46256 19766 46322
rect 19673 46154 19766 46220
tri 19673 46138 19689 46154 ne
rect 19689 46138 19766 46154
rect 19506 46039 19654 46121
rect 19394 46006 19471 46022
tri 19471 46006 19487 46022 sw
rect 19394 45940 19487 46006
rect 19523 45881 19637 46039
tri 19673 46006 19689 46022 se
rect 19689 46006 19766 46022
rect 19673 45940 19766 46006
rect 19394 45805 19766 45881
rect 19394 45680 19487 45746
rect 19394 45664 19471 45680
tri 19471 45664 19487 45680 nw
rect 19523 45647 19637 45805
rect 19673 45680 19766 45746
tri 19673 45664 19689 45680 ne
rect 19689 45664 19766 45680
rect 19506 45565 19654 45647
rect 19394 45532 19471 45548
tri 19471 45532 19487 45548 sw
rect 19394 45466 19487 45532
rect 19394 45364 19487 45430
rect 19394 45348 19471 45364
tri 19471 45348 19487 45364 nw
rect 19523 45331 19637 45565
tri 19673 45532 19689 45548 se
rect 19689 45532 19766 45548
rect 19673 45466 19766 45532
rect 19673 45364 19766 45430
tri 19673 45348 19689 45364 ne
rect 19689 45348 19766 45364
rect 19506 45249 19654 45331
rect 19394 45216 19471 45232
tri 19471 45216 19487 45232 sw
rect 19394 45150 19487 45216
rect 19523 45091 19637 45249
tri 19673 45216 19689 45232 se
rect 19689 45216 19766 45232
rect 19673 45150 19766 45216
rect 19394 45015 19766 45091
rect 19394 44890 19487 44956
rect 19394 44874 19471 44890
tri 19471 44874 19487 44890 nw
rect 19523 44857 19637 45015
rect 19673 44890 19766 44956
tri 19673 44874 19689 44890 ne
rect 19689 44874 19766 44890
rect 19506 44775 19654 44857
rect 19394 44742 19471 44758
tri 19471 44742 19487 44758 sw
rect 19394 44676 19487 44742
rect 19394 44574 19487 44640
rect 19394 44558 19471 44574
tri 19471 44558 19487 44574 nw
rect 19523 44541 19637 44775
tri 19673 44742 19689 44758 se
rect 19689 44742 19766 44758
rect 19673 44676 19766 44742
rect 19673 44574 19766 44640
tri 19673 44558 19689 44574 ne
rect 19689 44558 19766 44574
rect 19506 44459 19654 44541
rect 19394 44426 19471 44442
tri 19471 44426 19487 44442 sw
rect 19394 44360 19487 44426
rect 19523 44301 19637 44459
tri 19673 44426 19689 44442 se
rect 19689 44426 19766 44442
rect 19673 44360 19766 44426
rect 19394 44225 19766 44301
rect 19394 44100 19487 44166
rect 19394 44084 19471 44100
tri 19471 44084 19487 44100 nw
rect 19523 44067 19637 44225
rect 19673 44100 19766 44166
tri 19673 44084 19689 44100 ne
rect 19689 44084 19766 44100
rect 19506 43985 19654 44067
rect 19394 43952 19471 43968
tri 19471 43952 19487 43968 sw
rect 19394 43886 19487 43952
rect 19394 43784 19487 43850
rect 19394 43768 19471 43784
tri 19471 43768 19487 43784 nw
rect 19523 43751 19637 43985
tri 19673 43952 19689 43968 se
rect 19689 43952 19766 43968
rect 19673 43886 19766 43952
rect 19673 43784 19766 43850
tri 19673 43768 19689 43784 ne
rect 19689 43768 19766 43784
rect 19506 43669 19654 43751
rect 19394 43636 19471 43652
tri 19471 43636 19487 43652 sw
rect 19394 43570 19487 43636
rect 19523 43511 19637 43669
tri 19673 43636 19689 43652 se
rect 19689 43636 19766 43652
rect 19673 43570 19766 43636
rect 19394 43435 19766 43511
rect 19394 43310 19487 43376
rect 19394 43294 19471 43310
tri 19471 43294 19487 43310 nw
rect 19523 43277 19637 43435
rect 19673 43310 19766 43376
tri 19673 43294 19689 43310 ne
rect 19689 43294 19766 43310
rect 19506 43195 19654 43277
rect 19394 43162 19471 43178
tri 19471 43162 19487 43178 sw
rect 19394 43096 19487 43162
rect 19394 42994 19487 43060
rect 19394 42978 19471 42994
tri 19471 42978 19487 42994 nw
rect 19523 42961 19637 43195
tri 19673 43162 19689 43178 se
rect 19689 43162 19766 43178
rect 19673 43096 19766 43162
rect 19673 42994 19766 43060
tri 19673 42978 19689 42994 ne
rect 19689 42978 19766 42994
rect 19506 42879 19654 42961
rect 19394 42846 19471 42862
tri 19471 42846 19487 42862 sw
rect 19394 42780 19487 42846
rect 19523 42721 19637 42879
tri 19673 42846 19689 42862 se
rect 19689 42846 19766 42862
rect 19673 42780 19766 42846
rect 19394 42645 19766 42721
rect 19394 42520 19487 42586
rect 19394 42504 19471 42520
tri 19471 42504 19487 42520 nw
rect 19523 42487 19637 42645
rect 19673 42520 19766 42586
tri 19673 42504 19689 42520 ne
rect 19689 42504 19766 42520
rect 19506 42405 19654 42487
rect 19394 42372 19471 42388
tri 19471 42372 19487 42388 sw
rect 19394 42306 19487 42372
rect 19394 42204 19487 42270
rect 19394 42188 19471 42204
tri 19471 42188 19487 42204 nw
rect 19523 42171 19637 42405
tri 19673 42372 19689 42388 se
rect 19689 42372 19766 42388
rect 19673 42306 19766 42372
rect 19673 42204 19766 42270
tri 19673 42188 19689 42204 ne
rect 19689 42188 19766 42204
rect 19506 42089 19654 42171
rect 19394 42056 19471 42072
tri 19471 42056 19487 42072 sw
rect 19394 41990 19487 42056
rect 19523 41931 19637 42089
tri 19673 42056 19689 42072 se
rect 19689 42056 19766 42072
rect 19673 41990 19766 42056
rect 19394 41855 19766 41931
rect 19394 41730 19487 41796
rect 19394 41714 19471 41730
tri 19471 41714 19487 41730 nw
rect 19523 41697 19637 41855
rect 19673 41730 19766 41796
tri 19673 41714 19689 41730 ne
rect 19689 41714 19766 41730
rect 19506 41615 19654 41697
rect 19394 41582 19471 41598
tri 19471 41582 19487 41598 sw
rect 19394 41516 19487 41582
rect 19394 41414 19487 41480
rect 19394 41398 19471 41414
tri 19471 41398 19487 41414 nw
rect 19523 41381 19637 41615
tri 19673 41582 19689 41598 se
rect 19689 41582 19766 41598
rect 19673 41516 19766 41582
rect 19673 41414 19766 41480
tri 19673 41398 19689 41414 ne
rect 19689 41398 19766 41414
rect 19506 41299 19654 41381
rect 19394 41266 19471 41282
tri 19471 41266 19487 41282 sw
rect 19394 41200 19487 41266
rect 19523 41141 19637 41299
tri 19673 41266 19689 41282 se
rect 19689 41266 19766 41282
rect 19673 41200 19766 41266
rect 19394 41065 19766 41141
rect 19394 40940 19487 41006
rect 19394 40924 19471 40940
tri 19471 40924 19487 40940 nw
rect 19523 40907 19637 41065
rect 19673 40940 19766 41006
tri 19673 40924 19689 40940 ne
rect 19689 40924 19766 40940
rect 19506 40825 19654 40907
rect 19394 40792 19471 40808
tri 19471 40792 19487 40808 sw
rect 19394 40726 19487 40792
rect 19394 40624 19487 40690
rect 19394 40608 19471 40624
tri 19471 40608 19487 40624 nw
rect 19523 40591 19637 40825
tri 19673 40792 19689 40808 se
rect 19689 40792 19766 40808
rect 19673 40726 19766 40792
rect 19673 40624 19766 40690
tri 19673 40608 19689 40624 ne
rect 19689 40608 19766 40624
rect 19506 40509 19654 40591
rect 19394 40476 19471 40492
tri 19471 40476 19487 40492 sw
rect 19394 40410 19487 40476
rect 19523 40351 19637 40509
tri 19673 40476 19689 40492 se
rect 19689 40476 19766 40492
rect 19673 40410 19766 40476
rect 19394 40275 19766 40351
rect 19394 40150 19487 40216
rect 19394 40134 19471 40150
tri 19471 40134 19487 40150 nw
rect 19523 40117 19637 40275
rect 19673 40150 19766 40216
tri 19673 40134 19689 40150 ne
rect 19689 40134 19766 40150
rect 19506 40035 19654 40117
rect 19394 40002 19471 40018
tri 19471 40002 19487 40018 sw
rect 19394 39936 19487 40002
rect 19394 39834 19487 39900
rect 19394 39818 19471 39834
tri 19471 39818 19487 39834 nw
rect 19523 39801 19637 40035
tri 19673 40002 19689 40018 se
rect 19689 40002 19766 40018
rect 19673 39936 19766 40002
rect 19673 39834 19766 39900
tri 19673 39818 19689 39834 ne
rect 19689 39818 19766 39834
rect 19506 39719 19654 39801
rect 19394 39686 19471 39702
tri 19471 39686 19487 39702 sw
rect 19394 39620 19487 39686
rect 19523 39561 19637 39719
tri 19673 39686 19689 39702 se
rect 19689 39686 19766 39702
rect 19673 39620 19766 39686
rect 19394 39485 19766 39561
rect 19394 39360 19487 39426
rect 19394 39344 19471 39360
tri 19471 39344 19487 39360 nw
rect 19523 39327 19637 39485
rect 19673 39360 19766 39426
tri 19673 39344 19689 39360 ne
rect 19689 39344 19766 39360
rect 19506 39245 19654 39327
rect 19394 39212 19471 39228
tri 19471 39212 19487 39228 sw
rect 19394 39146 19487 39212
rect 19394 39044 19487 39110
rect 19394 39028 19471 39044
tri 19471 39028 19487 39044 nw
rect 19523 39011 19637 39245
tri 19673 39212 19689 39228 se
rect 19689 39212 19766 39228
rect 19673 39146 19766 39212
rect 19673 39044 19766 39110
tri 19673 39028 19689 39044 ne
rect 19689 39028 19766 39044
rect 19506 38929 19654 39011
rect 19394 38896 19471 38912
tri 19471 38896 19487 38912 sw
rect 19394 38830 19487 38896
rect 19523 38771 19637 38929
tri 19673 38896 19689 38912 se
rect 19689 38896 19766 38912
rect 19673 38830 19766 38896
rect 19394 38695 19766 38771
rect 19394 38570 19487 38636
rect 19394 38554 19471 38570
tri 19471 38554 19487 38570 nw
rect 19523 38537 19637 38695
rect 19673 38570 19766 38636
tri 19673 38554 19689 38570 ne
rect 19689 38554 19766 38570
rect 19506 38455 19654 38537
rect 19394 38422 19471 38438
tri 19471 38422 19487 38438 sw
rect 19394 38356 19487 38422
rect 19394 38254 19487 38320
rect 19394 38238 19471 38254
tri 19471 38238 19487 38254 nw
rect 19523 38221 19637 38455
tri 19673 38422 19689 38438 se
rect 19689 38422 19766 38438
rect 19673 38356 19766 38422
rect 19673 38254 19766 38320
tri 19673 38238 19689 38254 ne
rect 19689 38238 19766 38254
rect 19506 38139 19654 38221
rect 19394 38106 19471 38122
tri 19471 38106 19487 38122 sw
rect 19394 38040 19487 38106
rect 19523 37981 19637 38139
tri 19673 38106 19689 38122 se
rect 19689 38106 19766 38122
rect 19673 38040 19766 38106
rect 19394 37905 19766 37981
rect 19394 37780 19487 37846
rect 19394 37764 19471 37780
tri 19471 37764 19487 37780 nw
rect 19523 37747 19637 37905
rect 19673 37780 19766 37846
tri 19673 37764 19689 37780 ne
rect 19689 37764 19766 37780
rect 19506 37665 19654 37747
rect 19394 37632 19471 37648
tri 19471 37632 19487 37648 sw
rect 19394 37566 19487 37632
rect 19394 37464 19487 37530
rect 19394 37448 19471 37464
tri 19471 37448 19487 37464 nw
rect 19523 37431 19637 37665
tri 19673 37632 19689 37648 se
rect 19689 37632 19766 37648
rect 19673 37566 19766 37632
rect 19673 37464 19766 37530
tri 19673 37448 19689 37464 ne
rect 19689 37448 19766 37464
rect 19506 37349 19654 37431
rect 19394 37316 19471 37332
tri 19471 37316 19487 37332 sw
rect 19394 37250 19487 37316
rect 19523 37191 19637 37349
tri 19673 37316 19689 37332 se
rect 19689 37316 19766 37332
rect 19673 37250 19766 37316
rect 19394 37115 19766 37191
rect 19394 36990 19487 37056
rect 19394 36974 19471 36990
tri 19471 36974 19487 36990 nw
rect 19523 36957 19637 37115
rect 19673 36990 19766 37056
tri 19673 36974 19689 36990 ne
rect 19689 36974 19766 36990
rect 19506 36875 19654 36957
rect 19394 36842 19471 36858
tri 19471 36842 19487 36858 sw
rect 19394 36776 19487 36842
rect 19394 36674 19487 36740
rect 19394 36658 19471 36674
tri 19471 36658 19487 36674 nw
rect 19523 36641 19637 36875
tri 19673 36842 19689 36858 se
rect 19689 36842 19766 36858
rect 19673 36776 19766 36842
rect 19673 36674 19766 36740
tri 19673 36658 19689 36674 ne
rect 19689 36658 19766 36674
rect 19506 36559 19654 36641
rect 19394 36526 19471 36542
tri 19471 36526 19487 36542 sw
rect 19394 36460 19487 36526
rect 19523 36401 19637 36559
tri 19673 36526 19689 36542 se
rect 19689 36526 19766 36542
rect 19673 36460 19766 36526
rect 19394 36325 19766 36401
rect 19394 36200 19487 36266
rect 19394 36184 19471 36200
tri 19471 36184 19487 36200 nw
rect 19523 36167 19637 36325
rect 19673 36200 19766 36266
tri 19673 36184 19689 36200 ne
rect 19689 36184 19766 36200
rect 19506 36085 19654 36167
rect 19394 36052 19471 36068
tri 19471 36052 19487 36068 sw
rect 19394 35986 19487 36052
rect 19394 35884 19487 35950
rect 19394 35868 19471 35884
tri 19471 35868 19487 35884 nw
rect 19523 35851 19637 36085
tri 19673 36052 19689 36068 se
rect 19689 36052 19766 36068
rect 19673 35986 19766 36052
rect 19673 35884 19766 35950
tri 19673 35868 19689 35884 ne
rect 19689 35868 19766 35884
rect 19506 35769 19654 35851
rect 19394 35736 19471 35752
tri 19471 35736 19487 35752 sw
rect 19394 35670 19487 35736
rect 19523 35611 19637 35769
tri 19673 35736 19689 35752 se
rect 19689 35736 19766 35752
rect 19673 35670 19766 35736
rect 19394 35535 19766 35611
rect 19394 35410 19487 35476
rect 19394 35394 19471 35410
tri 19471 35394 19487 35410 nw
rect 19523 35377 19637 35535
rect 19673 35410 19766 35476
tri 19673 35394 19689 35410 ne
rect 19689 35394 19766 35410
rect 19506 35295 19654 35377
rect 19394 35262 19471 35278
tri 19471 35262 19487 35278 sw
rect 19394 35196 19487 35262
rect 19394 35094 19487 35160
rect 19394 35078 19471 35094
tri 19471 35078 19487 35094 nw
rect 19523 35061 19637 35295
tri 19673 35262 19689 35278 se
rect 19689 35262 19766 35278
rect 19673 35196 19766 35262
rect 19673 35094 19766 35160
tri 19673 35078 19689 35094 ne
rect 19689 35078 19766 35094
rect 19506 34979 19654 35061
rect 19394 34946 19471 34962
tri 19471 34946 19487 34962 sw
rect 19394 34880 19487 34946
rect 19523 34821 19637 34979
tri 19673 34946 19689 34962 se
rect 19689 34946 19766 34962
rect 19673 34880 19766 34946
rect 19394 34745 19766 34821
rect 19394 34620 19487 34686
rect 19394 34604 19471 34620
tri 19471 34604 19487 34620 nw
rect 19523 34587 19637 34745
rect 19673 34620 19766 34686
tri 19673 34604 19689 34620 ne
rect 19689 34604 19766 34620
rect 19506 34505 19654 34587
rect 19394 34472 19471 34488
tri 19471 34472 19487 34488 sw
rect 19394 34406 19487 34472
rect 19394 34304 19487 34370
rect 19394 34288 19471 34304
tri 19471 34288 19487 34304 nw
rect 19523 34271 19637 34505
tri 19673 34472 19689 34488 se
rect 19689 34472 19766 34488
rect 19673 34406 19766 34472
rect 19673 34304 19766 34370
tri 19673 34288 19689 34304 ne
rect 19689 34288 19766 34304
rect 19506 34189 19654 34271
rect 19394 34156 19471 34172
tri 19471 34156 19487 34172 sw
rect 19394 34090 19487 34156
rect 19523 34031 19637 34189
tri 19673 34156 19689 34172 se
rect 19689 34156 19766 34172
rect 19673 34090 19766 34156
rect 19394 33955 19766 34031
rect 19394 33830 19487 33896
rect 19394 33814 19471 33830
tri 19471 33814 19487 33830 nw
rect 19523 33797 19637 33955
rect 19673 33830 19766 33896
tri 19673 33814 19689 33830 ne
rect 19689 33814 19766 33830
rect 19506 33715 19654 33797
rect 19394 33682 19471 33698
tri 19471 33682 19487 33698 sw
rect 19394 33616 19487 33682
rect 19394 33514 19487 33580
rect 19394 33498 19471 33514
tri 19471 33498 19487 33514 nw
rect 19523 33481 19637 33715
tri 19673 33682 19689 33698 se
rect 19689 33682 19766 33698
rect 19673 33616 19766 33682
rect 19673 33514 19766 33580
tri 19673 33498 19689 33514 ne
rect 19689 33498 19766 33514
rect 19506 33399 19654 33481
rect 19394 33366 19471 33382
tri 19471 33366 19487 33382 sw
rect 19394 33300 19487 33366
rect 19523 33241 19637 33399
tri 19673 33366 19689 33382 se
rect 19689 33366 19766 33382
rect 19673 33300 19766 33366
rect 19394 33165 19766 33241
rect 19394 33040 19487 33106
rect 19394 33024 19471 33040
tri 19471 33024 19487 33040 nw
rect 19523 33007 19637 33165
rect 19673 33040 19766 33106
tri 19673 33024 19689 33040 ne
rect 19689 33024 19766 33040
rect 19506 32925 19654 33007
rect 19394 32892 19471 32908
tri 19471 32892 19487 32908 sw
rect 19394 32826 19487 32892
rect 19394 32724 19487 32790
rect 19394 32708 19471 32724
tri 19471 32708 19487 32724 nw
rect 19523 32691 19637 32925
tri 19673 32892 19689 32908 se
rect 19689 32892 19766 32908
rect 19673 32826 19766 32892
rect 19673 32724 19766 32790
tri 19673 32708 19689 32724 ne
rect 19689 32708 19766 32724
rect 19506 32609 19654 32691
rect 19394 32576 19471 32592
tri 19471 32576 19487 32592 sw
rect 19394 32510 19487 32576
rect 19523 32451 19637 32609
tri 19673 32576 19689 32592 se
rect 19689 32576 19766 32592
rect 19673 32510 19766 32576
rect 19394 32375 19766 32451
rect 19394 32250 19487 32316
rect 19394 32234 19471 32250
tri 19471 32234 19487 32250 nw
rect 19523 32217 19637 32375
rect 19673 32250 19766 32316
tri 19673 32234 19689 32250 ne
rect 19689 32234 19766 32250
rect 19506 32135 19654 32217
rect 19394 32102 19471 32118
tri 19471 32102 19487 32118 sw
rect 19394 32036 19487 32102
rect 19394 31934 19487 32000
rect 19394 31918 19471 31934
tri 19471 31918 19487 31934 nw
rect 19523 31901 19637 32135
tri 19673 32102 19689 32118 se
rect 19689 32102 19766 32118
rect 19673 32036 19766 32102
rect 19673 31934 19766 32000
tri 19673 31918 19689 31934 ne
rect 19689 31918 19766 31934
rect 19506 31819 19654 31901
rect 19394 31786 19471 31802
tri 19471 31786 19487 31802 sw
rect 19394 31720 19487 31786
rect 19523 31661 19637 31819
tri 19673 31786 19689 31802 se
rect 19689 31786 19766 31802
rect 19673 31720 19766 31786
rect 19394 31585 19766 31661
rect 19394 31460 19487 31526
rect 19394 31444 19471 31460
tri 19471 31444 19487 31460 nw
rect 19523 31427 19637 31585
rect 19673 31460 19766 31526
tri 19673 31444 19689 31460 ne
rect 19689 31444 19766 31460
rect 19506 31345 19654 31427
rect 19394 31312 19471 31328
tri 19471 31312 19487 31328 sw
rect 19394 31246 19487 31312
rect 19394 31144 19487 31210
rect 19394 31128 19471 31144
tri 19471 31128 19487 31144 nw
rect 19523 31111 19637 31345
tri 19673 31312 19689 31328 se
rect 19689 31312 19766 31328
rect 19673 31246 19766 31312
rect 19673 31144 19766 31210
tri 19673 31128 19689 31144 ne
rect 19689 31128 19766 31144
rect 19506 31029 19654 31111
rect 19394 30996 19471 31012
tri 19471 30996 19487 31012 sw
rect 19394 30930 19487 30996
rect 19523 30871 19637 31029
tri 19673 30996 19689 31012 se
rect 19689 30996 19766 31012
rect 19673 30930 19766 30996
rect 19394 30795 19766 30871
rect 19394 30670 19487 30736
rect 19394 30654 19471 30670
tri 19471 30654 19487 30670 nw
rect 19523 30637 19637 30795
rect 19673 30670 19766 30736
tri 19673 30654 19689 30670 ne
rect 19689 30654 19766 30670
rect 19506 30555 19654 30637
rect 19394 30522 19471 30538
tri 19471 30522 19487 30538 sw
rect 19394 30456 19487 30522
rect 19394 30354 19487 30420
rect 19394 30338 19471 30354
tri 19471 30338 19487 30354 nw
rect 19523 30321 19637 30555
tri 19673 30522 19689 30538 se
rect 19689 30522 19766 30538
rect 19673 30456 19766 30522
rect 19673 30354 19766 30420
tri 19673 30338 19689 30354 ne
rect 19689 30338 19766 30354
rect 19506 30239 19654 30321
rect 19394 30206 19471 30222
tri 19471 30206 19487 30222 sw
rect 19394 30140 19487 30206
rect 19523 30081 19637 30239
tri 19673 30206 19689 30222 se
rect 19689 30206 19766 30222
rect 19673 30140 19766 30206
rect 19394 30005 19766 30081
rect 19394 29880 19487 29946
rect 19394 29864 19471 29880
tri 19471 29864 19487 29880 nw
rect 19523 29847 19637 30005
rect 19673 29880 19766 29946
tri 19673 29864 19689 29880 ne
rect 19689 29864 19766 29880
rect 19506 29765 19654 29847
rect 19394 29732 19471 29748
tri 19471 29732 19487 29748 sw
rect 19394 29666 19487 29732
rect 19394 29564 19487 29630
rect 19394 29548 19471 29564
tri 19471 29548 19487 29564 nw
rect 19523 29531 19637 29765
tri 19673 29732 19689 29748 se
rect 19689 29732 19766 29748
rect 19673 29666 19766 29732
rect 19673 29564 19766 29630
tri 19673 29548 19689 29564 ne
rect 19689 29548 19766 29564
rect 19506 29449 19654 29531
rect 19394 29416 19471 29432
tri 19471 29416 19487 29432 sw
rect 19394 29350 19487 29416
rect 19523 29291 19637 29449
tri 19673 29416 19689 29432 se
rect 19689 29416 19766 29432
rect 19673 29350 19766 29416
rect 19394 29215 19766 29291
rect 19394 29090 19487 29156
rect 19394 29074 19471 29090
tri 19471 29074 19487 29090 nw
rect 19523 29057 19637 29215
rect 19673 29090 19766 29156
tri 19673 29074 19689 29090 ne
rect 19689 29074 19766 29090
rect 19506 28975 19654 29057
rect 19394 28942 19471 28958
tri 19471 28942 19487 28958 sw
rect 19394 28876 19487 28942
rect 19523 28833 19637 28975
tri 19673 28942 19689 28958 se
rect 19689 28942 19766 28958
rect 19673 28876 19766 28942
rect 19802 28463 19838 80603
rect 19874 28463 19910 80603
rect 19946 80445 19982 80603
rect 19938 80303 19990 80445
rect 19946 28763 19982 80303
rect 19938 28621 19990 28763
rect 19946 28463 19982 28621
rect 20018 28463 20054 80603
rect 20090 28463 20126 80603
rect 20162 28833 20246 80233
rect 20282 28463 20318 80603
rect 20354 28463 20390 80603
rect 20426 80445 20462 80603
rect 20418 80303 20470 80445
rect 20426 28763 20462 80303
rect 20418 28621 20470 28763
rect 20426 28463 20462 28621
rect 20498 28463 20534 80603
rect 20570 28463 20606 80603
rect 20642 80124 20735 80190
rect 20642 80108 20719 80124
tri 20719 80108 20735 80124 nw
rect 20771 80091 20885 80233
rect 20921 80124 21014 80190
tri 20921 80108 20937 80124 ne
rect 20937 80108 21014 80124
rect 20754 80009 20902 80091
rect 20642 79976 20719 79992
tri 20719 79976 20735 79992 sw
rect 20642 79910 20735 79976
rect 20771 79851 20885 80009
tri 20921 79976 20937 79992 se
rect 20937 79976 21014 79992
rect 20921 79910 21014 79976
rect 20642 79775 21014 79851
rect 20642 79650 20735 79716
rect 20642 79634 20719 79650
tri 20719 79634 20735 79650 nw
rect 20771 79617 20885 79775
rect 20921 79650 21014 79716
tri 20921 79634 20937 79650 ne
rect 20937 79634 21014 79650
rect 20754 79535 20902 79617
rect 20642 79502 20719 79518
tri 20719 79502 20735 79518 sw
rect 20642 79436 20735 79502
rect 20642 79334 20735 79400
rect 20642 79318 20719 79334
tri 20719 79318 20735 79334 nw
rect 20771 79301 20885 79535
tri 20921 79502 20937 79518 se
rect 20937 79502 21014 79518
rect 20921 79436 21014 79502
rect 20921 79334 21014 79400
tri 20921 79318 20937 79334 ne
rect 20937 79318 21014 79334
rect 20754 79219 20902 79301
rect 20642 79186 20719 79202
tri 20719 79186 20735 79202 sw
rect 20642 79120 20735 79186
rect 20771 79061 20885 79219
tri 20921 79186 20937 79202 se
rect 20937 79186 21014 79202
rect 20921 79120 21014 79186
rect 20642 78985 21014 79061
rect 20642 78860 20735 78926
rect 20642 78844 20719 78860
tri 20719 78844 20735 78860 nw
rect 20771 78827 20885 78985
rect 20921 78860 21014 78926
tri 20921 78844 20937 78860 ne
rect 20937 78844 21014 78860
rect 20754 78745 20902 78827
rect 20642 78712 20719 78728
tri 20719 78712 20735 78728 sw
rect 20642 78646 20735 78712
rect 20642 78544 20735 78610
rect 20642 78528 20719 78544
tri 20719 78528 20735 78544 nw
rect 20771 78511 20885 78745
tri 20921 78712 20937 78728 se
rect 20937 78712 21014 78728
rect 20921 78646 21014 78712
rect 20921 78544 21014 78610
tri 20921 78528 20937 78544 ne
rect 20937 78528 21014 78544
rect 20754 78429 20902 78511
rect 20642 78396 20719 78412
tri 20719 78396 20735 78412 sw
rect 20642 78330 20735 78396
rect 20771 78271 20885 78429
tri 20921 78396 20937 78412 se
rect 20937 78396 21014 78412
rect 20921 78330 21014 78396
rect 20642 78195 21014 78271
rect 20642 78070 20735 78136
rect 20642 78054 20719 78070
tri 20719 78054 20735 78070 nw
rect 20771 78037 20885 78195
rect 20921 78070 21014 78136
tri 20921 78054 20937 78070 ne
rect 20937 78054 21014 78070
rect 20754 77955 20902 78037
rect 20642 77922 20719 77938
tri 20719 77922 20735 77938 sw
rect 20642 77856 20735 77922
rect 20642 77754 20735 77820
rect 20642 77738 20719 77754
tri 20719 77738 20735 77754 nw
rect 20771 77721 20885 77955
tri 20921 77922 20937 77938 se
rect 20937 77922 21014 77938
rect 20921 77856 21014 77922
rect 20921 77754 21014 77820
tri 20921 77738 20937 77754 ne
rect 20937 77738 21014 77754
rect 20754 77639 20902 77721
rect 20642 77606 20719 77622
tri 20719 77606 20735 77622 sw
rect 20642 77540 20735 77606
rect 20771 77481 20885 77639
tri 20921 77606 20937 77622 se
rect 20937 77606 21014 77622
rect 20921 77540 21014 77606
rect 20642 77405 21014 77481
rect 20642 77280 20735 77346
rect 20642 77264 20719 77280
tri 20719 77264 20735 77280 nw
rect 20771 77247 20885 77405
rect 20921 77280 21014 77346
tri 20921 77264 20937 77280 ne
rect 20937 77264 21014 77280
rect 20754 77165 20902 77247
rect 20642 77132 20719 77148
tri 20719 77132 20735 77148 sw
rect 20642 77066 20735 77132
rect 20642 76964 20735 77030
rect 20642 76948 20719 76964
tri 20719 76948 20735 76964 nw
rect 20771 76931 20885 77165
tri 20921 77132 20937 77148 se
rect 20937 77132 21014 77148
rect 20921 77066 21014 77132
rect 20921 76964 21014 77030
tri 20921 76948 20937 76964 ne
rect 20937 76948 21014 76964
rect 20754 76849 20902 76931
rect 20642 76816 20719 76832
tri 20719 76816 20735 76832 sw
rect 20642 76750 20735 76816
rect 20771 76691 20885 76849
tri 20921 76816 20937 76832 se
rect 20937 76816 21014 76832
rect 20921 76750 21014 76816
rect 20642 76615 21014 76691
rect 20642 76490 20735 76556
rect 20642 76474 20719 76490
tri 20719 76474 20735 76490 nw
rect 20771 76457 20885 76615
rect 20921 76490 21014 76556
tri 20921 76474 20937 76490 ne
rect 20937 76474 21014 76490
rect 20754 76375 20902 76457
rect 20642 76342 20719 76358
tri 20719 76342 20735 76358 sw
rect 20642 76276 20735 76342
rect 20642 76174 20735 76240
rect 20642 76158 20719 76174
tri 20719 76158 20735 76174 nw
rect 20771 76141 20885 76375
tri 20921 76342 20937 76358 se
rect 20937 76342 21014 76358
rect 20921 76276 21014 76342
rect 20921 76174 21014 76240
tri 20921 76158 20937 76174 ne
rect 20937 76158 21014 76174
rect 20754 76059 20902 76141
rect 20642 76026 20719 76042
tri 20719 76026 20735 76042 sw
rect 20642 75960 20735 76026
rect 20771 75901 20885 76059
tri 20921 76026 20937 76042 se
rect 20937 76026 21014 76042
rect 20921 75960 21014 76026
rect 20642 75825 21014 75901
rect 20642 75700 20735 75766
rect 20642 75684 20719 75700
tri 20719 75684 20735 75700 nw
rect 20771 75667 20885 75825
rect 20921 75700 21014 75766
tri 20921 75684 20937 75700 ne
rect 20937 75684 21014 75700
rect 20754 75585 20902 75667
rect 20642 75552 20719 75568
tri 20719 75552 20735 75568 sw
rect 20642 75486 20735 75552
rect 20642 75384 20735 75450
rect 20642 75368 20719 75384
tri 20719 75368 20735 75384 nw
rect 20771 75351 20885 75585
tri 20921 75552 20937 75568 se
rect 20937 75552 21014 75568
rect 20921 75486 21014 75552
rect 20921 75384 21014 75450
tri 20921 75368 20937 75384 ne
rect 20937 75368 21014 75384
rect 20754 75269 20902 75351
rect 20642 75236 20719 75252
tri 20719 75236 20735 75252 sw
rect 20642 75170 20735 75236
rect 20771 75111 20885 75269
tri 20921 75236 20937 75252 se
rect 20937 75236 21014 75252
rect 20921 75170 21014 75236
rect 20642 75035 21014 75111
rect 20642 74910 20735 74976
rect 20642 74894 20719 74910
tri 20719 74894 20735 74910 nw
rect 20771 74877 20885 75035
rect 20921 74910 21014 74976
tri 20921 74894 20937 74910 ne
rect 20937 74894 21014 74910
rect 20754 74795 20902 74877
rect 20642 74762 20719 74778
tri 20719 74762 20735 74778 sw
rect 20642 74696 20735 74762
rect 20642 74594 20735 74660
rect 20642 74578 20719 74594
tri 20719 74578 20735 74594 nw
rect 20771 74561 20885 74795
tri 20921 74762 20937 74778 se
rect 20937 74762 21014 74778
rect 20921 74696 21014 74762
rect 20921 74594 21014 74660
tri 20921 74578 20937 74594 ne
rect 20937 74578 21014 74594
rect 20754 74479 20902 74561
rect 20642 74446 20719 74462
tri 20719 74446 20735 74462 sw
rect 20642 74380 20735 74446
rect 20771 74321 20885 74479
tri 20921 74446 20937 74462 se
rect 20937 74446 21014 74462
rect 20921 74380 21014 74446
rect 20642 74245 21014 74321
rect 20642 74120 20735 74186
rect 20642 74104 20719 74120
tri 20719 74104 20735 74120 nw
rect 20771 74087 20885 74245
rect 20921 74120 21014 74186
tri 20921 74104 20937 74120 ne
rect 20937 74104 21014 74120
rect 20754 74005 20902 74087
rect 20642 73972 20719 73988
tri 20719 73972 20735 73988 sw
rect 20642 73906 20735 73972
rect 20642 73804 20735 73870
rect 20642 73788 20719 73804
tri 20719 73788 20735 73804 nw
rect 20771 73771 20885 74005
tri 20921 73972 20937 73988 se
rect 20937 73972 21014 73988
rect 20921 73906 21014 73972
rect 20921 73804 21014 73870
tri 20921 73788 20937 73804 ne
rect 20937 73788 21014 73804
rect 20754 73689 20902 73771
rect 20642 73656 20719 73672
tri 20719 73656 20735 73672 sw
rect 20642 73590 20735 73656
rect 20771 73531 20885 73689
tri 20921 73656 20937 73672 se
rect 20937 73656 21014 73672
rect 20921 73590 21014 73656
rect 20642 73455 21014 73531
rect 20642 73330 20735 73396
rect 20642 73314 20719 73330
tri 20719 73314 20735 73330 nw
rect 20771 73297 20885 73455
rect 20921 73330 21014 73396
tri 20921 73314 20937 73330 ne
rect 20937 73314 21014 73330
rect 20754 73215 20902 73297
rect 20642 73182 20719 73198
tri 20719 73182 20735 73198 sw
rect 20642 73116 20735 73182
rect 20642 73014 20735 73080
rect 20642 72998 20719 73014
tri 20719 72998 20735 73014 nw
rect 20771 72981 20885 73215
tri 20921 73182 20937 73198 se
rect 20937 73182 21014 73198
rect 20921 73116 21014 73182
rect 20921 73014 21014 73080
tri 20921 72998 20937 73014 ne
rect 20937 72998 21014 73014
rect 20754 72899 20902 72981
rect 20642 72866 20719 72882
tri 20719 72866 20735 72882 sw
rect 20642 72800 20735 72866
rect 20771 72741 20885 72899
tri 20921 72866 20937 72882 se
rect 20937 72866 21014 72882
rect 20921 72800 21014 72866
rect 20642 72665 21014 72741
rect 20642 72540 20735 72606
rect 20642 72524 20719 72540
tri 20719 72524 20735 72540 nw
rect 20771 72507 20885 72665
rect 20921 72540 21014 72606
tri 20921 72524 20937 72540 ne
rect 20937 72524 21014 72540
rect 20754 72425 20902 72507
rect 20642 72392 20719 72408
tri 20719 72392 20735 72408 sw
rect 20642 72326 20735 72392
rect 20642 72224 20735 72290
rect 20642 72208 20719 72224
tri 20719 72208 20735 72224 nw
rect 20771 72191 20885 72425
tri 20921 72392 20937 72408 se
rect 20937 72392 21014 72408
rect 20921 72326 21014 72392
rect 20921 72224 21014 72290
tri 20921 72208 20937 72224 ne
rect 20937 72208 21014 72224
rect 20754 72109 20902 72191
rect 20642 72076 20719 72092
tri 20719 72076 20735 72092 sw
rect 20642 72010 20735 72076
rect 20771 71951 20885 72109
tri 20921 72076 20937 72092 se
rect 20937 72076 21014 72092
rect 20921 72010 21014 72076
rect 20642 71875 21014 71951
rect 20642 71750 20735 71816
rect 20642 71734 20719 71750
tri 20719 71734 20735 71750 nw
rect 20771 71717 20885 71875
rect 20921 71750 21014 71816
tri 20921 71734 20937 71750 ne
rect 20937 71734 21014 71750
rect 20754 71635 20902 71717
rect 20642 71602 20719 71618
tri 20719 71602 20735 71618 sw
rect 20642 71536 20735 71602
rect 20642 71434 20735 71500
rect 20642 71418 20719 71434
tri 20719 71418 20735 71434 nw
rect 20771 71401 20885 71635
tri 20921 71602 20937 71618 se
rect 20937 71602 21014 71618
rect 20921 71536 21014 71602
rect 20921 71434 21014 71500
tri 20921 71418 20937 71434 ne
rect 20937 71418 21014 71434
rect 20754 71319 20902 71401
rect 20642 71286 20719 71302
tri 20719 71286 20735 71302 sw
rect 20642 71220 20735 71286
rect 20771 71161 20885 71319
tri 20921 71286 20937 71302 se
rect 20937 71286 21014 71302
rect 20921 71220 21014 71286
rect 20642 71085 21014 71161
rect 20642 70960 20735 71026
rect 20642 70944 20719 70960
tri 20719 70944 20735 70960 nw
rect 20771 70927 20885 71085
rect 20921 70960 21014 71026
tri 20921 70944 20937 70960 ne
rect 20937 70944 21014 70960
rect 20754 70845 20902 70927
rect 20642 70812 20719 70828
tri 20719 70812 20735 70828 sw
rect 20642 70746 20735 70812
rect 20642 70644 20735 70710
rect 20642 70628 20719 70644
tri 20719 70628 20735 70644 nw
rect 20771 70611 20885 70845
tri 20921 70812 20937 70828 se
rect 20937 70812 21014 70828
rect 20921 70746 21014 70812
rect 20921 70644 21014 70710
tri 20921 70628 20937 70644 ne
rect 20937 70628 21014 70644
rect 20754 70529 20902 70611
rect 20642 70496 20719 70512
tri 20719 70496 20735 70512 sw
rect 20642 70430 20735 70496
rect 20771 70371 20885 70529
tri 20921 70496 20937 70512 se
rect 20937 70496 21014 70512
rect 20921 70430 21014 70496
rect 20642 70295 21014 70371
rect 20642 70170 20735 70236
rect 20642 70154 20719 70170
tri 20719 70154 20735 70170 nw
rect 20771 70137 20885 70295
rect 20921 70170 21014 70236
tri 20921 70154 20937 70170 ne
rect 20937 70154 21014 70170
rect 20754 70055 20902 70137
rect 20642 70022 20719 70038
tri 20719 70022 20735 70038 sw
rect 20642 69956 20735 70022
rect 20642 69854 20735 69920
rect 20642 69838 20719 69854
tri 20719 69838 20735 69854 nw
rect 20771 69821 20885 70055
tri 20921 70022 20937 70038 se
rect 20937 70022 21014 70038
rect 20921 69956 21014 70022
rect 20921 69854 21014 69920
tri 20921 69838 20937 69854 ne
rect 20937 69838 21014 69854
rect 20754 69739 20902 69821
rect 20642 69706 20719 69722
tri 20719 69706 20735 69722 sw
rect 20642 69640 20735 69706
rect 20771 69581 20885 69739
tri 20921 69706 20937 69722 se
rect 20937 69706 21014 69722
rect 20921 69640 21014 69706
rect 20642 69505 21014 69581
rect 20642 69380 20735 69446
rect 20642 69364 20719 69380
tri 20719 69364 20735 69380 nw
rect 20771 69347 20885 69505
rect 20921 69380 21014 69446
tri 20921 69364 20937 69380 ne
rect 20937 69364 21014 69380
rect 20754 69265 20902 69347
rect 20642 69232 20719 69248
tri 20719 69232 20735 69248 sw
rect 20642 69166 20735 69232
rect 20642 69064 20735 69130
rect 20642 69048 20719 69064
tri 20719 69048 20735 69064 nw
rect 20771 69031 20885 69265
tri 20921 69232 20937 69248 se
rect 20937 69232 21014 69248
rect 20921 69166 21014 69232
rect 20921 69064 21014 69130
tri 20921 69048 20937 69064 ne
rect 20937 69048 21014 69064
rect 20754 68949 20902 69031
rect 20642 68916 20719 68932
tri 20719 68916 20735 68932 sw
rect 20642 68850 20735 68916
rect 20771 68791 20885 68949
tri 20921 68916 20937 68932 se
rect 20937 68916 21014 68932
rect 20921 68850 21014 68916
rect 20642 68715 21014 68791
rect 20642 68590 20735 68656
rect 20642 68574 20719 68590
tri 20719 68574 20735 68590 nw
rect 20771 68557 20885 68715
rect 20921 68590 21014 68656
tri 20921 68574 20937 68590 ne
rect 20937 68574 21014 68590
rect 20754 68475 20902 68557
rect 20642 68442 20719 68458
tri 20719 68442 20735 68458 sw
rect 20642 68376 20735 68442
rect 20642 68274 20735 68340
rect 20642 68258 20719 68274
tri 20719 68258 20735 68274 nw
rect 20771 68241 20885 68475
tri 20921 68442 20937 68458 se
rect 20937 68442 21014 68458
rect 20921 68376 21014 68442
rect 20921 68274 21014 68340
tri 20921 68258 20937 68274 ne
rect 20937 68258 21014 68274
rect 20754 68159 20902 68241
rect 20642 68126 20719 68142
tri 20719 68126 20735 68142 sw
rect 20642 68060 20735 68126
rect 20771 68001 20885 68159
tri 20921 68126 20937 68142 se
rect 20937 68126 21014 68142
rect 20921 68060 21014 68126
rect 20642 67925 21014 68001
rect 20642 67800 20735 67866
rect 20642 67784 20719 67800
tri 20719 67784 20735 67800 nw
rect 20771 67767 20885 67925
rect 20921 67800 21014 67866
tri 20921 67784 20937 67800 ne
rect 20937 67784 21014 67800
rect 20754 67685 20902 67767
rect 20642 67652 20719 67668
tri 20719 67652 20735 67668 sw
rect 20642 67586 20735 67652
rect 20642 67484 20735 67550
rect 20642 67468 20719 67484
tri 20719 67468 20735 67484 nw
rect 20771 67451 20885 67685
tri 20921 67652 20937 67668 se
rect 20937 67652 21014 67668
rect 20921 67586 21014 67652
rect 20921 67484 21014 67550
tri 20921 67468 20937 67484 ne
rect 20937 67468 21014 67484
rect 20754 67369 20902 67451
rect 20642 67336 20719 67352
tri 20719 67336 20735 67352 sw
rect 20642 67270 20735 67336
rect 20771 67211 20885 67369
tri 20921 67336 20937 67352 se
rect 20937 67336 21014 67352
rect 20921 67270 21014 67336
rect 20642 67135 21014 67211
rect 20642 67010 20735 67076
rect 20642 66994 20719 67010
tri 20719 66994 20735 67010 nw
rect 20771 66977 20885 67135
rect 20921 67010 21014 67076
tri 20921 66994 20937 67010 ne
rect 20937 66994 21014 67010
rect 20754 66895 20902 66977
rect 20642 66862 20719 66878
tri 20719 66862 20735 66878 sw
rect 20642 66796 20735 66862
rect 20642 66694 20735 66760
rect 20642 66678 20719 66694
tri 20719 66678 20735 66694 nw
rect 20771 66661 20885 66895
tri 20921 66862 20937 66878 se
rect 20937 66862 21014 66878
rect 20921 66796 21014 66862
rect 20921 66694 21014 66760
tri 20921 66678 20937 66694 ne
rect 20937 66678 21014 66694
rect 20754 66579 20902 66661
rect 20642 66546 20719 66562
tri 20719 66546 20735 66562 sw
rect 20642 66480 20735 66546
rect 20771 66421 20885 66579
tri 20921 66546 20937 66562 se
rect 20937 66546 21014 66562
rect 20921 66480 21014 66546
rect 20642 66345 21014 66421
rect 20642 66220 20735 66286
rect 20642 66204 20719 66220
tri 20719 66204 20735 66220 nw
rect 20771 66187 20885 66345
rect 20921 66220 21014 66286
tri 20921 66204 20937 66220 ne
rect 20937 66204 21014 66220
rect 20754 66105 20902 66187
rect 20642 66072 20719 66088
tri 20719 66072 20735 66088 sw
rect 20642 66006 20735 66072
rect 20642 65904 20735 65970
rect 20642 65888 20719 65904
tri 20719 65888 20735 65904 nw
rect 20771 65871 20885 66105
tri 20921 66072 20937 66088 se
rect 20937 66072 21014 66088
rect 20921 66006 21014 66072
rect 20921 65904 21014 65970
tri 20921 65888 20937 65904 ne
rect 20937 65888 21014 65904
rect 20754 65789 20902 65871
rect 20642 65756 20719 65772
tri 20719 65756 20735 65772 sw
rect 20642 65690 20735 65756
rect 20771 65631 20885 65789
tri 20921 65756 20937 65772 se
rect 20937 65756 21014 65772
rect 20921 65690 21014 65756
rect 20642 65555 21014 65631
rect 20642 65430 20735 65496
rect 20642 65414 20719 65430
tri 20719 65414 20735 65430 nw
rect 20771 65397 20885 65555
rect 20921 65430 21014 65496
tri 20921 65414 20937 65430 ne
rect 20937 65414 21014 65430
rect 20754 65315 20902 65397
rect 20642 65282 20719 65298
tri 20719 65282 20735 65298 sw
rect 20642 65216 20735 65282
rect 20642 65114 20735 65180
rect 20642 65098 20719 65114
tri 20719 65098 20735 65114 nw
rect 20771 65081 20885 65315
tri 20921 65282 20937 65298 se
rect 20937 65282 21014 65298
rect 20921 65216 21014 65282
rect 20921 65114 21014 65180
tri 20921 65098 20937 65114 ne
rect 20937 65098 21014 65114
rect 20754 64999 20902 65081
rect 20642 64966 20719 64982
tri 20719 64966 20735 64982 sw
rect 20642 64900 20735 64966
rect 20771 64841 20885 64999
tri 20921 64966 20937 64982 se
rect 20937 64966 21014 64982
rect 20921 64900 21014 64966
rect 20642 64765 21014 64841
rect 20642 64640 20735 64706
rect 20642 64624 20719 64640
tri 20719 64624 20735 64640 nw
rect 20771 64607 20885 64765
rect 20921 64640 21014 64706
tri 20921 64624 20937 64640 ne
rect 20937 64624 21014 64640
rect 20754 64525 20902 64607
rect 20642 64492 20719 64508
tri 20719 64492 20735 64508 sw
rect 20642 64426 20735 64492
rect 20642 64324 20735 64390
rect 20642 64308 20719 64324
tri 20719 64308 20735 64324 nw
rect 20771 64291 20885 64525
tri 20921 64492 20937 64508 se
rect 20937 64492 21014 64508
rect 20921 64426 21014 64492
rect 20921 64324 21014 64390
tri 20921 64308 20937 64324 ne
rect 20937 64308 21014 64324
rect 20754 64209 20902 64291
rect 20642 64176 20719 64192
tri 20719 64176 20735 64192 sw
rect 20642 64110 20735 64176
rect 20771 64051 20885 64209
tri 20921 64176 20937 64192 se
rect 20937 64176 21014 64192
rect 20921 64110 21014 64176
rect 20642 63975 21014 64051
rect 20642 63850 20735 63916
rect 20642 63834 20719 63850
tri 20719 63834 20735 63850 nw
rect 20771 63817 20885 63975
rect 20921 63850 21014 63916
tri 20921 63834 20937 63850 ne
rect 20937 63834 21014 63850
rect 20754 63735 20902 63817
rect 20642 63702 20719 63718
tri 20719 63702 20735 63718 sw
rect 20642 63636 20735 63702
rect 20642 63534 20735 63600
rect 20642 63518 20719 63534
tri 20719 63518 20735 63534 nw
rect 20771 63501 20885 63735
tri 20921 63702 20937 63718 se
rect 20937 63702 21014 63718
rect 20921 63636 21014 63702
rect 20921 63534 21014 63600
tri 20921 63518 20937 63534 ne
rect 20937 63518 21014 63534
rect 20754 63419 20902 63501
rect 20642 63386 20719 63402
tri 20719 63386 20735 63402 sw
rect 20642 63320 20735 63386
rect 20771 63261 20885 63419
tri 20921 63386 20937 63402 se
rect 20937 63386 21014 63402
rect 20921 63320 21014 63386
rect 20642 63185 21014 63261
rect 20642 63060 20735 63126
rect 20642 63044 20719 63060
tri 20719 63044 20735 63060 nw
rect 20771 63027 20885 63185
rect 20921 63060 21014 63126
tri 20921 63044 20937 63060 ne
rect 20937 63044 21014 63060
rect 20754 62945 20902 63027
rect 20642 62912 20719 62928
tri 20719 62912 20735 62928 sw
rect 20642 62846 20735 62912
rect 20642 62744 20735 62810
rect 20642 62728 20719 62744
tri 20719 62728 20735 62744 nw
rect 20771 62711 20885 62945
tri 20921 62912 20937 62928 se
rect 20937 62912 21014 62928
rect 20921 62846 21014 62912
rect 20921 62744 21014 62810
tri 20921 62728 20937 62744 ne
rect 20937 62728 21014 62744
rect 20754 62629 20902 62711
rect 20642 62596 20719 62612
tri 20719 62596 20735 62612 sw
rect 20642 62530 20735 62596
rect 20771 62471 20885 62629
tri 20921 62596 20937 62612 se
rect 20937 62596 21014 62612
rect 20921 62530 21014 62596
rect 20642 62395 21014 62471
rect 20642 62270 20735 62336
rect 20642 62254 20719 62270
tri 20719 62254 20735 62270 nw
rect 20771 62237 20885 62395
rect 20921 62270 21014 62336
tri 20921 62254 20937 62270 ne
rect 20937 62254 21014 62270
rect 20754 62155 20902 62237
rect 20642 62122 20719 62138
tri 20719 62122 20735 62138 sw
rect 20642 62056 20735 62122
rect 20642 61954 20735 62020
rect 20642 61938 20719 61954
tri 20719 61938 20735 61954 nw
rect 20771 61921 20885 62155
tri 20921 62122 20937 62138 se
rect 20937 62122 21014 62138
rect 20921 62056 21014 62122
rect 20921 61954 21014 62020
tri 20921 61938 20937 61954 ne
rect 20937 61938 21014 61954
rect 20754 61839 20902 61921
rect 20642 61806 20719 61822
tri 20719 61806 20735 61822 sw
rect 20642 61740 20735 61806
rect 20771 61681 20885 61839
tri 20921 61806 20937 61822 se
rect 20937 61806 21014 61822
rect 20921 61740 21014 61806
rect 20642 61605 21014 61681
rect 20642 61480 20735 61546
rect 20642 61464 20719 61480
tri 20719 61464 20735 61480 nw
rect 20771 61447 20885 61605
rect 20921 61480 21014 61546
tri 20921 61464 20937 61480 ne
rect 20937 61464 21014 61480
rect 20754 61365 20902 61447
rect 20642 61332 20719 61348
tri 20719 61332 20735 61348 sw
rect 20642 61266 20735 61332
rect 20642 61164 20735 61230
rect 20642 61148 20719 61164
tri 20719 61148 20735 61164 nw
rect 20771 61131 20885 61365
tri 20921 61332 20937 61348 se
rect 20937 61332 21014 61348
rect 20921 61266 21014 61332
rect 20921 61164 21014 61230
tri 20921 61148 20937 61164 ne
rect 20937 61148 21014 61164
rect 20754 61049 20902 61131
rect 20642 61016 20719 61032
tri 20719 61016 20735 61032 sw
rect 20642 60950 20735 61016
rect 20771 60891 20885 61049
tri 20921 61016 20937 61032 se
rect 20937 61016 21014 61032
rect 20921 60950 21014 61016
rect 20642 60815 21014 60891
rect 20642 60690 20735 60756
rect 20642 60674 20719 60690
tri 20719 60674 20735 60690 nw
rect 20771 60657 20885 60815
rect 20921 60690 21014 60756
tri 20921 60674 20937 60690 ne
rect 20937 60674 21014 60690
rect 20754 60575 20902 60657
rect 20642 60542 20719 60558
tri 20719 60542 20735 60558 sw
rect 20642 60476 20735 60542
rect 20642 60374 20735 60440
rect 20642 60358 20719 60374
tri 20719 60358 20735 60374 nw
rect 20771 60341 20885 60575
tri 20921 60542 20937 60558 se
rect 20937 60542 21014 60558
rect 20921 60476 21014 60542
rect 20921 60374 21014 60440
tri 20921 60358 20937 60374 ne
rect 20937 60358 21014 60374
rect 20754 60259 20902 60341
rect 20642 60226 20719 60242
tri 20719 60226 20735 60242 sw
rect 20642 60160 20735 60226
rect 20771 60101 20885 60259
tri 20921 60226 20937 60242 se
rect 20937 60226 21014 60242
rect 20921 60160 21014 60226
rect 20642 60025 21014 60101
rect 20642 59900 20735 59966
rect 20642 59884 20719 59900
tri 20719 59884 20735 59900 nw
rect 20771 59867 20885 60025
rect 20921 59900 21014 59966
tri 20921 59884 20937 59900 ne
rect 20937 59884 21014 59900
rect 20754 59785 20902 59867
rect 20642 59752 20719 59768
tri 20719 59752 20735 59768 sw
rect 20642 59686 20735 59752
rect 20642 59584 20735 59650
rect 20642 59568 20719 59584
tri 20719 59568 20735 59584 nw
rect 20771 59551 20885 59785
tri 20921 59752 20937 59768 se
rect 20937 59752 21014 59768
rect 20921 59686 21014 59752
rect 20921 59584 21014 59650
tri 20921 59568 20937 59584 ne
rect 20937 59568 21014 59584
rect 20754 59469 20902 59551
rect 20642 59436 20719 59452
tri 20719 59436 20735 59452 sw
rect 20642 59370 20735 59436
rect 20771 59311 20885 59469
tri 20921 59436 20937 59452 se
rect 20937 59436 21014 59452
rect 20921 59370 21014 59436
rect 20642 59235 21014 59311
rect 20642 59110 20735 59176
rect 20642 59094 20719 59110
tri 20719 59094 20735 59110 nw
rect 20771 59077 20885 59235
rect 20921 59110 21014 59176
tri 20921 59094 20937 59110 ne
rect 20937 59094 21014 59110
rect 20754 58995 20902 59077
rect 20642 58962 20719 58978
tri 20719 58962 20735 58978 sw
rect 20642 58896 20735 58962
rect 20642 58794 20735 58860
rect 20642 58778 20719 58794
tri 20719 58778 20735 58794 nw
rect 20771 58761 20885 58995
tri 20921 58962 20937 58978 se
rect 20937 58962 21014 58978
rect 20921 58896 21014 58962
rect 20921 58794 21014 58860
tri 20921 58778 20937 58794 ne
rect 20937 58778 21014 58794
rect 20754 58679 20902 58761
rect 20642 58646 20719 58662
tri 20719 58646 20735 58662 sw
rect 20642 58580 20735 58646
rect 20771 58521 20885 58679
tri 20921 58646 20937 58662 se
rect 20937 58646 21014 58662
rect 20921 58580 21014 58646
rect 20642 58445 21014 58521
rect 20642 58320 20735 58386
rect 20642 58304 20719 58320
tri 20719 58304 20735 58320 nw
rect 20771 58287 20885 58445
rect 20921 58320 21014 58386
tri 20921 58304 20937 58320 ne
rect 20937 58304 21014 58320
rect 20754 58205 20902 58287
rect 20642 58172 20719 58188
tri 20719 58172 20735 58188 sw
rect 20642 58106 20735 58172
rect 20642 58004 20735 58070
rect 20642 57988 20719 58004
tri 20719 57988 20735 58004 nw
rect 20771 57971 20885 58205
tri 20921 58172 20937 58188 se
rect 20937 58172 21014 58188
rect 20921 58106 21014 58172
rect 20921 58004 21014 58070
tri 20921 57988 20937 58004 ne
rect 20937 57988 21014 58004
rect 20754 57889 20902 57971
rect 20642 57856 20719 57872
tri 20719 57856 20735 57872 sw
rect 20642 57790 20735 57856
rect 20771 57731 20885 57889
tri 20921 57856 20937 57872 se
rect 20937 57856 21014 57872
rect 20921 57790 21014 57856
rect 20642 57655 21014 57731
rect 20642 57530 20735 57596
rect 20642 57514 20719 57530
tri 20719 57514 20735 57530 nw
rect 20771 57497 20885 57655
rect 20921 57530 21014 57596
tri 20921 57514 20937 57530 ne
rect 20937 57514 21014 57530
rect 20754 57415 20902 57497
rect 20642 57382 20719 57398
tri 20719 57382 20735 57398 sw
rect 20642 57316 20735 57382
rect 20642 57214 20735 57280
rect 20642 57198 20719 57214
tri 20719 57198 20735 57214 nw
rect 20771 57181 20885 57415
tri 20921 57382 20937 57398 se
rect 20937 57382 21014 57398
rect 20921 57316 21014 57382
rect 20921 57214 21014 57280
tri 20921 57198 20937 57214 ne
rect 20937 57198 21014 57214
rect 20754 57099 20902 57181
rect 20642 57066 20719 57082
tri 20719 57066 20735 57082 sw
rect 20642 57000 20735 57066
rect 20771 56941 20885 57099
tri 20921 57066 20937 57082 se
rect 20937 57066 21014 57082
rect 20921 57000 21014 57066
rect 20642 56865 21014 56941
rect 20642 56740 20735 56806
rect 20642 56724 20719 56740
tri 20719 56724 20735 56740 nw
rect 20771 56707 20885 56865
rect 20921 56740 21014 56806
tri 20921 56724 20937 56740 ne
rect 20937 56724 21014 56740
rect 20754 56625 20902 56707
rect 20642 56592 20719 56608
tri 20719 56592 20735 56608 sw
rect 20642 56526 20735 56592
rect 20642 56424 20735 56490
rect 20642 56408 20719 56424
tri 20719 56408 20735 56424 nw
rect 20771 56391 20885 56625
tri 20921 56592 20937 56608 se
rect 20937 56592 21014 56608
rect 20921 56526 21014 56592
rect 20921 56424 21014 56490
tri 20921 56408 20937 56424 ne
rect 20937 56408 21014 56424
rect 20754 56309 20902 56391
rect 20642 56276 20719 56292
tri 20719 56276 20735 56292 sw
rect 20642 56210 20735 56276
rect 20771 56151 20885 56309
tri 20921 56276 20937 56292 se
rect 20937 56276 21014 56292
rect 20921 56210 21014 56276
rect 20642 56075 21014 56151
rect 20642 55950 20735 56016
rect 20642 55934 20719 55950
tri 20719 55934 20735 55950 nw
rect 20771 55917 20885 56075
rect 20921 55950 21014 56016
tri 20921 55934 20937 55950 ne
rect 20937 55934 21014 55950
rect 20754 55835 20902 55917
rect 20642 55802 20719 55818
tri 20719 55802 20735 55818 sw
rect 20642 55736 20735 55802
rect 20642 55634 20735 55700
rect 20642 55618 20719 55634
tri 20719 55618 20735 55634 nw
rect 20771 55601 20885 55835
tri 20921 55802 20937 55818 se
rect 20937 55802 21014 55818
rect 20921 55736 21014 55802
rect 20921 55634 21014 55700
tri 20921 55618 20937 55634 ne
rect 20937 55618 21014 55634
rect 20754 55519 20902 55601
rect 20642 55486 20719 55502
tri 20719 55486 20735 55502 sw
rect 20642 55420 20735 55486
rect 20771 55361 20885 55519
tri 20921 55486 20937 55502 se
rect 20937 55486 21014 55502
rect 20921 55420 21014 55486
rect 20642 55285 21014 55361
rect 20642 55160 20735 55226
rect 20642 55144 20719 55160
tri 20719 55144 20735 55160 nw
rect 20771 55127 20885 55285
rect 20921 55160 21014 55226
tri 20921 55144 20937 55160 ne
rect 20937 55144 21014 55160
rect 20754 55045 20902 55127
rect 20642 55012 20719 55028
tri 20719 55012 20735 55028 sw
rect 20642 54946 20735 55012
rect 20642 54844 20735 54910
rect 20642 54828 20719 54844
tri 20719 54828 20735 54844 nw
rect 20771 54811 20885 55045
tri 20921 55012 20937 55028 se
rect 20937 55012 21014 55028
rect 20921 54946 21014 55012
rect 20921 54844 21014 54910
tri 20921 54828 20937 54844 ne
rect 20937 54828 21014 54844
rect 20754 54729 20902 54811
rect 20642 54696 20719 54712
tri 20719 54696 20735 54712 sw
rect 20642 54630 20735 54696
rect 20771 54571 20885 54729
tri 20921 54696 20937 54712 se
rect 20937 54696 21014 54712
rect 20921 54630 21014 54696
rect 20642 54495 21014 54571
rect 20642 54370 20735 54436
rect 20642 54354 20719 54370
tri 20719 54354 20735 54370 nw
rect 20771 54337 20885 54495
rect 20921 54370 21014 54436
tri 20921 54354 20937 54370 ne
rect 20937 54354 21014 54370
rect 20754 54255 20902 54337
rect 20642 54222 20719 54238
tri 20719 54222 20735 54238 sw
rect 20642 54156 20735 54222
rect 20642 54054 20735 54120
rect 20642 54038 20719 54054
tri 20719 54038 20735 54054 nw
rect 20771 54021 20885 54255
tri 20921 54222 20937 54238 se
rect 20937 54222 21014 54238
rect 20921 54156 21014 54222
rect 20921 54054 21014 54120
tri 20921 54038 20937 54054 ne
rect 20937 54038 21014 54054
rect 20754 53939 20902 54021
rect 20642 53906 20719 53922
tri 20719 53906 20735 53922 sw
rect 20642 53840 20735 53906
rect 20771 53781 20885 53939
tri 20921 53906 20937 53922 se
rect 20937 53906 21014 53922
rect 20921 53840 21014 53906
rect 20642 53705 21014 53781
rect 20642 53580 20735 53646
rect 20642 53564 20719 53580
tri 20719 53564 20735 53580 nw
rect 20771 53547 20885 53705
rect 20921 53580 21014 53646
tri 20921 53564 20937 53580 ne
rect 20937 53564 21014 53580
rect 20754 53465 20902 53547
rect 20642 53432 20719 53448
tri 20719 53432 20735 53448 sw
rect 20642 53366 20735 53432
rect 20642 53264 20735 53330
rect 20642 53248 20719 53264
tri 20719 53248 20735 53264 nw
rect 20771 53231 20885 53465
tri 20921 53432 20937 53448 se
rect 20937 53432 21014 53448
rect 20921 53366 21014 53432
rect 20921 53264 21014 53330
tri 20921 53248 20937 53264 ne
rect 20937 53248 21014 53264
rect 20754 53149 20902 53231
rect 20642 53116 20719 53132
tri 20719 53116 20735 53132 sw
rect 20642 53050 20735 53116
rect 20771 52991 20885 53149
tri 20921 53116 20937 53132 se
rect 20937 53116 21014 53132
rect 20921 53050 21014 53116
rect 20642 52915 21014 52991
rect 20642 52790 20735 52856
rect 20642 52774 20719 52790
tri 20719 52774 20735 52790 nw
rect 20771 52757 20885 52915
rect 20921 52790 21014 52856
tri 20921 52774 20937 52790 ne
rect 20937 52774 21014 52790
rect 20754 52675 20902 52757
rect 20642 52642 20719 52658
tri 20719 52642 20735 52658 sw
rect 20642 52576 20735 52642
rect 20642 52474 20735 52540
rect 20642 52458 20719 52474
tri 20719 52458 20735 52474 nw
rect 20771 52441 20885 52675
tri 20921 52642 20937 52658 se
rect 20937 52642 21014 52658
rect 20921 52576 21014 52642
rect 20921 52474 21014 52540
tri 20921 52458 20937 52474 ne
rect 20937 52458 21014 52474
rect 20754 52359 20902 52441
rect 20642 52326 20719 52342
tri 20719 52326 20735 52342 sw
rect 20642 52260 20735 52326
rect 20771 52201 20885 52359
tri 20921 52326 20937 52342 se
rect 20937 52326 21014 52342
rect 20921 52260 21014 52326
rect 20642 52125 21014 52201
rect 20642 52000 20735 52066
rect 20642 51984 20719 52000
tri 20719 51984 20735 52000 nw
rect 20771 51967 20885 52125
rect 20921 52000 21014 52066
tri 20921 51984 20937 52000 ne
rect 20937 51984 21014 52000
rect 20754 51885 20902 51967
rect 20642 51852 20719 51868
tri 20719 51852 20735 51868 sw
rect 20642 51786 20735 51852
rect 20642 51684 20735 51750
rect 20642 51668 20719 51684
tri 20719 51668 20735 51684 nw
rect 20771 51651 20885 51885
tri 20921 51852 20937 51868 se
rect 20937 51852 21014 51868
rect 20921 51786 21014 51852
rect 20921 51684 21014 51750
tri 20921 51668 20937 51684 ne
rect 20937 51668 21014 51684
rect 20754 51569 20902 51651
rect 20642 51536 20719 51552
tri 20719 51536 20735 51552 sw
rect 20642 51470 20735 51536
rect 20771 51411 20885 51569
tri 20921 51536 20937 51552 se
rect 20937 51536 21014 51552
rect 20921 51470 21014 51536
rect 20642 51335 21014 51411
rect 20642 51210 20735 51276
rect 20642 51194 20719 51210
tri 20719 51194 20735 51210 nw
rect 20771 51177 20885 51335
rect 20921 51210 21014 51276
tri 20921 51194 20937 51210 ne
rect 20937 51194 21014 51210
rect 20754 51095 20902 51177
rect 20642 51062 20719 51078
tri 20719 51062 20735 51078 sw
rect 20642 50996 20735 51062
rect 20642 50894 20735 50960
rect 20642 50878 20719 50894
tri 20719 50878 20735 50894 nw
rect 20771 50861 20885 51095
tri 20921 51062 20937 51078 se
rect 20937 51062 21014 51078
rect 20921 50996 21014 51062
rect 20921 50894 21014 50960
tri 20921 50878 20937 50894 ne
rect 20937 50878 21014 50894
rect 20754 50779 20902 50861
rect 20642 50746 20719 50762
tri 20719 50746 20735 50762 sw
rect 20642 50680 20735 50746
rect 20771 50621 20885 50779
tri 20921 50746 20937 50762 se
rect 20937 50746 21014 50762
rect 20921 50680 21014 50746
rect 20642 50545 21014 50621
rect 20642 50420 20735 50486
rect 20642 50404 20719 50420
tri 20719 50404 20735 50420 nw
rect 20771 50387 20885 50545
rect 20921 50420 21014 50486
tri 20921 50404 20937 50420 ne
rect 20937 50404 21014 50420
rect 20754 50305 20902 50387
rect 20642 50272 20719 50288
tri 20719 50272 20735 50288 sw
rect 20642 50206 20735 50272
rect 20642 50104 20735 50170
rect 20642 50088 20719 50104
tri 20719 50088 20735 50104 nw
rect 20771 50071 20885 50305
tri 20921 50272 20937 50288 se
rect 20937 50272 21014 50288
rect 20921 50206 21014 50272
rect 20921 50104 21014 50170
tri 20921 50088 20937 50104 ne
rect 20937 50088 21014 50104
rect 20754 49989 20902 50071
rect 20642 49956 20719 49972
tri 20719 49956 20735 49972 sw
rect 20642 49890 20735 49956
rect 20771 49831 20885 49989
tri 20921 49956 20937 49972 se
rect 20937 49956 21014 49972
rect 20921 49890 21014 49956
rect 20642 49755 21014 49831
rect 20642 49630 20735 49696
rect 20642 49614 20719 49630
tri 20719 49614 20735 49630 nw
rect 20771 49597 20885 49755
rect 20921 49630 21014 49696
tri 20921 49614 20937 49630 ne
rect 20937 49614 21014 49630
rect 20754 49515 20902 49597
rect 20642 49482 20719 49498
tri 20719 49482 20735 49498 sw
rect 20642 49416 20735 49482
rect 20642 49314 20735 49380
rect 20642 49298 20719 49314
tri 20719 49298 20735 49314 nw
rect 20771 49281 20885 49515
tri 20921 49482 20937 49498 se
rect 20937 49482 21014 49498
rect 20921 49416 21014 49482
rect 20921 49314 21014 49380
tri 20921 49298 20937 49314 ne
rect 20937 49298 21014 49314
rect 20754 49199 20902 49281
rect 20642 49166 20719 49182
tri 20719 49166 20735 49182 sw
rect 20642 49100 20735 49166
rect 20771 49041 20885 49199
tri 20921 49166 20937 49182 se
rect 20937 49166 21014 49182
rect 20921 49100 21014 49166
rect 20642 48965 21014 49041
rect 20642 48840 20735 48906
rect 20642 48824 20719 48840
tri 20719 48824 20735 48840 nw
rect 20771 48807 20885 48965
rect 20921 48840 21014 48906
tri 20921 48824 20937 48840 ne
rect 20937 48824 21014 48840
rect 20754 48725 20902 48807
rect 20642 48692 20719 48708
tri 20719 48692 20735 48708 sw
rect 20642 48626 20735 48692
rect 20642 48524 20735 48590
rect 20642 48508 20719 48524
tri 20719 48508 20735 48524 nw
rect 20771 48491 20885 48725
tri 20921 48692 20937 48708 se
rect 20937 48692 21014 48708
rect 20921 48626 21014 48692
rect 20921 48524 21014 48590
tri 20921 48508 20937 48524 ne
rect 20937 48508 21014 48524
rect 20754 48409 20902 48491
rect 20642 48376 20719 48392
tri 20719 48376 20735 48392 sw
rect 20642 48310 20735 48376
rect 20771 48251 20885 48409
tri 20921 48376 20937 48392 se
rect 20937 48376 21014 48392
rect 20921 48310 21014 48376
rect 20642 48175 21014 48251
rect 20642 48050 20735 48116
rect 20642 48034 20719 48050
tri 20719 48034 20735 48050 nw
rect 20771 48017 20885 48175
rect 20921 48050 21014 48116
tri 20921 48034 20937 48050 ne
rect 20937 48034 21014 48050
rect 20754 47935 20902 48017
rect 20642 47902 20719 47918
tri 20719 47902 20735 47918 sw
rect 20642 47836 20735 47902
rect 20642 47734 20735 47800
rect 20642 47718 20719 47734
tri 20719 47718 20735 47734 nw
rect 20771 47701 20885 47935
tri 20921 47902 20937 47918 se
rect 20937 47902 21014 47918
rect 20921 47836 21014 47902
rect 20921 47734 21014 47800
tri 20921 47718 20937 47734 ne
rect 20937 47718 21014 47734
rect 20754 47619 20902 47701
rect 20642 47586 20719 47602
tri 20719 47586 20735 47602 sw
rect 20642 47520 20735 47586
rect 20771 47461 20885 47619
tri 20921 47586 20937 47602 se
rect 20937 47586 21014 47602
rect 20921 47520 21014 47586
rect 20642 47385 21014 47461
rect 20642 47260 20735 47326
rect 20642 47244 20719 47260
tri 20719 47244 20735 47260 nw
rect 20771 47227 20885 47385
rect 20921 47260 21014 47326
tri 20921 47244 20937 47260 ne
rect 20937 47244 21014 47260
rect 20754 47145 20902 47227
rect 20642 47112 20719 47128
tri 20719 47112 20735 47128 sw
rect 20642 47046 20735 47112
rect 20642 46944 20735 47010
rect 20642 46928 20719 46944
tri 20719 46928 20735 46944 nw
rect 20771 46911 20885 47145
tri 20921 47112 20937 47128 se
rect 20937 47112 21014 47128
rect 20921 47046 21014 47112
rect 20921 46944 21014 47010
tri 20921 46928 20937 46944 ne
rect 20937 46928 21014 46944
rect 20754 46829 20902 46911
rect 20642 46796 20719 46812
tri 20719 46796 20735 46812 sw
rect 20642 46730 20735 46796
rect 20771 46671 20885 46829
tri 20921 46796 20937 46812 se
rect 20937 46796 21014 46812
rect 20921 46730 21014 46796
rect 20642 46595 21014 46671
rect 20642 46470 20735 46536
rect 20642 46454 20719 46470
tri 20719 46454 20735 46470 nw
rect 20771 46437 20885 46595
rect 20921 46470 21014 46536
tri 20921 46454 20937 46470 ne
rect 20937 46454 21014 46470
rect 20754 46355 20902 46437
rect 20642 46322 20719 46338
tri 20719 46322 20735 46338 sw
rect 20642 46256 20735 46322
rect 20642 46154 20735 46220
rect 20642 46138 20719 46154
tri 20719 46138 20735 46154 nw
rect 20771 46121 20885 46355
tri 20921 46322 20937 46338 se
rect 20937 46322 21014 46338
rect 20921 46256 21014 46322
rect 20921 46154 21014 46220
tri 20921 46138 20937 46154 ne
rect 20937 46138 21014 46154
rect 20754 46039 20902 46121
rect 20642 46006 20719 46022
tri 20719 46006 20735 46022 sw
rect 20642 45940 20735 46006
rect 20771 45881 20885 46039
tri 20921 46006 20937 46022 se
rect 20937 46006 21014 46022
rect 20921 45940 21014 46006
rect 20642 45805 21014 45881
rect 20642 45680 20735 45746
rect 20642 45664 20719 45680
tri 20719 45664 20735 45680 nw
rect 20771 45647 20885 45805
rect 20921 45680 21014 45746
tri 20921 45664 20937 45680 ne
rect 20937 45664 21014 45680
rect 20754 45565 20902 45647
rect 20642 45532 20719 45548
tri 20719 45532 20735 45548 sw
rect 20642 45466 20735 45532
rect 20642 45364 20735 45430
rect 20642 45348 20719 45364
tri 20719 45348 20735 45364 nw
rect 20771 45331 20885 45565
tri 20921 45532 20937 45548 se
rect 20937 45532 21014 45548
rect 20921 45466 21014 45532
rect 20921 45364 21014 45430
tri 20921 45348 20937 45364 ne
rect 20937 45348 21014 45364
rect 20754 45249 20902 45331
rect 20642 45216 20719 45232
tri 20719 45216 20735 45232 sw
rect 20642 45150 20735 45216
rect 20771 45091 20885 45249
tri 20921 45216 20937 45232 se
rect 20937 45216 21014 45232
rect 20921 45150 21014 45216
rect 20642 45015 21014 45091
rect 20642 44890 20735 44956
rect 20642 44874 20719 44890
tri 20719 44874 20735 44890 nw
rect 20771 44857 20885 45015
rect 20921 44890 21014 44956
tri 20921 44874 20937 44890 ne
rect 20937 44874 21014 44890
rect 20754 44775 20902 44857
rect 20642 44742 20719 44758
tri 20719 44742 20735 44758 sw
rect 20642 44676 20735 44742
rect 20642 44574 20735 44640
rect 20642 44558 20719 44574
tri 20719 44558 20735 44574 nw
rect 20771 44541 20885 44775
tri 20921 44742 20937 44758 se
rect 20937 44742 21014 44758
rect 20921 44676 21014 44742
rect 20921 44574 21014 44640
tri 20921 44558 20937 44574 ne
rect 20937 44558 21014 44574
rect 20754 44459 20902 44541
rect 20642 44426 20719 44442
tri 20719 44426 20735 44442 sw
rect 20642 44360 20735 44426
rect 20771 44301 20885 44459
tri 20921 44426 20937 44442 se
rect 20937 44426 21014 44442
rect 20921 44360 21014 44426
rect 20642 44225 21014 44301
rect 20642 44100 20735 44166
rect 20642 44084 20719 44100
tri 20719 44084 20735 44100 nw
rect 20771 44067 20885 44225
rect 20921 44100 21014 44166
tri 20921 44084 20937 44100 ne
rect 20937 44084 21014 44100
rect 20754 43985 20902 44067
rect 20642 43952 20719 43968
tri 20719 43952 20735 43968 sw
rect 20642 43886 20735 43952
rect 20642 43784 20735 43850
rect 20642 43768 20719 43784
tri 20719 43768 20735 43784 nw
rect 20771 43751 20885 43985
tri 20921 43952 20937 43968 se
rect 20937 43952 21014 43968
rect 20921 43886 21014 43952
rect 20921 43784 21014 43850
tri 20921 43768 20937 43784 ne
rect 20937 43768 21014 43784
rect 20754 43669 20902 43751
rect 20642 43636 20719 43652
tri 20719 43636 20735 43652 sw
rect 20642 43570 20735 43636
rect 20771 43511 20885 43669
tri 20921 43636 20937 43652 se
rect 20937 43636 21014 43652
rect 20921 43570 21014 43636
rect 20642 43435 21014 43511
rect 20642 43310 20735 43376
rect 20642 43294 20719 43310
tri 20719 43294 20735 43310 nw
rect 20771 43277 20885 43435
rect 20921 43310 21014 43376
tri 20921 43294 20937 43310 ne
rect 20937 43294 21014 43310
rect 20754 43195 20902 43277
rect 20642 43162 20719 43178
tri 20719 43162 20735 43178 sw
rect 20642 43096 20735 43162
rect 20642 42994 20735 43060
rect 20642 42978 20719 42994
tri 20719 42978 20735 42994 nw
rect 20771 42961 20885 43195
tri 20921 43162 20937 43178 se
rect 20937 43162 21014 43178
rect 20921 43096 21014 43162
rect 20921 42994 21014 43060
tri 20921 42978 20937 42994 ne
rect 20937 42978 21014 42994
rect 20754 42879 20902 42961
rect 20642 42846 20719 42862
tri 20719 42846 20735 42862 sw
rect 20642 42780 20735 42846
rect 20771 42721 20885 42879
tri 20921 42846 20937 42862 se
rect 20937 42846 21014 42862
rect 20921 42780 21014 42846
rect 20642 42645 21014 42721
rect 20642 42520 20735 42586
rect 20642 42504 20719 42520
tri 20719 42504 20735 42520 nw
rect 20771 42487 20885 42645
rect 20921 42520 21014 42586
tri 20921 42504 20937 42520 ne
rect 20937 42504 21014 42520
rect 20754 42405 20902 42487
rect 20642 42372 20719 42388
tri 20719 42372 20735 42388 sw
rect 20642 42306 20735 42372
rect 20642 42204 20735 42270
rect 20642 42188 20719 42204
tri 20719 42188 20735 42204 nw
rect 20771 42171 20885 42405
tri 20921 42372 20937 42388 se
rect 20937 42372 21014 42388
rect 20921 42306 21014 42372
rect 20921 42204 21014 42270
tri 20921 42188 20937 42204 ne
rect 20937 42188 21014 42204
rect 20754 42089 20902 42171
rect 20642 42056 20719 42072
tri 20719 42056 20735 42072 sw
rect 20642 41990 20735 42056
rect 20771 41931 20885 42089
tri 20921 42056 20937 42072 se
rect 20937 42056 21014 42072
rect 20921 41990 21014 42056
rect 20642 41855 21014 41931
rect 20642 41730 20735 41796
rect 20642 41714 20719 41730
tri 20719 41714 20735 41730 nw
rect 20771 41697 20885 41855
rect 20921 41730 21014 41796
tri 20921 41714 20937 41730 ne
rect 20937 41714 21014 41730
rect 20754 41615 20902 41697
rect 20642 41582 20719 41598
tri 20719 41582 20735 41598 sw
rect 20642 41516 20735 41582
rect 20642 41414 20735 41480
rect 20642 41398 20719 41414
tri 20719 41398 20735 41414 nw
rect 20771 41381 20885 41615
tri 20921 41582 20937 41598 se
rect 20937 41582 21014 41598
rect 20921 41516 21014 41582
rect 20921 41414 21014 41480
tri 20921 41398 20937 41414 ne
rect 20937 41398 21014 41414
rect 20754 41299 20902 41381
rect 20642 41266 20719 41282
tri 20719 41266 20735 41282 sw
rect 20642 41200 20735 41266
rect 20771 41141 20885 41299
tri 20921 41266 20937 41282 se
rect 20937 41266 21014 41282
rect 20921 41200 21014 41266
rect 20642 41065 21014 41141
rect 20642 40940 20735 41006
rect 20642 40924 20719 40940
tri 20719 40924 20735 40940 nw
rect 20771 40907 20885 41065
rect 20921 40940 21014 41006
tri 20921 40924 20937 40940 ne
rect 20937 40924 21014 40940
rect 20754 40825 20902 40907
rect 20642 40792 20719 40808
tri 20719 40792 20735 40808 sw
rect 20642 40726 20735 40792
rect 20642 40624 20735 40690
rect 20642 40608 20719 40624
tri 20719 40608 20735 40624 nw
rect 20771 40591 20885 40825
tri 20921 40792 20937 40808 se
rect 20937 40792 21014 40808
rect 20921 40726 21014 40792
rect 20921 40624 21014 40690
tri 20921 40608 20937 40624 ne
rect 20937 40608 21014 40624
rect 20754 40509 20902 40591
rect 20642 40476 20719 40492
tri 20719 40476 20735 40492 sw
rect 20642 40410 20735 40476
rect 20771 40351 20885 40509
tri 20921 40476 20937 40492 se
rect 20937 40476 21014 40492
rect 20921 40410 21014 40476
rect 20642 40275 21014 40351
rect 20642 40150 20735 40216
rect 20642 40134 20719 40150
tri 20719 40134 20735 40150 nw
rect 20771 40117 20885 40275
rect 20921 40150 21014 40216
tri 20921 40134 20937 40150 ne
rect 20937 40134 21014 40150
rect 20754 40035 20902 40117
rect 20642 40002 20719 40018
tri 20719 40002 20735 40018 sw
rect 20642 39936 20735 40002
rect 20642 39834 20735 39900
rect 20642 39818 20719 39834
tri 20719 39818 20735 39834 nw
rect 20771 39801 20885 40035
tri 20921 40002 20937 40018 se
rect 20937 40002 21014 40018
rect 20921 39936 21014 40002
rect 20921 39834 21014 39900
tri 20921 39818 20937 39834 ne
rect 20937 39818 21014 39834
rect 20754 39719 20902 39801
rect 20642 39686 20719 39702
tri 20719 39686 20735 39702 sw
rect 20642 39620 20735 39686
rect 20771 39561 20885 39719
tri 20921 39686 20937 39702 se
rect 20937 39686 21014 39702
rect 20921 39620 21014 39686
rect 20642 39485 21014 39561
rect 20642 39360 20735 39426
rect 20642 39344 20719 39360
tri 20719 39344 20735 39360 nw
rect 20771 39327 20885 39485
rect 20921 39360 21014 39426
tri 20921 39344 20937 39360 ne
rect 20937 39344 21014 39360
rect 20754 39245 20902 39327
rect 20642 39212 20719 39228
tri 20719 39212 20735 39228 sw
rect 20642 39146 20735 39212
rect 20642 39044 20735 39110
rect 20642 39028 20719 39044
tri 20719 39028 20735 39044 nw
rect 20771 39011 20885 39245
tri 20921 39212 20937 39228 se
rect 20937 39212 21014 39228
rect 20921 39146 21014 39212
rect 20921 39044 21014 39110
tri 20921 39028 20937 39044 ne
rect 20937 39028 21014 39044
rect 20754 38929 20902 39011
rect 20642 38896 20719 38912
tri 20719 38896 20735 38912 sw
rect 20642 38830 20735 38896
rect 20771 38771 20885 38929
tri 20921 38896 20937 38912 se
rect 20937 38896 21014 38912
rect 20921 38830 21014 38896
rect 20642 38695 21014 38771
rect 20642 38570 20735 38636
rect 20642 38554 20719 38570
tri 20719 38554 20735 38570 nw
rect 20771 38537 20885 38695
rect 20921 38570 21014 38636
tri 20921 38554 20937 38570 ne
rect 20937 38554 21014 38570
rect 20754 38455 20902 38537
rect 20642 38422 20719 38438
tri 20719 38422 20735 38438 sw
rect 20642 38356 20735 38422
rect 20642 38254 20735 38320
rect 20642 38238 20719 38254
tri 20719 38238 20735 38254 nw
rect 20771 38221 20885 38455
tri 20921 38422 20937 38438 se
rect 20937 38422 21014 38438
rect 20921 38356 21014 38422
rect 20921 38254 21014 38320
tri 20921 38238 20937 38254 ne
rect 20937 38238 21014 38254
rect 20754 38139 20902 38221
rect 20642 38106 20719 38122
tri 20719 38106 20735 38122 sw
rect 20642 38040 20735 38106
rect 20771 37981 20885 38139
tri 20921 38106 20937 38122 se
rect 20937 38106 21014 38122
rect 20921 38040 21014 38106
rect 20642 37905 21014 37981
rect 20642 37780 20735 37846
rect 20642 37764 20719 37780
tri 20719 37764 20735 37780 nw
rect 20771 37747 20885 37905
rect 20921 37780 21014 37846
tri 20921 37764 20937 37780 ne
rect 20937 37764 21014 37780
rect 20754 37665 20902 37747
rect 20642 37632 20719 37648
tri 20719 37632 20735 37648 sw
rect 20642 37566 20735 37632
rect 20642 37464 20735 37530
rect 20642 37448 20719 37464
tri 20719 37448 20735 37464 nw
rect 20771 37431 20885 37665
tri 20921 37632 20937 37648 se
rect 20937 37632 21014 37648
rect 20921 37566 21014 37632
rect 20921 37464 21014 37530
tri 20921 37448 20937 37464 ne
rect 20937 37448 21014 37464
rect 20754 37349 20902 37431
rect 20642 37316 20719 37332
tri 20719 37316 20735 37332 sw
rect 20642 37250 20735 37316
rect 20771 37191 20885 37349
tri 20921 37316 20937 37332 se
rect 20937 37316 21014 37332
rect 20921 37250 21014 37316
rect 20642 37115 21014 37191
rect 20642 36990 20735 37056
rect 20642 36974 20719 36990
tri 20719 36974 20735 36990 nw
rect 20771 36957 20885 37115
rect 20921 36990 21014 37056
tri 20921 36974 20937 36990 ne
rect 20937 36974 21014 36990
rect 20754 36875 20902 36957
rect 20642 36842 20719 36858
tri 20719 36842 20735 36858 sw
rect 20642 36776 20735 36842
rect 20642 36674 20735 36740
rect 20642 36658 20719 36674
tri 20719 36658 20735 36674 nw
rect 20771 36641 20885 36875
tri 20921 36842 20937 36858 se
rect 20937 36842 21014 36858
rect 20921 36776 21014 36842
rect 20921 36674 21014 36740
tri 20921 36658 20937 36674 ne
rect 20937 36658 21014 36674
rect 20754 36559 20902 36641
rect 20642 36526 20719 36542
tri 20719 36526 20735 36542 sw
rect 20642 36460 20735 36526
rect 20771 36401 20885 36559
tri 20921 36526 20937 36542 se
rect 20937 36526 21014 36542
rect 20921 36460 21014 36526
rect 20642 36325 21014 36401
rect 20642 36200 20735 36266
rect 20642 36184 20719 36200
tri 20719 36184 20735 36200 nw
rect 20771 36167 20885 36325
rect 20921 36200 21014 36266
tri 20921 36184 20937 36200 ne
rect 20937 36184 21014 36200
rect 20754 36085 20902 36167
rect 20642 36052 20719 36068
tri 20719 36052 20735 36068 sw
rect 20642 35986 20735 36052
rect 20642 35884 20735 35950
rect 20642 35868 20719 35884
tri 20719 35868 20735 35884 nw
rect 20771 35851 20885 36085
tri 20921 36052 20937 36068 se
rect 20937 36052 21014 36068
rect 20921 35986 21014 36052
rect 20921 35884 21014 35950
tri 20921 35868 20937 35884 ne
rect 20937 35868 21014 35884
rect 20754 35769 20902 35851
rect 20642 35736 20719 35752
tri 20719 35736 20735 35752 sw
rect 20642 35670 20735 35736
rect 20771 35611 20885 35769
tri 20921 35736 20937 35752 se
rect 20937 35736 21014 35752
rect 20921 35670 21014 35736
rect 20642 35535 21014 35611
rect 20642 35410 20735 35476
rect 20642 35394 20719 35410
tri 20719 35394 20735 35410 nw
rect 20771 35377 20885 35535
rect 20921 35410 21014 35476
tri 20921 35394 20937 35410 ne
rect 20937 35394 21014 35410
rect 20754 35295 20902 35377
rect 20642 35262 20719 35278
tri 20719 35262 20735 35278 sw
rect 20642 35196 20735 35262
rect 20642 35094 20735 35160
rect 20642 35078 20719 35094
tri 20719 35078 20735 35094 nw
rect 20771 35061 20885 35295
tri 20921 35262 20937 35278 se
rect 20937 35262 21014 35278
rect 20921 35196 21014 35262
rect 20921 35094 21014 35160
tri 20921 35078 20937 35094 ne
rect 20937 35078 21014 35094
rect 20754 34979 20902 35061
rect 20642 34946 20719 34962
tri 20719 34946 20735 34962 sw
rect 20642 34880 20735 34946
rect 20771 34821 20885 34979
tri 20921 34946 20937 34962 se
rect 20937 34946 21014 34962
rect 20921 34880 21014 34946
rect 20642 34745 21014 34821
rect 20642 34620 20735 34686
rect 20642 34604 20719 34620
tri 20719 34604 20735 34620 nw
rect 20771 34587 20885 34745
rect 20921 34620 21014 34686
tri 20921 34604 20937 34620 ne
rect 20937 34604 21014 34620
rect 20754 34505 20902 34587
rect 20642 34472 20719 34488
tri 20719 34472 20735 34488 sw
rect 20642 34406 20735 34472
rect 20642 34304 20735 34370
rect 20642 34288 20719 34304
tri 20719 34288 20735 34304 nw
rect 20771 34271 20885 34505
tri 20921 34472 20937 34488 se
rect 20937 34472 21014 34488
rect 20921 34406 21014 34472
rect 20921 34304 21014 34370
tri 20921 34288 20937 34304 ne
rect 20937 34288 21014 34304
rect 20754 34189 20902 34271
rect 20642 34156 20719 34172
tri 20719 34156 20735 34172 sw
rect 20642 34090 20735 34156
rect 20771 34031 20885 34189
tri 20921 34156 20937 34172 se
rect 20937 34156 21014 34172
rect 20921 34090 21014 34156
rect 20642 33955 21014 34031
rect 20642 33830 20735 33896
rect 20642 33814 20719 33830
tri 20719 33814 20735 33830 nw
rect 20771 33797 20885 33955
rect 20921 33830 21014 33896
tri 20921 33814 20937 33830 ne
rect 20937 33814 21014 33830
rect 20754 33715 20902 33797
rect 20642 33682 20719 33698
tri 20719 33682 20735 33698 sw
rect 20642 33616 20735 33682
rect 20642 33514 20735 33580
rect 20642 33498 20719 33514
tri 20719 33498 20735 33514 nw
rect 20771 33481 20885 33715
tri 20921 33682 20937 33698 se
rect 20937 33682 21014 33698
rect 20921 33616 21014 33682
rect 20921 33514 21014 33580
tri 20921 33498 20937 33514 ne
rect 20937 33498 21014 33514
rect 20754 33399 20902 33481
rect 20642 33366 20719 33382
tri 20719 33366 20735 33382 sw
rect 20642 33300 20735 33366
rect 20771 33241 20885 33399
tri 20921 33366 20937 33382 se
rect 20937 33366 21014 33382
rect 20921 33300 21014 33366
rect 20642 33165 21014 33241
rect 20642 33040 20735 33106
rect 20642 33024 20719 33040
tri 20719 33024 20735 33040 nw
rect 20771 33007 20885 33165
rect 20921 33040 21014 33106
tri 20921 33024 20937 33040 ne
rect 20937 33024 21014 33040
rect 20754 32925 20902 33007
rect 20642 32892 20719 32908
tri 20719 32892 20735 32908 sw
rect 20642 32826 20735 32892
rect 20642 32724 20735 32790
rect 20642 32708 20719 32724
tri 20719 32708 20735 32724 nw
rect 20771 32691 20885 32925
tri 20921 32892 20937 32908 se
rect 20937 32892 21014 32908
rect 20921 32826 21014 32892
rect 20921 32724 21014 32790
tri 20921 32708 20937 32724 ne
rect 20937 32708 21014 32724
rect 20754 32609 20902 32691
rect 20642 32576 20719 32592
tri 20719 32576 20735 32592 sw
rect 20642 32510 20735 32576
rect 20771 32451 20885 32609
tri 20921 32576 20937 32592 se
rect 20937 32576 21014 32592
rect 20921 32510 21014 32576
rect 20642 32375 21014 32451
rect 20642 32250 20735 32316
rect 20642 32234 20719 32250
tri 20719 32234 20735 32250 nw
rect 20771 32217 20885 32375
rect 20921 32250 21014 32316
tri 20921 32234 20937 32250 ne
rect 20937 32234 21014 32250
rect 20754 32135 20902 32217
rect 20642 32102 20719 32118
tri 20719 32102 20735 32118 sw
rect 20642 32036 20735 32102
rect 20642 31934 20735 32000
rect 20642 31918 20719 31934
tri 20719 31918 20735 31934 nw
rect 20771 31901 20885 32135
tri 20921 32102 20937 32118 se
rect 20937 32102 21014 32118
rect 20921 32036 21014 32102
rect 20921 31934 21014 32000
tri 20921 31918 20937 31934 ne
rect 20937 31918 21014 31934
rect 20754 31819 20902 31901
rect 20642 31786 20719 31802
tri 20719 31786 20735 31802 sw
rect 20642 31720 20735 31786
rect 20771 31661 20885 31819
tri 20921 31786 20937 31802 se
rect 20937 31786 21014 31802
rect 20921 31720 21014 31786
rect 20642 31585 21014 31661
rect 20642 31460 20735 31526
rect 20642 31444 20719 31460
tri 20719 31444 20735 31460 nw
rect 20771 31427 20885 31585
rect 20921 31460 21014 31526
tri 20921 31444 20937 31460 ne
rect 20937 31444 21014 31460
rect 20754 31345 20902 31427
rect 20642 31312 20719 31328
tri 20719 31312 20735 31328 sw
rect 20642 31246 20735 31312
rect 20642 31144 20735 31210
rect 20642 31128 20719 31144
tri 20719 31128 20735 31144 nw
rect 20771 31111 20885 31345
tri 20921 31312 20937 31328 se
rect 20937 31312 21014 31328
rect 20921 31246 21014 31312
rect 20921 31144 21014 31210
tri 20921 31128 20937 31144 ne
rect 20937 31128 21014 31144
rect 20754 31029 20902 31111
rect 20642 30996 20719 31012
tri 20719 30996 20735 31012 sw
rect 20642 30930 20735 30996
rect 20771 30871 20885 31029
tri 20921 30996 20937 31012 se
rect 20937 30996 21014 31012
rect 20921 30930 21014 30996
rect 20642 30795 21014 30871
rect 20642 30670 20735 30736
rect 20642 30654 20719 30670
tri 20719 30654 20735 30670 nw
rect 20771 30637 20885 30795
rect 20921 30670 21014 30736
tri 20921 30654 20937 30670 ne
rect 20937 30654 21014 30670
rect 20754 30555 20902 30637
rect 20642 30522 20719 30538
tri 20719 30522 20735 30538 sw
rect 20642 30456 20735 30522
rect 20642 30354 20735 30420
rect 20642 30338 20719 30354
tri 20719 30338 20735 30354 nw
rect 20771 30321 20885 30555
tri 20921 30522 20937 30538 se
rect 20937 30522 21014 30538
rect 20921 30456 21014 30522
rect 20921 30354 21014 30420
tri 20921 30338 20937 30354 ne
rect 20937 30338 21014 30354
rect 20754 30239 20902 30321
rect 20642 30206 20719 30222
tri 20719 30206 20735 30222 sw
rect 20642 30140 20735 30206
rect 20771 30081 20885 30239
tri 20921 30206 20937 30222 se
rect 20937 30206 21014 30222
rect 20921 30140 21014 30206
rect 20642 30005 21014 30081
rect 20642 29880 20735 29946
rect 20642 29864 20719 29880
tri 20719 29864 20735 29880 nw
rect 20771 29847 20885 30005
rect 20921 29880 21014 29946
tri 20921 29864 20937 29880 ne
rect 20937 29864 21014 29880
rect 20754 29765 20902 29847
rect 20642 29732 20719 29748
tri 20719 29732 20735 29748 sw
rect 20642 29666 20735 29732
rect 20642 29564 20735 29630
rect 20642 29548 20719 29564
tri 20719 29548 20735 29564 nw
rect 20771 29531 20885 29765
tri 20921 29732 20937 29748 se
rect 20937 29732 21014 29748
rect 20921 29666 21014 29732
rect 20921 29564 21014 29630
tri 20921 29548 20937 29564 ne
rect 20937 29548 21014 29564
rect 20754 29449 20902 29531
rect 20642 29416 20719 29432
tri 20719 29416 20735 29432 sw
rect 20642 29350 20735 29416
rect 20771 29291 20885 29449
tri 20921 29416 20937 29432 se
rect 20937 29416 21014 29432
rect 20921 29350 21014 29416
rect 20642 29215 21014 29291
rect 20642 29090 20735 29156
rect 20642 29074 20719 29090
tri 20719 29074 20735 29090 nw
rect 20771 29057 20885 29215
rect 20921 29090 21014 29156
tri 20921 29074 20937 29090 ne
rect 20937 29074 21014 29090
rect 20754 28975 20902 29057
rect 20642 28942 20719 28958
tri 20719 28942 20735 28958 sw
rect 20642 28876 20735 28942
rect 20771 28833 20885 28975
tri 20921 28942 20937 28958 se
rect 20937 28942 21014 28958
rect 20921 28876 21014 28942
rect 21050 28463 21086 80603
rect 21122 28463 21158 80603
rect 21194 80445 21230 80603
rect 21186 80303 21238 80445
rect 21194 28763 21230 80303
rect 21186 28621 21238 28763
rect 21194 28463 21230 28621
rect 21266 28463 21302 80603
rect 21338 28463 21374 80603
rect 21410 28833 21494 80233
rect 21530 28463 21566 80603
rect 21602 28463 21638 80603
rect 21674 80445 21710 80603
rect 21666 80303 21718 80445
rect 21674 28763 21710 80303
rect 21666 28621 21718 28763
rect 21674 28463 21710 28621
rect 21746 28463 21782 80603
rect 21818 28463 21854 80603
rect 21890 80124 21983 80190
rect 21890 80108 21967 80124
tri 21967 80108 21983 80124 nw
rect 22019 80091 22133 80233
rect 22169 80124 22262 80190
tri 22169 80108 22185 80124 ne
rect 22185 80108 22262 80124
rect 22002 80009 22150 80091
rect 21890 79976 21967 79992
tri 21967 79976 21983 79992 sw
rect 21890 79910 21983 79976
rect 22019 79851 22133 80009
tri 22169 79976 22185 79992 se
rect 22185 79976 22262 79992
rect 22169 79910 22262 79976
rect 21890 79775 22262 79851
rect 21890 79650 21983 79716
rect 21890 79634 21967 79650
tri 21967 79634 21983 79650 nw
rect 22019 79617 22133 79775
rect 22169 79650 22262 79716
tri 22169 79634 22185 79650 ne
rect 22185 79634 22262 79650
rect 22002 79535 22150 79617
rect 21890 79502 21967 79518
tri 21967 79502 21983 79518 sw
rect 21890 79436 21983 79502
rect 21890 79334 21983 79400
rect 21890 79318 21967 79334
tri 21967 79318 21983 79334 nw
rect 22019 79301 22133 79535
tri 22169 79502 22185 79518 se
rect 22185 79502 22262 79518
rect 22169 79436 22262 79502
rect 22169 79334 22262 79400
tri 22169 79318 22185 79334 ne
rect 22185 79318 22262 79334
rect 22002 79219 22150 79301
rect 21890 79186 21967 79202
tri 21967 79186 21983 79202 sw
rect 21890 79120 21983 79186
rect 22019 79061 22133 79219
tri 22169 79186 22185 79202 se
rect 22185 79186 22262 79202
rect 22169 79120 22262 79186
rect 21890 78985 22262 79061
rect 21890 78860 21983 78926
rect 21890 78844 21967 78860
tri 21967 78844 21983 78860 nw
rect 22019 78827 22133 78985
rect 22169 78860 22262 78926
tri 22169 78844 22185 78860 ne
rect 22185 78844 22262 78860
rect 22002 78745 22150 78827
rect 21890 78712 21967 78728
tri 21967 78712 21983 78728 sw
rect 21890 78646 21983 78712
rect 21890 78544 21983 78610
rect 21890 78528 21967 78544
tri 21967 78528 21983 78544 nw
rect 22019 78511 22133 78745
tri 22169 78712 22185 78728 se
rect 22185 78712 22262 78728
rect 22169 78646 22262 78712
rect 22169 78544 22262 78610
tri 22169 78528 22185 78544 ne
rect 22185 78528 22262 78544
rect 22002 78429 22150 78511
rect 21890 78396 21967 78412
tri 21967 78396 21983 78412 sw
rect 21890 78330 21983 78396
rect 22019 78271 22133 78429
tri 22169 78396 22185 78412 se
rect 22185 78396 22262 78412
rect 22169 78330 22262 78396
rect 21890 78195 22262 78271
rect 21890 78070 21983 78136
rect 21890 78054 21967 78070
tri 21967 78054 21983 78070 nw
rect 22019 78037 22133 78195
rect 22169 78070 22262 78136
tri 22169 78054 22185 78070 ne
rect 22185 78054 22262 78070
rect 22002 77955 22150 78037
rect 21890 77922 21967 77938
tri 21967 77922 21983 77938 sw
rect 21890 77856 21983 77922
rect 21890 77754 21983 77820
rect 21890 77738 21967 77754
tri 21967 77738 21983 77754 nw
rect 22019 77721 22133 77955
tri 22169 77922 22185 77938 se
rect 22185 77922 22262 77938
rect 22169 77856 22262 77922
rect 22169 77754 22262 77820
tri 22169 77738 22185 77754 ne
rect 22185 77738 22262 77754
rect 22002 77639 22150 77721
rect 21890 77606 21967 77622
tri 21967 77606 21983 77622 sw
rect 21890 77540 21983 77606
rect 22019 77481 22133 77639
tri 22169 77606 22185 77622 se
rect 22185 77606 22262 77622
rect 22169 77540 22262 77606
rect 21890 77405 22262 77481
rect 21890 77280 21983 77346
rect 21890 77264 21967 77280
tri 21967 77264 21983 77280 nw
rect 22019 77247 22133 77405
rect 22169 77280 22262 77346
tri 22169 77264 22185 77280 ne
rect 22185 77264 22262 77280
rect 22002 77165 22150 77247
rect 21890 77132 21967 77148
tri 21967 77132 21983 77148 sw
rect 21890 77066 21983 77132
rect 21890 76964 21983 77030
rect 21890 76948 21967 76964
tri 21967 76948 21983 76964 nw
rect 22019 76931 22133 77165
tri 22169 77132 22185 77148 se
rect 22185 77132 22262 77148
rect 22169 77066 22262 77132
rect 22169 76964 22262 77030
tri 22169 76948 22185 76964 ne
rect 22185 76948 22262 76964
rect 22002 76849 22150 76931
rect 21890 76816 21967 76832
tri 21967 76816 21983 76832 sw
rect 21890 76750 21983 76816
rect 22019 76691 22133 76849
tri 22169 76816 22185 76832 se
rect 22185 76816 22262 76832
rect 22169 76750 22262 76816
rect 21890 76615 22262 76691
rect 21890 76490 21983 76556
rect 21890 76474 21967 76490
tri 21967 76474 21983 76490 nw
rect 22019 76457 22133 76615
rect 22169 76490 22262 76556
tri 22169 76474 22185 76490 ne
rect 22185 76474 22262 76490
rect 22002 76375 22150 76457
rect 21890 76342 21967 76358
tri 21967 76342 21983 76358 sw
rect 21890 76276 21983 76342
rect 21890 76174 21983 76240
rect 21890 76158 21967 76174
tri 21967 76158 21983 76174 nw
rect 22019 76141 22133 76375
tri 22169 76342 22185 76358 se
rect 22185 76342 22262 76358
rect 22169 76276 22262 76342
rect 22169 76174 22262 76240
tri 22169 76158 22185 76174 ne
rect 22185 76158 22262 76174
rect 22002 76059 22150 76141
rect 21890 76026 21967 76042
tri 21967 76026 21983 76042 sw
rect 21890 75960 21983 76026
rect 22019 75901 22133 76059
tri 22169 76026 22185 76042 se
rect 22185 76026 22262 76042
rect 22169 75960 22262 76026
rect 21890 75825 22262 75901
rect 21890 75700 21983 75766
rect 21890 75684 21967 75700
tri 21967 75684 21983 75700 nw
rect 22019 75667 22133 75825
rect 22169 75700 22262 75766
tri 22169 75684 22185 75700 ne
rect 22185 75684 22262 75700
rect 22002 75585 22150 75667
rect 21890 75552 21967 75568
tri 21967 75552 21983 75568 sw
rect 21890 75486 21983 75552
rect 21890 75384 21983 75450
rect 21890 75368 21967 75384
tri 21967 75368 21983 75384 nw
rect 22019 75351 22133 75585
tri 22169 75552 22185 75568 se
rect 22185 75552 22262 75568
rect 22169 75486 22262 75552
rect 22169 75384 22262 75450
tri 22169 75368 22185 75384 ne
rect 22185 75368 22262 75384
rect 22002 75269 22150 75351
rect 21890 75236 21967 75252
tri 21967 75236 21983 75252 sw
rect 21890 75170 21983 75236
rect 22019 75111 22133 75269
tri 22169 75236 22185 75252 se
rect 22185 75236 22262 75252
rect 22169 75170 22262 75236
rect 21890 75035 22262 75111
rect 21890 74910 21983 74976
rect 21890 74894 21967 74910
tri 21967 74894 21983 74910 nw
rect 22019 74877 22133 75035
rect 22169 74910 22262 74976
tri 22169 74894 22185 74910 ne
rect 22185 74894 22262 74910
rect 22002 74795 22150 74877
rect 21890 74762 21967 74778
tri 21967 74762 21983 74778 sw
rect 21890 74696 21983 74762
rect 21890 74594 21983 74660
rect 21890 74578 21967 74594
tri 21967 74578 21983 74594 nw
rect 22019 74561 22133 74795
tri 22169 74762 22185 74778 se
rect 22185 74762 22262 74778
rect 22169 74696 22262 74762
rect 22169 74594 22262 74660
tri 22169 74578 22185 74594 ne
rect 22185 74578 22262 74594
rect 22002 74479 22150 74561
rect 21890 74446 21967 74462
tri 21967 74446 21983 74462 sw
rect 21890 74380 21983 74446
rect 22019 74321 22133 74479
tri 22169 74446 22185 74462 se
rect 22185 74446 22262 74462
rect 22169 74380 22262 74446
rect 21890 74245 22262 74321
rect 21890 74120 21983 74186
rect 21890 74104 21967 74120
tri 21967 74104 21983 74120 nw
rect 22019 74087 22133 74245
rect 22169 74120 22262 74186
tri 22169 74104 22185 74120 ne
rect 22185 74104 22262 74120
rect 22002 74005 22150 74087
rect 21890 73972 21967 73988
tri 21967 73972 21983 73988 sw
rect 21890 73906 21983 73972
rect 21890 73804 21983 73870
rect 21890 73788 21967 73804
tri 21967 73788 21983 73804 nw
rect 22019 73771 22133 74005
tri 22169 73972 22185 73988 se
rect 22185 73972 22262 73988
rect 22169 73906 22262 73972
rect 22169 73804 22262 73870
tri 22169 73788 22185 73804 ne
rect 22185 73788 22262 73804
rect 22002 73689 22150 73771
rect 21890 73656 21967 73672
tri 21967 73656 21983 73672 sw
rect 21890 73590 21983 73656
rect 22019 73531 22133 73689
tri 22169 73656 22185 73672 se
rect 22185 73656 22262 73672
rect 22169 73590 22262 73656
rect 21890 73455 22262 73531
rect 21890 73330 21983 73396
rect 21890 73314 21967 73330
tri 21967 73314 21983 73330 nw
rect 22019 73297 22133 73455
rect 22169 73330 22262 73396
tri 22169 73314 22185 73330 ne
rect 22185 73314 22262 73330
rect 22002 73215 22150 73297
rect 21890 73182 21967 73198
tri 21967 73182 21983 73198 sw
rect 21890 73116 21983 73182
rect 21890 73014 21983 73080
rect 21890 72998 21967 73014
tri 21967 72998 21983 73014 nw
rect 22019 72981 22133 73215
tri 22169 73182 22185 73198 se
rect 22185 73182 22262 73198
rect 22169 73116 22262 73182
rect 22169 73014 22262 73080
tri 22169 72998 22185 73014 ne
rect 22185 72998 22262 73014
rect 22002 72899 22150 72981
rect 21890 72866 21967 72882
tri 21967 72866 21983 72882 sw
rect 21890 72800 21983 72866
rect 22019 72741 22133 72899
tri 22169 72866 22185 72882 se
rect 22185 72866 22262 72882
rect 22169 72800 22262 72866
rect 21890 72665 22262 72741
rect 21890 72540 21983 72606
rect 21890 72524 21967 72540
tri 21967 72524 21983 72540 nw
rect 22019 72507 22133 72665
rect 22169 72540 22262 72606
tri 22169 72524 22185 72540 ne
rect 22185 72524 22262 72540
rect 22002 72425 22150 72507
rect 21890 72392 21967 72408
tri 21967 72392 21983 72408 sw
rect 21890 72326 21983 72392
rect 21890 72224 21983 72290
rect 21890 72208 21967 72224
tri 21967 72208 21983 72224 nw
rect 22019 72191 22133 72425
tri 22169 72392 22185 72408 se
rect 22185 72392 22262 72408
rect 22169 72326 22262 72392
rect 22169 72224 22262 72290
tri 22169 72208 22185 72224 ne
rect 22185 72208 22262 72224
rect 22002 72109 22150 72191
rect 21890 72076 21967 72092
tri 21967 72076 21983 72092 sw
rect 21890 72010 21983 72076
rect 22019 71951 22133 72109
tri 22169 72076 22185 72092 se
rect 22185 72076 22262 72092
rect 22169 72010 22262 72076
rect 21890 71875 22262 71951
rect 21890 71750 21983 71816
rect 21890 71734 21967 71750
tri 21967 71734 21983 71750 nw
rect 22019 71717 22133 71875
rect 22169 71750 22262 71816
tri 22169 71734 22185 71750 ne
rect 22185 71734 22262 71750
rect 22002 71635 22150 71717
rect 21890 71602 21967 71618
tri 21967 71602 21983 71618 sw
rect 21890 71536 21983 71602
rect 21890 71434 21983 71500
rect 21890 71418 21967 71434
tri 21967 71418 21983 71434 nw
rect 22019 71401 22133 71635
tri 22169 71602 22185 71618 se
rect 22185 71602 22262 71618
rect 22169 71536 22262 71602
rect 22169 71434 22262 71500
tri 22169 71418 22185 71434 ne
rect 22185 71418 22262 71434
rect 22002 71319 22150 71401
rect 21890 71286 21967 71302
tri 21967 71286 21983 71302 sw
rect 21890 71220 21983 71286
rect 22019 71161 22133 71319
tri 22169 71286 22185 71302 se
rect 22185 71286 22262 71302
rect 22169 71220 22262 71286
rect 21890 71085 22262 71161
rect 21890 70960 21983 71026
rect 21890 70944 21967 70960
tri 21967 70944 21983 70960 nw
rect 22019 70927 22133 71085
rect 22169 70960 22262 71026
tri 22169 70944 22185 70960 ne
rect 22185 70944 22262 70960
rect 22002 70845 22150 70927
rect 21890 70812 21967 70828
tri 21967 70812 21983 70828 sw
rect 21890 70746 21983 70812
rect 21890 70644 21983 70710
rect 21890 70628 21967 70644
tri 21967 70628 21983 70644 nw
rect 22019 70611 22133 70845
tri 22169 70812 22185 70828 se
rect 22185 70812 22262 70828
rect 22169 70746 22262 70812
rect 22169 70644 22262 70710
tri 22169 70628 22185 70644 ne
rect 22185 70628 22262 70644
rect 22002 70529 22150 70611
rect 21890 70496 21967 70512
tri 21967 70496 21983 70512 sw
rect 21890 70430 21983 70496
rect 22019 70371 22133 70529
tri 22169 70496 22185 70512 se
rect 22185 70496 22262 70512
rect 22169 70430 22262 70496
rect 21890 70295 22262 70371
rect 21890 70170 21983 70236
rect 21890 70154 21967 70170
tri 21967 70154 21983 70170 nw
rect 22019 70137 22133 70295
rect 22169 70170 22262 70236
tri 22169 70154 22185 70170 ne
rect 22185 70154 22262 70170
rect 22002 70055 22150 70137
rect 21890 70022 21967 70038
tri 21967 70022 21983 70038 sw
rect 21890 69956 21983 70022
rect 21890 69854 21983 69920
rect 21890 69838 21967 69854
tri 21967 69838 21983 69854 nw
rect 22019 69821 22133 70055
tri 22169 70022 22185 70038 se
rect 22185 70022 22262 70038
rect 22169 69956 22262 70022
rect 22169 69854 22262 69920
tri 22169 69838 22185 69854 ne
rect 22185 69838 22262 69854
rect 22002 69739 22150 69821
rect 21890 69706 21967 69722
tri 21967 69706 21983 69722 sw
rect 21890 69640 21983 69706
rect 22019 69581 22133 69739
tri 22169 69706 22185 69722 se
rect 22185 69706 22262 69722
rect 22169 69640 22262 69706
rect 21890 69505 22262 69581
rect 21890 69380 21983 69446
rect 21890 69364 21967 69380
tri 21967 69364 21983 69380 nw
rect 22019 69347 22133 69505
rect 22169 69380 22262 69446
tri 22169 69364 22185 69380 ne
rect 22185 69364 22262 69380
rect 22002 69265 22150 69347
rect 21890 69232 21967 69248
tri 21967 69232 21983 69248 sw
rect 21890 69166 21983 69232
rect 21890 69064 21983 69130
rect 21890 69048 21967 69064
tri 21967 69048 21983 69064 nw
rect 22019 69031 22133 69265
tri 22169 69232 22185 69248 se
rect 22185 69232 22262 69248
rect 22169 69166 22262 69232
rect 22169 69064 22262 69130
tri 22169 69048 22185 69064 ne
rect 22185 69048 22262 69064
rect 22002 68949 22150 69031
rect 21890 68916 21967 68932
tri 21967 68916 21983 68932 sw
rect 21890 68850 21983 68916
rect 22019 68791 22133 68949
tri 22169 68916 22185 68932 se
rect 22185 68916 22262 68932
rect 22169 68850 22262 68916
rect 21890 68715 22262 68791
rect 21890 68590 21983 68656
rect 21890 68574 21967 68590
tri 21967 68574 21983 68590 nw
rect 22019 68557 22133 68715
rect 22169 68590 22262 68656
tri 22169 68574 22185 68590 ne
rect 22185 68574 22262 68590
rect 22002 68475 22150 68557
rect 21890 68442 21967 68458
tri 21967 68442 21983 68458 sw
rect 21890 68376 21983 68442
rect 21890 68274 21983 68340
rect 21890 68258 21967 68274
tri 21967 68258 21983 68274 nw
rect 22019 68241 22133 68475
tri 22169 68442 22185 68458 se
rect 22185 68442 22262 68458
rect 22169 68376 22262 68442
rect 22169 68274 22262 68340
tri 22169 68258 22185 68274 ne
rect 22185 68258 22262 68274
rect 22002 68159 22150 68241
rect 21890 68126 21967 68142
tri 21967 68126 21983 68142 sw
rect 21890 68060 21983 68126
rect 22019 68001 22133 68159
tri 22169 68126 22185 68142 se
rect 22185 68126 22262 68142
rect 22169 68060 22262 68126
rect 21890 67925 22262 68001
rect 21890 67800 21983 67866
rect 21890 67784 21967 67800
tri 21967 67784 21983 67800 nw
rect 22019 67767 22133 67925
rect 22169 67800 22262 67866
tri 22169 67784 22185 67800 ne
rect 22185 67784 22262 67800
rect 22002 67685 22150 67767
rect 21890 67652 21967 67668
tri 21967 67652 21983 67668 sw
rect 21890 67586 21983 67652
rect 21890 67484 21983 67550
rect 21890 67468 21967 67484
tri 21967 67468 21983 67484 nw
rect 22019 67451 22133 67685
tri 22169 67652 22185 67668 se
rect 22185 67652 22262 67668
rect 22169 67586 22262 67652
rect 22169 67484 22262 67550
tri 22169 67468 22185 67484 ne
rect 22185 67468 22262 67484
rect 22002 67369 22150 67451
rect 21890 67336 21967 67352
tri 21967 67336 21983 67352 sw
rect 21890 67270 21983 67336
rect 22019 67211 22133 67369
tri 22169 67336 22185 67352 se
rect 22185 67336 22262 67352
rect 22169 67270 22262 67336
rect 21890 67135 22262 67211
rect 21890 67010 21983 67076
rect 21890 66994 21967 67010
tri 21967 66994 21983 67010 nw
rect 22019 66977 22133 67135
rect 22169 67010 22262 67076
tri 22169 66994 22185 67010 ne
rect 22185 66994 22262 67010
rect 22002 66895 22150 66977
rect 21890 66862 21967 66878
tri 21967 66862 21983 66878 sw
rect 21890 66796 21983 66862
rect 21890 66694 21983 66760
rect 21890 66678 21967 66694
tri 21967 66678 21983 66694 nw
rect 22019 66661 22133 66895
tri 22169 66862 22185 66878 se
rect 22185 66862 22262 66878
rect 22169 66796 22262 66862
rect 22169 66694 22262 66760
tri 22169 66678 22185 66694 ne
rect 22185 66678 22262 66694
rect 22002 66579 22150 66661
rect 21890 66546 21967 66562
tri 21967 66546 21983 66562 sw
rect 21890 66480 21983 66546
rect 22019 66421 22133 66579
tri 22169 66546 22185 66562 se
rect 22185 66546 22262 66562
rect 22169 66480 22262 66546
rect 21890 66345 22262 66421
rect 21890 66220 21983 66286
rect 21890 66204 21967 66220
tri 21967 66204 21983 66220 nw
rect 22019 66187 22133 66345
rect 22169 66220 22262 66286
tri 22169 66204 22185 66220 ne
rect 22185 66204 22262 66220
rect 22002 66105 22150 66187
rect 21890 66072 21967 66088
tri 21967 66072 21983 66088 sw
rect 21890 66006 21983 66072
rect 21890 65904 21983 65970
rect 21890 65888 21967 65904
tri 21967 65888 21983 65904 nw
rect 22019 65871 22133 66105
tri 22169 66072 22185 66088 se
rect 22185 66072 22262 66088
rect 22169 66006 22262 66072
rect 22169 65904 22262 65970
tri 22169 65888 22185 65904 ne
rect 22185 65888 22262 65904
rect 22002 65789 22150 65871
rect 21890 65756 21967 65772
tri 21967 65756 21983 65772 sw
rect 21890 65690 21983 65756
rect 22019 65631 22133 65789
tri 22169 65756 22185 65772 se
rect 22185 65756 22262 65772
rect 22169 65690 22262 65756
rect 21890 65555 22262 65631
rect 21890 65430 21983 65496
rect 21890 65414 21967 65430
tri 21967 65414 21983 65430 nw
rect 22019 65397 22133 65555
rect 22169 65430 22262 65496
tri 22169 65414 22185 65430 ne
rect 22185 65414 22262 65430
rect 22002 65315 22150 65397
rect 21890 65282 21967 65298
tri 21967 65282 21983 65298 sw
rect 21890 65216 21983 65282
rect 21890 65114 21983 65180
rect 21890 65098 21967 65114
tri 21967 65098 21983 65114 nw
rect 22019 65081 22133 65315
tri 22169 65282 22185 65298 se
rect 22185 65282 22262 65298
rect 22169 65216 22262 65282
rect 22169 65114 22262 65180
tri 22169 65098 22185 65114 ne
rect 22185 65098 22262 65114
rect 22002 64999 22150 65081
rect 21890 64966 21967 64982
tri 21967 64966 21983 64982 sw
rect 21890 64900 21983 64966
rect 22019 64841 22133 64999
tri 22169 64966 22185 64982 se
rect 22185 64966 22262 64982
rect 22169 64900 22262 64966
rect 21890 64765 22262 64841
rect 21890 64640 21983 64706
rect 21890 64624 21967 64640
tri 21967 64624 21983 64640 nw
rect 22019 64607 22133 64765
rect 22169 64640 22262 64706
tri 22169 64624 22185 64640 ne
rect 22185 64624 22262 64640
rect 22002 64525 22150 64607
rect 21890 64492 21967 64508
tri 21967 64492 21983 64508 sw
rect 21890 64426 21983 64492
rect 21890 64324 21983 64390
rect 21890 64308 21967 64324
tri 21967 64308 21983 64324 nw
rect 22019 64291 22133 64525
tri 22169 64492 22185 64508 se
rect 22185 64492 22262 64508
rect 22169 64426 22262 64492
rect 22169 64324 22262 64390
tri 22169 64308 22185 64324 ne
rect 22185 64308 22262 64324
rect 22002 64209 22150 64291
rect 21890 64176 21967 64192
tri 21967 64176 21983 64192 sw
rect 21890 64110 21983 64176
rect 22019 64051 22133 64209
tri 22169 64176 22185 64192 se
rect 22185 64176 22262 64192
rect 22169 64110 22262 64176
rect 21890 63975 22262 64051
rect 21890 63850 21983 63916
rect 21890 63834 21967 63850
tri 21967 63834 21983 63850 nw
rect 22019 63817 22133 63975
rect 22169 63850 22262 63916
tri 22169 63834 22185 63850 ne
rect 22185 63834 22262 63850
rect 22002 63735 22150 63817
rect 21890 63702 21967 63718
tri 21967 63702 21983 63718 sw
rect 21890 63636 21983 63702
rect 21890 63534 21983 63600
rect 21890 63518 21967 63534
tri 21967 63518 21983 63534 nw
rect 22019 63501 22133 63735
tri 22169 63702 22185 63718 se
rect 22185 63702 22262 63718
rect 22169 63636 22262 63702
rect 22169 63534 22262 63600
tri 22169 63518 22185 63534 ne
rect 22185 63518 22262 63534
rect 22002 63419 22150 63501
rect 21890 63386 21967 63402
tri 21967 63386 21983 63402 sw
rect 21890 63320 21983 63386
rect 22019 63261 22133 63419
tri 22169 63386 22185 63402 se
rect 22185 63386 22262 63402
rect 22169 63320 22262 63386
rect 21890 63185 22262 63261
rect 21890 63060 21983 63126
rect 21890 63044 21967 63060
tri 21967 63044 21983 63060 nw
rect 22019 63027 22133 63185
rect 22169 63060 22262 63126
tri 22169 63044 22185 63060 ne
rect 22185 63044 22262 63060
rect 22002 62945 22150 63027
rect 21890 62912 21967 62928
tri 21967 62912 21983 62928 sw
rect 21890 62846 21983 62912
rect 21890 62744 21983 62810
rect 21890 62728 21967 62744
tri 21967 62728 21983 62744 nw
rect 22019 62711 22133 62945
tri 22169 62912 22185 62928 se
rect 22185 62912 22262 62928
rect 22169 62846 22262 62912
rect 22169 62744 22262 62810
tri 22169 62728 22185 62744 ne
rect 22185 62728 22262 62744
rect 22002 62629 22150 62711
rect 21890 62596 21967 62612
tri 21967 62596 21983 62612 sw
rect 21890 62530 21983 62596
rect 22019 62471 22133 62629
tri 22169 62596 22185 62612 se
rect 22185 62596 22262 62612
rect 22169 62530 22262 62596
rect 21890 62395 22262 62471
rect 21890 62270 21983 62336
rect 21890 62254 21967 62270
tri 21967 62254 21983 62270 nw
rect 22019 62237 22133 62395
rect 22169 62270 22262 62336
tri 22169 62254 22185 62270 ne
rect 22185 62254 22262 62270
rect 22002 62155 22150 62237
rect 21890 62122 21967 62138
tri 21967 62122 21983 62138 sw
rect 21890 62056 21983 62122
rect 21890 61954 21983 62020
rect 21890 61938 21967 61954
tri 21967 61938 21983 61954 nw
rect 22019 61921 22133 62155
tri 22169 62122 22185 62138 se
rect 22185 62122 22262 62138
rect 22169 62056 22262 62122
rect 22169 61954 22262 62020
tri 22169 61938 22185 61954 ne
rect 22185 61938 22262 61954
rect 22002 61839 22150 61921
rect 21890 61806 21967 61822
tri 21967 61806 21983 61822 sw
rect 21890 61740 21983 61806
rect 22019 61681 22133 61839
tri 22169 61806 22185 61822 se
rect 22185 61806 22262 61822
rect 22169 61740 22262 61806
rect 21890 61605 22262 61681
rect 21890 61480 21983 61546
rect 21890 61464 21967 61480
tri 21967 61464 21983 61480 nw
rect 22019 61447 22133 61605
rect 22169 61480 22262 61546
tri 22169 61464 22185 61480 ne
rect 22185 61464 22262 61480
rect 22002 61365 22150 61447
rect 21890 61332 21967 61348
tri 21967 61332 21983 61348 sw
rect 21890 61266 21983 61332
rect 21890 61164 21983 61230
rect 21890 61148 21967 61164
tri 21967 61148 21983 61164 nw
rect 22019 61131 22133 61365
tri 22169 61332 22185 61348 se
rect 22185 61332 22262 61348
rect 22169 61266 22262 61332
rect 22169 61164 22262 61230
tri 22169 61148 22185 61164 ne
rect 22185 61148 22262 61164
rect 22002 61049 22150 61131
rect 21890 61016 21967 61032
tri 21967 61016 21983 61032 sw
rect 21890 60950 21983 61016
rect 22019 60891 22133 61049
tri 22169 61016 22185 61032 se
rect 22185 61016 22262 61032
rect 22169 60950 22262 61016
rect 21890 60815 22262 60891
rect 21890 60690 21983 60756
rect 21890 60674 21967 60690
tri 21967 60674 21983 60690 nw
rect 22019 60657 22133 60815
rect 22169 60690 22262 60756
tri 22169 60674 22185 60690 ne
rect 22185 60674 22262 60690
rect 22002 60575 22150 60657
rect 21890 60542 21967 60558
tri 21967 60542 21983 60558 sw
rect 21890 60476 21983 60542
rect 21890 60374 21983 60440
rect 21890 60358 21967 60374
tri 21967 60358 21983 60374 nw
rect 22019 60341 22133 60575
tri 22169 60542 22185 60558 se
rect 22185 60542 22262 60558
rect 22169 60476 22262 60542
rect 22169 60374 22262 60440
tri 22169 60358 22185 60374 ne
rect 22185 60358 22262 60374
rect 22002 60259 22150 60341
rect 21890 60226 21967 60242
tri 21967 60226 21983 60242 sw
rect 21890 60160 21983 60226
rect 22019 60101 22133 60259
tri 22169 60226 22185 60242 se
rect 22185 60226 22262 60242
rect 22169 60160 22262 60226
rect 21890 60025 22262 60101
rect 21890 59900 21983 59966
rect 21890 59884 21967 59900
tri 21967 59884 21983 59900 nw
rect 22019 59867 22133 60025
rect 22169 59900 22262 59966
tri 22169 59884 22185 59900 ne
rect 22185 59884 22262 59900
rect 22002 59785 22150 59867
rect 21890 59752 21967 59768
tri 21967 59752 21983 59768 sw
rect 21890 59686 21983 59752
rect 21890 59584 21983 59650
rect 21890 59568 21967 59584
tri 21967 59568 21983 59584 nw
rect 22019 59551 22133 59785
tri 22169 59752 22185 59768 se
rect 22185 59752 22262 59768
rect 22169 59686 22262 59752
rect 22169 59584 22262 59650
tri 22169 59568 22185 59584 ne
rect 22185 59568 22262 59584
rect 22002 59469 22150 59551
rect 21890 59436 21967 59452
tri 21967 59436 21983 59452 sw
rect 21890 59370 21983 59436
rect 22019 59311 22133 59469
tri 22169 59436 22185 59452 se
rect 22185 59436 22262 59452
rect 22169 59370 22262 59436
rect 21890 59235 22262 59311
rect 21890 59110 21983 59176
rect 21890 59094 21967 59110
tri 21967 59094 21983 59110 nw
rect 22019 59077 22133 59235
rect 22169 59110 22262 59176
tri 22169 59094 22185 59110 ne
rect 22185 59094 22262 59110
rect 22002 58995 22150 59077
rect 21890 58962 21967 58978
tri 21967 58962 21983 58978 sw
rect 21890 58896 21983 58962
rect 21890 58794 21983 58860
rect 21890 58778 21967 58794
tri 21967 58778 21983 58794 nw
rect 22019 58761 22133 58995
tri 22169 58962 22185 58978 se
rect 22185 58962 22262 58978
rect 22169 58896 22262 58962
rect 22169 58794 22262 58860
tri 22169 58778 22185 58794 ne
rect 22185 58778 22262 58794
rect 22002 58679 22150 58761
rect 21890 58646 21967 58662
tri 21967 58646 21983 58662 sw
rect 21890 58580 21983 58646
rect 22019 58521 22133 58679
tri 22169 58646 22185 58662 se
rect 22185 58646 22262 58662
rect 22169 58580 22262 58646
rect 21890 58445 22262 58521
rect 21890 58320 21983 58386
rect 21890 58304 21967 58320
tri 21967 58304 21983 58320 nw
rect 22019 58287 22133 58445
rect 22169 58320 22262 58386
tri 22169 58304 22185 58320 ne
rect 22185 58304 22262 58320
rect 22002 58205 22150 58287
rect 21890 58172 21967 58188
tri 21967 58172 21983 58188 sw
rect 21890 58106 21983 58172
rect 21890 58004 21983 58070
rect 21890 57988 21967 58004
tri 21967 57988 21983 58004 nw
rect 22019 57971 22133 58205
tri 22169 58172 22185 58188 se
rect 22185 58172 22262 58188
rect 22169 58106 22262 58172
rect 22169 58004 22262 58070
tri 22169 57988 22185 58004 ne
rect 22185 57988 22262 58004
rect 22002 57889 22150 57971
rect 21890 57856 21967 57872
tri 21967 57856 21983 57872 sw
rect 21890 57790 21983 57856
rect 22019 57731 22133 57889
tri 22169 57856 22185 57872 se
rect 22185 57856 22262 57872
rect 22169 57790 22262 57856
rect 21890 57655 22262 57731
rect 21890 57530 21983 57596
rect 21890 57514 21967 57530
tri 21967 57514 21983 57530 nw
rect 22019 57497 22133 57655
rect 22169 57530 22262 57596
tri 22169 57514 22185 57530 ne
rect 22185 57514 22262 57530
rect 22002 57415 22150 57497
rect 21890 57382 21967 57398
tri 21967 57382 21983 57398 sw
rect 21890 57316 21983 57382
rect 21890 57214 21983 57280
rect 21890 57198 21967 57214
tri 21967 57198 21983 57214 nw
rect 22019 57181 22133 57415
tri 22169 57382 22185 57398 se
rect 22185 57382 22262 57398
rect 22169 57316 22262 57382
rect 22169 57214 22262 57280
tri 22169 57198 22185 57214 ne
rect 22185 57198 22262 57214
rect 22002 57099 22150 57181
rect 21890 57066 21967 57082
tri 21967 57066 21983 57082 sw
rect 21890 57000 21983 57066
rect 22019 56941 22133 57099
tri 22169 57066 22185 57082 se
rect 22185 57066 22262 57082
rect 22169 57000 22262 57066
rect 21890 56865 22262 56941
rect 21890 56740 21983 56806
rect 21890 56724 21967 56740
tri 21967 56724 21983 56740 nw
rect 22019 56707 22133 56865
rect 22169 56740 22262 56806
tri 22169 56724 22185 56740 ne
rect 22185 56724 22262 56740
rect 22002 56625 22150 56707
rect 21890 56592 21967 56608
tri 21967 56592 21983 56608 sw
rect 21890 56526 21983 56592
rect 21890 56424 21983 56490
rect 21890 56408 21967 56424
tri 21967 56408 21983 56424 nw
rect 22019 56391 22133 56625
tri 22169 56592 22185 56608 se
rect 22185 56592 22262 56608
rect 22169 56526 22262 56592
rect 22169 56424 22262 56490
tri 22169 56408 22185 56424 ne
rect 22185 56408 22262 56424
rect 22002 56309 22150 56391
rect 21890 56276 21967 56292
tri 21967 56276 21983 56292 sw
rect 21890 56210 21983 56276
rect 22019 56151 22133 56309
tri 22169 56276 22185 56292 se
rect 22185 56276 22262 56292
rect 22169 56210 22262 56276
rect 21890 56075 22262 56151
rect 21890 55950 21983 56016
rect 21890 55934 21967 55950
tri 21967 55934 21983 55950 nw
rect 22019 55917 22133 56075
rect 22169 55950 22262 56016
tri 22169 55934 22185 55950 ne
rect 22185 55934 22262 55950
rect 22002 55835 22150 55917
rect 21890 55802 21967 55818
tri 21967 55802 21983 55818 sw
rect 21890 55736 21983 55802
rect 21890 55634 21983 55700
rect 21890 55618 21967 55634
tri 21967 55618 21983 55634 nw
rect 22019 55601 22133 55835
tri 22169 55802 22185 55818 se
rect 22185 55802 22262 55818
rect 22169 55736 22262 55802
rect 22169 55634 22262 55700
tri 22169 55618 22185 55634 ne
rect 22185 55618 22262 55634
rect 22002 55519 22150 55601
rect 21890 55486 21967 55502
tri 21967 55486 21983 55502 sw
rect 21890 55420 21983 55486
rect 22019 55361 22133 55519
tri 22169 55486 22185 55502 se
rect 22185 55486 22262 55502
rect 22169 55420 22262 55486
rect 21890 55285 22262 55361
rect 21890 55160 21983 55226
rect 21890 55144 21967 55160
tri 21967 55144 21983 55160 nw
rect 22019 55127 22133 55285
rect 22169 55160 22262 55226
tri 22169 55144 22185 55160 ne
rect 22185 55144 22262 55160
rect 22002 55045 22150 55127
rect 21890 55012 21967 55028
tri 21967 55012 21983 55028 sw
rect 21890 54946 21983 55012
rect 21890 54844 21983 54910
rect 21890 54828 21967 54844
tri 21967 54828 21983 54844 nw
rect 22019 54811 22133 55045
tri 22169 55012 22185 55028 se
rect 22185 55012 22262 55028
rect 22169 54946 22262 55012
rect 22169 54844 22262 54910
tri 22169 54828 22185 54844 ne
rect 22185 54828 22262 54844
rect 22002 54729 22150 54811
rect 21890 54696 21967 54712
tri 21967 54696 21983 54712 sw
rect 21890 54630 21983 54696
rect 22019 54571 22133 54729
tri 22169 54696 22185 54712 se
rect 22185 54696 22262 54712
rect 22169 54630 22262 54696
rect 21890 54495 22262 54571
rect 21890 54370 21983 54436
rect 21890 54354 21967 54370
tri 21967 54354 21983 54370 nw
rect 22019 54337 22133 54495
rect 22169 54370 22262 54436
tri 22169 54354 22185 54370 ne
rect 22185 54354 22262 54370
rect 22002 54255 22150 54337
rect 21890 54222 21967 54238
tri 21967 54222 21983 54238 sw
rect 21890 54156 21983 54222
rect 21890 54054 21983 54120
rect 21890 54038 21967 54054
tri 21967 54038 21983 54054 nw
rect 22019 54021 22133 54255
tri 22169 54222 22185 54238 se
rect 22185 54222 22262 54238
rect 22169 54156 22262 54222
rect 22169 54054 22262 54120
tri 22169 54038 22185 54054 ne
rect 22185 54038 22262 54054
rect 22002 53939 22150 54021
rect 21890 53906 21967 53922
tri 21967 53906 21983 53922 sw
rect 21890 53840 21983 53906
rect 22019 53781 22133 53939
tri 22169 53906 22185 53922 se
rect 22185 53906 22262 53922
rect 22169 53840 22262 53906
rect 21890 53705 22262 53781
rect 21890 53580 21983 53646
rect 21890 53564 21967 53580
tri 21967 53564 21983 53580 nw
rect 22019 53547 22133 53705
rect 22169 53580 22262 53646
tri 22169 53564 22185 53580 ne
rect 22185 53564 22262 53580
rect 22002 53465 22150 53547
rect 21890 53432 21967 53448
tri 21967 53432 21983 53448 sw
rect 21890 53366 21983 53432
rect 21890 53264 21983 53330
rect 21890 53248 21967 53264
tri 21967 53248 21983 53264 nw
rect 22019 53231 22133 53465
tri 22169 53432 22185 53448 se
rect 22185 53432 22262 53448
rect 22169 53366 22262 53432
rect 22169 53264 22262 53330
tri 22169 53248 22185 53264 ne
rect 22185 53248 22262 53264
rect 22002 53149 22150 53231
rect 21890 53116 21967 53132
tri 21967 53116 21983 53132 sw
rect 21890 53050 21983 53116
rect 22019 52991 22133 53149
tri 22169 53116 22185 53132 se
rect 22185 53116 22262 53132
rect 22169 53050 22262 53116
rect 21890 52915 22262 52991
rect 21890 52790 21983 52856
rect 21890 52774 21967 52790
tri 21967 52774 21983 52790 nw
rect 22019 52757 22133 52915
rect 22169 52790 22262 52856
tri 22169 52774 22185 52790 ne
rect 22185 52774 22262 52790
rect 22002 52675 22150 52757
rect 21890 52642 21967 52658
tri 21967 52642 21983 52658 sw
rect 21890 52576 21983 52642
rect 21890 52474 21983 52540
rect 21890 52458 21967 52474
tri 21967 52458 21983 52474 nw
rect 22019 52441 22133 52675
tri 22169 52642 22185 52658 se
rect 22185 52642 22262 52658
rect 22169 52576 22262 52642
rect 22169 52474 22262 52540
tri 22169 52458 22185 52474 ne
rect 22185 52458 22262 52474
rect 22002 52359 22150 52441
rect 21890 52326 21967 52342
tri 21967 52326 21983 52342 sw
rect 21890 52260 21983 52326
rect 22019 52201 22133 52359
tri 22169 52326 22185 52342 se
rect 22185 52326 22262 52342
rect 22169 52260 22262 52326
rect 21890 52125 22262 52201
rect 21890 52000 21983 52066
rect 21890 51984 21967 52000
tri 21967 51984 21983 52000 nw
rect 22019 51967 22133 52125
rect 22169 52000 22262 52066
tri 22169 51984 22185 52000 ne
rect 22185 51984 22262 52000
rect 22002 51885 22150 51967
rect 21890 51852 21967 51868
tri 21967 51852 21983 51868 sw
rect 21890 51786 21983 51852
rect 21890 51684 21983 51750
rect 21890 51668 21967 51684
tri 21967 51668 21983 51684 nw
rect 22019 51651 22133 51885
tri 22169 51852 22185 51868 se
rect 22185 51852 22262 51868
rect 22169 51786 22262 51852
rect 22169 51684 22262 51750
tri 22169 51668 22185 51684 ne
rect 22185 51668 22262 51684
rect 22002 51569 22150 51651
rect 21890 51536 21967 51552
tri 21967 51536 21983 51552 sw
rect 21890 51470 21983 51536
rect 22019 51411 22133 51569
tri 22169 51536 22185 51552 se
rect 22185 51536 22262 51552
rect 22169 51470 22262 51536
rect 21890 51335 22262 51411
rect 21890 51210 21983 51276
rect 21890 51194 21967 51210
tri 21967 51194 21983 51210 nw
rect 22019 51177 22133 51335
rect 22169 51210 22262 51276
tri 22169 51194 22185 51210 ne
rect 22185 51194 22262 51210
rect 22002 51095 22150 51177
rect 21890 51062 21967 51078
tri 21967 51062 21983 51078 sw
rect 21890 50996 21983 51062
rect 21890 50894 21983 50960
rect 21890 50878 21967 50894
tri 21967 50878 21983 50894 nw
rect 22019 50861 22133 51095
tri 22169 51062 22185 51078 se
rect 22185 51062 22262 51078
rect 22169 50996 22262 51062
rect 22169 50894 22262 50960
tri 22169 50878 22185 50894 ne
rect 22185 50878 22262 50894
rect 22002 50779 22150 50861
rect 21890 50746 21967 50762
tri 21967 50746 21983 50762 sw
rect 21890 50680 21983 50746
rect 22019 50621 22133 50779
tri 22169 50746 22185 50762 se
rect 22185 50746 22262 50762
rect 22169 50680 22262 50746
rect 21890 50545 22262 50621
rect 21890 50420 21983 50486
rect 21890 50404 21967 50420
tri 21967 50404 21983 50420 nw
rect 22019 50387 22133 50545
rect 22169 50420 22262 50486
tri 22169 50404 22185 50420 ne
rect 22185 50404 22262 50420
rect 22002 50305 22150 50387
rect 21890 50272 21967 50288
tri 21967 50272 21983 50288 sw
rect 21890 50206 21983 50272
rect 21890 50104 21983 50170
rect 21890 50088 21967 50104
tri 21967 50088 21983 50104 nw
rect 22019 50071 22133 50305
tri 22169 50272 22185 50288 se
rect 22185 50272 22262 50288
rect 22169 50206 22262 50272
rect 22169 50104 22262 50170
tri 22169 50088 22185 50104 ne
rect 22185 50088 22262 50104
rect 22002 49989 22150 50071
rect 21890 49956 21967 49972
tri 21967 49956 21983 49972 sw
rect 21890 49890 21983 49956
rect 22019 49831 22133 49989
tri 22169 49956 22185 49972 se
rect 22185 49956 22262 49972
rect 22169 49890 22262 49956
rect 21890 49755 22262 49831
rect 21890 49630 21983 49696
rect 21890 49614 21967 49630
tri 21967 49614 21983 49630 nw
rect 22019 49597 22133 49755
rect 22169 49630 22262 49696
tri 22169 49614 22185 49630 ne
rect 22185 49614 22262 49630
rect 22002 49515 22150 49597
rect 21890 49482 21967 49498
tri 21967 49482 21983 49498 sw
rect 21890 49416 21983 49482
rect 21890 49314 21983 49380
rect 21890 49298 21967 49314
tri 21967 49298 21983 49314 nw
rect 22019 49281 22133 49515
tri 22169 49482 22185 49498 se
rect 22185 49482 22262 49498
rect 22169 49416 22262 49482
rect 22169 49314 22262 49380
tri 22169 49298 22185 49314 ne
rect 22185 49298 22262 49314
rect 22002 49199 22150 49281
rect 21890 49166 21967 49182
tri 21967 49166 21983 49182 sw
rect 21890 49100 21983 49166
rect 22019 49041 22133 49199
tri 22169 49166 22185 49182 se
rect 22185 49166 22262 49182
rect 22169 49100 22262 49166
rect 21890 48965 22262 49041
rect 21890 48840 21983 48906
rect 21890 48824 21967 48840
tri 21967 48824 21983 48840 nw
rect 22019 48807 22133 48965
rect 22169 48840 22262 48906
tri 22169 48824 22185 48840 ne
rect 22185 48824 22262 48840
rect 22002 48725 22150 48807
rect 21890 48692 21967 48708
tri 21967 48692 21983 48708 sw
rect 21890 48626 21983 48692
rect 21890 48524 21983 48590
rect 21890 48508 21967 48524
tri 21967 48508 21983 48524 nw
rect 22019 48491 22133 48725
tri 22169 48692 22185 48708 se
rect 22185 48692 22262 48708
rect 22169 48626 22262 48692
rect 22169 48524 22262 48590
tri 22169 48508 22185 48524 ne
rect 22185 48508 22262 48524
rect 22002 48409 22150 48491
rect 21890 48376 21967 48392
tri 21967 48376 21983 48392 sw
rect 21890 48310 21983 48376
rect 22019 48251 22133 48409
tri 22169 48376 22185 48392 se
rect 22185 48376 22262 48392
rect 22169 48310 22262 48376
rect 21890 48175 22262 48251
rect 21890 48050 21983 48116
rect 21890 48034 21967 48050
tri 21967 48034 21983 48050 nw
rect 22019 48017 22133 48175
rect 22169 48050 22262 48116
tri 22169 48034 22185 48050 ne
rect 22185 48034 22262 48050
rect 22002 47935 22150 48017
rect 21890 47902 21967 47918
tri 21967 47902 21983 47918 sw
rect 21890 47836 21983 47902
rect 21890 47734 21983 47800
rect 21890 47718 21967 47734
tri 21967 47718 21983 47734 nw
rect 22019 47701 22133 47935
tri 22169 47902 22185 47918 se
rect 22185 47902 22262 47918
rect 22169 47836 22262 47902
rect 22169 47734 22262 47800
tri 22169 47718 22185 47734 ne
rect 22185 47718 22262 47734
rect 22002 47619 22150 47701
rect 21890 47586 21967 47602
tri 21967 47586 21983 47602 sw
rect 21890 47520 21983 47586
rect 22019 47461 22133 47619
tri 22169 47586 22185 47602 se
rect 22185 47586 22262 47602
rect 22169 47520 22262 47586
rect 21890 47385 22262 47461
rect 21890 47260 21983 47326
rect 21890 47244 21967 47260
tri 21967 47244 21983 47260 nw
rect 22019 47227 22133 47385
rect 22169 47260 22262 47326
tri 22169 47244 22185 47260 ne
rect 22185 47244 22262 47260
rect 22002 47145 22150 47227
rect 21890 47112 21967 47128
tri 21967 47112 21983 47128 sw
rect 21890 47046 21983 47112
rect 21890 46944 21983 47010
rect 21890 46928 21967 46944
tri 21967 46928 21983 46944 nw
rect 22019 46911 22133 47145
tri 22169 47112 22185 47128 se
rect 22185 47112 22262 47128
rect 22169 47046 22262 47112
rect 22169 46944 22262 47010
tri 22169 46928 22185 46944 ne
rect 22185 46928 22262 46944
rect 22002 46829 22150 46911
rect 21890 46796 21967 46812
tri 21967 46796 21983 46812 sw
rect 21890 46730 21983 46796
rect 22019 46671 22133 46829
tri 22169 46796 22185 46812 se
rect 22185 46796 22262 46812
rect 22169 46730 22262 46796
rect 21890 46595 22262 46671
rect 21890 46470 21983 46536
rect 21890 46454 21967 46470
tri 21967 46454 21983 46470 nw
rect 22019 46437 22133 46595
rect 22169 46470 22262 46536
tri 22169 46454 22185 46470 ne
rect 22185 46454 22262 46470
rect 22002 46355 22150 46437
rect 21890 46322 21967 46338
tri 21967 46322 21983 46338 sw
rect 21890 46256 21983 46322
rect 21890 46154 21983 46220
rect 21890 46138 21967 46154
tri 21967 46138 21983 46154 nw
rect 22019 46121 22133 46355
tri 22169 46322 22185 46338 se
rect 22185 46322 22262 46338
rect 22169 46256 22262 46322
rect 22169 46154 22262 46220
tri 22169 46138 22185 46154 ne
rect 22185 46138 22262 46154
rect 22002 46039 22150 46121
rect 21890 46006 21967 46022
tri 21967 46006 21983 46022 sw
rect 21890 45940 21983 46006
rect 22019 45881 22133 46039
tri 22169 46006 22185 46022 se
rect 22185 46006 22262 46022
rect 22169 45940 22262 46006
rect 21890 45805 22262 45881
rect 21890 45680 21983 45746
rect 21890 45664 21967 45680
tri 21967 45664 21983 45680 nw
rect 22019 45647 22133 45805
rect 22169 45680 22262 45746
tri 22169 45664 22185 45680 ne
rect 22185 45664 22262 45680
rect 22002 45565 22150 45647
rect 21890 45532 21967 45548
tri 21967 45532 21983 45548 sw
rect 21890 45466 21983 45532
rect 21890 45364 21983 45430
rect 21890 45348 21967 45364
tri 21967 45348 21983 45364 nw
rect 22019 45331 22133 45565
tri 22169 45532 22185 45548 se
rect 22185 45532 22262 45548
rect 22169 45466 22262 45532
rect 22169 45364 22262 45430
tri 22169 45348 22185 45364 ne
rect 22185 45348 22262 45364
rect 22002 45249 22150 45331
rect 21890 45216 21967 45232
tri 21967 45216 21983 45232 sw
rect 21890 45150 21983 45216
rect 22019 45091 22133 45249
tri 22169 45216 22185 45232 se
rect 22185 45216 22262 45232
rect 22169 45150 22262 45216
rect 21890 45015 22262 45091
rect 21890 44890 21983 44956
rect 21890 44874 21967 44890
tri 21967 44874 21983 44890 nw
rect 22019 44857 22133 45015
rect 22169 44890 22262 44956
tri 22169 44874 22185 44890 ne
rect 22185 44874 22262 44890
rect 22002 44775 22150 44857
rect 21890 44742 21967 44758
tri 21967 44742 21983 44758 sw
rect 21890 44676 21983 44742
rect 21890 44574 21983 44640
rect 21890 44558 21967 44574
tri 21967 44558 21983 44574 nw
rect 22019 44541 22133 44775
tri 22169 44742 22185 44758 se
rect 22185 44742 22262 44758
rect 22169 44676 22262 44742
rect 22169 44574 22262 44640
tri 22169 44558 22185 44574 ne
rect 22185 44558 22262 44574
rect 22002 44459 22150 44541
rect 21890 44426 21967 44442
tri 21967 44426 21983 44442 sw
rect 21890 44360 21983 44426
rect 22019 44301 22133 44459
tri 22169 44426 22185 44442 se
rect 22185 44426 22262 44442
rect 22169 44360 22262 44426
rect 21890 44225 22262 44301
rect 21890 44100 21983 44166
rect 21890 44084 21967 44100
tri 21967 44084 21983 44100 nw
rect 22019 44067 22133 44225
rect 22169 44100 22262 44166
tri 22169 44084 22185 44100 ne
rect 22185 44084 22262 44100
rect 22002 43985 22150 44067
rect 21890 43952 21967 43968
tri 21967 43952 21983 43968 sw
rect 21890 43886 21983 43952
rect 21890 43784 21983 43850
rect 21890 43768 21967 43784
tri 21967 43768 21983 43784 nw
rect 22019 43751 22133 43985
tri 22169 43952 22185 43968 se
rect 22185 43952 22262 43968
rect 22169 43886 22262 43952
rect 22169 43784 22262 43850
tri 22169 43768 22185 43784 ne
rect 22185 43768 22262 43784
rect 22002 43669 22150 43751
rect 21890 43636 21967 43652
tri 21967 43636 21983 43652 sw
rect 21890 43570 21983 43636
rect 22019 43511 22133 43669
tri 22169 43636 22185 43652 se
rect 22185 43636 22262 43652
rect 22169 43570 22262 43636
rect 21890 43435 22262 43511
rect 21890 43310 21983 43376
rect 21890 43294 21967 43310
tri 21967 43294 21983 43310 nw
rect 22019 43277 22133 43435
rect 22169 43310 22262 43376
tri 22169 43294 22185 43310 ne
rect 22185 43294 22262 43310
rect 22002 43195 22150 43277
rect 21890 43162 21967 43178
tri 21967 43162 21983 43178 sw
rect 21890 43096 21983 43162
rect 21890 42994 21983 43060
rect 21890 42978 21967 42994
tri 21967 42978 21983 42994 nw
rect 22019 42961 22133 43195
tri 22169 43162 22185 43178 se
rect 22185 43162 22262 43178
rect 22169 43096 22262 43162
rect 22169 42994 22262 43060
tri 22169 42978 22185 42994 ne
rect 22185 42978 22262 42994
rect 22002 42879 22150 42961
rect 21890 42846 21967 42862
tri 21967 42846 21983 42862 sw
rect 21890 42780 21983 42846
rect 22019 42721 22133 42879
tri 22169 42846 22185 42862 se
rect 22185 42846 22262 42862
rect 22169 42780 22262 42846
rect 21890 42645 22262 42721
rect 21890 42520 21983 42586
rect 21890 42504 21967 42520
tri 21967 42504 21983 42520 nw
rect 22019 42487 22133 42645
rect 22169 42520 22262 42586
tri 22169 42504 22185 42520 ne
rect 22185 42504 22262 42520
rect 22002 42405 22150 42487
rect 21890 42372 21967 42388
tri 21967 42372 21983 42388 sw
rect 21890 42306 21983 42372
rect 21890 42204 21983 42270
rect 21890 42188 21967 42204
tri 21967 42188 21983 42204 nw
rect 22019 42171 22133 42405
tri 22169 42372 22185 42388 se
rect 22185 42372 22262 42388
rect 22169 42306 22262 42372
rect 22169 42204 22262 42270
tri 22169 42188 22185 42204 ne
rect 22185 42188 22262 42204
rect 22002 42089 22150 42171
rect 21890 42056 21967 42072
tri 21967 42056 21983 42072 sw
rect 21890 41990 21983 42056
rect 22019 41931 22133 42089
tri 22169 42056 22185 42072 se
rect 22185 42056 22262 42072
rect 22169 41990 22262 42056
rect 21890 41855 22262 41931
rect 21890 41730 21983 41796
rect 21890 41714 21967 41730
tri 21967 41714 21983 41730 nw
rect 22019 41697 22133 41855
rect 22169 41730 22262 41796
tri 22169 41714 22185 41730 ne
rect 22185 41714 22262 41730
rect 22002 41615 22150 41697
rect 21890 41582 21967 41598
tri 21967 41582 21983 41598 sw
rect 21890 41516 21983 41582
rect 21890 41414 21983 41480
rect 21890 41398 21967 41414
tri 21967 41398 21983 41414 nw
rect 22019 41381 22133 41615
tri 22169 41582 22185 41598 se
rect 22185 41582 22262 41598
rect 22169 41516 22262 41582
rect 22169 41414 22262 41480
tri 22169 41398 22185 41414 ne
rect 22185 41398 22262 41414
rect 22002 41299 22150 41381
rect 21890 41266 21967 41282
tri 21967 41266 21983 41282 sw
rect 21890 41200 21983 41266
rect 22019 41141 22133 41299
tri 22169 41266 22185 41282 se
rect 22185 41266 22262 41282
rect 22169 41200 22262 41266
rect 21890 41065 22262 41141
rect 21890 40940 21983 41006
rect 21890 40924 21967 40940
tri 21967 40924 21983 40940 nw
rect 22019 40907 22133 41065
rect 22169 40940 22262 41006
tri 22169 40924 22185 40940 ne
rect 22185 40924 22262 40940
rect 22002 40825 22150 40907
rect 21890 40792 21967 40808
tri 21967 40792 21983 40808 sw
rect 21890 40726 21983 40792
rect 21890 40624 21983 40690
rect 21890 40608 21967 40624
tri 21967 40608 21983 40624 nw
rect 22019 40591 22133 40825
tri 22169 40792 22185 40808 se
rect 22185 40792 22262 40808
rect 22169 40726 22262 40792
rect 22169 40624 22262 40690
tri 22169 40608 22185 40624 ne
rect 22185 40608 22262 40624
rect 22002 40509 22150 40591
rect 21890 40476 21967 40492
tri 21967 40476 21983 40492 sw
rect 21890 40410 21983 40476
rect 22019 40351 22133 40509
tri 22169 40476 22185 40492 se
rect 22185 40476 22262 40492
rect 22169 40410 22262 40476
rect 21890 40275 22262 40351
rect 21890 40150 21983 40216
rect 21890 40134 21967 40150
tri 21967 40134 21983 40150 nw
rect 22019 40117 22133 40275
rect 22169 40150 22262 40216
tri 22169 40134 22185 40150 ne
rect 22185 40134 22262 40150
rect 22002 40035 22150 40117
rect 21890 40002 21967 40018
tri 21967 40002 21983 40018 sw
rect 21890 39936 21983 40002
rect 21890 39834 21983 39900
rect 21890 39818 21967 39834
tri 21967 39818 21983 39834 nw
rect 22019 39801 22133 40035
tri 22169 40002 22185 40018 se
rect 22185 40002 22262 40018
rect 22169 39936 22262 40002
rect 22169 39834 22262 39900
tri 22169 39818 22185 39834 ne
rect 22185 39818 22262 39834
rect 22002 39719 22150 39801
rect 21890 39686 21967 39702
tri 21967 39686 21983 39702 sw
rect 21890 39620 21983 39686
rect 22019 39561 22133 39719
tri 22169 39686 22185 39702 se
rect 22185 39686 22262 39702
rect 22169 39620 22262 39686
rect 21890 39485 22262 39561
rect 21890 39360 21983 39426
rect 21890 39344 21967 39360
tri 21967 39344 21983 39360 nw
rect 22019 39327 22133 39485
rect 22169 39360 22262 39426
tri 22169 39344 22185 39360 ne
rect 22185 39344 22262 39360
rect 22002 39245 22150 39327
rect 21890 39212 21967 39228
tri 21967 39212 21983 39228 sw
rect 21890 39146 21983 39212
rect 21890 39044 21983 39110
rect 21890 39028 21967 39044
tri 21967 39028 21983 39044 nw
rect 22019 39011 22133 39245
tri 22169 39212 22185 39228 se
rect 22185 39212 22262 39228
rect 22169 39146 22262 39212
rect 22169 39044 22262 39110
tri 22169 39028 22185 39044 ne
rect 22185 39028 22262 39044
rect 22002 38929 22150 39011
rect 21890 38896 21967 38912
tri 21967 38896 21983 38912 sw
rect 21890 38830 21983 38896
rect 22019 38771 22133 38929
tri 22169 38896 22185 38912 se
rect 22185 38896 22262 38912
rect 22169 38830 22262 38896
rect 21890 38695 22262 38771
rect 21890 38570 21983 38636
rect 21890 38554 21967 38570
tri 21967 38554 21983 38570 nw
rect 22019 38537 22133 38695
rect 22169 38570 22262 38636
tri 22169 38554 22185 38570 ne
rect 22185 38554 22262 38570
rect 22002 38455 22150 38537
rect 21890 38422 21967 38438
tri 21967 38422 21983 38438 sw
rect 21890 38356 21983 38422
rect 21890 38254 21983 38320
rect 21890 38238 21967 38254
tri 21967 38238 21983 38254 nw
rect 22019 38221 22133 38455
tri 22169 38422 22185 38438 se
rect 22185 38422 22262 38438
rect 22169 38356 22262 38422
rect 22169 38254 22262 38320
tri 22169 38238 22185 38254 ne
rect 22185 38238 22262 38254
rect 22002 38139 22150 38221
rect 21890 38106 21967 38122
tri 21967 38106 21983 38122 sw
rect 21890 38040 21983 38106
rect 22019 37981 22133 38139
tri 22169 38106 22185 38122 se
rect 22185 38106 22262 38122
rect 22169 38040 22262 38106
rect 21890 37905 22262 37981
rect 21890 37780 21983 37846
rect 21890 37764 21967 37780
tri 21967 37764 21983 37780 nw
rect 22019 37747 22133 37905
rect 22169 37780 22262 37846
tri 22169 37764 22185 37780 ne
rect 22185 37764 22262 37780
rect 22002 37665 22150 37747
rect 21890 37632 21967 37648
tri 21967 37632 21983 37648 sw
rect 21890 37566 21983 37632
rect 21890 37464 21983 37530
rect 21890 37448 21967 37464
tri 21967 37448 21983 37464 nw
rect 22019 37431 22133 37665
tri 22169 37632 22185 37648 se
rect 22185 37632 22262 37648
rect 22169 37566 22262 37632
rect 22169 37464 22262 37530
tri 22169 37448 22185 37464 ne
rect 22185 37448 22262 37464
rect 22002 37349 22150 37431
rect 21890 37316 21967 37332
tri 21967 37316 21983 37332 sw
rect 21890 37250 21983 37316
rect 22019 37191 22133 37349
tri 22169 37316 22185 37332 se
rect 22185 37316 22262 37332
rect 22169 37250 22262 37316
rect 21890 37115 22262 37191
rect 21890 36990 21983 37056
rect 21890 36974 21967 36990
tri 21967 36974 21983 36990 nw
rect 22019 36957 22133 37115
rect 22169 36990 22262 37056
tri 22169 36974 22185 36990 ne
rect 22185 36974 22262 36990
rect 22002 36875 22150 36957
rect 21890 36842 21967 36858
tri 21967 36842 21983 36858 sw
rect 21890 36776 21983 36842
rect 21890 36674 21983 36740
rect 21890 36658 21967 36674
tri 21967 36658 21983 36674 nw
rect 22019 36641 22133 36875
tri 22169 36842 22185 36858 se
rect 22185 36842 22262 36858
rect 22169 36776 22262 36842
rect 22169 36674 22262 36740
tri 22169 36658 22185 36674 ne
rect 22185 36658 22262 36674
rect 22002 36559 22150 36641
rect 21890 36526 21967 36542
tri 21967 36526 21983 36542 sw
rect 21890 36460 21983 36526
rect 22019 36401 22133 36559
tri 22169 36526 22185 36542 se
rect 22185 36526 22262 36542
rect 22169 36460 22262 36526
rect 21890 36325 22262 36401
rect 21890 36200 21983 36266
rect 21890 36184 21967 36200
tri 21967 36184 21983 36200 nw
rect 22019 36167 22133 36325
rect 22169 36200 22262 36266
tri 22169 36184 22185 36200 ne
rect 22185 36184 22262 36200
rect 22002 36085 22150 36167
rect 21890 36052 21967 36068
tri 21967 36052 21983 36068 sw
rect 21890 35986 21983 36052
rect 21890 35884 21983 35950
rect 21890 35868 21967 35884
tri 21967 35868 21983 35884 nw
rect 22019 35851 22133 36085
tri 22169 36052 22185 36068 se
rect 22185 36052 22262 36068
rect 22169 35986 22262 36052
rect 22169 35884 22262 35950
tri 22169 35868 22185 35884 ne
rect 22185 35868 22262 35884
rect 22002 35769 22150 35851
rect 21890 35736 21967 35752
tri 21967 35736 21983 35752 sw
rect 21890 35670 21983 35736
rect 22019 35611 22133 35769
tri 22169 35736 22185 35752 se
rect 22185 35736 22262 35752
rect 22169 35670 22262 35736
rect 21890 35535 22262 35611
rect 21890 35410 21983 35476
rect 21890 35394 21967 35410
tri 21967 35394 21983 35410 nw
rect 22019 35377 22133 35535
rect 22169 35410 22262 35476
tri 22169 35394 22185 35410 ne
rect 22185 35394 22262 35410
rect 22002 35295 22150 35377
rect 21890 35262 21967 35278
tri 21967 35262 21983 35278 sw
rect 21890 35196 21983 35262
rect 21890 35094 21983 35160
rect 21890 35078 21967 35094
tri 21967 35078 21983 35094 nw
rect 22019 35061 22133 35295
tri 22169 35262 22185 35278 se
rect 22185 35262 22262 35278
rect 22169 35196 22262 35262
rect 22169 35094 22262 35160
tri 22169 35078 22185 35094 ne
rect 22185 35078 22262 35094
rect 22002 34979 22150 35061
rect 21890 34946 21967 34962
tri 21967 34946 21983 34962 sw
rect 21890 34880 21983 34946
rect 22019 34821 22133 34979
tri 22169 34946 22185 34962 se
rect 22185 34946 22262 34962
rect 22169 34880 22262 34946
rect 21890 34745 22262 34821
rect 21890 34620 21983 34686
rect 21890 34604 21967 34620
tri 21967 34604 21983 34620 nw
rect 22019 34587 22133 34745
rect 22169 34620 22262 34686
tri 22169 34604 22185 34620 ne
rect 22185 34604 22262 34620
rect 22002 34505 22150 34587
rect 21890 34472 21967 34488
tri 21967 34472 21983 34488 sw
rect 21890 34406 21983 34472
rect 21890 34304 21983 34370
rect 21890 34288 21967 34304
tri 21967 34288 21983 34304 nw
rect 22019 34271 22133 34505
tri 22169 34472 22185 34488 se
rect 22185 34472 22262 34488
rect 22169 34406 22262 34472
rect 22169 34304 22262 34370
tri 22169 34288 22185 34304 ne
rect 22185 34288 22262 34304
rect 22002 34189 22150 34271
rect 21890 34156 21967 34172
tri 21967 34156 21983 34172 sw
rect 21890 34090 21983 34156
rect 22019 34031 22133 34189
tri 22169 34156 22185 34172 se
rect 22185 34156 22262 34172
rect 22169 34090 22262 34156
rect 21890 33955 22262 34031
rect 21890 33830 21983 33896
rect 21890 33814 21967 33830
tri 21967 33814 21983 33830 nw
rect 22019 33797 22133 33955
rect 22169 33830 22262 33896
tri 22169 33814 22185 33830 ne
rect 22185 33814 22262 33830
rect 22002 33715 22150 33797
rect 21890 33682 21967 33698
tri 21967 33682 21983 33698 sw
rect 21890 33616 21983 33682
rect 21890 33514 21983 33580
rect 21890 33498 21967 33514
tri 21967 33498 21983 33514 nw
rect 22019 33481 22133 33715
tri 22169 33682 22185 33698 se
rect 22185 33682 22262 33698
rect 22169 33616 22262 33682
rect 22169 33514 22262 33580
tri 22169 33498 22185 33514 ne
rect 22185 33498 22262 33514
rect 22002 33399 22150 33481
rect 21890 33366 21967 33382
tri 21967 33366 21983 33382 sw
rect 21890 33300 21983 33366
rect 22019 33241 22133 33399
tri 22169 33366 22185 33382 se
rect 22185 33366 22262 33382
rect 22169 33300 22262 33366
rect 21890 33165 22262 33241
rect 21890 33040 21983 33106
rect 21890 33024 21967 33040
tri 21967 33024 21983 33040 nw
rect 22019 33007 22133 33165
rect 22169 33040 22262 33106
tri 22169 33024 22185 33040 ne
rect 22185 33024 22262 33040
rect 22002 32925 22150 33007
rect 21890 32892 21967 32908
tri 21967 32892 21983 32908 sw
rect 21890 32826 21983 32892
rect 21890 32724 21983 32790
rect 21890 32708 21967 32724
tri 21967 32708 21983 32724 nw
rect 22019 32691 22133 32925
tri 22169 32892 22185 32908 se
rect 22185 32892 22262 32908
rect 22169 32826 22262 32892
rect 22169 32724 22262 32790
tri 22169 32708 22185 32724 ne
rect 22185 32708 22262 32724
rect 22002 32609 22150 32691
rect 21890 32576 21967 32592
tri 21967 32576 21983 32592 sw
rect 21890 32510 21983 32576
rect 22019 32451 22133 32609
tri 22169 32576 22185 32592 se
rect 22185 32576 22262 32592
rect 22169 32510 22262 32576
rect 21890 32375 22262 32451
rect 21890 32250 21983 32316
rect 21890 32234 21967 32250
tri 21967 32234 21983 32250 nw
rect 22019 32217 22133 32375
rect 22169 32250 22262 32316
tri 22169 32234 22185 32250 ne
rect 22185 32234 22262 32250
rect 22002 32135 22150 32217
rect 21890 32102 21967 32118
tri 21967 32102 21983 32118 sw
rect 21890 32036 21983 32102
rect 21890 31934 21983 32000
rect 21890 31918 21967 31934
tri 21967 31918 21983 31934 nw
rect 22019 31901 22133 32135
tri 22169 32102 22185 32118 se
rect 22185 32102 22262 32118
rect 22169 32036 22262 32102
rect 22169 31934 22262 32000
tri 22169 31918 22185 31934 ne
rect 22185 31918 22262 31934
rect 22002 31819 22150 31901
rect 21890 31786 21967 31802
tri 21967 31786 21983 31802 sw
rect 21890 31720 21983 31786
rect 22019 31661 22133 31819
tri 22169 31786 22185 31802 se
rect 22185 31786 22262 31802
rect 22169 31720 22262 31786
rect 21890 31585 22262 31661
rect 21890 31460 21983 31526
rect 21890 31444 21967 31460
tri 21967 31444 21983 31460 nw
rect 22019 31427 22133 31585
rect 22169 31460 22262 31526
tri 22169 31444 22185 31460 ne
rect 22185 31444 22262 31460
rect 22002 31345 22150 31427
rect 21890 31312 21967 31328
tri 21967 31312 21983 31328 sw
rect 21890 31246 21983 31312
rect 21890 31144 21983 31210
rect 21890 31128 21967 31144
tri 21967 31128 21983 31144 nw
rect 22019 31111 22133 31345
tri 22169 31312 22185 31328 se
rect 22185 31312 22262 31328
rect 22169 31246 22262 31312
rect 22169 31144 22262 31210
tri 22169 31128 22185 31144 ne
rect 22185 31128 22262 31144
rect 22002 31029 22150 31111
rect 21890 30996 21967 31012
tri 21967 30996 21983 31012 sw
rect 21890 30930 21983 30996
rect 22019 30871 22133 31029
tri 22169 30996 22185 31012 se
rect 22185 30996 22262 31012
rect 22169 30930 22262 30996
rect 21890 30795 22262 30871
rect 21890 30670 21983 30736
rect 21890 30654 21967 30670
tri 21967 30654 21983 30670 nw
rect 22019 30637 22133 30795
rect 22169 30670 22262 30736
tri 22169 30654 22185 30670 ne
rect 22185 30654 22262 30670
rect 22002 30555 22150 30637
rect 21890 30522 21967 30538
tri 21967 30522 21983 30538 sw
rect 21890 30456 21983 30522
rect 21890 30354 21983 30420
rect 21890 30338 21967 30354
tri 21967 30338 21983 30354 nw
rect 22019 30321 22133 30555
tri 22169 30522 22185 30538 se
rect 22185 30522 22262 30538
rect 22169 30456 22262 30522
rect 22169 30354 22262 30420
tri 22169 30338 22185 30354 ne
rect 22185 30338 22262 30354
rect 22002 30239 22150 30321
rect 21890 30206 21967 30222
tri 21967 30206 21983 30222 sw
rect 21890 30140 21983 30206
rect 22019 30081 22133 30239
tri 22169 30206 22185 30222 se
rect 22185 30206 22262 30222
rect 22169 30140 22262 30206
rect 21890 30005 22262 30081
rect 21890 29880 21983 29946
rect 21890 29864 21967 29880
tri 21967 29864 21983 29880 nw
rect 22019 29847 22133 30005
rect 22169 29880 22262 29946
tri 22169 29864 22185 29880 ne
rect 22185 29864 22262 29880
rect 22002 29765 22150 29847
rect 21890 29732 21967 29748
tri 21967 29732 21983 29748 sw
rect 21890 29666 21983 29732
rect 21890 29564 21983 29630
rect 21890 29548 21967 29564
tri 21967 29548 21983 29564 nw
rect 22019 29531 22133 29765
tri 22169 29732 22185 29748 se
rect 22185 29732 22262 29748
rect 22169 29666 22262 29732
rect 22169 29564 22262 29630
tri 22169 29548 22185 29564 ne
rect 22185 29548 22262 29564
rect 22002 29449 22150 29531
rect 21890 29416 21967 29432
tri 21967 29416 21983 29432 sw
rect 21890 29350 21983 29416
rect 22019 29291 22133 29449
tri 22169 29416 22185 29432 se
rect 22185 29416 22262 29432
rect 22169 29350 22262 29416
rect 21890 29215 22262 29291
rect 21890 29090 21983 29156
rect 21890 29074 21967 29090
tri 21967 29074 21983 29090 nw
rect 22019 29057 22133 29215
rect 22169 29090 22262 29156
tri 22169 29074 22185 29090 ne
rect 22185 29074 22262 29090
rect 22002 28975 22150 29057
rect 21890 28942 21967 28958
tri 21967 28942 21983 28958 sw
rect 21890 28876 21983 28942
rect 22019 28833 22133 28975
tri 22169 28942 22185 28958 se
rect 22185 28942 22262 28958
rect 22169 28876 22262 28942
rect 22298 28463 22334 80603
rect 22370 28463 22406 80603
rect 22442 80445 22478 80603
rect 22434 80303 22486 80445
rect 22442 28763 22478 80303
rect 22434 28621 22486 28763
rect 22442 28463 22478 28621
rect 22514 28463 22550 80603
rect 22586 28463 22622 80603
rect 22658 28833 22742 80233
rect 22778 28463 22814 80603
rect 22850 28463 22886 80603
rect 22922 80445 22958 80603
rect 22914 80303 22966 80445
rect 22922 28763 22958 80303
rect 22914 28621 22966 28763
rect 22922 28463 22958 28621
rect 22994 28463 23030 80603
rect 23066 28463 23102 80603
rect 23138 80124 23231 80190
rect 23138 80108 23215 80124
tri 23215 80108 23231 80124 nw
rect 23267 80091 23381 80233
rect 23417 80124 23510 80190
tri 23417 80108 23433 80124 ne
rect 23433 80108 23510 80124
rect 23250 80009 23398 80091
rect 23138 79976 23215 79992
tri 23215 79976 23231 79992 sw
rect 23138 79910 23231 79976
rect 23267 79851 23381 80009
tri 23417 79976 23433 79992 se
rect 23433 79976 23510 79992
rect 23417 79910 23510 79976
rect 23138 79775 23510 79851
rect 23138 79650 23231 79716
rect 23138 79634 23215 79650
tri 23215 79634 23231 79650 nw
rect 23267 79617 23381 79775
rect 23417 79650 23510 79716
tri 23417 79634 23433 79650 ne
rect 23433 79634 23510 79650
rect 23250 79535 23398 79617
rect 23138 79502 23215 79518
tri 23215 79502 23231 79518 sw
rect 23138 79436 23231 79502
rect 23138 79334 23231 79400
rect 23138 79318 23215 79334
tri 23215 79318 23231 79334 nw
rect 23267 79301 23381 79535
tri 23417 79502 23433 79518 se
rect 23433 79502 23510 79518
rect 23417 79436 23510 79502
rect 23417 79334 23510 79400
tri 23417 79318 23433 79334 ne
rect 23433 79318 23510 79334
rect 23250 79219 23398 79301
rect 23138 79186 23215 79202
tri 23215 79186 23231 79202 sw
rect 23138 79120 23231 79186
rect 23267 79061 23381 79219
tri 23417 79186 23433 79202 se
rect 23433 79186 23510 79202
rect 23417 79120 23510 79186
rect 23138 78985 23510 79061
rect 23138 78860 23231 78926
rect 23138 78844 23215 78860
tri 23215 78844 23231 78860 nw
rect 23267 78827 23381 78985
rect 23417 78860 23510 78926
tri 23417 78844 23433 78860 ne
rect 23433 78844 23510 78860
rect 23250 78745 23398 78827
rect 23138 78712 23215 78728
tri 23215 78712 23231 78728 sw
rect 23138 78646 23231 78712
rect 23138 78544 23231 78610
rect 23138 78528 23215 78544
tri 23215 78528 23231 78544 nw
rect 23267 78511 23381 78745
tri 23417 78712 23433 78728 se
rect 23433 78712 23510 78728
rect 23417 78646 23510 78712
rect 23417 78544 23510 78610
tri 23417 78528 23433 78544 ne
rect 23433 78528 23510 78544
rect 23250 78429 23398 78511
rect 23138 78396 23215 78412
tri 23215 78396 23231 78412 sw
rect 23138 78330 23231 78396
rect 23267 78271 23381 78429
tri 23417 78396 23433 78412 se
rect 23433 78396 23510 78412
rect 23417 78330 23510 78396
rect 23138 78195 23510 78271
rect 23138 78070 23231 78136
rect 23138 78054 23215 78070
tri 23215 78054 23231 78070 nw
rect 23267 78037 23381 78195
rect 23417 78070 23510 78136
tri 23417 78054 23433 78070 ne
rect 23433 78054 23510 78070
rect 23250 77955 23398 78037
rect 23138 77922 23215 77938
tri 23215 77922 23231 77938 sw
rect 23138 77856 23231 77922
rect 23138 77754 23231 77820
rect 23138 77738 23215 77754
tri 23215 77738 23231 77754 nw
rect 23267 77721 23381 77955
tri 23417 77922 23433 77938 se
rect 23433 77922 23510 77938
rect 23417 77856 23510 77922
rect 23417 77754 23510 77820
tri 23417 77738 23433 77754 ne
rect 23433 77738 23510 77754
rect 23250 77639 23398 77721
rect 23138 77606 23215 77622
tri 23215 77606 23231 77622 sw
rect 23138 77540 23231 77606
rect 23267 77481 23381 77639
tri 23417 77606 23433 77622 se
rect 23433 77606 23510 77622
rect 23417 77540 23510 77606
rect 23138 77405 23510 77481
rect 23138 77280 23231 77346
rect 23138 77264 23215 77280
tri 23215 77264 23231 77280 nw
rect 23267 77247 23381 77405
rect 23417 77280 23510 77346
tri 23417 77264 23433 77280 ne
rect 23433 77264 23510 77280
rect 23250 77165 23398 77247
rect 23138 77132 23215 77148
tri 23215 77132 23231 77148 sw
rect 23138 77066 23231 77132
rect 23138 76964 23231 77030
rect 23138 76948 23215 76964
tri 23215 76948 23231 76964 nw
rect 23267 76931 23381 77165
tri 23417 77132 23433 77148 se
rect 23433 77132 23510 77148
rect 23417 77066 23510 77132
rect 23417 76964 23510 77030
tri 23417 76948 23433 76964 ne
rect 23433 76948 23510 76964
rect 23250 76849 23398 76931
rect 23138 76816 23215 76832
tri 23215 76816 23231 76832 sw
rect 23138 76750 23231 76816
rect 23267 76691 23381 76849
tri 23417 76816 23433 76832 se
rect 23433 76816 23510 76832
rect 23417 76750 23510 76816
rect 23138 76615 23510 76691
rect 23138 76490 23231 76556
rect 23138 76474 23215 76490
tri 23215 76474 23231 76490 nw
rect 23267 76457 23381 76615
rect 23417 76490 23510 76556
tri 23417 76474 23433 76490 ne
rect 23433 76474 23510 76490
rect 23250 76375 23398 76457
rect 23138 76342 23215 76358
tri 23215 76342 23231 76358 sw
rect 23138 76276 23231 76342
rect 23138 76174 23231 76240
rect 23138 76158 23215 76174
tri 23215 76158 23231 76174 nw
rect 23267 76141 23381 76375
tri 23417 76342 23433 76358 se
rect 23433 76342 23510 76358
rect 23417 76276 23510 76342
rect 23417 76174 23510 76240
tri 23417 76158 23433 76174 ne
rect 23433 76158 23510 76174
rect 23250 76059 23398 76141
rect 23138 76026 23215 76042
tri 23215 76026 23231 76042 sw
rect 23138 75960 23231 76026
rect 23267 75901 23381 76059
tri 23417 76026 23433 76042 se
rect 23433 76026 23510 76042
rect 23417 75960 23510 76026
rect 23138 75825 23510 75901
rect 23138 75700 23231 75766
rect 23138 75684 23215 75700
tri 23215 75684 23231 75700 nw
rect 23267 75667 23381 75825
rect 23417 75700 23510 75766
tri 23417 75684 23433 75700 ne
rect 23433 75684 23510 75700
rect 23250 75585 23398 75667
rect 23138 75552 23215 75568
tri 23215 75552 23231 75568 sw
rect 23138 75486 23231 75552
rect 23138 75384 23231 75450
rect 23138 75368 23215 75384
tri 23215 75368 23231 75384 nw
rect 23267 75351 23381 75585
tri 23417 75552 23433 75568 se
rect 23433 75552 23510 75568
rect 23417 75486 23510 75552
rect 23417 75384 23510 75450
tri 23417 75368 23433 75384 ne
rect 23433 75368 23510 75384
rect 23250 75269 23398 75351
rect 23138 75236 23215 75252
tri 23215 75236 23231 75252 sw
rect 23138 75170 23231 75236
rect 23267 75111 23381 75269
tri 23417 75236 23433 75252 se
rect 23433 75236 23510 75252
rect 23417 75170 23510 75236
rect 23138 75035 23510 75111
rect 23138 74910 23231 74976
rect 23138 74894 23215 74910
tri 23215 74894 23231 74910 nw
rect 23267 74877 23381 75035
rect 23417 74910 23510 74976
tri 23417 74894 23433 74910 ne
rect 23433 74894 23510 74910
rect 23250 74795 23398 74877
rect 23138 74762 23215 74778
tri 23215 74762 23231 74778 sw
rect 23138 74696 23231 74762
rect 23138 74594 23231 74660
rect 23138 74578 23215 74594
tri 23215 74578 23231 74594 nw
rect 23267 74561 23381 74795
tri 23417 74762 23433 74778 se
rect 23433 74762 23510 74778
rect 23417 74696 23510 74762
rect 23417 74594 23510 74660
tri 23417 74578 23433 74594 ne
rect 23433 74578 23510 74594
rect 23250 74479 23398 74561
rect 23138 74446 23215 74462
tri 23215 74446 23231 74462 sw
rect 23138 74380 23231 74446
rect 23267 74321 23381 74479
tri 23417 74446 23433 74462 se
rect 23433 74446 23510 74462
rect 23417 74380 23510 74446
rect 23138 74245 23510 74321
rect 23138 74120 23231 74186
rect 23138 74104 23215 74120
tri 23215 74104 23231 74120 nw
rect 23267 74087 23381 74245
rect 23417 74120 23510 74186
tri 23417 74104 23433 74120 ne
rect 23433 74104 23510 74120
rect 23250 74005 23398 74087
rect 23138 73972 23215 73988
tri 23215 73972 23231 73988 sw
rect 23138 73906 23231 73972
rect 23138 73804 23231 73870
rect 23138 73788 23215 73804
tri 23215 73788 23231 73804 nw
rect 23267 73771 23381 74005
tri 23417 73972 23433 73988 se
rect 23433 73972 23510 73988
rect 23417 73906 23510 73972
rect 23417 73804 23510 73870
tri 23417 73788 23433 73804 ne
rect 23433 73788 23510 73804
rect 23250 73689 23398 73771
rect 23138 73656 23215 73672
tri 23215 73656 23231 73672 sw
rect 23138 73590 23231 73656
rect 23267 73531 23381 73689
tri 23417 73656 23433 73672 se
rect 23433 73656 23510 73672
rect 23417 73590 23510 73656
rect 23138 73455 23510 73531
rect 23138 73330 23231 73396
rect 23138 73314 23215 73330
tri 23215 73314 23231 73330 nw
rect 23267 73297 23381 73455
rect 23417 73330 23510 73396
tri 23417 73314 23433 73330 ne
rect 23433 73314 23510 73330
rect 23250 73215 23398 73297
rect 23138 73182 23215 73198
tri 23215 73182 23231 73198 sw
rect 23138 73116 23231 73182
rect 23138 73014 23231 73080
rect 23138 72998 23215 73014
tri 23215 72998 23231 73014 nw
rect 23267 72981 23381 73215
tri 23417 73182 23433 73198 se
rect 23433 73182 23510 73198
rect 23417 73116 23510 73182
rect 23417 73014 23510 73080
tri 23417 72998 23433 73014 ne
rect 23433 72998 23510 73014
rect 23250 72899 23398 72981
rect 23138 72866 23215 72882
tri 23215 72866 23231 72882 sw
rect 23138 72800 23231 72866
rect 23267 72741 23381 72899
tri 23417 72866 23433 72882 se
rect 23433 72866 23510 72882
rect 23417 72800 23510 72866
rect 23138 72665 23510 72741
rect 23138 72540 23231 72606
rect 23138 72524 23215 72540
tri 23215 72524 23231 72540 nw
rect 23267 72507 23381 72665
rect 23417 72540 23510 72606
tri 23417 72524 23433 72540 ne
rect 23433 72524 23510 72540
rect 23250 72425 23398 72507
rect 23138 72392 23215 72408
tri 23215 72392 23231 72408 sw
rect 23138 72326 23231 72392
rect 23138 72224 23231 72290
rect 23138 72208 23215 72224
tri 23215 72208 23231 72224 nw
rect 23267 72191 23381 72425
tri 23417 72392 23433 72408 se
rect 23433 72392 23510 72408
rect 23417 72326 23510 72392
rect 23417 72224 23510 72290
tri 23417 72208 23433 72224 ne
rect 23433 72208 23510 72224
rect 23250 72109 23398 72191
rect 23138 72076 23215 72092
tri 23215 72076 23231 72092 sw
rect 23138 72010 23231 72076
rect 23267 71951 23381 72109
tri 23417 72076 23433 72092 se
rect 23433 72076 23510 72092
rect 23417 72010 23510 72076
rect 23138 71875 23510 71951
rect 23138 71750 23231 71816
rect 23138 71734 23215 71750
tri 23215 71734 23231 71750 nw
rect 23267 71717 23381 71875
rect 23417 71750 23510 71816
tri 23417 71734 23433 71750 ne
rect 23433 71734 23510 71750
rect 23250 71635 23398 71717
rect 23138 71602 23215 71618
tri 23215 71602 23231 71618 sw
rect 23138 71536 23231 71602
rect 23138 71434 23231 71500
rect 23138 71418 23215 71434
tri 23215 71418 23231 71434 nw
rect 23267 71401 23381 71635
tri 23417 71602 23433 71618 se
rect 23433 71602 23510 71618
rect 23417 71536 23510 71602
rect 23417 71434 23510 71500
tri 23417 71418 23433 71434 ne
rect 23433 71418 23510 71434
rect 23250 71319 23398 71401
rect 23138 71286 23215 71302
tri 23215 71286 23231 71302 sw
rect 23138 71220 23231 71286
rect 23267 71161 23381 71319
tri 23417 71286 23433 71302 se
rect 23433 71286 23510 71302
rect 23417 71220 23510 71286
rect 23138 71085 23510 71161
rect 23138 70960 23231 71026
rect 23138 70944 23215 70960
tri 23215 70944 23231 70960 nw
rect 23267 70927 23381 71085
rect 23417 70960 23510 71026
tri 23417 70944 23433 70960 ne
rect 23433 70944 23510 70960
rect 23250 70845 23398 70927
rect 23138 70812 23215 70828
tri 23215 70812 23231 70828 sw
rect 23138 70746 23231 70812
rect 23138 70644 23231 70710
rect 23138 70628 23215 70644
tri 23215 70628 23231 70644 nw
rect 23267 70611 23381 70845
tri 23417 70812 23433 70828 se
rect 23433 70812 23510 70828
rect 23417 70746 23510 70812
rect 23417 70644 23510 70710
tri 23417 70628 23433 70644 ne
rect 23433 70628 23510 70644
rect 23250 70529 23398 70611
rect 23138 70496 23215 70512
tri 23215 70496 23231 70512 sw
rect 23138 70430 23231 70496
rect 23267 70371 23381 70529
tri 23417 70496 23433 70512 se
rect 23433 70496 23510 70512
rect 23417 70430 23510 70496
rect 23138 70295 23510 70371
rect 23138 70170 23231 70236
rect 23138 70154 23215 70170
tri 23215 70154 23231 70170 nw
rect 23267 70137 23381 70295
rect 23417 70170 23510 70236
tri 23417 70154 23433 70170 ne
rect 23433 70154 23510 70170
rect 23250 70055 23398 70137
rect 23138 70022 23215 70038
tri 23215 70022 23231 70038 sw
rect 23138 69956 23231 70022
rect 23138 69854 23231 69920
rect 23138 69838 23215 69854
tri 23215 69838 23231 69854 nw
rect 23267 69821 23381 70055
tri 23417 70022 23433 70038 se
rect 23433 70022 23510 70038
rect 23417 69956 23510 70022
rect 23417 69854 23510 69920
tri 23417 69838 23433 69854 ne
rect 23433 69838 23510 69854
rect 23250 69739 23398 69821
rect 23138 69706 23215 69722
tri 23215 69706 23231 69722 sw
rect 23138 69640 23231 69706
rect 23267 69581 23381 69739
tri 23417 69706 23433 69722 se
rect 23433 69706 23510 69722
rect 23417 69640 23510 69706
rect 23138 69505 23510 69581
rect 23138 69380 23231 69446
rect 23138 69364 23215 69380
tri 23215 69364 23231 69380 nw
rect 23267 69347 23381 69505
rect 23417 69380 23510 69446
tri 23417 69364 23433 69380 ne
rect 23433 69364 23510 69380
rect 23250 69265 23398 69347
rect 23138 69232 23215 69248
tri 23215 69232 23231 69248 sw
rect 23138 69166 23231 69232
rect 23138 69064 23231 69130
rect 23138 69048 23215 69064
tri 23215 69048 23231 69064 nw
rect 23267 69031 23381 69265
tri 23417 69232 23433 69248 se
rect 23433 69232 23510 69248
rect 23417 69166 23510 69232
rect 23417 69064 23510 69130
tri 23417 69048 23433 69064 ne
rect 23433 69048 23510 69064
rect 23250 68949 23398 69031
rect 23138 68916 23215 68932
tri 23215 68916 23231 68932 sw
rect 23138 68850 23231 68916
rect 23267 68791 23381 68949
tri 23417 68916 23433 68932 se
rect 23433 68916 23510 68932
rect 23417 68850 23510 68916
rect 23138 68715 23510 68791
rect 23138 68590 23231 68656
rect 23138 68574 23215 68590
tri 23215 68574 23231 68590 nw
rect 23267 68557 23381 68715
rect 23417 68590 23510 68656
tri 23417 68574 23433 68590 ne
rect 23433 68574 23510 68590
rect 23250 68475 23398 68557
rect 23138 68442 23215 68458
tri 23215 68442 23231 68458 sw
rect 23138 68376 23231 68442
rect 23138 68274 23231 68340
rect 23138 68258 23215 68274
tri 23215 68258 23231 68274 nw
rect 23267 68241 23381 68475
tri 23417 68442 23433 68458 se
rect 23433 68442 23510 68458
rect 23417 68376 23510 68442
rect 23417 68274 23510 68340
tri 23417 68258 23433 68274 ne
rect 23433 68258 23510 68274
rect 23250 68159 23398 68241
rect 23138 68126 23215 68142
tri 23215 68126 23231 68142 sw
rect 23138 68060 23231 68126
rect 23267 68001 23381 68159
tri 23417 68126 23433 68142 se
rect 23433 68126 23510 68142
rect 23417 68060 23510 68126
rect 23138 67925 23510 68001
rect 23138 67800 23231 67866
rect 23138 67784 23215 67800
tri 23215 67784 23231 67800 nw
rect 23267 67767 23381 67925
rect 23417 67800 23510 67866
tri 23417 67784 23433 67800 ne
rect 23433 67784 23510 67800
rect 23250 67685 23398 67767
rect 23138 67652 23215 67668
tri 23215 67652 23231 67668 sw
rect 23138 67586 23231 67652
rect 23138 67484 23231 67550
rect 23138 67468 23215 67484
tri 23215 67468 23231 67484 nw
rect 23267 67451 23381 67685
tri 23417 67652 23433 67668 se
rect 23433 67652 23510 67668
rect 23417 67586 23510 67652
rect 23417 67484 23510 67550
tri 23417 67468 23433 67484 ne
rect 23433 67468 23510 67484
rect 23250 67369 23398 67451
rect 23138 67336 23215 67352
tri 23215 67336 23231 67352 sw
rect 23138 67270 23231 67336
rect 23267 67211 23381 67369
tri 23417 67336 23433 67352 se
rect 23433 67336 23510 67352
rect 23417 67270 23510 67336
rect 23138 67135 23510 67211
rect 23138 67010 23231 67076
rect 23138 66994 23215 67010
tri 23215 66994 23231 67010 nw
rect 23267 66977 23381 67135
rect 23417 67010 23510 67076
tri 23417 66994 23433 67010 ne
rect 23433 66994 23510 67010
rect 23250 66895 23398 66977
rect 23138 66862 23215 66878
tri 23215 66862 23231 66878 sw
rect 23138 66796 23231 66862
rect 23138 66694 23231 66760
rect 23138 66678 23215 66694
tri 23215 66678 23231 66694 nw
rect 23267 66661 23381 66895
tri 23417 66862 23433 66878 se
rect 23433 66862 23510 66878
rect 23417 66796 23510 66862
rect 23417 66694 23510 66760
tri 23417 66678 23433 66694 ne
rect 23433 66678 23510 66694
rect 23250 66579 23398 66661
rect 23138 66546 23215 66562
tri 23215 66546 23231 66562 sw
rect 23138 66480 23231 66546
rect 23267 66421 23381 66579
tri 23417 66546 23433 66562 se
rect 23433 66546 23510 66562
rect 23417 66480 23510 66546
rect 23138 66345 23510 66421
rect 23138 66220 23231 66286
rect 23138 66204 23215 66220
tri 23215 66204 23231 66220 nw
rect 23267 66187 23381 66345
rect 23417 66220 23510 66286
tri 23417 66204 23433 66220 ne
rect 23433 66204 23510 66220
rect 23250 66105 23398 66187
rect 23138 66072 23215 66088
tri 23215 66072 23231 66088 sw
rect 23138 66006 23231 66072
rect 23138 65904 23231 65970
rect 23138 65888 23215 65904
tri 23215 65888 23231 65904 nw
rect 23267 65871 23381 66105
tri 23417 66072 23433 66088 se
rect 23433 66072 23510 66088
rect 23417 66006 23510 66072
rect 23417 65904 23510 65970
tri 23417 65888 23433 65904 ne
rect 23433 65888 23510 65904
rect 23250 65789 23398 65871
rect 23138 65756 23215 65772
tri 23215 65756 23231 65772 sw
rect 23138 65690 23231 65756
rect 23267 65631 23381 65789
tri 23417 65756 23433 65772 se
rect 23433 65756 23510 65772
rect 23417 65690 23510 65756
rect 23138 65555 23510 65631
rect 23138 65430 23231 65496
rect 23138 65414 23215 65430
tri 23215 65414 23231 65430 nw
rect 23267 65397 23381 65555
rect 23417 65430 23510 65496
tri 23417 65414 23433 65430 ne
rect 23433 65414 23510 65430
rect 23250 65315 23398 65397
rect 23138 65282 23215 65298
tri 23215 65282 23231 65298 sw
rect 23138 65216 23231 65282
rect 23138 65114 23231 65180
rect 23138 65098 23215 65114
tri 23215 65098 23231 65114 nw
rect 23267 65081 23381 65315
tri 23417 65282 23433 65298 se
rect 23433 65282 23510 65298
rect 23417 65216 23510 65282
rect 23417 65114 23510 65180
tri 23417 65098 23433 65114 ne
rect 23433 65098 23510 65114
rect 23250 64999 23398 65081
rect 23138 64966 23215 64982
tri 23215 64966 23231 64982 sw
rect 23138 64900 23231 64966
rect 23267 64841 23381 64999
tri 23417 64966 23433 64982 se
rect 23433 64966 23510 64982
rect 23417 64900 23510 64966
rect 23138 64765 23510 64841
rect 23138 64640 23231 64706
rect 23138 64624 23215 64640
tri 23215 64624 23231 64640 nw
rect 23267 64607 23381 64765
rect 23417 64640 23510 64706
tri 23417 64624 23433 64640 ne
rect 23433 64624 23510 64640
rect 23250 64525 23398 64607
rect 23138 64492 23215 64508
tri 23215 64492 23231 64508 sw
rect 23138 64426 23231 64492
rect 23138 64324 23231 64390
rect 23138 64308 23215 64324
tri 23215 64308 23231 64324 nw
rect 23267 64291 23381 64525
tri 23417 64492 23433 64508 se
rect 23433 64492 23510 64508
rect 23417 64426 23510 64492
rect 23417 64324 23510 64390
tri 23417 64308 23433 64324 ne
rect 23433 64308 23510 64324
rect 23250 64209 23398 64291
rect 23138 64176 23215 64192
tri 23215 64176 23231 64192 sw
rect 23138 64110 23231 64176
rect 23267 64051 23381 64209
tri 23417 64176 23433 64192 se
rect 23433 64176 23510 64192
rect 23417 64110 23510 64176
rect 23138 63975 23510 64051
rect 23138 63850 23231 63916
rect 23138 63834 23215 63850
tri 23215 63834 23231 63850 nw
rect 23267 63817 23381 63975
rect 23417 63850 23510 63916
tri 23417 63834 23433 63850 ne
rect 23433 63834 23510 63850
rect 23250 63735 23398 63817
rect 23138 63702 23215 63718
tri 23215 63702 23231 63718 sw
rect 23138 63636 23231 63702
rect 23138 63534 23231 63600
rect 23138 63518 23215 63534
tri 23215 63518 23231 63534 nw
rect 23267 63501 23381 63735
tri 23417 63702 23433 63718 se
rect 23433 63702 23510 63718
rect 23417 63636 23510 63702
rect 23417 63534 23510 63600
tri 23417 63518 23433 63534 ne
rect 23433 63518 23510 63534
rect 23250 63419 23398 63501
rect 23138 63386 23215 63402
tri 23215 63386 23231 63402 sw
rect 23138 63320 23231 63386
rect 23267 63261 23381 63419
tri 23417 63386 23433 63402 se
rect 23433 63386 23510 63402
rect 23417 63320 23510 63386
rect 23138 63185 23510 63261
rect 23138 63060 23231 63126
rect 23138 63044 23215 63060
tri 23215 63044 23231 63060 nw
rect 23267 63027 23381 63185
rect 23417 63060 23510 63126
tri 23417 63044 23433 63060 ne
rect 23433 63044 23510 63060
rect 23250 62945 23398 63027
rect 23138 62912 23215 62928
tri 23215 62912 23231 62928 sw
rect 23138 62846 23231 62912
rect 23138 62744 23231 62810
rect 23138 62728 23215 62744
tri 23215 62728 23231 62744 nw
rect 23267 62711 23381 62945
tri 23417 62912 23433 62928 se
rect 23433 62912 23510 62928
rect 23417 62846 23510 62912
rect 23417 62744 23510 62810
tri 23417 62728 23433 62744 ne
rect 23433 62728 23510 62744
rect 23250 62629 23398 62711
rect 23138 62596 23215 62612
tri 23215 62596 23231 62612 sw
rect 23138 62530 23231 62596
rect 23267 62471 23381 62629
tri 23417 62596 23433 62612 se
rect 23433 62596 23510 62612
rect 23417 62530 23510 62596
rect 23138 62395 23510 62471
rect 23138 62270 23231 62336
rect 23138 62254 23215 62270
tri 23215 62254 23231 62270 nw
rect 23267 62237 23381 62395
rect 23417 62270 23510 62336
tri 23417 62254 23433 62270 ne
rect 23433 62254 23510 62270
rect 23250 62155 23398 62237
rect 23138 62122 23215 62138
tri 23215 62122 23231 62138 sw
rect 23138 62056 23231 62122
rect 23138 61954 23231 62020
rect 23138 61938 23215 61954
tri 23215 61938 23231 61954 nw
rect 23267 61921 23381 62155
tri 23417 62122 23433 62138 se
rect 23433 62122 23510 62138
rect 23417 62056 23510 62122
rect 23417 61954 23510 62020
tri 23417 61938 23433 61954 ne
rect 23433 61938 23510 61954
rect 23250 61839 23398 61921
rect 23138 61806 23215 61822
tri 23215 61806 23231 61822 sw
rect 23138 61740 23231 61806
rect 23267 61681 23381 61839
tri 23417 61806 23433 61822 se
rect 23433 61806 23510 61822
rect 23417 61740 23510 61806
rect 23138 61605 23510 61681
rect 23138 61480 23231 61546
rect 23138 61464 23215 61480
tri 23215 61464 23231 61480 nw
rect 23267 61447 23381 61605
rect 23417 61480 23510 61546
tri 23417 61464 23433 61480 ne
rect 23433 61464 23510 61480
rect 23250 61365 23398 61447
rect 23138 61332 23215 61348
tri 23215 61332 23231 61348 sw
rect 23138 61266 23231 61332
rect 23138 61164 23231 61230
rect 23138 61148 23215 61164
tri 23215 61148 23231 61164 nw
rect 23267 61131 23381 61365
tri 23417 61332 23433 61348 se
rect 23433 61332 23510 61348
rect 23417 61266 23510 61332
rect 23417 61164 23510 61230
tri 23417 61148 23433 61164 ne
rect 23433 61148 23510 61164
rect 23250 61049 23398 61131
rect 23138 61016 23215 61032
tri 23215 61016 23231 61032 sw
rect 23138 60950 23231 61016
rect 23267 60891 23381 61049
tri 23417 61016 23433 61032 se
rect 23433 61016 23510 61032
rect 23417 60950 23510 61016
rect 23138 60815 23510 60891
rect 23138 60690 23231 60756
rect 23138 60674 23215 60690
tri 23215 60674 23231 60690 nw
rect 23267 60657 23381 60815
rect 23417 60690 23510 60756
tri 23417 60674 23433 60690 ne
rect 23433 60674 23510 60690
rect 23250 60575 23398 60657
rect 23138 60542 23215 60558
tri 23215 60542 23231 60558 sw
rect 23138 60476 23231 60542
rect 23138 60374 23231 60440
rect 23138 60358 23215 60374
tri 23215 60358 23231 60374 nw
rect 23267 60341 23381 60575
tri 23417 60542 23433 60558 se
rect 23433 60542 23510 60558
rect 23417 60476 23510 60542
rect 23417 60374 23510 60440
tri 23417 60358 23433 60374 ne
rect 23433 60358 23510 60374
rect 23250 60259 23398 60341
rect 23138 60226 23215 60242
tri 23215 60226 23231 60242 sw
rect 23138 60160 23231 60226
rect 23267 60101 23381 60259
tri 23417 60226 23433 60242 se
rect 23433 60226 23510 60242
rect 23417 60160 23510 60226
rect 23138 60025 23510 60101
rect 23138 59900 23231 59966
rect 23138 59884 23215 59900
tri 23215 59884 23231 59900 nw
rect 23267 59867 23381 60025
rect 23417 59900 23510 59966
tri 23417 59884 23433 59900 ne
rect 23433 59884 23510 59900
rect 23250 59785 23398 59867
rect 23138 59752 23215 59768
tri 23215 59752 23231 59768 sw
rect 23138 59686 23231 59752
rect 23138 59584 23231 59650
rect 23138 59568 23215 59584
tri 23215 59568 23231 59584 nw
rect 23267 59551 23381 59785
tri 23417 59752 23433 59768 se
rect 23433 59752 23510 59768
rect 23417 59686 23510 59752
rect 23417 59584 23510 59650
tri 23417 59568 23433 59584 ne
rect 23433 59568 23510 59584
rect 23250 59469 23398 59551
rect 23138 59436 23215 59452
tri 23215 59436 23231 59452 sw
rect 23138 59370 23231 59436
rect 23267 59311 23381 59469
tri 23417 59436 23433 59452 se
rect 23433 59436 23510 59452
rect 23417 59370 23510 59436
rect 23138 59235 23510 59311
rect 23138 59110 23231 59176
rect 23138 59094 23215 59110
tri 23215 59094 23231 59110 nw
rect 23267 59077 23381 59235
rect 23417 59110 23510 59176
tri 23417 59094 23433 59110 ne
rect 23433 59094 23510 59110
rect 23250 58995 23398 59077
rect 23138 58962 23215 58978
tri 23215 58962 23231 58978 sw
rect 23138 58896 23231 58962
rect 23138 58794 23231 58860
rect 23138 58778 23215 58794
tri 23215 58778 23231 58794 nw
rect 23267 58761 23381 58995
tri 23417 58962 23433 58978 se
rect 23433 58962 23510 58978
rect 23417 58896 23510 58962
rect 23417 58794 23510 58860
tri 23417 58778 23433 58794 ne
rect 23433 58778 23510 58794
rect 23250 58679 23398 58761
rect 23138 58646 23215 58662
tri 23215 58646 23231 58662 sw
rect 23138 58580 23231 58646
rect 23267 58521 23381 58679
tri 23417 58646 23433 58662 se
rect 23433 58646 23510 58662
rect 23417 58580 23510 58646
rect 23138 58445 23510 58521
rect 23138 58320 23231 58386
rect 23138 58304 23215 58320
tri 23215 58304 23231 58320 nw
rect 23267 58287 23381 58445
rect 23417 58320 23510 58386
tri 23417 58304 23433 58320 ne
rect 23433 58304 23510 58320
rect 23250 58205 23398 58287
rect 23138 58172 23215 58188
tri 23215 58172 23231 58188 sw
rect 23138 58106 23231 58172
rect 23138 58004 23231 58070
rect 23138 57988 23215 58004
tri 23215 57988 23231 58004 nw
rect 23267 57971 23381 58205
tri 23417 58172 23433 58188 se
rect 23433 58172 23510 58188
rect 23417 58106 23510 58172
rect 23417 58004 23510 58070
tri 23417 57988 23433 58004 ne
rect 23433 57988 23510 58004
rect 23250 57889 23398 57971
rect 23138 57856 23215 57872
tri 23215 57856 23231 57872 sw
rect 23138 57790 23231 57856
rect 23267 57731 23381 57889
tri 23417 57856 23433 57872 se
rect 23433 57856 23510 57872
rect 23417 57790 23510 57856
rect 23138 57655 23510 57731
rect 23138 57530 23231 57596
rect 23138 57514 23215 57530
tri 23215 57514 23231 57530 nw
rect 23267 57497 23381 57655
rect 23417 57530 23510 57596
tri 23417 57514 23433 57530 ne
rect 23433 57514 23510 57530
rect 23250 57415 23398 57497
rect 23138 57382 23215 57398
tri 23215 57382 23231 57398 sw
rect 23138 57316 23231 57382
rect 23138 57214 23231 57280
rect 23138 57198 23215 57214
tri 23215 57198 23231 57214 nw
rect 23267 57181 23381 57415
tri 23417 57382 23433 57398 se
rect 23433 57382 23510 57398
rect 23417 57316 23510 57382
rect 23417 57214 23510 57280
tri 23417 57198 23433 57214 ne
rect 23433 57198 23510 57214
rect 23250 57099 23398 57181
rect 23138 57066 23215 57082
tri 23215 57066 23231 57082 sw
rect 23138 57000 23231 57066
rect 23267 56941 23381 57099
tri 23417 57066 23433 57082 se
rect 23433 57066 23510 57082
rect 23417 57000 23510 57066
rect 23138 56865 23510 56941
rect 23138 56740 23231 56806
rect 23138 56724 23215 56740
tri 23215 56724 23231 56740 nw
rect 23267 56707 23381 56865
rect 23417 56740 23510 56806
tri 23417 56724 23433 56740 ne
rect 23433 56724 23510 56740
rect 23250 56625 23398 56707
rect 23138 56592 23215 56608
tri 23215 56592 23231 56608 sw
rect 23138 56526 23231 56592
rect 23138 56424 23231 56490
rect 23138 56408 23215 56424
tri 23215 56408 23231 56424 nw
rect 23267 56391 23381 56625
tri 23417 56592 23433 56608 se
rect 23433 56592 23510 56608
rect 23417 56526 23510 56592
rect 23417 56424 23510 56490
tri 23417 56408 23433 56424 ne
rect 23433 56408 23510 56424
rect 23250 56309 23398 56391
rect 23138 56276 23215 56292
tri 23215 56276 23231 56292 sw
rect 23138 56210 23231 56276
rect 23267 56151 23381 56309
tri 23417 56276 23433 56292 se
rect 23433 56276 23510 56292
rect 23417 56210 23510 56276
rect 23138 56075 23510 56151
rect 23138 55950 23231 56016
rect 23138 55934 23215 55950
tri 23215 55934 23231 55950 nw
rect 23267 55917 23381 56075
rect 23417 55950 23510 56016
tri 23417 55934 23433 55950 ne
rect 23433 55934 23510 55950
rect 23250 55835 23398 55917
rect 23138 55802 23215 55818
tri 23215 55802 23231 55818 sw
rect 23138 55736 23231 55802
rect 23138 55634 23231 55700
rect 23138 55618 23215 55634
tri 23215 55618 23231 55634 nw
rect 23267 55601 23381 55835
tri 23417 55802 23433 55818 se
rect 23433 55802 23510 55818
rect 23417 55736 23510 55802
rect 23417 55634 23510 55700
tri 23417 55618 23433 55634 ne
rect 23433 55618 23510 55634
rect 23250 55519 23398 55601
rect 23138 55486 23215 55502
tri 23215 55486 23231 55502 sw
rect 23138 55420 23231 55486
rect 23267 55361 23381 55519
tri 23417 55486 23433 55502 se
rect 23433 55486 23510 55502
rect 23417 55420 23510 55486
rect 23138 55285 23510 55361
rect 23138 55160 23231 55226
rect 23138 55144 23215 55160
tri 23215 55144 23231 55160 nw
rect 23267 55127 23381 55285
rect 23417 55160 23510 55226
tri 23417 55144 23433 55160 ne
rect 23433 55144 23510 55160
rect 23250 55045 23398 55127
rect 23138 55012 23215 55028
tri 23215 55012 23231 55028 sw
rect 23138 54946 23231 55012
rect 23138 54844 23231 54910
rect 23138 54828 23215 54844
tri 23215 54828 23231 54844 nw
rect 23267 54811 23381 55045
tri 23417 55012 23433 55028 se
rect 23433 55012 23510 55028
rect 23417 54946 23510 55012
rect 23417 54844 23510 54910
tri 23417 54828 23433 54844 ne
rect 23433 54828 23510 54844
rect 23250 54729 23398 54811
rect 23138 54696 23215 54712
tri 23215 54696 23231 54712 sw
rect 23138 54630 23231 54696
rect 23267 54571 23381 54729
tri 23417 54696 23433 54712 se
rect 23433 54696 23510 54712
rect 23417 54630 23510 54696
rect 23138 54495 23510 54571
rect 23138 54370 23231 54436
rect 23138 54354 23215 54370
tri 23215 54354 23231 54370 nw
rect 23267 54337 23381 54495
rect 23417 54370 23510 54436
tri 23417 54354 23433 54370 ne
rect 23433 54354 23510 54370
rect 23250 54255 23398 54337
rect 23138 54222 23215 54238
tri 23215 54222 23231 54238 sw
rect 23138 54156 23231 54222
rect 23138 54054 23231 54120
rect 23138 54038 23215 54054
tri 23215 54038 23231 54054 nw
rect 23267 54021 23381 54255
tri 23417 54222 23433 54238 se
rect 23433 54222 23510 54238
rect 23417 54156 23510 54222
rect 23417 54054 23510 54120
tri 23417 54038 23433 54054 ne
rect 23433 54038 23510 54054
rect 23250 53939 23398 54021
rect 23138 53906 23215 53922
tri 23215 53906 23231 53922 sw
rect 23138 53840 23231 53906
rect 23267 53781 23381 53939
tri 23417 53906 23433 53922 se
rect 23433 53906 23510 53922
rect 23417 53840 23510 53906
rect 23138 53705 23510 53781
rect 23138 53580 23231 53646
rect 23138 53564 23215 53580
tri 23215 53564 23231 53580 nw
rect 23267 53547 23381 53705
rect 23417 53580 23510 53646
tri 23417 53564 23433 53580 ne
rect 23433 53564 23510 53580
rect 23250 53465 23398 53547
rect 23138 53432 23215 53448
tri 23215 53432 23231 53448 sw
rect 23138 53366 23231 53432
rect 23138 53264 23231 53330
rect 23138 53248 23215 53264
tri 23215 53248 23231 53264 nw
rect 23267 53231 23381 53465
tri 23417 53432 23433 53448 se
rect 23433 53432 23510 53448
rect 23417 53366 23510 53432
rect 23417 53264 23510 53330
tri 23417 53248 23433 53264 ne
rect 23433 53248 23510 53264
rect 23250 53149 23398 53231
rect 23138 53116 23215 53132
tri 23215 53116 23231 53132 sw
rect 23138 53050 23231 53116
rect 23267 52991 23381 53149
tri 23417 53116 23433 53132 se
rect 23433 53116 23510 53132
rect 23417 53050 23510 53116
rect 23138 52915 23510 52991
rect 23138 52790 23231 52856
rect 23138 52774 23215 52790
tri 23215 52774 23231 52790 nw
rect 23267 52757 23381 52915
rect 23417 52790 23510 52856
tri 23417 52774 23433 52790 ne
rect 23433 52774 23510 52790
rect 23250 52675 23398 52757
rect 23138 52642 23215 52658
tri 23215 52642 23231 52658 sw
rect 23138 52576 23231 52642
rect 23138 52474 23231 52540
rect 23138 52458 23215 52474
tri 23215 52458 23231 52474 nw
rect 23267 52441 23381 52675
tri 23417 52642 23433 52658 se
rect 23433 52642 23510 52658
rect 23417 52576 23510 52642
rect 23417 52474 23510 52540
tri 23417 52458 23433 52474 ne
rect 23433 52458 23510 52474
rect 23250 52359 23398 52441
rect 23138 52326 23215 52342
tri 23215 52326 23231 52342 sw
rect 23138 52260 23231 52326
rect 23267 52201 23381 52359
tri 23417 52326 23433 52342 se
rect 23433 52326 23510 52342
rect 23417 52260 23510 52326
rect 23138 52125 23510 52201
rect 23138 52000 23231 52066
rect 23138 51984 23215 52000
tri 23215 51984 23231 52000 nw
rect 23267 51967 23381 52125
rect 23417 52000 23510 52066
tri 23417 51984 23433 52000 ne
rect 23433 51984 23510 52000
rect 23250 51885 23398 51967
rect 23138 51852 23215 51868
tri 23215 51852 23231 51868 sw
rect 23138 51786 23231 51852
rect 23138 51684 23231 51750
rect 23138 51668 23215 51684
tri 23215 51668 23231 51684 nw
rect 23267 51651 23381 51885
tri 23417 51852 23433 51868 se
rect 23433 51852 23510 51868
rect 23417 51786 23510 51852
rect 23417 51684 23510 51750
tri 23417 51668 23433 51684 ne
rect 23433 51668 23510 51684
rect 23250 51569 23398 51651
rect 23138 51536 23215 51552
tri 23215 51536 23231 51552 sw
rect 23138 51470 23231 51536
rect 23267 51411 23381 51569
tri 23417 51536 23433 51552 se
rect 23433 51536 23510 51552
rect 23417 51470 23510 51536
rect 23138 51335 23510 51411
rect 23138 51210 23231 51276
rect 23138 51194 23215 51210
tri 23215 51194 23231 51210 nw
rect 23267 51177 23381 51335
rect 23417 51210 23510 51276
tri 23417 51194 23433 51210 ne
rect 23433 51194 23510 51210
rect 23250 51095 23398 51177
rect 23138 51062 23215 51078
tri 23215 51062 23231 51078 sw
rect 23138 50996 23231 51062
rect 23138 50894 23231 50960
rect 23138 50878 23215 50894
tri 23215 50878 23231 50894 nw
rect 23267 50861 23381 51095
tri 23417 51062 23433 51078 se
rect 23433 51062 23510 51078
rect 23417 50996 23510 51062
rect 23417 50894 23510 50960
tri 23417 50878 23433 50894 ne
rect 23433 50878 23510 50894
rect 23250 50779 23398 50861
rect 23138 50746 23215 50762
tri 23215 50746 23231 50762 sw
rect 23138 50680 23231 50746
rect 23267 50621 23381 50779
tri 23417 50746 23433 50762 se
rect 23433 50746 23510 50762
rect 23417 50680 23510 50746
rect 23138 50545 23510 50621
rect 23138 50420 23231 50486
rect 23138 50404 23215 50420
tri 23215 50404 23231 50420 nw
rect 23267 50387 23381 50545
rect 23417 50420 23510 50486
tri 23417 50404 23433 50420 ne
rect 23433 50404 23510 50420
rect 23250 50305 23398 50387
rect 23138 50272 23215 50288
tri 23215 50272 23231 50288 sw
rect 23138 50206 23231 50272
rect 23138 50104 23231 50170
rect 23138 50088 23215 50104
tri 23215 50088 23231 50104 nw
rect 23267 50071 23381 50305
tri 23417 50272 23433 50288 se
rect 23433 50272 23510 50288
rect 23417 50206 23510 50272
rect 23417 50104 23510 50170
tri 23417 50088 23433 50104 ne
rect 23433 50088 23510 50104
rect 23250 49989 23398 50071
rect 23138 49956 23215 49972
tri 23215 49956 23231 49972 sw
rect 23138 49890 23231 49956
rect 23267 49831 23381 49989
tri 23417 49956 23433 49972 se
rect 23433 49956 23510 49972
rect 23417 49890 23510 49956
rect 23138 49755 23510 49831
rect 23138 49630 23231 49696
rect 23138 49614 23215 49630
tri 23215 49614 23231 49630 nw
rect 23267 49597 23381 49755
rect 23417 49630 23510 49696
tri 23417 49614 23433 49630 ne
rect 23433 49614 23510 49630
rect 23250 49515 23398 49597
rect 23138 49482 23215 49498
tri 23215 49482 23231 49498 sw
rect 23138 49416 23231 49482
rect 23138 49314 23231 49380
rect 23138 49298 23215 49314
tri 23215 49298 23231 49314 nw
rect 23267 49281 23381 49515
tri 23417 49482 23433 49498 se
rect 23433 49482 23510 49498
rect 23417 49416 23510 49482
rect 23417 49314 23510 49380
tri 23417 49298 23433 49314 ne
rect 23433 49298 23510 49314
rect 23250 49199 23398 49281
rect 23138 49166 23215 49182
tri 23215 49166 23231 49182 sw
rect 23138 49100 23231 49166
rect 23267 49041 23381 49199
tri 23417 49166 23433 49182 se
rect 23433 49166 23510 49182
rect 23417 49100 23510 49166
rect 23138 48965 23510 49041
rect 23138 48840 23231 48906
rect 23138 48824 23215 48840
tri 23215 48824 23231 48840 nw
rect 23267 48807 23381 48965
rect 23417 48840 23510 48906
tri 23417 48824 23433 48840 ne
rect 23433 48824 23510 48840
rect 23250 48725 23398 48807
rect 23138 48692 23215 48708
tri 23215 48692 23231 48708 sw
rect 23138 48626 23231 48692
rect 23138 48524 23231 48590
rect 23138 48508 23215 48524
tri 23215 48508 23231 48524 nw
rect 23267 48491 23381 48725
tri 23417 48692 23433 48708 se
rect 23433 48692 23510 48708
rect 23417 48626 23510 48692
rect 23417 48524 23510 48590
tri 23417 48508 23433 48524 ne
rect 23433 48508 23510 48524
rect 23250 48409 23398 48491
rect 23138 48376 23215 48392
tri 23215 48376 23231 48392 sw
rect 23138 48310 23231 48376
rect 23267 48251 23381 48409
tri 23417 48376 23433 48392 se
rect 23433 48376 23510 48392
rect 23417 48310 23510 48376
rect 23138 48175 23510 48251
rect 23138 48050 23231 48116
rect 23138 48034 23215 48050
tri 23215 48034 23231 48050 nw
rect 23267 48017 23381 48175
rect 23417 48050 23510 48116
tri 23417 48034 23433 48050 ne
rect 23433 48034 23510 48050
rect 23250 47935 23398 48017
rect 23138 47902 23215 47918
tri 23215 47902 23231 47918 sw
rect 23138 47836 23231 47902
rect 23138 47734 23231 47800
rect 23138 47718 23215 47734
tri 23215 47718 23231 47734 nw
rect 23267 47701 23381 47935
tri 23417 47902 23433 47918 se
rect 23433 47902 23510 47918
rect 23417 47836 23510 47902
rect 23417 47734 23510 47800
tri 23417 47718 23433 47734 ne
rect 23433 47718 23510 47734
rect 23250 47619 23398 47701
rect 23138 47586 23215 47602
tri 23215 47586 23231 47602 sw
rect 23138 47520 23231 47586
rect 23267 47461 23381 47619
tri 23417 47586 23433 47602 se
rect 23433 47586 23510 47602
rect 23417 47520 23510 47586
rect 23138 47385 23510 47461
rect 23138 47260 23231 47326
rect 23138 47244 23215 47260
tri 23215 47244 23231 47260 nw
rect 23267 47227 23381 47385
rect 23417 47260 23510 47326
tri 23417 47244 23433 47260 ne
rect 23433 47244 23510 47260
rect 23250 47145 23398 47227
rect 23138 47112 23215 47128
tri 23215 47112 23231 47128 sw
rect 23138 47046 23231 47112
rect 23138 46944 23231 47010
rect 23138 46928 23215 46944
tri 23215 46928 23231 46944 nw
rect 23267 46911 23381 47145
tri 23417 47112 23433 47128 se
rect 23433 47112 23510 47128
rect 23417 47046 23510 47112
rect 23417 46944 23510 47010
tri 23417 46928 23433 46944 ne
rect 23433 46928 23510 46944
rect 23250 46829 23398 46911
rect 23138 46796 23215 46812
tri 23215 46796 23231 46812 sw
rect 23138 46730 23231 46796
rect 23267 46671 23381 46829
tri 23417 46796 23433 46812 se
rect 23433 46796 23510 46812
rect 23417 46730 23510 46796
rect 23138 46595 23510 46671
rect 23138 46470 23231 46536
rect 23138 46454 23215 46470
tri 23215 46454 23231 46470 nw
rect 23267 46437 23381 46595
rect 23417 46470 23510 46536
tri 23417 46454 23433 46470 ne
rect 23433 46454 23510 46470
rect 23250 46355 23398 46437
rect 23138 46322 23215 46338
tri 23215 46322 23231 46338 sw
rect 23138 46256 23231 46322
rect 23138 46154 23231 46220
rect 23138 46138 23215 46154
tri 23215 46138 23231 46154 nw
rect 23267 46121 23381 46355
tri 23417 46322 23433 46338 se
rect 23433 46322 23510 46338
rect 23417 46256 23510 46322
rect 23417 46154 23510 46220
tri 23417 46138 23433 46154 ne
rect 23433 46138 23510 46154
rect 23250 46039 23398 46121
rect 23138 46006 23215 46022
tri 23215 46006 23231 46022 sw
rect 23138 45940 23231 46006
rect 23267 45881 23381 46039
tri 23417 46006 23433 46022 se
rect 23433 46006 23510 46022
rect 23417 45940 23510 46006
rect 23138 45805 23510 45881
rect 23138 45680 23231 45746
rect 23138 45664 23215 45680
tri 23215 45664 23231 45680 nw
rect 23267 45647 23381 45805
rect 23417 45680 23510 45746
tri 23417 45664 23433 45680 ne
rect 23433 45664 23510 45680
rect 23250 45565 23398 45647
rect 23138 45532 23215 45548
tri 23215 45532 23231 45548 sw
rect 23138 45466 23231 45532
rect 23138 45364 23231 45430
rect 23138 45348 23215 45364
tri 23215 45348 23231 45364 nw
rect 23267 45331 23381 45565
tri 23417 45532 23433 45548 se
rect 23433 45532 23510 45548
rect 23417 45466 23510 45532
rect 23417 45364 23510 45430
tri 23417 45348 23433 45364 ne
rect 23433 45348 23510 45364
rect 23250 45249 23398 45331
rect 23138 45216 23215 45232
tri 23215 45216 23231 45232 sw
rect 23138 45150 23231 45216
rect 23267 45091 23381 45249
tri 23417 45216 23433 45232 se
rect 23433 45216 23510 45232
rect 23417 45150 23510 45216
rect 23138 45015 23510 45091
rect 23138 44890 23231 44956
rect 23138 44874 23215 44890
tri 23215 44874 23231 44890 nw
rect 23267 44857 23381 45015
rect 23417 44890 23510 44956
tri 23417 44874 23433 44890 ne
rect 23433 44874 23510 44890
rect 23250 44775 23398 44857
rect 23138 44742 23215 44758
tri 23215 44742 23231 44758 sw
rect 23138 44676 23231 44742
rect 23138 44574 23231 44640
rect 23138 44558 23215 44574
tri 23215 44558 23231 44574 nw
rect 23267 44541 23381 44775
tri 23417 44742 23433 44758 se
rect 23433 44742 23510 44758
rect 23417 44676 23510 44742
rect 23417 44574 23510 44640
tri 23417 44558 23433 44574 ne
rect 23433 44558 23510 44574
rect 23250 44459 23398 44541
rect 23138 44426 23215 44442
tri 23215 44426 23231 44442 sw
rect 23138 44360 23231 44426
rect 23267 44301 23381 44459
tri 23417 44426 23433 44442 se
rect 23433 44426 23510 44442
rect 23417 44360 23510 44426
rect 23138 44225 23510 44301
rect 23138 44100 23231 44166
rect 23138 44084 23215 44100
tri 23215 44084 23231 44100 nw
rect 23267 44067 23381 44225
rect 23417 44100 23510 44166
tri 23417 44084 23433 44100 ne
rect 23433 44084 23510 44100
rect 23250 43985 23398 44067
rect 23138 43952 23215 43968
tri 23215 43952 23231 43968 sw
rect 23138 43886 23231 43952
rect 23138 43784 23231 43850
rect 23138 43768 23215 43784
tri 23215 43768 23231 43784 nw
rect 23267 43751 23381 43985
tri 23417 43952 23433 43968 se
rect 23433 43952 23510 43968
rect 23417 43886 23510 43952
rect 23417 43784 23510 43850
tri 23417 43768 23433 43784 ne
rect 23433 43768 23510 43784
rect 23250 43669 23398 43751
rect 23138 43636 23215 43652
tri 23215 43636 23231 43652 sw
rect 23138 43570 23231 43636
rect 23267 43511 23381 43669
tri 23417 43636 23433 43652 se
rect 23433 43636 23510 43652
rect 23417 43570 23510 43636
rect 23138 43435 23510 43511
rect 23138 43310 23231 43376
rect 23138 43294 23215 43310
tri 23215 43294 23231 43310 nw
rect 23267 43277 23381 43435
rect 23417 43310 23510 43376
tri 23417 43294 23433 43310 ne
rect 23433 43294 23510 43310
rect 23250 43195 23398 43277
rect 23138 43162 23215 43178
tri 23215 43162 23231 43178 sw
rect 23138 43096 23231 43162
rect 23138 42994 23231 43060
rect 23138 42978 23215 42994
tri 23215 42978 23231 42994 nw
rect 23267 42961 23381 43195
tri 23417 43162 23433 43178 se
rect 23433 43162 23510 43178
rect 23417 43096 23510 43162
rect 23417 42994 23510 43060
tri 23417 42978 23433 42994 ne
rect 23433 42978 23510 42994
rect 23250 42879 23398 42961
rect 23138 42846 23215 42862
tri 23215 42846 23231 42862 sw
rect 23138 42780 23231 42846
rect 23267 42721 23381 42879
tri 23417 42846 23433 42862 se
rect 23433 42846 23510 42862
rect 23417 42780 23510 42846
rect 23138 42645 23510 42721
rect 23138 42520 23231 42586
rect 23138 42504 23215 42520
tri 23215 42504 23231 42520 nw
rect 23267 42487 23381 42645
rect 23417 42520 23510 42586
tri 23417 42504 23433 42520 ne
rect 23433 42504 23510 42520
rect 23250 42405 23398 42487
rect 23138 42372 23215 42388
tri 23215 42372 23231 42388 sw
rect 23138 42306 23231 42372
rect 23138 42204 23231 42270
rect 23138 42188 23215 42204
tri 23215 42188 23231 42204 nw
rect 23267 42171 23381 42405
tri 23417 42372 23433 42388 se
rect 23433 42372 23510 42388
rect 23417 42306 23510 42372
rect 23417 42204 23510 42270
tri 23417 42188 23433 42204 ne
rect 23433 42188 23510 42204
rect 23250 42089 23398 42171
rect 23138 42056 23215 42072
tri 23215 42056 23231 42072 sw
rect 23138 41990 23231 42056
rect 23267 41931 23381 42089
tri 23417 42056 23433 42072 se
rect 23433 42056 23510 42072
rect 23417 41990 23510 42056
rect 23138 41855 23510 41931
rect 23138 41730 23231 41796
rect 23138 41714 23215 41730
tri 23215 41714 23231 41730 nw
rect 23267 41697 23381 41855
rect 23417 41730 23510 41796
tri 23417 41714 23433 41730 ne
rect 23433 41714 23510 41730
rect 23250 41615 23398 41697
rect 23138 41582 23215 41598
tri 23215 41582 23231 41598 sw
rect 23138 41516 23231 41582
rect 23138 41414 23231 41480
rect 23138 41398 23215 41414
tri 23215 41398 23231 41414 nw
rect 23267 41381 23381 41615
tri 23417 41582 23433 41598 se
rect 23433 41582 23510 41598
rect 23417 41516 23510 41582
rect 23417 41414 23510 41480
tri 23417 41398 23433 41414 ne
rect 23433 41398 23510 41414
rect 23250 41299 23398 41381
rect 23138 41266 23215 41282
tri 23215 41266 23231 41282 sw
rect 23138 41200 23231 41266
rect 23267 41141 23381 41299
tri 23417 41266 23433 41282 se
rect 23433 41266 23510 41282
rect 23417 41200 23510 41266
rect 23138 41065 23510 41141
rect 23138 40940 23231 41006
rect 23138 40924 23215 40940
tri 23215 40924 23231 40940 nw
rect 23267 40907 23381 41065
rect 23417 40940 23510 41006
tri 23417 40924 23433 40940 ne
rect 23433 40924 23510 40940
rect 23250 40825 23398 40907
rect 23138 40792 23215 40808
tri 23215 40792 23231 40808 sw
rect 23138 40726 23231 40792
rect 23138 40624 23231 40690
rect 23138 40608 23215 40624
tri 23215 40608 23231 40624 nw
rect 23267 40591 23381 40825
tri 23417 40792 23433 40808 se
rect 23433 40792 23510 40808
rect 23417 40726 23510 40792
rect 23417 40624 23510 40690
tri 23417 40608 23433 40624 ne
rect 23433 40608 23510 40624
rect 23250 40509 23398 40591
rect 23138 40476 23215 40492
tri 23215 40476 23231 40492 sw
rect 23138 40410 23231 40476
rect 23267 40351 23381 40509
tri 23417 40476 23433 40492 se
rect 23433 40476 23510 40492
rect 23417 40410 23510 40476
rect 23138 40275 23510 40351
rect 23138 40150 23231 40216
rect 23138 40134 23215 40150
tri 23215 40134 23231 40150 nw
rect 23267 40117 23381 40275
rect 23417 40150 23510 40216
tri 23417 40134 23433 40150 ne
rect 23433 40134 23510 40150
rect 23250 40035 23398 40117
rect 23138 40002 23215 40018
tri 23215 40002 23231 40018 sw
rect 23138 39936 23231 40002
rect 23138 39834 23231 39900
rect 23138 39818 23215 39834
tri 23215 39818 23231 39834 nw
rect 23267 39801 23381 40035
tri 23417 40002 23433 40018 se
rect 23433 40002 23510 40018
rect 23417 39936 23510 40002
rect 23417 39834 23510 39900
tri 23417 39818 23433 39834 ne
rect 23433 39818 23510 39834
rect 23250 39719 23398 39801
rect 23138 39686 23215 39702
tri 23215 39686 23231 39702 sw
rect 23138 39620 23231 39686
rect 23267 39561 23381 39719
tri 23417 39686 23433 39702 se
rect 23433 39686 23510 39702
rect 23417 39620 23510 39686
rect 23138 39485 23510 39561
rect 23138 39360 23231 39426
rect 23138 39344 23215 39360
tri 23215 39344 23231 39360 nw
rect 23267 39327 23381 39485
rect 23417 39360 23510 39426
tri 23417 39344 23433 39360 ne
rect 23433 39344 23510 39360
rect 23250 39245 23398 39327
rect 23138 39212 23215 39228
tri 23215 39212 23231 39228 sw
rect 23138 39146 23231 39212
rect 23138 39044 23231 39110
rect 23138 39028 23215 39044
tri 23215 39028 23231 39044 nw
rect 23267 39011 23381 39245
tri 23417 39212 23433 39228 se
rect 23433 39212 23510 39228
rect 23417 39146 23510 39212
rect 23417 39044 23510 39110
tri 23417 39028 23433 39044 ne
rect 23433 39028 23510 39044
rect 23250 38929 23398 39011
rect 23138 38896 23215 38912
tri 23215 38896 23231 38912 sw
rect 23138 38830 23231 38896
rect 23267 38771 23381 38929
tri 23417 38896 23433 38912 se
rect 23433 38896 23510 38912
rect 23417 38830 23510 38896
rect 23138 38695 23510 38771
rect 23138 38570 23231 38636
rect 23138 38554 23215 38570
tri 23215 38554 23231 38570 nw
rect 23267 38537 23381 38695
rect 23417 38570 23510 38636
tri 23417 38554 23433 38570 ne
rect 23433 38554 23510 38570
rect 23250 38455 23398 38537
rect 23138 38422 23215 38438
tri 23215 38422 23231 38438 sw
rect 23138 38356 23231 38422
rect 23138 38254 23231 38320
rect 23138 38238 23215 38254
tri 23215 38238 23231 38254 nw
rect 23267 38221 23381 38455
tri 23417 38422 23433 38438 se
rect 23433 38422 23510 38438
rect 23417 38356 23510 38422
rect 23417 38254 23510 38320
tri 23417 38238 23433 38254 ne
rect 23433 38238 23510 38254
rect 23250 38139 23398 38221
rect 23138 38106 23215 38122
tri 23215 38106 23231 38122 sw
rect 23138 38040 23231 38106
rect 23267 37981 23381 38139
tri 23417 38106 23433 38122 se
rect 23433 38106 23510 38122
rect 23417 38040 23510 38106
rect 23138 37905 23510 37981
rect 23138 37780 23231 37846
rect 23138 37764 23215 37780
tri 23215 37764 23231 37780 nw
rect 23267 37747 23381 37905
rect 23417 37780 23510 37846
tri 23417 37764 23433 37780 ne
rect 23433 37764 23510 37780
rect 23250 37665 23398 37747
rect 23138 37632 23215 37648
tri 23215 37632 23231 37648 sw
rect 23138 37566 23231 37632
rect 23138 37464 23231 37530
rect 23138 37448 23215 37464
tri 23215 37448 23231 37464 nw
rect 23267 37431 23381 37665
tri 23417 37632 23433 37648 se
rect 23433 37632 23510 37648
rect 23417 37566 23510 37632
rect 23417 37464 23510 37530
tri 23417 37448 23433 37464 ne
rect 23433 37448 23510 37464
rect 23250 37349 23398 37431
rect 23138 37316 23215 37332
tri 23215 37316 23231 37332 sw
rect 23138 37250 23231 37316
rect 23267 37191 23381 37349
tri 23417 37316 23433 37332 se
rect 23433 37316 23510 37332
rect 23417 37250 23510 37316
rect 23138 37115 23510 37191
rect 23138 36990 23231 37056
rect 23138 36974 23215 36990
tri 23215 36974 23231 36990 nw
rect 23267 36957 23381 37115
rect 23417 36990 23510 37056
tri 23417 36974 23433 36990 ne
rect 23433 36974 23510 36990
rect 23250 36875 23398 36957
rect 23138 36842 23215 36858
tri 23215 36842 23231 36858 sw
rect 23138 36776 23231 36842
rect 23138 36674 23231 36740
rect 23138 36658 23215 36674
tri 23215 36658 23231 36674 nw
rect 23267 36641 23381 36875
tri 23417 36842 23433 36858 se
rect 23433 36842 23510 36858
rect 23417 36776 23510 36842
rect 23417 36674 23510 36740
tri 23417 36658 23433 36674 ne
rect 23433 36658 23510 36674
rect 23250 36559 23398 36641
rect 23138 36526 23215 36542
tri 23215 36526 23231 36542 sw
rect 23138 36460 23231 36526
rect 23267 36401 23381 36559
tri 23417 36526 23433 36542 se
rect 23433 36526 23510 36542
rect 23417 36460 23510 36526
rect 23138 36325 23510 36401
rect 23138 36200 23231 36266
rect 23138 36184 23215 36200
tri 23215 36184 23231 36200 nw
rect 23267 36167 23381 36325
rect 23417 36200 23510 36266
tri 23417 36184 23433 36200 ne
rect 23433 36184 23510 36200
rect 23250 36085 23398 36167
rect 23138 36052 23215 36068
tri 23215 36052 23231 36068 sw
rect 23138 35986 23231 36052
rect 23138 35884 23231 35950
rect 23138 35868 23215 35884
tri 23215 35868 23231 35884 nw
rect 23267 35851 23381 36085
tri 23417 36052 23433 36068 se
rect 23433 36052 23510 36068
rect 23417 35986 23510 36052
rect 23417 35884 23510 35950
tri 23417 35868 23433 35884 ne
rect 23433 35868 23510 35884
rect 23250 35769 23398 35851
rect 23138 35736 23215 35752
tri 23215 35736 23231 35752 sw
rect 23138 35670 23231 35736
rect 23267 35611 23381 35769
tri 23417 35736 23433 35752 se
rect 23433 35736 23510 35752
rect 23417 35670 23510 35736
rect 23138 35535 23510 35611
rect 23138 35410 23231 35476
rect 23138 35394 23215 35410
tri 23215 35394 23231 35410 nw
rect 23267 35377 23381 35535
rect 23417 35410 23510 35476
tri 23417 35394 23433 35410 ne
rect 23433 35394 23510 35410
rect 23250 35295 23398 35377
rect 23138 35262 23215 35278
tri 23215 35262 23231 35278 sw
rect 23138 35196 23231 35262
rect 23138 35094 23231 35160
rect 23138 35078 23215 35094
tri 23215 35078 23231 35094 nw
rect 23267 35061 23381 35295
tri 23417 35262 23433 35278 se
rect 23433 35262 23510 35278
rect 23417 35196 23510 35262
rect 23417 35094 23510 35160
tri 23417 35078 23433 35094 ne
rect 23433 35078 23510 35094
rect 23250 34979 23398 35061
rect 23138 34946 23215 34962
tri 23215 34946 23231 34962 sw
rect 23138 34880 23231 34946
rect 23267 34821 23381 34979
tri 23417 34946 23433 34962 se
rect 23433 34946 23510 34962
rect 23417 34880 23510 34946
rect 23138 34745 23510 34821
rect 23138 34620 23231 34686
rect 23138 34604 23215 34620
tri 23215 34604 23231 34620 nw
rect 23267 34587 23381 34745
rect 23417 34620 23510 34686
tri 23417 34604 23433 34620 ne
rect 23433 34604 23510 34620
rect 23250 34505 23398 34587
rect 23138 34472 23215 34488
tri 23215 34472 23231 34488 sw
rect 23138 34406 23231 34472
rect 23138 34304 23231 34370
rect 23138 34288 23215 34304
tri 23215 34288 23231 34304 nw
rect 23267 34271 23381 34505
tri 23417 34472 23433 34488 se
rect 23433 34472 23510 34488
rect 23417 34406 23510 34472
rect 23417 34304 23510 34370
tri 23417 34288 23433 34304 ne
rect 23433 34288 23510 34304
rect 23250 34189 23398 34271
rect 23138 34156 23215 34172
tri 23215 34156 23231 34172 sw
rect 23138 34090 23231 34156
rect 23267 34031 23381 34189
tri 23417 34156 23433 34172 se
rect 23433 34156 23510 34172
rect 23417 34090 23510 34156
rect 23138 33955 23510 34031
rect 23138 33830 23231 33896
rect 23138 33814 23215 33830
tri 23215 33814 23231 33830 nw
rect 23267 33797 23381 33955
rect 23417 33830 23510 33896
tri 23417 33814 23433 33830 ne
rect 23433 33814 23510 33830
rect 23250 33715 23398 33797
rect 23138 33682 23215 33698
tri 23215 33682 23231 33698 sw
rect 23138 33616 23231 33682
rect 23138 33514 23231 33580
rect 23138 33498 23215 33514
tri 23215 33498 23231 33514 nw
rect 23267 33481 23381 33715
tri 23417 33682 23433 33698 se
rect 23433 33682 23510 33698
rect 23417 33616 23510 33682
rect 23417 33514 23510 33580
tri 23417 33498 23433 33514 ne
rect 23433 33498 23510 33514
rect 23250 33399 23398 33481
rect 23138 33366 23215 33382
tri 23215 33366 23231 33382 sw
rect 23138 33300 23231 33366
rect 23267 33241 23381 33399
tri 23417 33366 23433 33382 se
rect 23433 33366 23510 33382
rect 23417 33300 23510 33366
rect 23138 33165 23510 33241
rect 23138 33040 23231 33106
rect 23138 33024 23215 33040
tri 23215 33024 23231 33040 nw
rect 23267 33007 23381 33165
rect 23417 33040 23510 33106
tri 23417 33024 23433 33040 ne
rect 23433 33024 23510 33040
rect 23250 32925 23398 33007
rect 23138 32892 23215 32908
tri 23215 32892 23231 32908 sw
rect 23138 32826 23231 32892
rect 23138 32724 23231 32790
rect 23138 32708 23215 32724
tri 23215 32708 23231 32724 nw
rect 23267 32691 23381 32925
tri 23417 32892 23433 32908 se
rect 23433 32892 23510 32908
rect 23417 32826 23510 32892
rect 23417 32724 23510 32790
tri 23417 32708 23433 32724 ne
rect 23433 32708 23510 32724
rect 23250 32609 23398 32691
rect 23138 32576 23215 32592
tri 23215 32576 23231 32592 sw
rect 23138 32510 23231 32576
rect 23267 32451 23381 32609
tri 23417 32576 23433 32592 se
rect 23433 32576 23510 32592
rect 23417 32510 23510 32576
rect 23138 32375 23510 32451
rect 23138 32250 23231 32316
rect 23138 32234 23215 32250
tri 23215 32234 23231 32250 nw
rect 23267 32217 23381 32375
rect 23417 32250 23510 32316
tri 23417 32234 23433 32250 ne
rect 23433 32234 23510 32250
rect 23250 32135 23398 32217
rect 23138 32102 23215 32118
tri 23215 32102 23231 32118 sw
rect 23138 32036 23231 32102
rect 23138 31934 23231 32000
rect 23138 31918 23215 31934
tri 23215 31918 23231 31934 nw
rect 23267 31901 23381 32135
tri 23417 32102 23433 32118 se
rect 23433 32102 23510 32118
rect 23417 32036 23510 32102
rect 23417 31934 23510 32000
tri 23417 31918 23433 31934 ne
rect 23433 31918 23510 31934
rect 23250 31819 23398 31901
rect 23138 31786 23215 31802
tri 23215 31786 23231 31802 sw
rect 23138 31720 23231 31786
rect 23267 31661 23381 31819
tri 23417 31786 23433 31802 se
rect 23433 31786 23510 31802
rect 23417 31720 23510 31786
rect 23138 31585 23510 31661
rect 23138 31460 23231 31526
rect 23138 31444 23215 31460
tri 23215 31444 23231 31460 nw
rect 23267 31427 23381 31585
rect 23417 31460 23510 31526
tri 23417 31444 23433 31460 ne
rect 23433 31444 23510 31460
rect 23250 31345 23398 31427
rect 23138 31312 23215 31328
tri 23215 31312 23231 31328 sw
rect 23138 31246 23231 31312
rect 23138 31144 23231 31210
rect 23138 31128 23215 31144
tri 23215 31128 23231 31144 nw
rect 23267 31111 23381 31345
tri 23417 31312 23433 31328 se
rect 23433 31312 23510 31328
rect 23417 31246 23510 31312
rect 23417 31144 23510 31210
tri 23417 31128 23433 31144 ne
rect 23433 31128 23510 31144
rect 23250 31029 23398 31111
rect 23138 30996 23215 31012
tri 23215 30996 23231 31012 sw
rect 23138 30930 23231 30996
rect 23267 30871 23381 31029
tri 23417 30996 23433 31012 se
rect 23433 30996 23510 31012
rect 23417 30930 23510 30996
rect 23138 30795 23510 30871
rect 23138 30670 23231 30736
rect 23138 30654 23215 30670
tri 23215 30654 23231 30670 nw
rect 23267 30637 23381 30795
rect 23417 30670 23510 30736
tri 23417 30654 23433 30670 ne
rect 23433 30654 23510 30670
rect 23250 30555 23398 30637
rect 23138 30522 23215 30538
tri 23215 30522 23231 30538 sw
rect 23138 30456 23231 30522
rect 23138 30354 23231 30420
rect 23138 30338 23215 30354
tri 23215 30338 23231 30354 nw
rect 23267 30321 23381 30555
tri 23417 30522 23433 30538 se
rect 23433 30522 23510 30538
rect 23417 30456 23510 30522
rect 23417 30354 23510 30420
tri 23417 30338 23433 30354 ne
rect 23433 30338 23510 30354
rect 23250 30239 23398 30321
rect 23138 30206 23215 30222
tri 23215 30206 23231 30222 sw
rect 23138 30140 23231 30206
rect 23267 30081 23381 30239
tri 23417 30206 23433 30222 se
rect 23433 30206 23510 30222
rect 23417 30140 23510 30206
rect 23138 30005 23510 30081
rect 23138 29880 23231 29946
rect 23138 29864 23215 29880
tri 23215 29864 23231 29880 nw
rect 23267 29847 23381 30005
rect 23417 29880 23510 29946
tri 23417 29864 23433 29880 ne
rect 23433 29864 23510 29880
rect 23250 29765 23398 29847
rect 23138 29732 23215 29748
tri 23215 29732 23231 29748 sw
rect 23138 29666 23231 29732
rect 23138 29564 23231 29630
rect 23138 29548 23215 29564
tri 23215 29548 23231 29564 nw
rect 23267 29531 23381 29765
tri 23417 29732 23433 29748 se
rect 23433 29732 23510 29748
rect 23417 29666 23510 29732
rect 23417 29564 23510 29630
tri 23417 29548 23433 29564 ne
rect 23433 29548 23510 29564
rect 23250 29449 23398 29531
rect 23138 29416 23215 29432
tri 23215 29416 23231 29432 sw
rect 23138 29350 23231 29416
rect 23267 29291 23381 29449
tri 23417 29416 23433 29432 se
rect 23433 29416 23510 29432
rect 23417 29350 23510 29416
rect 23138 29215 23510 29291
rect 23138 29090 23231 29156
rect 23138 29074 23215 29090
tri 23215 29074 23231 29090 nw
rect 23267 29057 23381 29215
rect 23417 29090 23510 29156
tri 23417 29074 23433 29090 ne
rect 23433 29074 23510 29090
rect 23250 28975 23398 29057
rect 23138 28942 23215 28958
tri 23215 28942 23231 28958 sw
rect 23138 28876 23231 28942
rect 23267 28833 23381 28975
tri 23417 28942 23433 28958 se
rect 23433 28942 23510 28958
rect 23417 28876 23510 28942
rect 23546 28463 23582 80603
rect 23618 28463 23654 80603
rect 23690 80445 23726 80603
rect 23682 80303 23734 80445
rect 23690 28763 23726 80303
rect 23682 28621 23734 28763
rect 23690 28463 23726 28621
rect 23762 28463 23798 80603
rect 23834 28463 23870 80603
rect 23906 28833 23990 80233
rect 24026 28463 24062 80603
rect 24098 28463 24134 80603
rect 24170 80445 24206 80603
rect 24162 80303 24214 80445
rect 24170 28763 24206 80303
rect 24162 28621 24214 28763
rect 24170 28463 24206 28621
rect 24242 28463 24278 80603
rect 24314 28463 24350 80603
rect 24386 80124 24479 80190
rect 24386 80108 24463 80124
tri 24463 80108 24479 80124 nw
rect 24515 80091 24629 80233
rect 24665 80124 24758 80190
tri 24665 80108 24681 80124 ne
rect 24681 80108 24758 80124
rect 24498 80009 24646 80091
rect 24386 79976 24463 79992
tri 24463 79976 24479 79992 sw
rect 24386 79910 24479 79976
rect 24515 79851 24629 80009
tri 24665 79976 24681 79992 se
rect 24681 79976 24758 79992
rect 24665 79910 24758 79976
rect 24386 79775 24758 79851
rect 24386 79650 24479 79716
rect 24386 79634 24463 79650
tri 24463 79634 24479 79650 nw
rect 24515 79617 24629 79775
rect 24665 79650 24758 79716
tri 24665 79634 24681 79650 ne
rect 24681 79634 24758 79650
rect 24498 79535 24646 79617
rect 24386 79502 24463 79518
tri 24463 79502 24479 79518 sw
rect 24386 79436 24479 79502
rect 24386 79334 24479 79400
rect 24386 79318 24463 79334
tri 24463 79318 24479 79334 nw
rect 24515 79301 24629 79535
tri 24665 79502 24681 79518 se
rect 24681 79502 24758 79518
rect 24665 79436 24758 79502
rect 24665 79334 24758 79400
tri 24665 79318 24681 79334 ne
rect 24681 79318 24758 79334
rect 24498 79219 24646 79301
rect 24386 79186 24463 79202
tri 24463 79186 24479 79202 sw
rect 24386 79120 24479 79186
rect 24515 79061 24629 79219
tri 24665 79186 24681 79202 se
rect 24681 79186 24758 79202
rect 24665 79120 24758 79186
rect 24386 78985 24758 79061
rect 24386 78860 24479 78926
rect 24386 78844 24463 78860
tri 24463 78844 24479 78860 nw
rect 24515 78827 24629 78985
rect 24665 78860 24758 78926
tri 24665 78844 24681 78860 ne
rect 24681 78844 24758 78860
rect 24498 78745 24646 78827
rect 24386 78712 24463 78728
tri 24463 78712 24479 78728 sw
rect 24386 78646 24479 78712
rect 24386 78544 24479 78610
rect 24386 78528 24463 78544
tri 24463 78528 24479 78544 nw
rect 24515 78511 24629 78745
tri 24665 78712 24681 78728 se
rect 24681 78712 24758 78728
rect 24665 78646 24758 78712
rect 24665 78544 24758 78610
tri 24665 78528 24681 78544 ne
rect 24681 78528 24758 78544
rect 24498 78429 24646 78511
rect 24386 78396 24463 78412
tri 24463 78396 24479 78412 sw
rect 24386 78330 24479 78396
rect 24515 78271 24629 78429
tri 24665 78396 24681 78412 se
rect 24681 78396 24758 78412
rect 24665 78330 24758 78396
rect 24386 78195 24758 78271
rect 24386 78070 24479 78136
rect 24386 78054 24463 78070
tri 24463 78054 24479 78070 nw
rect 24515 78037 24629 78195
rect 24665 78070 24758 78136
tri 24665 78054 24681 78070 ne
rect 24681 78054 24758 78070
rect 24498 77955 24646 78037
rect 24386 77922 24463 77938
tri 24463 77922 24479 77938 sw
rect 24386 77856 24479 77922
rect 24386 77754 24479 77820
rect 24386 77738 24463 77754
tri 24463 77738 24479 77754 nw
rect 24515 77721 24629 77955
tri 24665 77922 24681 77938 se
rect 24681 77922 24758 77938
rect 24665 77856 24758 77922
rect 24665 77754 24758 77820
tri 24665 77738 24681 77754 ne
rect 24681 77738 24758 77754
rect 24498 77639 24646 77721
rect 24386 77606 24463 77622
tri 24463 77606 24479 77622 sw
rect 24386 77540 24479 77606
rect 24515 77481 24629 77639
tri 24665 77606 24681 77622 se
rect 24681 77606 24758 77622
rect 24665 77540 24758 77606
rect 24386 77405 24758 77481
rect 24386 77280 24479 77346
rect 24386 77264 24463 77280
tri 24463 77264 24479 77280 nw
rect 24515 77247 24629 77405
rect 24665 77280 24758 77346
tri 24665 77264 24681 77280 ne
rect 24681 77264 24758 77280
rect 24498 77165 24646 77247
rect 24386 77132 24463 77148
tri 24463 77132 24479 77148 sw
rect 24386 77066 24479 77132
rect 24386 76964 24479 77030
rect 24386 76948 24463 76964
tri 24463 76948 24479 76964 nw
rect 24515 76931 24629 77165
tri 24665 77132 24681 77148 se
rect 24681 77132 24758 77148
rect 24665 77066 24758 77132
rect 24665 76964 24758 77030
tri 24665 76948 24681 76964 ne
rect 24681 76948 24758 76964
rect 24498 76849 24646 76931
rect 24386 76816 24463 76832
tri 24463 76816 24479 76832 sw
rect 24386 76750 24479 76816
rect 24515 76691 24629 76849
tri 24665 76816 24681 76832 se
rect 24681 76816 24758 76832
rect 24665 76750 24758 76816
rect 24386 76615 24758 76691
rect 24386 76490 24479 76556
rect 24386 76474 24463 76490
tri 24463 76474 24479 76490 nw
rect 24515 76457 24629 76615
rect 24665 76490 24758 76556
tri 24665 76474 24681 76490 ne
rect 24681 76474 24758 76490
rect 24498 76375 24646 76457
rect 24386 76342 24463 76358
tri 24463 76342 24479 76358 sw
rect 24386 76276 24479 76342
rect 24386 76174 24479 76240
rect 24386 76158 24463 76174
tri 24463 76158 24479 76174 nw
rect 24515 76141 24629 76375
tri 24665 76342 24681 76358 se
rect 24681 76342 24758 76358
rect 24665 76276 24758 76342
rect 24665 76174 24758 76240
tri 24665 76158 24681 76174 ne
rect 24681 76158 24758 76174
rect 24498 76059 24646 76141
rect 24386 76026 24463 76042
tri 24463 76026 24479 76042 sw
rect 24386 75960 24479 76026
rect 24515 75901 24629 76059
tri 24665 76026 24681 76042 se
rect 24681 76026 24758 76042
rect 24665 75960 24758 76026
rect 24386 75825 24758 75901
rect 24386 75700 24479 75766
rect 24386 75684 24463 75700
tri 24463 75684 24479 75700 nw
rect 24515 75667 24629 75825
rect 24665 75700 24758 75766
tri 24665 75684 24681 75700 ne
rect 24681 75684 24758 75700
rect 24498 75585 24646 75667
rect 24386 75552 24463 75568
tri 24463 75552 24479 75568 sw
rect 24386 75486 24479 75552
rect 24386 75384 24479 75450
rect 24386 75368 24463 75384
tri 24463 75368 24479 75384 nw
rect 24515 75351 24629 75585
tri 24665 75552 24681 75568 se
rect 24681 75552 24758 75568
rect 24665 75486 24758 75552
rect 24665 75384 24758 75450
tri 24665 75368 24681 75384 ne
rect 24681 75368 24758 75384
rect 24498 75269 24646 75351
rect 24386 75236 24463 75252
tri 24463 75236 24479 75252 sw
rect 24386 75170 24479 75236
rect 24515 75111 24629 75269
tri 24665 75236 24681 75252 se
rect 24681 75236 24758 75252
rect 24665 75170 24758 75236
rect 24386 75035 24758 75111
rect 24386 74910 24479 74976
rect 24386 74894 24463 74910
tri 24463 74894 24479 74910 nw
rect 24515 74877 24629 75035
rect 24665 74910 24758 74976
tri 24665 74894 24681 74910 ne
rect 24681 74894 24758 74910
rect 24498 74795 24646 74877
rect 24386 74762 24463 74778
tri 24463 74762 24479 74778 sw
rect 24386 74696 24479 74762
rect 24386 74594 24479 74660
rect 24386 74578 24463 74594
tri 24463 74578 24479 74594 nw
rect 24515 74561 24629 74795
tri 24665 74762 24681 74778 se
rect 24681 74762 24758 74778
rect 24665 74696 24758 74762
rect 24665 74594 24758 74660
tri 24665 74578 24681 74594 ne
rect 24681 74578 24758 74594
rect 24498 74479 24646 74561
rect 24386 74446 24463 74462
tri 24463 74446 24479 74462 sw
rect 24386 74380 24479 74446
rect 24515 74321 24629 74479
tri 24665 74446 24681 74462 se
rect 24681 74446 24758 74462
rect 24665 74380 24758 74446
rect 24386 74245 24758 74321
rect 24386 74120 24479 74186
rect 24386 74104 24463 74120
tri 24463 74104 24479 74120 nw
rect 24515 74087 24629 74245
rect 24665 74120 24758 74186
tri 24665 74104 24681 74120 ne
rect 24681 74104 24758 74120
rect 24498 74005 24646 74087
rect 24386 73972 24463 73988
tri 24463 73972 24479 73988 sw
rect 24386 73906 24479 73972
rect 24386 73804 24479 73870
rect 24386 73788 24463 73804
tri 24463 73788 24479 73804 nw
rect 24515 73771 24629 74005
tri 24665 73972 24681 73988 se
rect 24681 73972 24758 73988
rect 24665 73906 24758 73972
rect 24665 73804 24758 73870
tri 24665 73788 24681 73804 ne
rect 24681 73788 24758 73804
rect 24498 73689 24646 73771
rect 24386 73656 24463 73672
tri 24463 73656 24479 73672 sw
rect 24386 73590 24479 73656
rect 24515 73531 24629 73689
tri 24665 73656 24681 73672 se
rect 24681 73656 24758 73672
rect 24665 73590 24758 73656
rect 24386 73455 24758 73531
rect 24386 73330 24479 73396
rect 24386 73314 24463 73330
tri 24463 73314 24479 73330 nw
rect 24515 73297 24629 73455
rect 24665 73330 24758 73396
tri 24665 73314 24681 73330 ne
rect 24681 73314 24758 73330
rect 24498 73215 24646 73297
rect 24386 73182 24463 73198
tri 24463 73182 24479 73198 sw
rect 24386 73116 24479 73182
rect 24386 73014 24479 73080
rect 24386 72998 24463 73014
tri 24463 72998 24479 73014 nw
rect 24515 72981 24629 73215
tri 24665 73182 24681 73198 se
rect 24681 73182 24758 73198
rect 24665 73116 24758 73182
rect 24665 73014 24758 73080
tri 24665 72998 24681 73014 ne
rect 24681 72998 24758 73014
rect 24498 72899 24646 72981
rect 24386 72866 24463 72882
tri 24463 72866 24479 72882 sw
rect 24386 72800 24479 72866
rect 24515 72741 24629 72899
tri 24665 72866 24681 72882 se
rect 24681 72866 24758 72882
rect 24665 72800 24758 72866
rect 24386 72665 24758 72741
rect 24386 72540 24479 72606
rect 24386 72524 24463 72540
tri 24463 72524 24479 72540 nw
rect 24515 72507 24629 72665
rect 24665 72540 24758 72606
tri 24665 72524 24681 72540 ne
rect 24681 72524 24758 72540
rect 24498 72425 24646 72507
rect 24386 72392 24463 72408
tri 24463 72392 24479 72408 sw
rect 24386 72326 24479 72392
rect 24386 72224 24479 72290
rect 24386 72208 24463 72224
tri 24463 72208 24479 72224 nw
rect 24515 72191 24629 72425
tri 24665 72392 24681 72408 se
rect 24681 72392 24758 72408
rect 24665 72326 24758 72392
rect 24665 72224 24758 72290
tri 24665 72208 24681 72224 ne
rect 24681 72208 24758 72224
rect 24498 72109 24646 72191
rect 24386 72076 24463 72092
tri 24463 72076 24479 72092 sw
rect 24386 72010 24479 72076
rect 24515 71951 24629 72109
tri 24665 72076 24681 72092 se
rect 24681 72076 24758 72092
rect 24665 72010 24758 72076
rect 24386 71875 24758 71951
rect 24386 71750 24479 71816
rect 24386 71734 24463 71750
tri 24463 71734 24479 71750 nw
rect 24515 71717 24629 71875
rect 24665 71750 24758 71816
tri 24665 71734 24681 71750 ne
rect 24681 71734 24758 71750
rect 24498 71635 24646 71717
rect 24386 71602 24463 71618
tri 24463 71602 24479 71618 sw
rect 24386 71536 24479 71602
rect 24386 71434 24479 71500
rect 24386 71418 24463 71434
tri 24463 71418 24479 71434 nw
rect 24515 71401 24629 71635
tri 24665 71602 24681 71618 se
rect 24681 71602 24758 71618
rect 24665 71536 24758 71602
rect 24665 71434 24758 71500
tri 24665 71418 24681 71434 ne
rect 24681 71418 24758 71434
rect 24498 71319 24646 71401
rect 24386 71286 24463 71302
tri 24463 71286 24479 71302 sw
rect 24386 71220 24479 71286
rect 24515 71161 24629 71319
tri 24665 71286 24681 71302 se
rect 24681 71286 24758 71302
rect 24665 71220 24758 71286
rect 24386 71085 24758 71161
rect 24386 70960 24479 71026
rect 24386 70944 24463 70960
tri 24463 70944 24479 70960 nw
rect 24515 70927 24629 71085
rect 24665 70960 24758 71026
tri 24665 70944 24681 70960 ne
rect 24681 70944 24758 70960
rect 24498 70845 24646 70927
rect 24386 70812 24463 70828
tri 24463 70812 24479 70828 sw
rect 24386 70746 24479 70812
rect 24386 70644 24479 70710
rect 24386 70628 24463 70644
tri 24463 70628 24479 70644 nw
rect 24515 70611 24629 70845
tri 24665 70812 24681 70828 se
rect 24681 70812 24758 70828
rect 24665 70746 24758 70812
rect 24665 70644 24758 70710
tri 24665 70628 24681 70644 ne
rect 24681 70628 24758 70644
rect 24498 70529 24646 70611
rect 24386 70496 24463 70512
tri 24463 70496 24479 70512 sw
rect 24386 70430 24479 70496
rect 24515 70371 24629 70529
tri 24665 70496 24681 70512 se
rect 24681 70496 24758 70512
rect 24665 70430 24758 70496
rect 24386 70295 24758 70371
rect 24386 70170 24479 70236
rect 24386 70154 24463 70170
tri 24463 70154 24479 70170 nw
rect 24515 70137 24629 70295
rect 24665 70170 24758 70236
tri 24665 70154 24681 70170 ne
rect 24681 70154 24758 70170
rect 24498 70055 24646 70137
rect 24386 70022 24463 70038
tri 24463 70022 24479 70038 sw
rect 24386 69956 24479 70022
rect 24386 69854 24479 69920
rect 24386 69838 24463 69854
tri 24463 69838 24479 69854 nw
rect 24515 69821 24629 70055
tri 24665 70022 24681 70038 se
rect 24681 70022 24758 70038
rect 24665 69956 24758 70022
rect 24665 69854 24758 69920
tri 24665 69838 24681 69854 ne
rect 24681 69838 24758 69854
rect 24498 69739 24646 69821
rect 24386 69706 24463 69722
tri 24463 69706 24479 69722 sw
rect 24386 69640 24479 69706
rect 24515 69581 24629 69739
tri 24665 69706 24681 69722 se
rect 24681 69706 24758 69722
rect 24665 69640 24758 69706
rect 24386 69505 24758 69581
rect 24386 69380 24479 69446
rect 24386 69364 24463 69380
tri 24463 69364 24479 69380 nw
rect 24515 69347 24629 69505
rect 24665 69380 24758 69446
tri 24665 69364 24681 69380 ne
rect 24681 69364 24758 69380
rect 24498 69265 24646 69347
rect 24386 69232 24463 69248
tri 24463 69232 24479 69248 sw
rect 24386 69166 24479 69232
rect 24386 69064 24479 69130
rect 24386 69048 24463 69064
tri 24463 69048 24479 69064 nw
rect 24515 69031 24629 69265
tri 24665 69232 24681 69248 se
rect 24681 69232 24758 69248
rect 24665 69166 24758 69232
rect 24665 69064 24758 69130
tri 24665 69048 24681 69064 ne
rect 24681 69048 24758 69064
rect 24498 68949 24646 69031
rect 24386 68916 24463 68932
tri 24463 68916 24479 68932 sw
rect 24386 68850 24479 68916
rect 24515 68791 24629 68949
tri 24665 68916 24681 68932 se
rect 24681 68916 24758 68932
rect 24665 68850 24758 68916
rect 24386 68715 24758 68791
rect 24386 68590 24479 68656
rect 24386 68574 24463 68590
tri 24463 68574 24479 68590 nw
rect 24515 68557 24629 68715
rect 24665 68590 24758 68656
tri 24665 68574 24681 68590 ne
rect 24681 68574 24758 68590
rect 24498 68475 24646 68557
rect 24386 68442 24463 68458
tri 24463 68442 24479 68458 sw
rect 24386 68376 24479 68442
rect 24386 68274 24479 68340
rect 24386 68258 24463 68274
tri 24463 68258 24479 68274 nw
rect 24515 68241 24629 68475
tri 24665 68442 24681 68458 se
rect 24681 68442 24758 68458
rect 24665 68376 24758 68442
rect 24665 68274 24758 68340
tri 24665 68258 24681 68274 ne
rect 24681 68258 24758 68274
rect 24498 68159 24646 68241
rect 24386 68126 24463 68142
tri 24463 68126 24479 68142 sw
rect 24386 68060 24479 68126
rect 24515 68001 24629 68159
tri 24665 68126 24681 68142 se
rect 24681 68126 24758 68142
rect 24665 68060 24758 68126
rect 24386 67925 24758 68001
rect 24386 67800 24479 67866
rect 24386 67784 24463 67800
tri 24463 67784 24479 67800 nw
rect 24515 67767 24629 67925
rect 24665 67800 24758 67866
tri 24665 67784 24681 67800 ne
rect 24681 67784 24758 67800
rect 24498 67685 24646 67767
rect 24386 67652 24463 67668
tri 24463 67652 24479 67668 sw
rect 24386 67586 24479 67652
rect 24386 67484 24479 67550
rect 24386 67468 24463 67484
tri 24463 67468 24479 67484 nw
rect 24515 67451 24629 67685
tri 24665 67652 24681 67668 se
rect 24681 67652 24758 67668
rect 24665 67586 24758 67652
rect 24665 67484 24758 67550
tri 24665 67468 24681 67484 ne
rect 24681 67468 24758 67484
rect 24498 67369 24646 67451
rect 24386 67336 24463 67352
tri 24463 67336 24479 67352 sw
rect 24386 67270 24479 67336
rect 24515 67211 24629 67369
tri 24665 67336 24681 67352 se
rect 24681 67336 24758 67352
rect 24665 67270 24758 67336
rect 24386 67135 24758 67211
rect 24386 67010 24479 67076
rect 24386 66994 24463 67010
tri 24463 66994 24479 67010 nw
rect 24515 66977 24629 67135
rect 24665 67010 24758 67076
tri 24665 66994 24681 67010 ne
rect 24681 66994 24758 67010
rect 24498 66895 24646 66977
rect 24386 66862 24463 66878
tri 24463 66862 24479 66878 sw
rect 24386 66796 24479 66862
rect 24386 66694 24479 66760
rect 24386 66678 24463 66694
tri 24463 66678 24479 66694 nw
rect 24515 66661 24629 66895
tri 24665 66862 24681 66878 se
rect 24681 66862 24758 66878
rect 24665 66796 24758 66862
rect 24665 66694 24758 66760
tri 24665 66678 24681 66694 ne
rect 24681 66678 24758 66694
rect 24498 66579 24646 66661
rect 24386 66546 24463 66562
tri 24463 66546 24479 66562 sw
rect 24386 66480 24479 66546
rect 24515 66421 24629 66579
tri 24665 66546 24681 66562 se
rect 24681 66546 24758 66562
rect 24665 66480 24758 66546
rect 24386 66345 24758 66421
rect 24386 66220 24479 66286
rect 24386 66204 24463 66220
tri 24463 66204 24479 66220 nw
rect 24515 66187 24629 66345
rect 24665 66220 24758 66286
tri 24665 66204 24681 66220 ne
rect 24681 66204 24758 66220
rect 24498 66105 24646 66187
rect 24386 66072 24463 66088
tri 24463 66072 24479 66088 sw
rect 24386 66006 24479 66072
rect 24386 65904 24479 65970
rect 24386 65888 24463 65904
tri 24463 65888 24479 65904 nw
rect 24515 65871 24629 66105
tri 24665 66072 24681 66088 se
rect 24681 66072 24758 66088
rect 24665 66006 24758 66072
rect 24665 65904 24758 65970
tri 24665 65888 24681 65904 ne
rect 24681 65888 24758 65904
rect 24498 65789 24646 65871
rect 24386 65756 24463 65772
tri 24463 65756 24479 65772 sw
rect 24386 65690 24479 65756
rect 24515 65631 24629 65789
tri 24665 65756 24681 65772 se
rect 24681 65756 24758 65772
rect 24665 65690 24758 65756
rect 24386 65555 24758 65631
rect 24386 65430 24479 65496
rect 24386 65414 24463 65430
tri 24463 65414 24479 65430 nw
rect 24515 65397 24629 65555
rect 24665 65430 24758 65496
tri 24665 65414 24681 65430 ne
rect 24681 65414 24758 65430
rect 24498 65315 24646 65397
rect 24386 65282 24463 65298
tri 24463 65282 24479 65298 sw
rect 24386 65216 24479 65282
rect 24386 65114 24479 65180
rect 24386 65098 24463 65114
tri 24463 65098 24479 65114 nw
rect 24515 65081 24629 65315
tri 24665 65282 24681 65298 se
rect 24681 65282 24758 65298
rect 24665 65216 24758 65282
rect 24665 65114 24758 65180
tri 24665 65098 24681 65114 ne
rect 24681 65098 24758 65114
rect 24498 64999 24646 65081
rect 24386 64966 24463 64982
tri 24463 64966 24479 64982 sw
rect 24386 64900 24479 64966
rect 24515 64841 24629 64999
tri 24665 64966 24681 64982 se
rect 24681 64966 24758 64982
rect 24665 64900 24758 64966
rect 24386 64765 24758 64841
rect 24386 64640 24479 64706
rect 24386 64624 24463 64640
tri 24463 64624 24479 64640 nw
rect 24515 64607 24629 64765
rect 24665 64640 24758 64706
tri 24665 64624 24681 64640 ne
rect 24681 64624 24758 64640
rect 24498 64525 24646 64607
rect 24386 64492 24463 64508
tri 24463 64492 24479 64508 sw
rect 24386 64426 24479 64492
rect 24386 64324 24479 64390
rect 24386 64308 24463 64324
tri 24463 64308 24479 64324 nw
rect 24515 64291 24629 64525
tri 24665 64492 24681 64508 se
rect 24681 64492 24758 64508
rect 24665 64426 24758 64492
rect 24665 64324 24758 64390
tri 24665 64308 24681 64324 ne
rect 24681 64308 24758 64324
rect 24498 64209 24646 64291
rect 24386 64176 24463 64192
tri 24463 64176 24479 64192 sw
rect 24386 64110 24479 64176
rect 24515 64051 24629 64209
tri 24665 64176 24681 64192 se
rect 24681 64176 24758 64192
rect 24665 64110 24758 64176
rect 24386 63975 24758 64051
rect 24386 63850 24479 63916
rect 24386 63834 24463 63850
tri 24463 63834 24479 63850 nw
rect 24515 63817 24629 63975
rect 24665 63850 24758 63916
tri 24665 63834 24681 63850 ne
rect 24681 63834 24758 63850
rect 24498 63735 24646 63817
rect 24386 63702 24463 63718
tri 24463 63702 24479 63718 sw
rect 24386 63636 24479 63702
rect 24386 63534 24479 63600
rect 24386 63518 24463 63534
tri 24463 63518 24479 63534 nw
rect 24515 63501 24629 63735
tri 24665 63702 24681 63718 se
rect 24681 63702 24758 63718
rect 24665 63636 24758 63702
rect 24665 63534 24758 63600
tri 24665 63518 24681 63534 ne
rect 24681 63518 24758 63534
rect 24498 63419 24646 63501
rect 24386 63386 24463 63402
tri 24463 63386 24479 63402 sw
rect 24386 63320 24479 63386
rect 24515 63261 24629 63419
tri 24665 63386 24681 63402 se
rect 24681 63386 24758 63402
rect 24665 63320 24758 63386
rect 24386 63185 24758 63261
rect 24386 63060 24479 63126
rect 24386 63044 24463 63060
tri 24463 63044 24479 63060 nw
rect 24515 63027 24629 63185
rect 24665 63060 24758 63126
tri 24665 63044 24681 63060 ne
rect 24681 63044 24758 63060
rect 24498 62945 24646 63027
rect 24386 62912 24463 62928
tri 24463 62912 24479 62928 sw
rect 24386 62846 24479 62912
rect 24386 62744 24479 62810
rect 24386 62728 24463 62744
tri 24463 62728 24479 62744 nw
rect 24515 62711 24629 62945
tri 24665 62912 24681 62928 se
rect 24681 62912 24758 62928
rect 24665 62846 24758 62912
rect 24665 62744 24758 62810
tri 24665 62728 24681 62744 ne
rect 24681 62728 24758 62744
rect 24498 62629 24646 62711
rect 24386 62596 24463 62612
tri 24463 62596 24479 62612 sw
rect 24386 62530 24479 62596
rect 24515 62471 24629 62629
tri 24665 62596 24681 62612 se
rect 24681 62596 24758 62612
rect 24665 62530 24758 62596
rect 24386 62395 24758 62471
rect 24386 62270 24479 62336
rect 24386 62254 24463 62270
tri 24463 62254 24479 62270 nw
rect 24515 62237 24629 62395
rect 24665 62270 24758 62336
tri 24665 62254 24681 62270 ne
rect 24681 62254 24758 62270
rect 24498 62155 24646 62237
rect 24386 62122 24463 62138
tri 24463 62122 24479 62138 sw
rect 24386 62056 24479 62122
rect 24386 61954 24479 62020
rect 24386 61938 24463 61954
tri 24463 61938 24479 61954 nw
rect 24515 61921 24629 62155
tri 24665 62122 24681 62138 se
rect 24681 62122 24758 62138
rect 24665 62056 24758 62122
rect 24665 61954 24758 62020
tri 24665 61938 24681 61954 ne
rect 24681 61938 24758 61954
rect 24498 61839 24646 61921
rect 24386 61806 24463 61822
tri 24463 61806 24479 61822 sw
rect 24386 61740 24479 61806
rect 24515 61681 24629 61839
tri 24665 61806 24681 61822 se
rect 24681 61806 24758 61822
rect 24665 61740 24758 61806
rect 24386 61605 24758 61681
rect 24386 61480 24479 61546
rect 24386 61464 24463 61480
tri 24463 61464 24479 61480 nw
rect 24515 61447 24629 61605
rect 24665 61480 24758 61546
tri 24665 61464 24681 61480 ne
rect 24681 61464 24758 61480
rect 24498 61365 24646 61447
rect 24386 61332 24463 61348
tri 24463 61332 24479 61348 sw
rect 24386 61266 24479 61332
rect 24386 61164 24479 61230
rect 24386 61148 24463 61164
tri 24463 61148 24479 61164 nw
rect 24515 61131 24629 61365
tri 24665 61332 24681 61348 se
rect 24681 61332 24758 61348
rect 24665 61266 24758 61332
rect 24665 61164 24758 61230
tri 24665 61148 24681 61164 ne
rect 24681 61148 24758 61164
rect 24498 61049 24646 61131
rect 24386 61016 24463 61032
tri 24463 61016 24479 61032 sw
rect 24386 60950 24479 61016
rect 24515 60891 24629 61049
tri 24665 61016 24681 61032 se
rect 24681 61016 24758 61032
rect 24665 60950 24758 61016
rect 24386 60815 24758 60891
rect 24386 60690 24479 60756
rect 24386 60674 24463 60690
tri 24463 60674 24479 60690 nw
rect 24515 60657 24629 60815
rect 24665 60690 24758 60756
tri 24665 60674 24681 60690 ne
rect 24681 60674 24758 60690
rect 24498 60575 24646 60657
rect 24386 60542 24463 60558
tri 24463 60542 24479 60558 sw
rect 24386 60476 24479 60542
rect 24386 60374 24479 60440
rect 24386 60358 24463 60374
tri 24463 60358 24479 60374 nw
rect 24515 60341 24629 60575
tri 24665 60542 24681 60558 se
rect 24681 60542 24758 60558
rect 24665 60476 24758 60542
rect 24665 60374 24758 60440
tri 24665 60358 24681 60374 ne
rect 24681 60358 24758 60374
rect 24498 60259 24646 60341
rect 24386 60226 24463 60242
tri 24463 60226 24479 60242 sw
rect 24386 60160 24479 60226
rect 24515 60101 24629 60259
tri 24665 60226 24681 60242 se
rect 24681 60226 24758 60242
rect 24665 60160 24758 60226
rect 24386 60025 24758 60101
rect 24386 59900 24479 59966
rect 24386 59884 24463 59900
tri 24463 59884 24479 59900 nw
rect 24515 59867 24629 60025
rect 24665 59900 24758 59966
tri 24665 59884 24681 59900 ne
rect 24681 59884 24758 59900
rect 24498 59785 24646 59867
rect 24386 59752 24463 59768
tri 24463 59752 24479 59768 sw
rect 24386 59686 24479 59752
rect 24386 59584 24479 59650
rect 24386 59568 24463 59584
tri 24463 59568 24479 59584 nw
rect 24515 59551 24629 59785
tri 24665 59752 24681 59768 se
rect 24681 59752 24758 59768
rect 24665 59686 24758 59752
rect 24665 59584 24758 59650
tri 24665 59568 24681 59584 ne
rect 24681 59568 24758 59584
rect 24498 59469 24646 59551
rect 24386 59436 24463 59452
tri 24463 59436 24479 59452 sw
rect 24386 59370 24479 59436
rect 24515 59311 24629 59469
tri 24665 59436 24681 59452 se
rect 24681 59436 24758 59452
rect 24665 59370 24758 59436
rect 24386 59235 24758 59311
rect 24386 59110 24479 59176
rect 24386 59094 24463 59110
tri 24463 59094 24479 59110 nw
rect 24515 59077 24629 59235
rect 24665 59110 24758 59176
tri 24665 59094 24681 59110 ne
rect 24681 59094 24758 59110
rect 24498 58995 24646 59077
rect 24386 58962 24463 58978
tri 24463 58962 24479 58978 sw
rect 24386 58896 24479 58962
rect 24386 58794 24479 58860
rect 24386 58778 24463 58794
tri 24463 58778 24479 58794 nw
rect 24515 58761 24629 58995
tri 24665 58962 24681 58978 se
rect 24681 58962 24758 58978
rect 24665 58896 24758 58962
rect 24665 58794 24758 58860
tri 24665 58778 24681 58794 ne
rect 24681 58778 24758 58794
rect 24498 58679 24646 58761
rect 24386 58646 24463 58662
tri 24463 58646 24479 58662 sw
rect 24386 58580 24479 58646
rect 24515 58521 24629 58679
tri 24665 58646 24681 58662 se
rect 24681 58646 24758 58662
rect 24665 58580 24758 58646
rect 24386 58445 24758 58521
rect 24386 58320 24479 58386
rect 24386 58304 24463 58320
tri 24463 58304 24479 58320 nw
rect 24515 58287 24629 58445
rect 24665 58320 24758 58386
tri 24665 58304 24681 58320 ne
rect 24681 58304 24758 58320
rect 24498 58205 24646 58287
rect 24386 58172 24463 58188
tri 24463 58172 24479 58188 sw
rect 24386 58106 24479 58172
rect 24386 58004 24479 58070
rect 24386 57988 24463 58004
tri 24463 57988 24479 58004 nw
rect 24515 57971 24629 58205
tri 24665 58172 24681 58188 se
rect 24681 58172 24758 58188
rect 24665 58106 24758 58172
rect 24665 58004 24758 58070
tri 24665 57988 24681 58004 ne
rect 24681 57988 24758 58004
rect 24498 57889 24646 57971
rect 24386 57856 24463 57872
tri 24463 57856 24479 57872 sw
rect 24386 57790 24479 57856
rect 24515 57731 24629 57889
tri 24665 57856 24681 57872 se
rect 24681 57856 24758 57872
rect 24665 57790 24758 57856
rect 24386 57655 24758 57731
rect 24386 57530 24479 57596
rect 24386 57514 24463 57530
tri 24463 57514 24479 57530 nw
rect 24515 57497 24629 57655
rect 24665 57530 24758 57596
tri 24665 57514 24681 57530 ne
rect 24681 57514 24758 57530
rect 24498 57415 24646 57497
rect 24386 57382 24463 57398
tri 24463 57382 24479 57398 sw
rect 24386 57316 24479 57382
rect 24386 57214 24479 57280
rect 24386 57198 24463 57214
tri 24463 57198 24479 57214 nw
rect 24515 57181 24629 57415
tri 24665 57382 24681 57398 se
rect 24681 57382 24758 57398
rect 24665 57316 24758 57382
rect 24665 57214 24758 57280
tri 24665 57198 24681 57214 ne
rect 24681 57198 24758 57214
rect 24498 57099 24646 57181
rect 24386 57066 24463 57082
tri 24463 57066 24479 57082 sw
rect 24386 57000 24479 57066
rect 24515 56941 24629 57099
tri 24665 57066 24681 57082 se
rect 24681 57066 24758 57082
rect 24665 57000 24758 57066
rect 24386 56865 24758 56941
rect 24386 56740 24479 56806
rect 24386 56724 24463 56740
tri 24463 56724 24479 56740 nw
rect 24515 56707 24629 56865
rect 24665 56740 24758 56806
tri 24665 56724 24681 56740 ne
rect 24681 56724 24758 56740
rect 24498 56625 24646 56707
rect 24386 56592 24463 56608
tri 24463 56592 24479 56608 sw
rect 24386 56526 24479 56592
rect 24386 56424 24479 56490
rect 24386 56408 24463 56424
tri 24463 56408 24479 56424 nw
rect 24515 56391 24629 56625
tri 24665 56592 24681 56608 se
rect 24681 56592 24758 56608
rect 24665 56526 24758 56592
rect 24665 56424 24758 56490
tri 24665 56408 24681 56424 ne
rect 24681 56408 24758 56424
rect 24498 56309 24646 56391
rect 24386 56276 24463 56292
tri 24463 56276 24479 56292 sw
rect 24386 56210 24479 56276
rect 24515 56151 24629 56309
tri 24665 56276 24681 56292 se
rect 24681 56276 24758 56292
rect 24665 56210 24758 56276
rect 24386 56075 24758 56151
rect 24386 55950 24479 56016
rect 24386 55934 24463 55950
tri 24463 55934 24479 55950 nw
rect 24515 55917 24629 56075
rect 24665 55950 24758 56016
tri 24665 55934 24681 55950 ne
rect 24681 55934 24758 55950
rect 24498 55835 24646 55917
rect 24386 55802 24463 55818
tri 24463 55802 24479 55818 sw
rect 24386 55736 24479 55802
rect 24386 55634 24479 55700
rect 24386 55618 24463 55634
tri 24463 55618 24479 55634 nw
rect 24515 55601 24629 55835
tri 24665 55802 24681 55818 se
rect 24681 55802 24758 55818
rect 24665 55736 24758 55802
rect 24665 55634 24758 55700
tri 24665 55618 24681 55634 ne
rect 24681 55618 24758 55634
rect 24498 55519 24646 55601
rect 24386 55486 24463 55502
tri 24463 55486 24479 55502 sw
rect 24386 55420 24479 55486
rect 24515 55361 24629 55519
tri 24665 55486 24681 55502 se
rect 24681 55486 24758 55502
rect 24665 55420 24758 55486
rect 24386 55285 24758 55361
rect 24386 55160 24479 55226
rect 24386 55144 24463 55160
tri 24463 55144 24479 55160 nw
rect 24515 55127 24629 55285
rect 24665 55160 24758 55226
tri 24665 55144 24681 55160 ne
rect 24681 55144 24758 55160
rect 24498 55045 24646 55127
rect 24386 55012 24463 55028
tri 24463 55012 24479 55028 sw
rect 24386 54946 24479 55012
rect 24386 54844 24479 54910
rect 24386 54828 24463 54844
tri 24463 54828 24479 54844 nw
rect 24515 54811 24629 55045
tri 24665 55012 24681 55028 se
rect 24681 55012 24758 55028
rect 24665 54946 24758 55012
rect 24665 54844 24758 54910
tri 24665 54828 24681 54844 ne
rect 24681 54828 24758 54844
rect 24498 54729 24646 54811
rect 24386 54696 24463 54712
tri 24463 54696 24479 54712 sw
rect 24386 54630 24479 54696
rect 24515 54571 24629 54729
tri 24665 54696 24681 54712 se
rect 24681 54696 24758 54712
rect 24665 54630 24758 54696
rect 24386 54495 24758 54571
rect 24386 54370 24479 54436
rect 24386 54354 24463 54370
tri 24463 54354 24479 54370 nw
rect 24515 54337 24629 54495
rect 24665 54370 24758 54436
tri 24665 54354 24681 54370 ne
rect 24681 54354 24758 54370
rect 24498 54255 24646 54337
rect 24386 54222 24463 54238
tri 24463 54222 24479 54238 sw
rect 24386 54156 24479 54222
rect 24386 54054 24479 54120
rect 24386 54038 24463 54054
tri 24463 54038 24479 54054 nw
rect 24515 54021 24629 54255
tri 24665 54222 24681 54238 se
rect 24681 54222 24758 54238
rect 24665 54156 24758 54222
rect 24665 54054 24758 54120
tri 24665 54038 24681 54054 ne
rect 24681 54038 24758 54054
rect 24498 53939 24646 54021
rect 24386 53906 24463 53922
tri 24463 53906 24479 53922 sw
rect 24386 53840 24479 53906
rect 24515 53781 24629 53939
tri 24665 53906 24681 53922 se
rect 24681 53906 24758 53922
rect 24665 53840 24758 53906
rect 24386 53705 24758 53781
rect 24386 53580 24479 53646
rect 24386 53564 24463 53580
tri 24463 53564 24479 53580 nw
rect 24515 53547 24629 53705
rect 24665 53580 24758 53646
tri 24665 53564 24681 53580 ne
rect 24681 53564 24758 53580
rect 24498 53465 24646 53547
rect 24386 53432 24463 53448
tri 24463 53432 24479 53448 sw
rect 24386 53366 24479 53432
rect 24386 53264 24479 53330
rect 24386 53248 24463 53264
tri 24463 53248 24479 53264 nw
rect 24515 53231 24629 53465
tri 24665 53432 24681 53448 se
rect 24681 53432 24758 53448
rect 24665 53366 24758 53432
rect 24665 53264 24758 53330
tri 24665 53248 24681 53264 ne
rect 24681 53248 24758 53264
rect 24498 53149 24646 53231
rect 24386 53116 24463 53132
tri 24463 53116 24479 53132 sw
rect 24386 53050 24479 53116
rect 24515 52991 24629 53149
tri 24665 53116 24681 53132 se
rect 24681 53116 24758 53132
rect 24665 53050 24758 53116
rect 24386 52915 24758 52991
rect 24386 52790 24479 52856
rect 24386 52774 24463 52790
tri 24463 52774 24479 52790 nw
rect 24515 52757 24629 52915
rect 24665 52790 24758 52856
tri 24665 52774 24681 52790 ne
rect 24681 52774 24758 52790
rect 24498 52675 24646 52757
rect 24386 52642 24463 52658
tri 24463 52642 24479 52658 sw
rect 24386 52576 24479 52642
rect 24386 52474 24479 52540
rect 24386 52458 24463 52474
tri 24463 52458 24479 52474 nw
rect 24515 52441 24629 52675
tri 24665 52642 24681 52658 se
rect 24681 52642 24758 52658
rect 24665 52576 24758 52642
rect 24665 52474 24758 52540
tri 24665 52458 24681 52474 ne
rect 24681 52458 24758 52474
rect 24498 52359 24646 52441
rect 24386 52326 24463 52342
tri 24463 52326 24479 52342 sw
rect 24386 52260 24479 52326
rect 24515 52201 24629 52359
tri 24665 52326 24681 52342 se
rect 24681 52326 24758 52342
rect 24665 52260 24758 52326
rect 24386 52125 24758 52201
rect 24386 52000 24479 52066
rect 24386 51984 24463 52000
tri 24463 51984 24479 52000 nw
rect 24515 51967 24629 52125
rect 24665 52000 24758 52066
tri 24665 51984 24681 52000 ne
rect 24681 51984 24758 52000
rect 24498 51885 24646 51967
rect 24386 51852 24463 51868
tri 24463 51852 24479 51868 sw
rect 24386 51786 24479 51852
rect 24386 51684 24479 51750
rect 24386 51668 24463 51684
tri 24463 51668 24479 51684 nw
rect 24515 51651 24629 51885
tri 24665 51852 24681 51868 se
rect 24681 51852 24758 51868
rect 24665 51786 24758 51852
rect 24665 51684 24758 51750
tri 24665 51668 24681 51684 ne
rect 24681 51668 24758 51684
rect 24498 51569 24646 51651
rect 24386 51536 24463 51552
tri 24463 51536 24479 51552 sw
rect 24386 51470 24479 51536
rect 24515 51411 24629 51569
tri 24665 51536 24681 51552 se
rect 24681 51536 24758 51552
rect 24665 51470 24758 51536
rect 24386 51335 24758 51411
rect 24386 51210 24479 51276
rect 24386 51194 24463 51210
tri 24463 51194 24479 51210 nw
rect 24515 51177 24629 51335
rect 24665 51210 24758 51276
tri 24665 51194 24681 51210 ne
rect 24681 51194 24758 51210
rect 24498 51095 24646 51177
rect 24386 51062 24463 51078
tri 24463 51062 24479 51078 sw
rect 24386 50996 24479 51062
rect 24386 50894 24479 50960
rect 24386 50878 24463 50894
tri 24463 50878 24479 50894 nw
rect 24515 50861 24629 51095
tri 24665 51062 24681 51078 se
rect 24681 51062 24758 51078
rect 24665 50996 24758 51062
rect 24665 50894 24758 50960
tri 24665 50878 24681 50894 ne
rect 24681 50878 24758 50894
rect 24498 50779 24646 50861
rect 24386 50746 24463 50762
tri 24463 50746 24479 50762 sw
rect 24386 50680 24479 50746
rect 24515 50621 24629 50779
tri 24665 50746 24681 50762 se
rect 24681 50746 24758 50762
rect 24665 50680 24758 50746
rect 24386 50545 24758 50621
rect 24386 50420 24479 50486
rect 24386 50404 24463 50420
tri 24463 50404 24479 50420 nw
rect 24515 50387 24629 50545
rect 24665 50420 24758 50486
tri 24665 50404 24681 50420 ne
rect 24681 50404 24758 50420
rect 24498 50305 24646 50387
rect 24386 50272 24463 50288
tri 24463 50272 24479 50288 sw
rect 24386 50206 24479 50272
rect 24386 50104 24479 50170
rect 24386 50088 24463 50104
tri 24463 50088 24479 50104 nw
rect 24515 50071 24629 50305
tri 24665 50272 24681 50288 se
rect 24681 50272 24758 50288
rect 24665 50206 24758 50272
rect 24665 50104 24758 50170
tri 24665 50088 24681 50104 ne
rect 24681 50088 24758 50104
rect 24498 49989 24646 50071
rect 24386 49956 24463 49972
tri 24463 49956 24479 49972 sw
rect 24386 49890 24479 49956
rect 24515 49831 24629 49989
tri 24665 49956 24681 49972 se
rect 24681 49956 24758 49972
rect 24665 49890 24758 49956
rect 24386 49755 24758 49831
rect 24386 49630 24479 49696
rect 24386 49614 24463 49630
tri 24463 49614 24479 49630 nw
rect 24515 49597 24629 49755
rect 24665 49630 24758 49696
tri 24665 49614 24681 49630 ne
rect 24681 49614 24758 49630
rect 24498 49515 24646 49597
rect 24386 49482 24463 49498
tri 24463 49482 24479 49498 sw
rect 24386 49416 24479 49482
rect 24386 49314 24479 49380
rect 24386 49298 24463 49314
tri 24463 49298 24479 49314 nw
rect 24515 49281 24629 49515
tri 24665 49482 24681 49498 se
rect 24681 49482 24758 49498
rect 24665 49416 24758 49482
rect 24665 49314 24758 49380
tri 24665 49298 24681 49314 ne
rect 24681 49298 24758 49314
rect 24498 49199 24646 49281
rect 24386 49166 24463 49182
tri 24463 49166 24479 49182 sw
rect 24386 49100 24479 49166
rect 24515 49041 24629 49199
tri 24665 49166 24681 49182 se
rect 24681 49166 24758 49182
rect 24665 49100 24758 49166
rect 24386 48965 24758 49041
rect 24386 48840 24479 48906
rect 24386 48824 24463 48840
tri 24463 48824 24479 48840 nw
rect 24515 48807 24629 48965
rect 24665 48840 24758 48906
tri 24665 48824 24681 48840 ne
rect 24681 48824 24758 48840
rect 24498 48725 24646 48807
rect 24386 48692 24463 48708
tri 24463 48692 24479 48708 sw
rect 24386 48626 24479 48692
rect 24386 48524 24479 48590
rect 24386 48508 24463 48524
tri 24463 48508 24479 48524 nw
rect 24515 48491 24629 48725
tri 24665 48692 24681 48708 se
rect 24681 48692 24758 48708
rect 24665 48626 24758 48692
rect 24665 48524 24758 48590
tri 24665 48508 24681 48524 ne
rect 24681 48508 24758 48524
rect 24498 48409 24646 48491
rect 24386 48376 24463 48392
tri 24463 48376 24479 48392 sw
rect 24386 48310 24479 48376
rect 24515 48251 24629 48409
tri 24665 48376 24681 48392 se
rect 24681 48376 24758 48392
rect 24665 48310 24758 48376
rect 24386 48175 24758 48251
rect 24386 48050 24479 48116
rect 24386 48034 24463 48050
tri 24463 48034 24479 48050 nw
rect 24515 48017 24629 48175
rect 24665 48050 24758 48116
tri 24665 48034 24681 48050 ne
rect 24681 48034 24758 48050
rect 24498 47935 24646 48017
rect 24386 47902 24463 47918
tri 24463 47902 24479 47918 sw
rect 24386 47836 24479 47902
rect 24386 47734 24479 47800
rect 24386 47718 24463 47734
tri 24463 47718 24479 47734 nw
rect 24515 47701 24629 47935
tri 24665 47902 24681 47918 se
rect 24681 47902 24758 47918
rect 24665 47836 24758 47902
rect 24665 47734 24758 47800
tri 24665 47718 24681 47734 ne
rect 24681 47718 24758 47734
rect 24498 47619 24646 47701
rect 24386 47586 24463 47602
tri 24463 47586 24479 47602 sw
rect 24386 47520 24479 47586
rect 24515 47461 24629 47619
tri 24665 47586 24681 47602 se
rect 24681 47586 24758 47602
rect 24665 47520 24758 47586
rect 24386 47385 24758 47461
rect 24386 47260 24479 47326
rect 24386 47244 24463 47260
tri 24463 47244 24479 47260 nw
rect 24515 47227 24629 47385
rect 24665 47260 24758 47326
tri 24665 47244 24681 47260 ne
rect 24681 47244 24758 47260
rect 24498 47145 24646 47227
rect 24386 47112 24463 47128
tri 24463 47112 24479 47128 sw
rect 24386 47046 24479 47112
rect 24386 46944 24479 47010
rect 24386 46928 24463 46944
tri 24463 46928 24479 46944 nw
rect 24515 46911 24629 47145
tri 24665 47112 24681 47128 se
rect 24681 47112 24758 47128
rect 24665 47046 24758 47112
rect 24665 46944 24758 47010
tri 24665 46928 24681 46944 ne
rect 24681 46928 24758 46944
rect 24498 46829 24646 46911
rect 24386 46796 24463 46812
tri 24463 46796 24479 46812 sw
rect 24386 46730 24479 46796
rect 24515 46671 24629 46829
tri 24665 46796 24681 46812 se
rect 24681 46796 24758 46812
rect 24665 46730 24758 46796
rect 24386 46595 24758 46671
rect 24386 46470 24479 46536
rect 24386 46454 24463 46470
tri 24463 46454 24479 46470 nw
rect 24515 46437 24629 46595
rect 24665 46470 24758 46536
tri 24665 46454 24681 46470 ne
rect 24681 46454 24758 46470
rect 24498 46355 24646 46437
rect 24386 46322 24463 46338
tri 24463 46322 24479 46338 sw
rect 24386 46256 24479 46322
rect 24386 46154 24479 46220
rect 24386 46138 24463 46154
tri 24463 46138 24479 46154 nw
rect 24515 46121 24629 46355
tri 24665 46322 24681 46338 se
rect 24681 46322 24758 46338
rect 24665 46256 24758 46322
rect 24665 46154 24758 46220
tri 24665 46138 24681 46154 ne
rect 24681 46138 24758 46154
rect 24498 46039 24646 46121
rect 24386 46006 24463 46022
tri 24463 46006 24479 46022 sw
rect 24386 45940 24479 46006
rect 24515 45881 24629 46039
tri 24665 46006 24681 46022 se
rect 24681 46006 24758 46022
rect 24665 45940 24758 46006
rect 24386 45805 24758 45881
rect 24386 45680 24479 45746
rect 24386 45664 24463 45680
tri 24463 45664 24479 45680 nw
rect 24515 45647 24629 45805
rect 24665 45680 24758 45746
tri 24665 45664 24681 45680 ne
rect 24681 45664 24758 45680
rect 24498 45565 24646 45647
rect 24386 45532 24463 45548
tri 24463 45532 24479 45548 sw
rect 24386 45466 24479 45532
rect 24386 45364 24479 45430
rect 24386 45348 24463 45364
tri 24463 45348 24479 45364 nw
rect 24515 45331 24629 45565
tri 24665 45532 24681 45548 se
rect 24681 45532 24758 45548
rect 24665 45466 24758 45532
rect 24665 45364 24758 45430
tri 24665 45348 24681 45364 ne
rect 24681 45348 24758 45364
rect 24498 45249 24646 45331
rect 24386 45216 24463 45232
tri 24463 45216 24479 45232 sw
rect 24386 45150 24479 45216
rect 24515 45091 24629 45249
tri 24665 45216 24681 45232 se
rect 24681 45216 24758 45232
rect 24665 45150 24758 45216
rect 24386 45015 24758 45091
rect 24386 44890 24479 44956
rect 24386 44874 24463 44890
tri 24463 44874 24479 44890 nw
rect 24515 44857 24629 45015
rect 24665 44890 24758 44956
tri 24665 44874 24681 44890 ne
rect 24681 44874 24758 44890
rect 24498 44775 24646 44857
rect 24386 44742 24463 44758
tri 24463 44742 24479 44758 sw
rect 24386 44676 24479 44742
rect 24386 44574 24479 44640
rect 24386 44558 24463 44574
tri 24463 44558 24479 44574 nw
rect 24515 44541 24629 44775
tri 24665 44742 24681 44758 se
rect 24681 44742 24758 44758
rect 24665 44676 24758 44742
rect 24665 44574 24758 44640
tri 24665 44558 24681 44574 ne
rect 24681 44558 24758 44574
rect 24498 44459 24646 44541
rect 24386 44426 24463 44442
tri 24463 44426 24479 44442 sw
rect 24386 44360 24479 44426
rect 24515 44301 24629 44459
tri 24665 44426 24681 44442 se
rect 24681 44426 24758 44442
rect 24665 44360 24758 44426
rect 24386 44225 24758 44301
rect 24386 44100 24479 44166
rect 24386 44084 24463 44100
tri 24463 44084 24479 44100 nw
rect 24515 44067 24629 44225
rect 24665 44100 24758 44166
tri 24665 44084 24681 44100 ne
rect 24681 44084 24758 44100
rect 24498 43985 24646 44067
rect 24386 43952 24463 43968
tri 24463 43952 24479 43968 sw
rect 24386 43886 24479 43952
rect 24386 43784 24479 43850
rect 24386 43768 24463 43784
tri 24463 43768 24479 43784 nw
rect 24515 43751 24629 43985
tri 24665 43952 24681 43968 se
rect 24681 43952 24758 43968
rect 24665 43886 24758 43952
rect 24665 43784 24758 43850
tri 24665 43768 24681 43784 ne
rect 24681 43768 24758 43784
rect 24498 43669 24646 43751
rect 24386 43636 24463 43652
tri 24463 43636 24479 43652 sw
rect 24386 43570 24479 43636
rect 24515 43511 24629 43669
tri 24665 43636 24681 43652 se
rect 24681 43636 24758 43652
rect 24665 43570 24758 43636
rect 24386 43435 24758 43511
rect 24386 43310 24479 43376
rect 24386 43294 24463 43310
tri 24463 43294 24479 43310 nw
rect 24515 43277 24629 43435
rect 24665 43310 24758 43376
tri 24665 43294 24681 43310 ne
rect 24681 43294 24758 43310
rect 24498 43195 24646 43277
rect 24386 43162 24463 43178
tri 24463 43162 24479 43178 sw
rect 24386 43096 24479 43162
rect 24386 42994 24479 43060
rect 24386 42978 24463 42994
tri 24463 42978 24479 42994 nw
rect 24515 42961 24629 43195
tri 24665 43162 24681 43178 se
rect 24681 43162 24758 43178
rect 24665 43096 24758 43162
rect 24665 42994 24758 43060
tri 24665 42978 24681 42994 ne
rect 24681 42978 24758 42994
rect 24498 42879 24646 42961
rect 24386 42846 24463 42862
tri 24463 42846 24479 42862 sw
rect 24386 42780 24479 42846
rect 24515 42721 24629 42879
tri 24665 42846 24681 42862 se
rect 24681 42846 24758 42862
rect 24665 42780 24758 42846
rect 24386 42645 24758 42721
rect 24386 42520 24479 42586
rect 24386 42504 24463 42520
tri 24463 42504 24479 42520 nw
rect 24515 42487 24629 42645
rect 24665 42520 24758 42586
tri 24665 42504 24681 42520 ne
rect 24681 42504 24758 42520
rect 24498 42405 24646 42487
rect 24386 42372 24463 42388
tri 24463 42372 24479 42388 sw
rect 24386 42306 24479 42372
rect 24386 42204 24479 42270
rect 24386 42188 24463 42204
tri 24463 42188 24479 42204 nw
rect 24515 42171 24629 42405
tri 24665 42372 24681 42388 se
rect 24681 42372 24758 42388
rect 24665 42306 24758 42372
rect 24665 42204 24758 42270
tri 24665 42188 24681 42204 ne
rect 24681 42188 24758 42204
rect 24498 42089 24646 42171
rect 24386 42056 24463 42072
tri 24463 42056 24479 42072 sw
rect 24386 41990 24479 42056
rect 24515 41931 24629 42089
tri 24665 42056 24681 42072 se
rect 24681 42056 24758 42072
rect 24665 41990 24758 42056
rect 24386 41855 24758 41931
rect 24386 41730 24479 41796
rect 24386 41714 24463 41730
tri 24463 41714 24479 41730 nw
rect 24515 41697 24629 41855
rect 24665 41730 24758 41796
tri 24665 41714 24681 41730 ne
rect 24681 41714 24758 41730
rect 24498 41615 24646 41697
rect 24386 41582 24463 41598
tri 24463 41582 24479 41598 sw
rect 24386 41516 24479 41582
rect 24386 41414 24479 41480
rect 24386 41398 24463 41414
tri 24463 41398 24479 41414 nw
rect 24515 41381 24629 41615
tri 24665 41582 24681 41598 se
rect 24681 41582 24758 41598
rect 24665 41516 24758 41582
rect 24665 41414 24758 41480
tri 24665 41398 24681 41414 ne
rect 24681 41398 24758 41414
rect 24498 41299 24646 41381
rect 24386 41266 24463 41282
tri 24463 41266 24479 41282 sw
rect 24386 41200 24479 41266
rect 24515 41141 24629 41299
tri 24665 41266 24681 41282 se
rect 24681 41266 24758 41282
rect 24665 41200 24758 41266
rect 24386 41065 24758 41141
rect 24386 40940 24479 41006
rect 24386 40924 24463 40940
tri 24463 40924 24479 40940 nw
rect 24515 40907 24629 41065
rect 24665 40940 24758 41006
tri 24665 40924 24681 40940 ne
rect 24681 40924 24758 40940
rect 24498 40825 24646 40907
rect 24386 40792 24463 40808
tri 24463 40792 24479 40808 sw
rect 24386 40726 24479 40792
rect 24386 40624 24479 40690
rect 24386 40608 24463 40624
tri 24463 40608 24479 40624 nw
rect 24515 40591 24629 40825
tri 24665 40792 24681 40808 se
rect 24681 40792 24758 40808
rect 24665 40726 24758 40792
rect 24665 40624 24758 40690
tri 24665 40608 24681 40624 ne
rect 24681 40608 24758 40624
rect 24498 40509 24646 40591
rect 24386 40476 24463 40492
tri 24463 40476 24479 40492 sw
rect 24386 40410 24479 40476
rect 24515 40351 24629 40509
tri 24665 40476 24681 40492 se
rect 24681 40476 24758 40492
rect 24665 40410 24758 40476
rect 24386 40275 24758 40351
rect 24386 40150 24479 40216
rect 24386 40134 24463 40150
tri 24463 40134 24479 40150 nw
rect 24515 40117 24629 40275
rect 24665 40150 24758 40216
tri 24665 40134 24681 40150 ne
rect 24681 40134 24758 40150
rect 24498 40035 24646 40117
rect 24386 40002 24463 40018
tri 24463 40002 24479 40018 sw
rect 24386 39936 24479 40002
rect 24386 39834 24479 39900
rect 24386 39818 24463 39834
tri 24463 39818 24479 39834 nw
rect 24515 39801 24629 40035
tri 24665 40002 24681 40018 se
rect 24681 40002 24758 40018
rect 24665 39936 24758 40002
rect 24665 39834 24758 39900
tri 24665 39818 24681 39834 ne
rect 24681 39818 24758 39834
rect 24498 39719 24646 39801
rect 24386 39686 24463 39702
tri 24463 39686 24479 39702 sw
rect 24386 39620 24479 39686
rect 24515 39561 24629 39719
tri 24665 39686 24681 39702 se
rect 24681 39686 24758 39702
rect 24665 39620 24758 39686
rect 24386 39485 24758 39561
rect 24386 39360 24479 39426
rect 24386 39344 24463 39360
tri 24463 39344 24479 39360 nw
rect 24515 39327 24629 39485
rect 24665 39360 24758 39426
tri 24665 39344 24681 39360 ne
rect 24681 39344 24758 39360
rect 24498 39245 24646 39327
rect 24386 39212 24463 39228
tri 24463 39212 24479 39228 sw
rect 24386 39146 24479 39212
rect 24386 39044 24479 39110
rect 24386 39028 24463 39044
tri 24463 39028 24479 39044 nw
rect 24515 39011 24629 39245
tri 24665 39212 24681 39228 se
rect 24681 39212 24758 39228
rect 24665 39146 24758 39212
rect 24665 39044 24758 39110
tri 24665 39028 24681 39044 ne
rect 24681 39028 24758 39044
rect 24498 38929 24646 39011
rect 24386 38896 24463 38912
tri 24463 38896 24479 38912 sw
rect 24386 38830 24479 38896
rect 24515 38771 24629 38929
tri 24665 38896 24681 38912 se
rect 24681 38896 24758 38912
rect 24665 38830 24758 38896
rect 24386 38695 24758 38771
rect 24386 38570 24479 38636
rect 24386 38554 24463 38570
tri 24463 38554 24479 38570 nw
rect 24515 38537 24629 38695
rect 24665 38570 24758 38636
tri 24665 38554 24681 38570 ne
rect 24681 38554 24758 38570
rect 24498 38455 24646 38537
rect 24386 38422 24463 38438
tri 24463 38422 24479 38438 sw
rect 24386 38356 24479 38422
rect 24386 38254 24479 38320
rect 24386 38238 24463 38254
tri 24463 38238 24479 38254 nw
rect 24515 38221 24629 38455
tri 24665 38422 24681 38438 se
rect 24681 38422 24758 38438
rect 24665 38356 24758 38422
rect 24665 38254 24758 38320
tri 24665 38238 24681 38254 ne
rect 24681 38238 24758 38254
rect 24498 38139 24646 38221
rect 24386 38106 24463 38122
tri 24463 38106 24479 38122 sw
rect 24386 38040 24479 38106
rect 24515 37981 24629 38139
tri 24665 38106 24681 38122 se
rect 24681 38106 24758 38122
rect 24665 38040 24758 38106
rect 24386 37905 24758 37981
rect 24386 37780 24479 37846
rect 24386 37764 24463 37780
tri 24463 37764 24479 37780 nw
rect 24515 37747 24629 37905
rect 24665 37780 24758 37846
tri 24665 37764 24681 37780 ne
rect 24681 37764 24758 37780
rect 24498 37665 24646 37747
rect 24386 37632 24463 37648
tri 24463 37632 24479 37648 sw
rect 24386 37566 24479 37632
rect 24386 37464 24479 37530
rect 24386 37448 24463 37464
tri 24463 37448 24479 37464 nw
rect 24515 37431 24629 37665
tri 24665 37632 24681 37648 se
rect 24681 37632 24758 37648
rect 24665 37566 24758 37632
rect 24665 37464 24758 37530
tri 24665 37448 24681 37464 ne
rect 24681 37448 24758 37464
rect 24498 37349 24646 37431
rect 24386 37316 24463 37332
tri 24463 37316 24479 37332 sw
rect 24386 37250 24479 37316
rect 24515 37191 24629 37349
tri 24665 37316 24681 37332 se
rect 24681 37316 24758 37332
rect 24665 37250 24758 37316
rect 24386 37115 24758 37191
rect 24386 36990 24479 37056
rect 24386 36974 24463 36990
tri 24463 36974 24479 36990 nw
rect 24515 36957 24629 37115
rect 24665 36990 24758 37056
tri 24665 36974 24681 36990 ne
rect 24681 36974 24758 36990
rect 24498 36875 24646 36957
rect 24386 36842 24463 36858
tri 24463 36842 24479 36858 sw
rect 24386 36776 24479 36842
rect 24386 36674 24479 36740
rect 24386 36658 24463 36674
tri 24463 36658 24479 36674 nw
rect 24515 36641 24629 36875
tri 24665 36842 24681 36858 se
rect 24681 36842 24758 36858
rect 24665 36776 24758 36842
rect 24665 36674 24758 36740
tri 24665 36658 24681 36674 ne
rect 24681 36658 24758 36674
rect 24498 36559 24646 36641
rect 24386 36526 24463 36542
tri 24463 36526 24479 36542 sw
rect 24386 36460 24479 36526
rect 24515 36401 24629 36559
tri 24665 36526 24681 36542 se
rect 24681 36526 24758 36542
rect 24665 36460 24758 36526
rect 24386 36325 24758 36401
rect 24386 36200 24479 36266
rect 24386 36184 24463 36200
tri 24463 36184 24479 36200 nw
rect 24515 36167 24629 36325
rect 24665 36200 24758 36266
tri 24665 36184 24681 36200 ne
rect 24681 36184 24758 36200
rect 24498 36085 24646 36167
rect 24386 36052 24463 36068
tri 24463 36052 24479 36068 sw
rect 24386 35986 24479 36052
rect 24386 35884 24479 35950
rect 24386 35868 24463 35884
tri 24463 35868 24479 35884 nw
rect 24515 35851 24629 36085
tri 24665 36052 24681 36068 se
rect 24681 36052 24758 36068
rect 24665 35986 24758 36052
rect 24665 35884 24758 35950
tri 24665 35868 24681 35884 ne
rect 24681 35868 24758 35884
rect 24498 35769 24646 35851
rect 24386 35736 24463 35752
tri 24463 35736 24479 35752 sw
rect 24386 35670 24479 35736
rect 24515 35611 24629 35769
tri 24665 35736 24681 35752 se
rect 24681 35736 24758 35752
rect 24665 35670 24758 35736
rect 24386 35535 24758 35611
rect 24386 35410 24479 35476
rect 24386 35394 24463 35410
tri 24463 35394 24479 35410 nw
rect 24515 35377 24629 35535
rect 24665 35410 24758 35476
tri 24665 35394 24681 35410 ne
rect 24681 35394 24758 35410
rect 24498 35295 24646 35377
rect 24386 35262 24463 35278
tri 24463 35262 24479 35278 sw
rect 24386 35196 24479 35262
rect 24386 35094 24479 35160
rect 24386 35078 24463 35094
tri 24463 35078 24479 35094 nw
rect 24515 35061 24629 35295
tri 24665 35262 24681 35278 se
rect 24681 35262 24758 35278
rect 24665 35196 24758 35262
rect 24665 35094 24758 35160
tri 24665 35078 24681 35094 ne
rect 24681 35078 24758 35094
rect 24498 34979 24646 35061
rect 24386 34946 24463 34962
tri 24463 34946 24479 34962 sw
rect 24386 34880 24479 34946
rect 24515 34821 24629 34979
tri 24665 34946 24681 34962 se
rect 24681 34946 24758 34962
rect 24665 34880 24758 34946
rect 24386 34745 24758 34821
rect 24386 34620 24479 34686
rect 24386 34604 24463 34620
tri 24463 34604 24479 34620 nw
rect 24515 34587 24629 34745
rect 24665 34620 24758 34686
tri 24665 34604 24681 34620 ne
rect 24681 34604 24758 34620
rect 24498 34505 24646 34587
rect 24386 34472 24463 34488
tri 24463 34472 24479 34488 sw
rect 24386 34406 24479 34472
rect 24386 34304 24479 34370
rect 24386 34288 24463 34304
tri 24463 34288 24479 34304 nw
rect 24515 34271 24629 34505
tri 24665 34472 24681 34488 se
rect 24681 34472 24758 34488
rect 24665 34406 24758 34472
rect 24665 34304 24758 34370
tri 24665 34288 24681 34304 ne
rect 24681 34288 24758 34304
rect 24498 34189 24646 34271
rect 24386 34156 24463 34172
tri 24463 34156 24479 34172 sw
rect 24386 34090 24479 34156
rect 24515 34031 24629 34189
tri 24665 34156 24681 34172 se
rect 24681 34156 24758 34172
rect 24665 34090 24758 34156
rect 24386 33955 24758 34031
rect 24386 33830 24479 33896
rect 24386 33814 24463 33830
tri 24463 33814 24479 33830 nw
rect 24515 33797 24629 33955
rect 24665 33830 24758 33896
tri 24665 33814 24681 33830 ne
rect 24681 33814 24758 33830
rect 24498 33715 24646 33797
rect 24386 33682 24463 33698
tri 24463 33682 24479 33698 sw
rect 24386 33616 24479 33682
rect 24386 33514 24479 33580
rect 24386 33498 24463 33514
tri 24463 33498 24479 33514 nw
rect 24515 33481 24629 33715
tri 24665 33682 24681 33698 se
rect 24681 33682 24758 33698
rect 24665 33616 24758 33682
rect 24665 33514 24758 33580
tri 24665 33498 24681 33514 ne
rect 24681 33498 24758 33514
rect 24498 33399 24646 33481
rect 24386 33366 24463 33382
tri 24463 33366 24479 33382 sw
rect 24386 33300 24479 33366
rect 24515 33241 24629 33399
tri 24665 33366 24681 33382 se
rect 24681 33366 24758 33382
rect 24665 33300 24758 33366
rect 24386 33165 24758 33241
rect 24386 33040 24479 33106
rect 24386 33024 24463 33040
tri 24463 33024 24479 33040 nw
rect 24515 33007 24629 33165
rect 24665 33040 24758 33106
tri 24665 33024 24681 33040 ne
rect 24681 33024 24758 33040
rect 24498 32925 24646 33007
rect 24386 32892 24463 32908
tri 24463 32892 24479 32908 sw
rect 24386 32826 24479 32892
rect 24386 32724 24479 32790
rect 24386 32708 24463 32724
tri 24463 32708 24479 32724 nw
rect 24515 32691 24629 32925
tri 24665 32892 24681 32908 se
rect 24681 32892 24758 32908
rect 24665 32826 24758 32892
rect 24665 32724 24758 32790
tri 24665 32708 24681 32724 ne
rect 24681 32708 24758 32724
rect 24498 32609 24646 32691
rect 24386 32576 24463 32592
tri 24463 32576 24479 32592 sw
rect 24386 32510 24479 32576
rect 24515 32451 24629 32609
tri 24665 32576 24681 32592 se
rect 24681 32576 24758 32592
rect 24665 32510 24758 32576
rect 24386 32375 24758 32451
rect 24386 32250 24479 32316
rect 24386 32234 24463 32250
tri 24463 32234 24479 32250 nw
rect 24515 32217 24629 32375
rect 24665 32250 24758 32316
tri 24665 32234 24681 32250 ne
rect 24681 32234 24758 32250
rect 24498 32135 24646 32217
rect 24386 32102 24463 32118
tri 24463 32102 24479 32118 sw
rect 24386 32036 24479 32102
rect 24386 31934 24479 32000
rect 24386 31918 24463 31934
tri 24463 31918 24479 31934 nw
rect 24515 31901 24629 32135
tri 24665 32102 24681 32118 se
rect 24681 32102 24758 32118
rect 24665 32036 24758 32102
rect 24665 31934 24758 32000
tri 24665 31918 24681 31934 ne
rect 24681 31918 24758 31934
rect 24498 31819 24646 31901
rect 24386 31786 24463 31802
tri 24463 31786 24479 31802 sw
rect 24386 31720 24479 31786
rect 24515 31661 24629 31819
tri 24665 31786 24681 31802 se
rect 24681 31786 24758 31802
rect 24665 31720 24758 31786
rect 24386 31585 24758 31661
rect 24386 31460 24479 31526
rect 24386 31444 24463 31460
tri 24463 31444 24479 31460 nw
rect 24515 31427 24629 31585
rect 24665 31460 24758 31526
tri 24665 31444 24681 31460 ne
rect 24681 31444 24758 31460
rect 24498 31345 24646 31427
rect 24386 31312 24463 31328
tri 24463 31312 24479 31328 sw
rect 24386 31246 24479 31312
rect 24386 31144 24479 31210
rect 24386 31128 24463 31144
tri 24463 31128 24479 31144 nw
rect 24515 31111 24629 31345
tri 24665 31312 24681 31328 se
rect 24681 31312 24758 31328
rect 24665 31246 24758 31312
rect 24665 31144 24758 31210
tri 24665 31128 24681 31144 ne
rect 24681 31128 24758 31144
rect 24498 31029 24646 31111
rect 24386 30996 24463 31012
tri 24463 30996 24479 31012 sw
rect 24386 30930 24479 30996
rect 24515 30871 24629 31029
tri 24665 30996 24681 31012 se
rect 24681 30996 24758 31012
rect 24665 30930 24758 30996
rect 24386 30795 24758 30871
rect 24386 30670 24479 30736
rect 24386 30654 24463 30670
tri 24463 30654 24479 30670 nw
rect 24515 30637 24629 30795
rect 24665 30670 24758 30736
tri 24665 30654 24681 30670 ne
rect 24681 30654 24758 30670
rect 24498 30555 24646 30637
rect 24386 30522 24463 30538
tri 24463 30522 24479 30538 sw
rect 24386 30456 24479 30522
rect 24386 30354 24479 30420
rect 24386 30338 24463 30354
tri 24463 30338 24479 30354 nw
rect 24515 30321 24629 30555
tri 24665 30522 24681 30538 se
rect 24681 30522 24758 30538
rect 24665 30456 24758 30522
rect 24665 30354 24758 30420
tri 24665 30338 24681 30354 ne
rect 24681 30338 24758 30354
rect 24498 30239 24646 30321
rect 24386 30206 24463 30222
tri 24463 30206 24479 30222 sw
rect 24386 30140 24479 30206
rect 24515 30081 24629 30239
tri 24665 30206 24681 30222 se
rect 24681 30206 24758 30222
rect 24665 30140 24758 30206
rect 24386 30005 24758 30081
rect 24386 29880 24479 29946
rect 24386 29864 24463 29880
tri 24463 29864 24479 29880 nw
rect 24515 29847 24629 30005
rect 24665 29880 24758 29946
tri 24665 29864 24681 29880 ne
rect 24681 29864 24758 29880
rect 24498 29765 24646 29847
rect 24386 29732 24463 29748
tri 24463 29732 24479 29748 sw
rect 24386 29666 24479 29732
rect 24386 29564 24479 29630
rect 24386 29548 24463 29564
tri 24463 29548 24479 29564 nw
rect 24515 29531 24629 29765
tri 24665 29732 24681 29748 se
rect 24681 29732 24758 29748
rect 24665 29666 24758 29732
rect 24665 29564 24758 29630
tri 24665 29548 24681 29564 ne
rect 24681 29548 24758 29564
rect 24498 29449 24646 29531
rect 24386 29416 24463 29432
tri 24463 29416 24479 29432 sw
rect 24386 29350 24479 29416
rect 24515 29291 24629 29449
tri 24665 29416 24681 29432 se
rect 24681 29416 24758 29432
rect 24665 29350 24758 29416
rect 24386 29215 24758 29291
rect 24386 29090 24479 29156
rect 24386 29074 24463 29090
tri 24463 29074 24479 29090 nw
rect 24515 29057 24629 29215
rect 24665 29090 24758 29156
tri 24665 29074 24681 29090 ne
rect 24681 29074 24758 29090
rect 24498 28975 24646 29057
rect 24386 28942 24463 28958
tri 24463 28942 24479 28958 sw
rect 24386 28876 24479 28942
rect 24515 28833 24629 28975
tri 24665 28942 24681 28958 se
rect 24681 28942 24758 28958
rect 24665 28876 24758 28942
rect 24794 28463 24830 80603
rect 24866 28463 24902 80603
rect 24938 80445 24974 80603
rect 24930 80303 24982 80445
rect 24938 28763 24974 80303
rect 24930 28621 24982 28763
rect 24938 28463 24974 28621
rect 25010 28463 25046 80603
rect 25082 28463 25118 80603
rect 25154 28833 25238 80233
rect 25274 28463 25310 80603
rect 25346 28463 25382 80603
rect 25418 80445 25454 80603
rect 25410 80303 25462 80445
rect 25418 28763 25454 80303
rect 25410 28621 25462 28763
rect 25418 28463 25454 28621
rect 25490 28463 25526 80603
rect 25562 28463 25598 80603
rect 25634 80124 25727 80190
rect 25634 80108 25711 80124
tri 25711 80108 25727 80124 nw
rect 25763 80091 25877 80233
rect 25913 80124 26006 80190
tri 25913 80108 25929 80124 ne
rect 25929 80108 26006 80124
rect 25746 80009 25894 80091
rect 25634 79976 25711 79992
tri 25711 79976 25727 79992 sw
rect 25634 79910 25727 79976
rect 25763 79851 25877 80009
tri 25913 79976 25929 79992 se
rect 25929 79976 26006 79992
rect 25913 79910 26006 79976
rect 25634 79775 26006 79851
rect 25634 79650 25727 79716
rect 25634 79634 25711 79650
tri 25711 79634 25727 79650 nw
rect 25763 79617 25877 79775
rect 25913 79650 26006 79716
tri 25913 79634 25929 79650 ne
rect 25929 79634 26006 79650
rect 25746 79535 25894 79617
rect 25634 79502 25711 79518
tri 25711 79502 25727 79518 sw
rect 25634 79436 25727 79502
rect 25634 79334 25727 79400
rect 25634 79318 25711 79334
tri 25711 79318 25727 79334 nw
rect 25763 79301 25877 79535
tri 25913 79502 25929 79518 se
rect 25929 79502 26006 79518
rect 25913 79436 26006 79502
rect 25913 79334 26006 79400
tri 25913 79318 25929 79334 ne
rect 25929 79318 26006 79334
rect 25746 79219 25894 79301
rect 25634 79186 25711 79202
tri 25711 79186 25727 79202 sw
rect 25634 79120 25727 79186
rect 25763 79061 25877 79219
tri 25913 79186 25929 79202 se
rect 25929 79186 26006 79202
rect 25913 79120 26006 79186
rect 25634 78985 26006 79061
rect 25634 78860 25727 78926
rect 25634 78844 25711 78860
tri 25711 78844 25727 78860 nw
rect 25763 78827 25877 78985
rect 25913 78860 26006 78926
tri 25913 78844 25929 78860 ne
rect 25929 78844 26006 78860
rect 25746 78745 25894 78827
rect 25634 78712 25711 78728
tri 25711 78712 25727 78728 sw
rect 25634 78646 25727 78712
rect 25634 78544 25727 78610
rect 25634 78528 25711 78544
tri 25711 78528 25727 78544 nw
rect 25763 78511 25877 78745
tri 25913 78712 25929 78728 se
rect 25929 78712 26006 78728
rect 25913 78646 26006 78712
rect 25913 78544 26006 78610
tri 25913 78528 25929 78544 ne
rect 25929 78528 26006 78544
rect 25746 78429 25894 78511
rect 25634 78396 25711 78412
tri 25711 78396 25727 78412 sw
rect 25634 78330 25727 78396
rect 25763 78271 25877 78429
tri 25913 78396 25929 78412 se
rect 25929 78396 26006 78412
rect 25913 78330 26006 78396
rect 25634 78195 26006 78271
rect 25634 78070 25727 78136
rect 25634 78054 25711 78070
tri 25711 78054 25727 78070 nw
rect 25763 78037 25877 78195
rect 25913 78070 26006 78136
tri 25913 78054 25929 78070 ne
rect 25929 78054 26006 78070
rect 25746 77955 25894 78037
rect 25634 77922 25711 77938
tri 25711 77922 25727 77938 sw
rect 25634 77856 25727 77922
rect 25634 77754 25727 77820
rect 25634 77738 25711 77754
tri 25711 77738 25727 77754 nw
rect 25763 77721 25877 77955
tri 25913 77922 25929 77938 se
rect 25929 77922 26006 77938
rect 25913 77856 26006 77922
rect 25913 77754 26006 77820
tri 25913 77738 25929 77754 ne
rect 25929 77738 26006 77754
rect 25746 77639 25894 77721
rect 25634 77606 25711 77622
tri 25711 77606 25727 77622 sw
rect 25634 77540 25727 77606
rect 25763 77481 25877 77639
tri 25913 77606 25929 77622 se
rect 25929 77606 26006 77622
rect 25913 77540 26006 77606
rect 25634 77405 26006 77481
rect 25634 77280 25727 77346
rect 25634 77264 25711 77280
tri 25711 77264 25727 77280 nw
rect 25763 77247 25877 77405
rect 25913 77280 26006 77346
tri 25913 77264 25929 77280 ne
rect 25929 77264 26006 77280
rect 25746 77165 25894 77247
rect 25634 77132 25711 77148
tri 25711 77132 25727 77148 sw
rect 25634 77066 25727 77132
rect 25634 76964 25727 77030
rect 25634 76948 25711 76964
tri 25711 76948 25727 76964 nw
rect 25763 76931 25877 77165
tri 25913 77132 25929 77148 se
rect 25929 77132 26006 77148
rect 25913 77066 26006 77132
rect 25913 76964 26006 77030
tri 25913 76948 25929 76964 ne
rect 25929 76948 26006 76964
rect 25746 76849 25894 76931
rect 25634 76816 25711 76832
tri 25711 76816 25727 76832 sw
rect 25634 76750 25727 76816
rect 25763 76691 25877 76849
tri 25913 76816 25929 76832 se
rect 25929 76816 26006 76832
rect 25913 76750 26006 76816
rect 25634 76615 26006 76691
rect 25634 76490 25727 76556
rect 25634 76474 25711 76490
tri 25711 76474 25727 76490 nw
rect 25763 76457 25877 76615
rect 25913 76490 26006 76556
tri 25913 76474 25929 76490 ne
rect 25929 76474 26006 76490
rect 25746 76375 25894 76457
rect 25634 76342 25711 76358
tri 25711 76342 25727 76358 sw
rect 25634 76276 25727 76342
rect 25634 76174 25727 76240
rect 25634 76158 25711 76174
tri 25711 76158 25727 76174 nw
rect 25763 76141 25877 76375
tri 25913 76342 25929 76358 se
rect 25929 76342 26006 76358
rect 25913 76276 26006 76342
rect 25913 76174 26006 76240
tri 25913 76158 25929 76174 ne
rect 25929 76158 26006 76174
rect 25746 76059 25894 76141
rect 25634 76026 25711 76042
tri 25711 76026 25727 76042 sw
rect 25634 75960 25727 76026
rect 25763 75901 25877 76059
tri 25913 76026 25929 76042 se
rect 25929 76026 26006 76042
rect 25913 75960 26006 76026
rect 25634 75825 26006 75901
rect 25634 75700 25727 75766
rect 25634 75684 25711 75700
tri 25711 75684 25727 75700 nw
rect 25763 75667 25877 75825
rect 25913 75700 26006 75766
tri 25913 75684 25929 75700 ne
rect 25929 75684 26006 75700
rect 25746 75585 25894 75667
rect 25634 75552 25711 75568
tri 25711 75552 25727 75568 sw
rect 25634 75486 25727 75552
rect 25634 75384 25727 75450
rect 25634 75368 25711 75384
tri 25711 75368 25727 75384 nw
rect 25763 75351 25877 75585
tri 25913 75552 25929 75568 se
rect 25929 75552 26006 75568
rect 25913 75486 26006 75552
rect 25913 75384 26006 75450
tri 25913 75368 25929 75384 ne
rect 25929 75368 26006 75384
rect 25746 75269 25894 75351
rect 25634 75236 25711 75252
tri 25711 75236 25727 75252 sw
rect 25634 75170 25727 75236
rect 25763 75111 25877 75269
tri 25913 75236 25929 75252 se
rect 25929 75236 26006 75252
rect 25913 75170 26006 75236
rect 25634 75035 26006 75111
rect 25634 74910 25727 74976
rect 25634 74894 25711 74910
tri 25711 74894 25727 74910 nw
rect 25763 74877 25877 75035
rect 25913 74910 26006 74976
tri 25913 74894 25929 74910 ne
rect 25929 74894 26006 74910
rect 25746 74795 25894 74877
rect 25634 74762 25711 74778
tri 25711 74762 25727 74778 sw
rect 25634 74696 25727 74762
rect 25634 74594 25727 74660
rect 25634 74578 25711 74594
tri 25711 74578 25727 74594 nw
rect 25763 74561 25877 74795
tri 25913 74762 25929 74778 se
rect 25929 74762 26006 74778
rect 25913 74696 26006 74762
rect 25913 74594 26006 74660
tri 25913 74578 25929 74594 ne
rect 25929 74578 26006 74594
rect 25746 74479 25894 74561
rect 25634 74446 25711 74462
tri 25711 74446 25727 74462 sw
rect 25634 74380 25727 74446
rect 25763 74321 25877 74479
tri 25913 74446 25929 74462 se
rect 25929 74446 26006 74462
rect 25913 74380 26006 74446
rect 25634 74245 26006 74321
rect 25634 74120 25727 74186
rect 25634 74104 25711 74120
tri 25711 74104 25727 74120 nw
rect 25763 74087 25877 74245
rect 25913 74120 26006 74186
tri 25913 74104 25929 74120 ne
rect 25929 74104 26006 74120
rect 25746 74005 25894 74087
rect 25634 73972 25711 73988
tri 25711 73972 25727 73988 sw
rect 25634 73906 25727 73972
rect 25634 73804 25727 73870
rect 25634 73788 25711 73804
tri 25711 73788 25727 73804 nw
rect 25763 73771 25877 74005
tri 25913 73972 25929 73988 se
rect 25929 73972 26006 73988
rect 25913 73906 26006 73972
rect 25913 73804 26006 73870
tri 25913 73788 25929 73804 ne
rect 25929 73788 26006 73804
rect 25746 73689 25894 73771
rect 25634 73656 25711 73672
tri 25711 73656 25727 73672 sw
rect 25634 73590 25727 73656
rect 25763 73531 25877 73689
tri 25913 73656 25929 73672 se
rect 25929 73656 26006 73672
rect 25913 73590 26006 73656
rect 25634 73455 26006 73531
rect 25634 73330 25727 73396
rect 25634 73314 25711 73330
tri 25711 73314 25727 73330 nw
rect 25763 73297 25877 73455
rect 25913 73330 26006 73396
tri 25913 73314 25929 73330 ne
rect 25929 73314 26006 73330
rect 25746 73215 25894 73297
rect 25634 73182 25711 73198
tri 25711 73182 25727 73198 sw
rect 25634 73116 25727 73182
rect 25634 73014 25727 73080
rect 25634 72998 25711 73014
tri 25711 72998 25727 73014 nw
rect 25763 72981 25877 73215
tri 25913 73182 25929 73198 se
rect 25929 73182 26006 73198
rect 25913 73116 26006 73182
rect 25913 73014 26006 73080
tri 25913 72998 25929 73014 ne
rect 25929 72998 26006 73014
rect 25746 72899 25894 72981
rect 25634 72866 25711 72882
tri 25711 72866 25727 72882 sw
rect 25634 72800 25727 72866
rect 25763 72741 25877 72899
tri 25913 72866 25929 72882 se
rect 25929 72866 26006 72882
rect 25913 72800 26006 72866
rect 25634 72665 26006 72741
rect 25634 72540 25727 72606
rect 25634 72524 25711 72540
tri 25711 72524 25727 72540 nw
rect 25763 72507 25877 72665
rect 25913 72540 26006 72606
tri 25913 72524 25929 72540 ne
rect 25929 72524 26006 72540
rect 25746 72425 25894 72507
rect 25634 72392 25711 72408
tri 25711 72392 25727 72408 sw
rect 25634 72326 25727 72392
rect 25634 72224 25727 72290
rect 25634 72208 25711 72224
tri 25711 72208 25727 72224 nw
rect 25763 72191 25877 72425
tri 25913 72392 25929 72408 se
rect 25929 72392 26006 72408
rect 25913 72326 26006 72392
rect 25913 72224 26006 72290
tri 25913 72208 25929 72224 ne
rect 25929 72208 26006 72224
rect 25746 72109 25894 72191
rect 25634 72076 25711 72092
tri 25711 72076 25727 72092 sw
rect 25634 72010 25727 72076
rect 25763 71951 25877 72109
tri 25913 72076 25929 72092 se
rect 25929 72076 26006 72092
rect 25913 72010 26006 72076
rect 25634 71875 26006 71951
rect 25634 71750 25727 71816
rect 25634 71734 25711 71750
tri 25711 71734 25727 71750 nw
rect 25763 71717 25877 71875
rect 25913 71750 26006 71816
tri 25913 71734 25929 71750 ne
rect 25929 71734 26006 71750
rect 25746 71635 25894 71717
rect 25634 71602 25711 71618
tri 25711 71602 25727 71618 sw
rect 25634 71536 25727 71602
rect 25634 71434 25727 71500
rect 25634 71418 25711 71434
tri 25711 71418 25727 71434 nw
rect 25763 71401 25877 71635
tri 25913 71602 25929 71618 se
rect 25929 71602 26006 71618
rect 25913 71536 26006 71602
rect 25913 71434 26006 71500
tri 25913 71418 25929 71434 ne
rect 25929 71418 26006 71434
rect 25746 71319 25894 71401
rect 25634 71286 25711 71302
tri 25711 71286 25727 71302 sw
rect 25634 71220 25727 71286
rect 25763 71161 25877 71319
tri 25913 71286 25929 71302 se
rect 25929 71286 26006 71302
rect 25913 71220 26006 71286
rect 25634 71085 26006 71161
rect 25634 70960 25727 71026
rect 25634 70944 25711 70960
tri 25711 70944 25727 70960 nw
rect 25763 70927 25877 71085
rect 25913 70960 26006 71026
tri 25913 70944 25929 70960 ne
rect 25929 70944 26006 70960
rect 25746 70845 25894 70927
rect 25634 70812 25711 70828
tri 25711 70812 25727 70828 sw
rect 25634 70746 25727 70812
rect 25634 70644 25727 70710
rect 25634 70628 25711 70644
tri 25711 70628 25727 70644 nw
rect 25763 70611 25877 70845
tri 25913 70812 25929 70828 se
rect 25929 70812 26006 70828
rect 25913 70746 26006 70812
rect 25913 70644 26006 70710
tri 25913 70628 25929 70644 ne
rect 25929 70628 26006 70644
rect 25746 70529 25894 70611
rect 25634 70496 25711 70512
tri 25711 70496 25727 70512 sw
rect 25634 70430 25727 70496
rect 25763 70371 25877 70529
tri 25913 70496 25929 70512 se
rect 25929 70496 26006 70512
rect 25913 70430 26006 70496
rect 25634 70295 26006 70371
rect 25634 70170 25727 70236
rect 25634 70154 25711 70170
tri 25711 70154 25727 70170 nw
rect 25763 70137 25877 70295
rect 25913 70170 26006 70236
tri 25913 70154 25929 70170 ne
rect 25929 70154 26006 70170
rect 25746 70055 25894 70137
rect 25634 70022 25711 70038
tri 25711 70022 25727 70038 sw
rect 25634 69956 25727 70022
rect 25634 69854 25727 69920
rect 25634 69838 25711 69854
tri 25711 69838 25727 69854 nw
rect 25763 69821 25877 70055
tri 25913 70022 25929 70038 se
rect 25929 70022 26006 70038
rect 25913 69956 26006 70022
rect 25913 69854 26006 69920
tri 25913 69838 25929 69854 ne
rect 25929 69838 26006 69854
rect 25746 69739 25894 69821
rect 25634 69706 25711 69722
tri 25711 69706 25727 69722 sw
rect 25634 69640 25727 69706
rect 25763 69581 25877 69739
tri 25913 69706 25929 69722 se
rect 25929 69706 26006 69722
rect 25913 69640 26006 69706
rect 25634 69505 26006 69581
rect 25634 69380 25727 69446
rect 25634 69364 25711 69380
tri 25711 69364 25727 69380 nw
rect 25763 69347 25877 69505
rect 25913 69380 26006 69446
tri 25913 69364 25929 69380 ne
rect 25929 69364 26006 69380
rect 25746 69265 25894 69347
rect 25634 69232 25711 69248
tri 25711 69232 25727 69248 sw
rect 25634 69166 25727 69232
rect 25634 69064 25727 69130
rect 25634 69048 25711 69064
tri 25711 69048 25727 69064 nw
rect 25763 69031 25877 69265
tri 25913 69232 25929 69248 se
rect 25929 69232 26006 69248
rect 25913 69166 26006 69232
rect 25913 69064 26006 69130
tri 25913 69048 25929 69064 ne
rect 25929 69048 26006 69064
rect 25746 68949 25894 69031
rect 25634 68916 25711 68932
tri 25711 68916 25727 68932 sw
rect 25634 68850 25727 68916
rect 25763 68791 25877 68949
tri 25913 68916 25929 68932 se
rect 25929 68916 26006 68932
rect 25913 68850 26006 68916
rect 25634 68715 26006 68791
rect 25634 68590 25727 68656
rect 25634 68574 25711 68590
tri 25711 68574 25727 68590 nw
rect 25763 68557 25877 68715
rect 25913 68590 26006 68656
tri 25913 68574 25929 68590 ne
rect 25929 68574 26006 68590
rect 25746 68475 25894 68557
rect 25634 68442 25711 68458
tri 25711 68442 25727 68458 sw
rect 25634 68376 25727 68442
rect 25634 68274 25727 68340
rect 25634 68258 25711 68274
tri 25711 68258 25727 68274 nw
rect 25763 68241 25877 68475
tri 25913 68442 25929 68458 se
rect 25929 68442 26006 68458
rect 25913 68376 26006 68442
rect 25913 68274 26006 68340
tri 25913 68258 25929 68274 ne
rect 25929 68258 26006 68274
rect 25746 68159 25894 68241
rect 25634 68126 25711 68142
tri 25711 68126 25727 68142 sw
rect 25634 68060 25727 68126
rect 25763 68001 25877 68159
tri 25913 68126 25929 68142 se
rect 25929 68126 26006 68142
rect 25913 68060 26006 68126
rect 25634 67925 26006 68001
rect 25634 67800 25727 67866
rect 25634 67784 25711 67800
tri 25711 67784 25727 67800 nw
rect 25763 67767 25877 67925
rect 25913 67800 26006 67866
tri 25913 67784 25929 67800 ne
rect 25929 67784 26006 67800
rect 25746 67685 25894 67767
rect 25634 67652 25711 67668
tri 25711 67652 25727 67668 sw
rect 25634 67586 25727 67652
rect 25634 67484 25727 67550
rect 25634 67468 25711 67484
tri 25711 67468 25727 67484 nw
rect 25763 67451 25877 67685
tri 25913 67652 25929 67668 se
rect 25929 67652 26006 67668
rect 25913 67586 26006 67652
rect 25913 67484 26006 67550
tri 25913 67468 25929 67484 ne
rect 25929 67468 26006 67484
rect 25746 67369 25894 67451
rect 25634 67336 25711 67352
tri 25711 67336 25727 67352 sw
rect 25634 67270 25727 67336
rect 25763 67211 25877 67369
tri 25913 67336 25929 67352 se
rect 25929 67336 26006 67352
rect 25913 67270 26006 67336
rect 25634 67135 26006 67211
rect 25634 67010 25727 67076
rect 25634 66994 25711 67010
tri 25711 66994 25727 67010 nw
rect 25763 66977 25877 67135
rect 25913 67010 26006 67076
tri 25913 66994 25929 67010 ne
rect 25929 66994 26006 67010
rect 25746 66895 25894 66977
rect 25634 66862 25711 66878
tri 25711 66862 25727 66878 sw
rect 25634 66796 25727 66862
rect 25634 66694 25727 66760
rect 25634 66678 25711 66694
tri 25711 66678 25727 66694 nw
rect 25763 66661 25877 66895
tri 25913 66862 25929 66878 se
rect 25929 66862 26006 66878
rect 25913 66796 26006 66862
rect 25913 66694 26006 66760
tri 25913 66678 25929 66694 ne
rect 25929 66678 26006 66694
rect 25746 66579 25894 66661
rect 25634 66546 25711 66562
tri 25711 66546 25727 66562 sw
rect 25634 66480 25727 66546
rect 25763 66421 25877 66579
tri 25913 66546 25929 66562 se
rect 25929 66546 26006 66562
rect 25913 66480 26006 66546
rect 25634 66345 26006 66421
rect 25634 66220 25727 66286
rect 25634 66204 25711 66220
tri 25711 66204 25727 66220 nw
rect 25763 66187 25877 66345
rect 25913 66220 26006 66286
tri 25913 66204 25929 66220 ne
rect 25929 66204 26006 66220
rect 25746 66105 25894 66187
rect 25634 66072 25711 66088
tri 25711 66072 25727 66088 sw
rect 25634 66006 25727 66072
rect 25634 65904 25727 65970
rect 25634 65888 25711 65904
tri 25711 65888 25727 65904 nw
rect 25763 65871 25877 66105
tri 25913 66072 25929 66088 se
rect 25929 66072 26006 66088
rect 25913 66006 26006 66072
rect 25913 65904 26006 65970
tri 25913 65888 25929 65904 ne
rect 25929 65888 26006 65904
rect 25746 65789 25894 65871
rect 25634 65756 25711 65772
tri 25711 65756 25727 65772 sw
rect 25634 65690 25727 65756
rect 25763 65631 25877 65789
tri 25913 65756 25929 65772 se
rect 25929 65756 26006 65772
rect 25913 65690 26006 65756
rect 25634 65555 26006 65631
rect 25634 65430 25727 65496
rect 25634 65414 25711 65430
tri 25711 65414 25727 65430 nw
rect 25763 65397 25877 65555
rect 25913 65430 26006 65496
tri 25913 65414 25929 65430 ne
rect 25929 65414 26006 65430
rect 25746 65315 25894 65397
rect 25634 65282 25711 65298
tri 25711 65282 25727 65298 sw
rect 25634 65216 25727 65282
rect 25634 65114 25727 65180
rect 25634 65098 25711 65114
tri 25711 65098 25727 65114 nw
rect 25763 65081 25877 65315
tri 25913 65282 25929 65298 se
rect 25929 65282 26006 65298
rect 25913 65216 26006 65282
rect 25913 65114 26006 65180
tri 25913 65098 25929 65114 ne
rect 25929 65098 26006 65114
rect 25746 64999 25894 65081
rect 25634 64966 25711 64982
tri 25711 64966 25727 64982 sw
rect 25634 64900 25727 64966
rect 25763 64841 25877 64999
tri 25913 64966 25929 64982 se
rect 25929 64966 26006 64982
rect 25913 64900 26006 64966
rect 25634 64765 26006 64841
rect 25634 64640 25727 64706
rect 25634 64624 25711 64640
tri 25711 64624 25727 64640 nw
rect 25763 64607 25877 64765
rect 25913 64640 26006 64706
tri 25913 64624 25929 64640 ne
rect 25929 64624 26006 64640
rect 25746 64525 25894 64607
rect 25634 64492 25711 64508
tri 25711 64492 25727 64508 sw
rect 25634 64426 25727 64492
rect 25634 64324 25727 64390
rect 25634 64308 25711 64324
tri 25711 64308 25727 64324 nw
rect 25763 64291 25877 64525
tri 25913 64492 25929 64508 se
rect 25929 64492 26006 64508
rect 25913 64426 26006 64492
rect 25913 64324 26006 64390
tri 25913 64308 25929 64324 ne
rect 25929 64308 26006 64324
rect 25746 64209 25894 64291
rect 25634 64176 25711 64192
tri 25711 64176 25727 64192 sw
rect 25634 64110 25727 64176
rect 25763 64051 25877 64209
tri 25913 64176 25929 64192 se
rect 25929 64176 26006 64192
rect 25913 64110 26006 64176
rect 25634 63975 26006 64051
rect 25634 63850 25727 63916
rect 25634 63834 25711 63850
tri 25711 63834 25727 63850 nw
rect 25763 63817 25877 63975
rect 25913 63850 26006 63916
tri 25913 63834 25929 63850 ne
rect 25929 63834 26006 63850
rect 25746 63735 25894 63817
rect 25634 63702 25711 63718
tri 25711 63702 25727 63718 sw
rect 25634 63636 25727 63702
rect 25634 63534 25727 63600
rect 25634 63518 25711 63534
tri 25711 63518 25727 63534 nw
rect 25763 63501 25877 63735
tri 25913 63702 25929 63718 se
rect 25929 63702 26006 63718
rect 25913 63636 26006 63702
rect 25913 63534 26006 63600
tri 25913 63518 25929 63534 ne
rect 25929 63518 26006 63534
rect 25746 63419 25894 63501
rect 25634 63386 25711 63402
tri 25711 63386 25727 63402 sw
rect 25634 63320 25727 63386
rect 25763 63261 25877 63419
tri 25913 63386 25929 63402 se
rect 25929 63386 26006 63402
rect 25913 63320 26006 63386
rect 25634 63185 26006 63261
rect 25634 63060 25727 63126
rect 25634 63044 25711 63060
tri 25711 63044 25727 63060 nw
rect 25763 63027 25877 63185
rect 25913 63060 26006 63126
tri 25913 63044 25929 63060 ne
rect 25929 63044 26006 63060
rect 25746 62945 25894 63027
rect 25634 62912 25711 62928
tri 25711 62912 25727 62928 sw
rect 25634 62846 25727 62912
rect 25634 62744 25727 62810
rect 25634 62728 25711 62744
tri 25711 62728 25727 62744 nw
rect 25763 62711 25877 62945
tri 25913 62912 25929 62928 se
rect 25929 62912 26006 62928
rect 25913 62846 26006 62912
rect 25913 62744 26006 62810
tri 25913 62728 25929 62744 ne
rect 25929 62728 26006 62744
rect 25746 62629 25894 62711
rect 25634 62596 25711 62612
tri 25711 62596 25727 62612 sw
rect 25634 62530 25727 62596
rect 25763 62471 25877 62629
tri 25913 62596 25929 62612 se
rect 25929 62596 26006 62612
rect 25913 62530 26006 62596
rect 25634 62395 26006 62471
rect 25634 62270 25727 62336
rect 25634 62254 25711 62270
tri 25711 62254 25727 62270 nw
rect 25763 62237 25877 62395
rect 25913 62270 26006 62336
tri 25913 62254 25929 62270 ne
rect 25929 62254 26006 62270
rect 25746 62155 25894 62237
rect 25634 62122 25711 62138
tri 25711 62122 25727 62138 sw
rect 25634 62056 25727 62122
rect 25634 61954 25727 62020
rect 25634 61938 25711 61954
tri 25711 61938 25727 61954 nw
rect 25763 61921 25877 62155
tri 25913 62122 25929 62138 se
rect 25929 62122 26006 62138
rect 25913 62056 26006 62122
rect 25913 61954 26006 62020
tri 25913 61938 25929 61954 ne
rect 25929 61938 26006 61954
rect 25746 61839 25894 61921
rect 25634 61806 25711 61822
tri 25711 61806 25727 61822 sw
rect 25634 61740 25727 61806
rect 25763 61681 25877 61839
tri 25913 61806 25929 61822 se
rect 25929 61806 26006 61822
rect 25913 61740 26006 61806
rect 25634 61605 26006 61681
rect 25634 61480 25727 61546
rect 25634 61464 25711 61480
tri 25711 61464 25727 61480 nw
rect 25763 61447 25877 61605
rect 25913 61480 26006 61546
tri 25913 61464 25929 61480 ne
rect 25929 61464 26006 61480
rect 25746 61365 25894 61447
rect 25634 61332 25711 61348
tri 25711 61332 25727 61348 sw
rect 25634 61266 25727 61332
rect 25634 61164 25727 61230
rect 25634 61148 25711 61164
tri 25711 61148 25727 61164 nw
rect 25763 61131 25877 61365
tri 25913 61332 25929 61348 se
rect 25929 61332 26006 61348
rect 25913 61266 26006 61332
rect 25913 61164 26006 61230
tri 25913 61148 25929 61164 ne
rect 25929 61148 26006 61164
rect 25746 61049 25894 61131
rect 25634 61016 25711 61032
tri 25711 61016 25727 61032 sw
rect 25634 60950 25727 61016
rect 25763 60891 25877 61049
tri 25913 61016 25929 61032 se
rect 25929 61016 26006 61032
rect 25913 60950 26006 61016
rect 25634 60815 26006 60891
rect 25634 60690 25727 60756
rect 25634 60674 25711 60690
tri 25711 60674 25727 60690 nw
rect 25763 60657 25877 60815
rect 25913 60690 26006 60756
tri 25913 60674 25929 60690 ne
rect 25929 60674 26006 60690
rect 25746 60575 25894 60657
rect 25634 60542 25711 60558
tri 25711 60542 25727 60558 sw
rect 25634 60476 25727 60542
rect 25634 60374 25727 60440
rect 25634 60358 25711 60374
tri 25711 60358 25727 60374 nw
rect 25763 60341 25877 60575
tri 25913 60542 25929 60558 se
rect 25929 60542 26006 60558
rect 25913 60476 26006 60542
rect 25913 60374 26006 60440
tri 25913 60358 25929 60374 ne
rect 25929 60358 26006 60374
rect 25746 60259 25894 60341
rect 25634 60226 25711 60242
tri 25711 60226 25727 60242 sw
rect 25634 60160 25727 60226
rect 25763 60101 25877 60259
tri 25913 60226 25929 60242 se
rect 25929 60226 26006 60242
rect 25913 60160 26006 60226
rect 25634 60025 26006 60101
rect 25634 59900 25727 59966
rect 25634 59884 25711 59900
tri 25711 59884 25727 59900 nw
rect 25763 59867 25877 60025
rect 25913 59900 26006 59966
tri 25913 59884 25929 59900 ne
rect 25929 59884 26006 59900
rect 25746 59785 25894 59867
rect 25634 59752 25711 59768
tri 25711 59752 25727 59768 sw
rect 25634 59686 25727 59752
rect 25634 59584 25727 59650
rect 25634 59568 25711 59584
tri 25711 59568 25727 59584 nw
rect 25763 59551 25877 59785
tri 25913 59752 25929 59768 se
rect 25929 59752 26006 59768
rect 25913 59686 26006 59752
rect 25913 59584 26006 59650
tri 25913 59568 25929 59584 ne
rect 25929 59568 26006 59584
rect 25746 59469 25894 59551
rect 25634 59436 25711 59452
tri 25711 59436 25727 59452 sw
rect 25634 59370 25727 59436
rect 25763 59311 25877 59469
tri 25913 59436 25929 59452 se
rect 25929 59436 26006 59452
rect 25913 59370 26006 59436
rect 25634 59235 26006 59311
rect 25634 59110 25727 59176
rect 25634 59094 25711 59110
tri 25711 59094 25727 59110 nw
rect 25763 59077 25877 59235
rect 25913 59110 26006 59176
tri 25913 59094 25929 59110 ne
rect 25929 59094 26006 59110
rect 25746 58995 25894 59077
rect 25634 58962 25711 58978
tri 25711 58962 25727 58978 sw
rect 25634 58896 25727 58962
rect 25634 58794 25727 58860
rect 25634 58778 25711 58794
tri 25711 58778 25727 58794 nw
rect 25763 58761 25877 58995
tri 25913 58962 25929 58978 se
rect 25929 58962 26006 58978
rect 25913 58896 26006 58962
rect 25913 58794 26006 58860
tri 25913 58778 25929 58794 ne
rect 25929 58778 26006 58794
rect 25746 58679 25894 58761
rect 25634 58646 25711 58662
tri 25711 58646 25727 58662 sw
rect 25634 58580 25727 58646
rect 25763 58521 25877 58679
tri 25913 58646 25929 58662 se
rect 25929 58646 26006 58662
rect 25913 58580 26006 58646
rect 25634 58445 26006 58521
rect 25634 58320 25727 58386
rect 25634 58304 25711 58320
tri 25711 58304 25727 58320 nw
rect 25763 58287 25877 58445
rect 25913 58320 26006 58386
tri 25913 58304 25929 58320 ne
rect 25929 58304 26006 58320
rect 25746 58205 25894 58287
rect 25634 58172 25711 58188
tri 25711 58172 25727 58188 sw
rect 25634 58106 25727 58172
rect 25634 58004 25727 58070
rect 25634 57988 25711 58004
tri 25711 57988 25727 58004 nw
rect 25763 57971 25877 58205
tri 25913 58172 25929 58188 se
rect 25929 58172 26006 58188
rect 25913 58106 26006 58172
rect 25913 58004 26006 58070
tri 25913 57988 25929 58004 ne
rect 25929 57988 26006 58004
rect 25746 57889 25894 57971
rect 25634 57856 25711 57872
tri 25711 57856 25727 57872 sw
rect 25634 57790 25727 57856
rect 25763 57731 25877 57889
tri 25913 57856 25929 57872 se
rect 25929 57856 26006 57872
rect 25913 57790 26006 57856
rect 25634 57655 26006 57731
rect 25634 57530 25727 57596
rect 25634 57514 25711 57530
tri 25711 57514 25727 57530 nw
rect 25763 57497 25877 57655
rect 25913 57530 26006 57596
tri 25913 57514 25929 57530 ne
rect 25929 57514 26006 57530
rect 25746 57415 25894 57497
rect 25634 57382 25711 57398
tri 25711 57382 25727 57398 sw
rect 25634 57316 25727 57382
rect 25634 57214 25727 57280
rect 25634 57198 25711 57214
tri 25711 57198 25727 57214 nw
rect 25763 57181 25877 57415
tri 25913 57382 25929 57398 se
rect 25929 57382 26006 57398
rect 25913 57316 26006 57382
rect 25913 57214 26006 57280
tri 25913 57198 25929 57214 ne
rect 25929 57198 26006 57214
rect 25746 57099 25894 57181
rect 25634 57066 25711 57082
tri 25711 57066 25727 57082 sw
rect 25634 57000 25727 57066
rect 25763 56941 25877 57099
tri 25913 57066 25929 57082 se
rect 25929 57066 26006 57082
rect 25913 57000 26006 57066
rect 25634 56865 26006 56941
rect 25634 56740 25727 56806
rect 25634 56724 25711 56740
tri 25711 56724 25727 56740 nw
rect 25763 56707 25877 56865
rect 25913 56740 26006 56806
tri 25913 56724 25929 56740 ne
rect 25929 56724 26006 56740
rect 25746 56625 25894 56707
rect 25634 56592 25711 56608
tri 25711 56592 25727 56608 sw
rect 25634 56526 25727 56592
rect 25634 56424 25727 56490
rect 25634 56408 25711 56424
tri 25711 56408 25727 56424 nw
rect 25763 56391 25877 56625
tri 25913 56592 25929 56608 se
rect 25929 56592 26006 56608
rect 25913 56526 26006 56592
rect 25913 56424 26006 56490
tri 25913 56408 25929 56424 ne
rect 25929 56408 26006 56424
rect 25746 56309 25894 56391
rect 25634 56276 25711 56292
tri 25711 56276 25727 56292 sw
rect 25634 56210 25727 56276
rect 25763 56151 25877 56309
tri 25913 56276 25929 56292 se
rect 25929 56276 26006 56292
rect 25913 56210 26006 56276
rect 25634 56075 26006 56151
rect 25634 55950 25727 56016
rect 25634 55934 25711 55950
tri 25711 55934 25727 55950 nw
rect 25763 55917 25877 56075
rect 25913 55950 26006 56016
tri 25913 55934 25929 55950 ne
rect 25929 55934 26006 55950
rect 25746 55835 25894 55917
rect 25634 55802 25711 55818
tri 25711 55802 25727 55818 sw
rect 25634 55736 25727 55802
rect 25634 55634 25727 55700
rect 25634 55618 25711 55634
tri 25711 55618 25727 55634 nw
rect 25763 55601 25877 55835
tri 25913 55802 25929 55818 se
rect 25929 55802 26006 55818
rect 25913 55736 26006 55802
rect 25913 55634 26006 55700
tri 25913 55618 25929 55634 ne
rect 25929 55618 26006 55634
rect 25746 55519 25894 55601
rect 25634 55486 25711 55502
tri 25711 55486 25727 55502 sw
rect 25634 55420 25727 55486
rect 25763 55361 25877 55519
tri 25913 55486 25929 55502 se
rect 25929 55486 26006 55502
rect 25913 55420 26006 55486
rect 25634 55285 26006 55361
rect 25634 55160 25727 55226
rect 25634 55144 25711 55160
tri 25711 55144 25727 55160 nw
rect 25763 55127 25877 55285
rect 25913 55160 26006 55226
tri 25913 55144 25929 55160 ne
rect 25929 55144 26006 55160
rect 25746 55045 25894 55127
rect 25634 55012 25711 55028
tri 25711 55012 25727 55028 sw
rect 25634 54946 25727 55012
rect 25634 54844 25727 54910
rect 25634 54828 25711 54844
tri 25711 54828 25727 54844 nw
rect 25763 54811 25877 55045
tri 25913 55012 25929 55028 se
rect 25929 55012 26006 55028
rect 25913 54946 26006 55012
rect 25913 54844 26006 54910
tri 25913 54828 25929 54844 ne
rect 25929 54828 26006 54844
rect 25746 54729 25894 54811
rect 25634 54696 25711 54712
tri 25711 54696 25727 54712 sw
rect 25634 54630 25727 54696
rect 25763 54571 25877 54729
tri 25913 54696 25929 54712 se
rect 25929 54696 26006 54712
rect 25913 54630 26006 54696
rect 25634 54495 26006 54571
rect 25634 54370 25727 54436
rect 25634 54354 25711 54370
tri 25711 54354 25727 54370 nw
rect 25763 54337 25877 54495
rect 25913 54370 26006 54436
tri 25913 54354 25929 54370 ne
rect 25929 54354 26006 54370
rect 25746 54255 25894 54337
rect 25634 54222 25711 54238
tri 25711 54222 25727 54238 sw
rect 25634 54156 25727 54222
rect 25634 54054 25727 54120
rect 25634 54038 25711 54054
tri 25711 54038 25727 54054 nw
rect 25763 54021 25877 54255
tri 25913 54222 25929 54238 se
rect 25929 54222 26006 54238
rect 25913 54156 26006 54222
rect 25913 54054 26006 54120
tri 25913 54038 25929 54054 ne
rect 25929 54038 26006 54054
rect 25746 53939 25894 54021
rect 25634 53906 25711 53922
tri 25711 53906 25727 53922 sw
rect 25634 53840 25727 53906
rect 25763 53781 25877 53939
tri 25913 53906 25929 53922 se
rect 25929 53906 26006 53922
rect 25913 53840 26006 53906
rect 25634 53705 26006 53781
rect 25634 53580 25727 53646
rect 25634 53564 25711 53580
tri 25711 53564 25727 53580 nw
rect 25763 53547 25877 53705
rect 25913 53580 26006 53646
tri 25913 53564 25929 53580 ne
rect 25929 53564 26006 53580
rect 25746 53465 25894 53547
rect 25634 53432 25711 53448
tri 25711 53432 25727 53448 sw
rect 25634 53366 25727 53432
rect 25634 53264 25727 53330
rect 25634 53248 25711 53264
tri 25711 53248 25727 53264 nw
rect 25763 53231 25877 53465
tri 25913 53432 25929 53448 se
rect 25929 53432 26006 53448
rect 25913 53366 26006 53432
rect 25913 53264 26006 53330
tri 25913 53248 25929 53264 ne
rect 25929 53248 26006 53264
rect 25746 53149 25894 53231
rect 25634 53116 25711 53132
tri 25711 53116 25727 53132 sw
rect 25634 53050 25727 53116
rect 25763 52991 25877 53149
tri 25913 53116 25929 53132 se
rect 25929 53116 26006 53132
rect 25913 53050 26006 53116
rect 25634 52915 26006 52991
rect 25634 52790 25727 52856
rect 25634 52774 25711 52790
tri 25711 52774 25727 52790 nw
rect 25763 52757 25877 52915
rect 25913 52790 26006 52856
tri 25913 52774 25929 52790 ne
rect 25929 52774 26006 52790
rect 25746 52675 25894 52757
rect 25634 52642 25711 52658
tri 25711 52642 25727 52658 sw
rect 25634 52576 25727 52642
rect 25634 52474 25727 52540
rect 25634 52458 25711 52474
tri 25711 52458 25727 52474 nw
rect 25763 52441 25877 52675
tri 25913 52642 25929 52658 se
rect 25929 52642 26006 52658
rect 25913 52576 26006 52642
rect 25913 52474 26006 52540
tri 25913 52458 25929 52474 ne
rect 25929 52458 26006 52474
rect 25746 52359 25894 52441
rect 25634 52326 25711 52342
tri 25711 52326 25727 52342 sw
rect 25634 52260 25727 52326
rect 25763 52201 25877 52359
tri 25913 52326 25929 52342 se
rect 25929 52326 26006 52342
rect 25913 52260 26006 52326
rect 25634 52125 26006 52201
rect 25634 52000 25727 52066
rect 25634 51984 25711 52000
tri 25711 51984 25727 52000 nw
rect 25763 51967 25877 52125
rect 25913 52000 26006 52066
tri 25913 51984 25929 52000 ne
rect 25929 51984 26006 52000
rect 25746 51885 25894 51967
rect 25634 51852 25711 51868
tri 25711 51852 25727 51868 sw
rect 25634 51786 25727 51852
rect 25634 51684 25727 51750
rect 25634 51668 25711 51684
tri 25711 51668 25727 51684 nw
rect 25763 51651 25877 51885
tri 25913 51852 25929 51868 se
rect 25929 51852 26006 51868
rect 25913 51786 26006 51852
rect 25913 51684 26006 51750
tri 25913 51668 25929 51684 ne
rect 25929 51668 26006 51684
rect 25746 51569 25894 51651
rect 25634 51536 25711 51552
tri 25711 51536 25727 51552 sw
rect 25634 51470 25727 51536
rect 25763 51411 25877 51569
tri 25913 51536 25929 51552 se
rect 25929 51536 26006 51552
rect 25913 51470 26006 51536
rect 25634 51335 26006 51411
rect 25634 51210 25727 51276
rect 25634 51194 25711 51210
tri 25711 51194 25727 51210 nw
rect 25763 51177 25877 51335
rect 25913 51210 26006 51276
tri 25913 51194 25929 51210 ne
rect 25929 51194 26006 51210
rect 25746 51095 25894 51177
rect 25634 51062 25711 51078
tri 25711 51062 25727 51078 sw
rect 25634 50996 25727 51062
rect 25634 50894 25727 50960
rect 25634 50878 25711 50894
tri 25711 50878 25727 50894 nw
rect 25763 50861 25877 51095
tri 25913 51062 25929 51078 se
rect 25929 51062 26006 51078
rect 25913 50996 26006 51062
rect 25913 50894 26006 50960
tri 25913 50878 25929 50894 ne
rect 25929 50878 26006 50894
rect 25746 50779 25894 50861
rect 25634 50746 25711 50762
tri 25711 50746 25727 50762 sw
rect 25634 50680 25727 50746
rect 25763 50621 25877 50779
tri 25913 50746 25929 50762 se
rect 25929 50746 26006 50762
rect 25913 50680 26006 50746
rect 25634 50545 26006 50621
rect 25634 50420 25727 50486
rect 25634 50404 25711 50420
tri 25711 50404 25727 50420 nw
rect 25763 50387 25877 50545
rect 25913 50420 26006 50486
tri 25913 50404 25929 50420 ne
rect 25929 50404 26006 50420
rect 25746 50305 25894 50387
rect 25634 50272 25711 50288
tri 25711 50272 25727 50288 sw
rect 25634 50206 25727 50272
rect 25634 50104 25727 50170
rect 25634 50088 25711 50104
tri 25711 50088 25727 50104 nw
rect 25763 50071 25877 50305
tri 25913 50272 25929 50288 se
rect 25929 50272 26006 50288
rect 25913 50206 26006 50272
rect 25913 50104 26006 50170
tri 25913 50088 25929 50104 ne
rect 25929 50088 26006 50104
rect 25746 49989 25894 50071
rect 25634 49956 25711 49972
tri 25711 49956 25727 49972 sw
rect 25634 49890 25727 49956
rect 25763 49831 25877 49989
tri 25913 49956 25929 49972 se
rect 25929 49956 26006 49972
rect 25913 49890 26006 49956
rect 25634 49755 26006 49831
rect 25634 49630 25727 49696
rect 25634 49614 25711 49630
tri 25711 49614 25727 49630 nw
rect 25763 49597 25877 49755
rect 25913 49630 26006 49696
tri 25913 49614 25929 49630 ne
rect 25929 49614 26006 49630
rect 25746 49515 25894 49597
rect 25634 49482 25711 49498
tri 25711 49482 25727 49498 sw
rect 25634 49416 25727 49482
rect 25634 49314 25727 49380
rect 25634 49298 25711 49314
tri 25711 49298 25727 49314 nw
rect 25763 49281 25877 49515
tri 25913 49482 25929 49498 se
rect 25929 49482 26006 49498
rect 25913 49416 26006 49482
rect 25913 49314 26006 49380
tri 25913 49298 25929 49314 ne
rect 25929 49298 26006 49314
rect 25746 49199 25894 49281
rect 25634 49166 25711 49182
tri 25711 49166 25727 49182 sw
rect 25634 49100 25727 49166
rect 25763 49041 25877 49199
tri 25913 49166 25929 49182 se
rect 25929 49166 26006 49182
rect 25913 49100 26006 49166
rect 25634 48965 26006 49041
rect 25634 48840 25727 48906
rect 25634 48824 25711 48840
tri 25711 48824 25727 48840 nw
rect 25763 48807 25877 48965
rect 25913 48840 26006 48906
tri 25913 48824 25929 48840 ne
rect 25929 48824 26006 48840
rect 25746 48725 25894 48807
rect 25634 48692 25711 48708
tri 25711 48692 25727 48708 sw
rect 25634 48626 25727 48692
rect 25634 48524 25727 48590
rect 25634 48508 25711 48524
tri 25711 48508 25727 48524 nw
rect 25763 48491 25877 48725
tri 25913 48692 25929 48708 se
rect 25929 48692 26006 48708
rect 25913 48626 26006 48692
rect 25913 48524 26006 48590
tri 25913 48508 25929 48524 ne
rect 25929 48508 26006 48524
rect 25746 48409 25894 48491
rect 25634 48376 25711 48392
tri 25711 48376 25727 48392 sw
rect 25634 48310 25727 48376
rect 25763 48251 25877 48409
tri 25913 48376 25929 48392 se
rect 25929 48376 26006 48392
rect 25913 48310 26006 48376
rect 25634 48175 26006 48251
rect 25634 48050 25727 48116
rect 25634 48034 25711 48050
tri 25711 48034 25727 48050 nw
rect 25763 48017 25877 48175
rect 25913 48050 26006 48116
tri 25913 48034 25929 48050 ne
rect 25929 48034 26006 48050
rect 25746 47935 25894 48017
rect 25634 47902 25711 47918
tri 25711 47902 25727 47918 sw
rect 25634 47836 25727 47902
rect 25634 47734 25727 47800
rect 25634 47718 25711 47734
tri 25711 47718 25727 47734 nw
rect 25763 47701 25877 47935
tri 25913 47902 25929 47918 se
rect 25929 47902 26006 47918
rect 25913 47836 26006 47902
rect 25913 47734 26006 47800
tri 25913 47718 25929 47734 ne
rect 25929 47718 26006 47734
rect 25746 47619 25894 47701
rect 25634 47586 25711 47602
tri 25711 47586 25727 47602 sw
rect 25634 47520 25727 47586
rect 25763 47461 25877 47619
tri 25913 47586 25929 47602 se
rect 25929 47586 26006 47602
rect 25913 47520 26006 47586
rect 25634 47385 26006 47461
rect 25634 47260 25727 47326
rect 25634 47244 25711 47260
tri 25711 47244 25727 47260 nw
rect 25763 47227 25877 47385
rect 25913 47260 26006 47326
tri 25913 47244 25929 47260 ne
rect 25929 47244 26006 47260
rect 25746 47145 25894 47227
rect 25634 47112 25711 47128
tri 25711 47112 25727 47128 sw
rect 25634 47046 25727 47112
rect 25634 46944 25727 47010
rect 25634 46928 25711 46944
tri 25711 46928 25727 46944 nw
rect 25763 46911 25877 47145
tri 25913 47112 25929 47128 se
rect 25929 47112 26006 47128
rect 25913 47046 26006 47112
rect 25913 46944 26006 47010
tri 25913 46928 25929 46944 ne
rect 25929 46928 26006 46944
rect 25746 46829 25894 46911
rect 25634 46796 25711 46812
tri 25711 46796 25727 46812 sw
rect 25634 46730 25727 46796
rect 25763 46671 25877 46829
tri 25913 46796 25929 46812 se
rect 25929 46796 26006 46812
rect 25913 46730 26006 46796
rect 25634 46595 26006 46671
rect 25634 46470 25727 46536
rect 25634 46454 25711 46470
tri 25711 46454 25727 46470 nw
rect 25763 46437 25877 46595
rect 25913 46470 26006 46536
tri 25913 46454 25929 46470 ne
rect 25929 46454 26006 46470
rect 25746 46355 25894 46437
rect 25634 46322 25711 46338
tri 25711 46322 25727 46338 sw
rect 25634 46256 25727 46322
rect 25634 46154 25727 46220
rect 25634 46138 25711 46154
tri 25711 46138 25727 46154 nw
rect 25763 46121 25877 46355
tri 25913 46322 25929 46338 se
rect 25929 46322 26006 46338
rect 25913 46256 26006 46322
rect 25913 46154 26006 46220
tri 25913 46138 25929 46154 ne
rect 25929 46138 26006 46154
rect 25746 46039 25894 46121
rect 25634 46006 25711 46022
tri 25711 46006 25727 46022 sw
rect 25634 45940 25727 46006
rect 25763 45881 25877 46039
tri 25913 46006 25929 46022 se
rect 25929 46006 26006 46022
rect 25913 45940 26006 46006
rect 25634 45805 26006 45881
rect 25634 45680 25727 45746
rect 25634 45664 25711 45680
tri 25711 45664 25727 45680 nw
rect 25763 45647 25877 45805
rect 25913 45680 26006 45746
tri 25913 45664 25929 45680 ne
rect 25929 45664 26006 45680
rect 25746 45565 25894 45647
rect 25634 45532 25711 45548
tri 25711 45532 25727 45548 sw
rect 25634 45466 25727 45532
rect 25634 45364 25727 45430
rect 25634 45348 25711 45364
tri 25711 45348 25727 45364 nw
rect 25763 45331 25877 45565
tri 25913 45532 25929 45548 se
rect 25929 45532 26006 45548
rect 25913 45466 26006 45532
rect 25913 45364 26006 45430
tri 25913 45348 25929 45364 ne
rect 25929 45348 26006 45364
rect 25746 45249 25894 45331
rect 25634 45216 25711 45232
tri 25711 45216 25727 45232 sw
rect 25634 45150 25727 45216
rect 25763 45091 25877 45249
tri 25913 45216 25929 45232 se
rect 25929 45216 26006 45232
rect 25913 45150 26006 45216
rect 25634 45015 26006 45091
rect 25634 44890 25727 44956
rect 25634 44874 25711 44890
tri 25711 44874 25727 44890 nw
rect 25763 44857 25877 45015
rect 25913 44890 26006 44956
tri 25913 44874 25929 44890 ne
rect 25929 44874 26006 44890
rect 25746 44775 25894 44857
rect 25634 44742 25711 44758
tri 25711 44742 25727 44758 sw
rect 25634 44676 25727 44742
rect 25634 44574 25727 44640
rect 25634 44558 25711 44574
tri 25711 44558 25727 44574 nw
rect 25763 44541 25877 44775
tri 25913 44742 25929 44758 se
rect 25929 44742 26006 44758
rect 25913 44676 26006 44742
rect 25913 44574 26006 44640
tri 25913 44558 25929 44574 ne
rect 25929 44558 26006 44574
rect 25746 44459 25894 44541
rect 25634 44426 25711 44442
tri 25711 44426 25727 44442 sw
rect 25634 44360 25727 44426
rect 25763 44301 25877 44459
tri 25913 44426 25929 44442 se
rect 25929 44426 26006 44442
rect 25913 44360 26006 44426
rect 25634 44225 26006 44301
rect 25634 44100 25727 44166
rect 25634 44084 25711 44100
tri 25711 44084 25727 44100 nw
rect 25763 44067 25877 44225
rect 25913 44100 26006 44166
tri 25913 44084 25929 44100 ne
rect 25929 44084 26006 44100
rect 25746 43985 25894 44067
rect 25634 43952 25711 43968
tri 25711 43952 25727 43968 sw
rect 25634 43886 25727 43952
rect 25634 43784 25727 43850
rect 25634 43768 25711 43784
tri 25711 43768 25727 43784 nw
rect 25763 43751 25877 43985
tri 25913 43952 25929 43968 se
rect 25929 43952 26006 43968
rect 25913 43886 26006 43952
rect 25913 43784 26006 43850
tri 25913 43768 25929 43784 ne
rect 25929 43768 26006 43784
rect 25746 43669 25894 43751
rect 25634 43636 25711 43652
tri 25711 43636 25727 43652 sw
rect 25634 43570 25727 43636
rect 25763 43511 25877 43669
tri 25913 43636 25929 43652 se
rect 25929 43636 26006 43652
rect 25913 43570 26006 43636
rect 25634 43435 26006 43511
rect 25634 43310 25727 43376
rect 25634 43294 25711 43310
tri 25711 43294 25727 43310 nw
rect 25763 43277 25877 43435
rect 25913 43310 26006 43376
tri 25913 43294 25929 43310 ne
rect 25929 43294 26006 43310
rect 25746 43195 25894 43277
rect 25634 43162 25711 43178
tri 25711 43162 25727 43178 sw
rect 25634 43096 25727 43162
rect 25634 42994 25727 43060
rect 25634 42978 25711 42994
tri 25711 42978 25727 42994 nw
rect 25763 42961 25877 43195
tri 25913 43162 25929 43178 se
rect 25929 43162 26006 43178
rect 25913 43096 26006 43162
rect 25913 42994 26006 43060
tri 25913 42978 25929 42994 ne
rect 25929 42978 26006 42994
rect 25746 42879 25894 42961
rect 25634 42846 25711 42862
tri 25711 42846 25727 42862 sw
rect 25634 42780 25727 42846
rect 25763 42721 25877 42879
tri 25913 42846 25929 42862 se
rect 25929 42846 26006 42862
rect 25913 42780 26006 42846
rect 25634 42645 26006 42721
rect 25634 42520 25727 42586
rect 25634 42504 25711 42520
tri 25711 42504 25727 42520 nw
rect 25763 42487 25877 42645
rect 25913 42520 26006 42586
tri 25913 42504 25929 42520 ne
rect 25929 42504 26006 42520
rect 25746 42405 25894 42487
rect 25634 42372 25711 42388
tri 25711 42372 25727 42388 sw
rect 25634 42306 25727 42372
rect 25634 42204 25727 42270
rect 25634 42188 25711 42204
tri 25711 42188 25727 42204 nw
rect 25763 42171 25877 42405
tri 25913 42372 25929 42388 se
rect 25929 42372 26006 42388
rect 25913 42306 26006 42372
rect 25913 42204 26006 42270
tri 25913 42188 25929 42204 ne
rect 25929 42188 26006 42204
rect 25746 42089 25894 42171
rect 25634 42056 25711 42072
tri 25711 42056 25727 42072 sw
rect 25634 41990 25727 42056
rect 25763 41931 25877 42089
tri 25913 42056 25929 42072 se
rect 25929 42056 26006 42072
rect 25913 41990 26006 42056
rect 25634 41855 26006 41931
rect 25634 41730 25727 41796
rect 25634 41714 25711 41730
tri 25711 41714 25727 41730 nw
rect 25763 41697 25877 41855
rect 25913 41730 26006 41796
tri 25913 41714 25929 41730 ne
rect 25929 41714 26006 41730
rect 25746 41615 25894 41697
rect 25634 41582 25711 41598
tri 25711 41582 25727 41598 sw
rect 25634 41516 25727 41582
rect 25634 41414 25727 41480
rect 25634 41398 25711 41414
tri 25711 41398 25727 41414 nw
rect 25763 41381 25877 41615
tri 25913 41582 25929 41598 se
rect 25929 41582 26006 41598
rect 25913 41516 26006 41582
rect 25913 41414 26006 41480
tri 25913 41398 25929 41414 ne
rect 25929 41398 26006 41414
rect 25746 41299 25894 41381
rect 25634 41266 25711 41282
tri 25711 41266 25727 41282 sw
rect 25634 41200 25727 41266
rect 25763 41141 25877 41299
tri 25913 41266 25929 41282 se
rect 25929 41266 26006 41282
rect 25913 41200 26006 41266
rect 25634 41065 26006 41141
rect 25634 40940 25727 41006
rect 25634 40924 25711 40940
tri 25711 40924 25727 40940 nw
rect 25763 40907 25877 41065
rect 25913 40940 26006 41006
tri 25913 40924 25929 40940 ne
rect 25929 40924 26006 40940
rect 25746 40825 25894 40907
rect 25634 40792 25711 40808
tri 25711 40792 25727 40808 sw
rect 25634 40726 25727 40792
rect 25634 40624 25727 40690
rect 25634 40608 25711 40624
tri 25711 40608 25727 40624 nw
rect 25763 40591 25877 40825
tri 25913 40792 25929 40808 se
rect 25929 40792 26006 40808
rect 25913 40726 26006 40792
rect 25913 40624 26006 40690
tri 25913 40608 25929 40624 ne
rect 25929 40608 26006 40624
rect 25746 40509 25894 40591
rect 25634 40476 25711 40492
tri 25711 40476 25727 40492 sw
rect 25634 40410 25727 40476
rect 25763 40351 25877 40509
tri 25913 40476 25929 40492 se
rect 25929 40476 26006 40492
rect 25913 40410 26006 40476
rect 25634 40275 26006 40351
rect 25634 40150 25727 40216
rect 25634 40134 25711 40150
tri 25711 40134 25727 40150 nw
rect 25763 40117 25877 40275
rect 25913 40150 26006 40216
tri 25913 40134 25929 40150 ne
rect 25929 40134 26006 40150
rect 25746 40035 25894 40117
rect 25634 40002 25711 40018
tri 25711 40002 25727 40018 sw
rect 25634 39936 25727 40002
rect 25634 39834 25727 39900
rect 25634 39818 25711 39834
tri 25711 39818 25727 39834 nw
rect 25763 39801 25877 40035
tri 25913 40002 25929 40018 se
rect 25929 40002 26006 40018
rect 25913 39936 26006 40002
rect 25913 39834 26006 39900
tri 25913 39818 25929 39834 ne
rect 25929 39818 26006 39834
rect 25746 39719 25894 39801
rect 25634 39686 25711 39702
tri 25711 39686 25727 39702 sw
rect 25634 39620 25727 39686
rect 25763 39561 25877 39719
tri 25913 39686 25929 39702 se
rect 25929 39686 26006 39702
rect 25913 39620 26006 39686
rect 25634 39485 26006 39561
rect 25634 39360 25727 39426
rect 25634 39344 25711 39360
tri 25711 39344 25727 39360 nw
rect 25763 39327 25877 39485
rect 25913 39360 26006 39426
tri 25913 39344 25929 39360 ne
rect 25929 39344 26006 39360
rect 25746 39245 25894 39327
rect 25634 39212 25711 39228
tri 25711 39212 25727 39228 sw
rect 25634 39146 25727 39212
rect 25634 39044 25727 39110
rect 25634 39028 25711 39044
tri 25711 39028 25727 39044 nw
rect 25763 39011 25877 39245
tri 25913 39212 25929 39228 se
rect 25929 39212 26006 39228
rect 25913 39146 26006 39212
rect 25913 39044 26006 39110
tri 25913 39028 25929 39044 ne
rect 25929 39028 26006 39044
rect 25746 38929 25894 39011
rect 25634 38896 25711 38912
tri 25711 38896 25727 38912 sw
rect 25634 38830 25727 38896
rect 25763 38771 25877 38929
tri 25913 38896 25929 38912 se
rect 25929 38896 26006 38912
rect 25913 38830 26006 38896
rect 25634 38695 26006 38771
rect 25634 38570 25727 38636
rect 25634 38554 25711 38570
tri 25711 38554 25727 38570 nw
rect 25763 38537 25877 38695
rect 25913 38570 26006 38636
tri 25913 38554 25929 38570 ne
rect 25929 38554 26006 38570
rect 25746 38455 25894 38537
rect 25634 38422 25711 38438
tri 25711 38422 25727 38438 sw
rect 25634 38356 25727 38422
rect 25634 38254 25727 38320
rect 25634 38238 25711 38254
tri 25711 38238 25727 38254 nw
rect 25763 38221 25877 38455
tri 25913 38422 25929 38438 se
rect 25929 38422 26006 38438
rect 25913 38356 26006 38422
rect 25913 38254 26006 38320
tri 25913 38238 25929 38254 ne
rect 25929 38238 26006 38254
rect 25746 38139 25894 38221
rect 25634 38106 25711 38122
tri 25711 38106 25727 38122 sw
rect 25634 38040 25727 38106
rect 25763 37981 25877 38139
tri 25913 38106 25929 38122 se
rect 25929 38106 26006 38122
rect 25913 38040 26006 38106
rect 25634 37905 26006 37981
rect 25634 37780 25727 37846
rect 25634 37764 25711 37780
tri 25711 37764 25727 37780 nw
rect 25763 37747 25877 37905
rect 25913 37780 26006 37846
tri 25913 37764 25929 37780 ne
rect 25929 37764 26006 37780
rect 25746 37665 25894 37747
rect 25634 37632 25711 37648
tri 25711 37632 25727 37648 sw
rect 25634 37566 25727 37632
rect 25634 37464 25727 37530
rect 25634 37448 25711 37464
tri 25711 37448 25727 37464 nw
rect 25763 37431 25877 37665
tri 25913 37632 25929 37648 se
rect 25929 37632 26006 37648
rect 25913 37566 26006 37632
rect 25913 37464 26006 37530
tri 25913 37448 25929 37464 ne
rect 25929 37448 26006 37464
rect 25746 37349 25894 37431
rect 25634 37316 25711 37332
tri 25711 37316 25727 37332 sw
rect 25634 37250 25727 37316
rect 25763 37191 25877 37349
tri 25913 37316 25929 37332 se
rect 25929 37316 26006 37332
rect 25913 37250 26006 37316
rect 25634 37115 26006 37191
rect 25634 36990 25727 37056
rect 25634 36974 25711 36990
tri 25711 36974 25727 36990 nw
rect 25763 36957 25877 37115
rect 25913 36990 26006 37056
tri 25913 36974 25929 36990 ne
rect 25929 36974 26006 36990
rect 25746 36875 25894 36957
rect 25634 36842 25711 36858
tri 25711 36842 25727 36858 sw
rect 25634 36776 25727 36842
rect 25634 36674 25727 36740
rect 25634 36658 25711 36674
tri 25711 36658 25727 36674 nw
rect 25763 36641 25877 36875
tri 25913 36842 25929 36858 se
rect 25929 36842 26006 36858
rect 25913 36776 26006 36842
rect 25913 36674 26006 36740
tri 25913 36658 25929 36674 ne
rect 25929 36658 26006 36674
rect 25746 36559 25894 36641
rect 25634 36526 25711 36542
tri 25711 36526 25727 36542 sw
rect 25634 36460 25727 36526
rect 25763 36401 25877 36559
tri 25913 36526 25929 36542 se
rect 25929 36526 26006 36542
rect 25913 36460 26006 36526
rect 25634 36325 26006 36401
rect 25634 36200 25727 36266
rect 25634 36184 25711 36200
tri 25711 36184 25727 36200 nw
rect 25763 36167 25877 36325
rect 25913 36200 26006 36266
tri 25913 36184 25929 36200 ne
rect 25929 36184 26006 36200
rect 25746 36085 25894 36167
rect 25634 36052 25711 36068
tri 25711 36052 25727 36068 sw
rect 25634 35986 25727 36052
rect 25634 35884 25727 35950
rect 25634 35868 25711 35884
tri 25711 35868 25727 35884 nw
rect 25763 35851 25877 36085
tri 25913 36052 25929 36068 se
rect 25929 36052 26006 36068
rect 25913 35986 26006 36052
rect 25913 35884 26006 35950
tri 25913 35868 25929 35884 ne
rect 25929 35868 26006 35884
rect 25746 35769 25894 35851
rect 25634 35736 25711 35752
tri 25711 35736 25727 35752 sw
rect 25634 35670 25727 35736
rect 25763 35611 25877 35769
tri 25913 35736 25929 35752 se
rect 25929 35736 26006 35752
rect 25913 35670 26006 35736
rect 25634 35535 26006 35611
rect 25634 35410 25727 35476
rect 25634 35394 25711 35410
tri 25711 35394 25727 35410 nw
rect 25763 35377 25877 35535
rect 25913 35410 26006 35476
tri 25913 35394 25929 35410 ne
rect 25929 35394 26006 35410
rect 25746 35295 25894 35377
rect 25634 35262 25711 35278
tri 25711 35262 25727 35278 sw
rect 25634 35196 25727 35262
rect 25634 35094 25727 35160
rect 25634 35078 25711 35094
tri 25711 35078 25727 35094 nw
rect 25763 35061 25877 35295
tri 25913 35262 25929 35278 se
rect 25929 35262 26006 35278
rect 25913 35196 26006 35262
rect 25913 35094 26006 35160
tri 25913 35078 25929 35094 ne
rect 25929 35078 26006 35094
rect 25746 34979 25894 35061
rect 25634 34946 25711 34962
tri 25711 34946 25727 34962 sw
rect 25634 34880 25727 34946
rect 25763 34821 25877 34979
tri 25913 34946 25929 34962 se
rect 25929 34946 26006 34962
rect 25913 34880 26006 34946
rect 25634 34745 26006 34821
rect 25634 34620 25727 34686
rect 25634 34604 25711 34620
tri 25711 34604 25727 34620 nw
rect 25763 34587 25877 34745
rect 25913 34620 26006 34686
tri 25913 34604 25929 34620 ne
rect 25929 34604 26006 34620
rect 25746 34505 25894 34587
rect 25634 34472 25711 34488
tri 25711 34472 25727 34488 sw
rect 25634 34406 25727 34472
rect 25634 34304 25727 34370
rect 25634 34288 25711 34304
tri 25711 34288 25727 34304 nw
rect 25763 34271 25877 34505
tri 25913 34472 25929 34488 se
rect 25929 34472 26006 34488
rect 25913 34406 26006 34472
rect 25913 34304 26006 34370
tri 25913 34288 25929 34304 ne
rect 25929 34288 26006 34304
rect 25746 34189 25894 34271
rect 25634 34156 25711 34172
tri 25711 34156 25727 34172 sw
rect 25634 34090 25727 34156
rect 25763 34031 25877 34189
tri 25913 34156 25929 34172 se
rect 25929 34156 26006 34172
rect 25913 34090 26006 34156
rect 25634 33955 26006 34031
rect 25634 33830 25727 33896
rect 25634 33814 25711 33830
tri 25711 33814 25727 33830 nw
rect 25763 33797 25877 33955
rect 25913 33830 26006 33896
tri 25913 33814 25929 33830 ne
rect 25929 33814 26006 33830
rect 25746 33715 25894 33797
rect 25634 33682 25711 33698
tri 25711 33682 25727 33698 sw
rect 25634 33616 25727 33682
rect 25634 33514 25727 33580
rect 25634 33498 25711 33514
tri 25711 33498 25727 33514 nw
rect 25763 33481 25877 33715
tri 25913 33682 25929 33698 se
rect 25929 33682 26006 33698
rect 25913 33616 26006 33682
rect 25913 33514 26006 33580
tri 25913 33498 25929 33514 ne
rect 25929 33498 26006 33514
rect 25746 33399 25894 33481
rect 25634 33366 25711 33382
tri 25711 33366 25727 33382 sw
rect 25634 33300 25727 33366
rect 25763 33241 25877 33399
tri 25913 33366 25929 33382 se
rect 25929 33366 26006 33382
rect 25913 33300 26006 33366
rect 25634 33165 26006 33241
rect 25634 33040 25727 33106
rect 25634 33024 25711 33040
tri 25711 33024 25727 33040 nw
rect 25763 33007 25877 33165
rect 25913 33040 26006 33106
tri 25913 33024 25929 33040 ne
rect 25929 33024 26006 33040
rect 25746 32925 25894 33007
rect 25634 32892 25711 32908
tri 25711 32892 25727 32908 sw
rect 25634 32826 25727 32892
rect 25634 32724 25727 32790
rect 25634 32708 25711 32724
tri 25711 32708 25727 32724 nw
rect 25763 32691 25877 32925
tri 25913 32892 25929 32908 se
rect 25929 32892 26006 32908
rect 25913 32826 26006 32892
rect 25913 32724 26006 32790
tri 25913 32708 25929 32724 ne
rect 25929 32708 26006 32724
rect 25746 32609 25894 32691
rect 25634 32576 25711 32592
tri 25711 32576 25727 32592 sw
rect 25634 32510 25727 32576
rect 25763 32451 25877 32609
tri 25913 32576 25929 32592 se
rect 25929 32576 26006 32592
rect 25913 32510 26006 32576
rect 25634 32375 26006 32451
rect 25634 32250 25727 32316
rect 25634 32234 25711 32250
tri 25711 32234 25727 32250 nw
rect 25763 32217 25877 32375
rect 25913 32250 26006 32316
tri 25913 32234 25929 32250 ne
rect 25929 32234 26006 32250
rect 25746 32135 25894 32217
rect 25634 32102 25711 32118
tri 25711 32102 25727 32118 sw
rect 25634 32036 25727 32102
rect 25634 31934 25727 32000
rect 25634 31918 25711 31934
tri 25711 31918 25727 31934 nw
rect 25763 31901 25877 32135
tri 25913 32102 25929 32118 se
rect 25929 32102 26006 32118
rect 25913 32036 26006 32102
rect 25913 31934 26006 32000
tri 25913 31918 25929 31934 ne
rect 25929 31918 26006 31934
rect 25746 31819 25894 31901
rect 25634 31786 25711 31802
tri 25711 31786 25727 31802 sw
rect 25634 31720 25727 31786
rect 25763 31661 25877 31819
tri 25913 31786 25929 31802 se
rect 25929 31786 26006 31802
rect 25913 31720 26006 31786
rect 25634 31585 26006 31661
rect 25634 31460 25727 31526
rect 25634 31444 25711 31460
tri 25711 31444 25727 31460 nw
rect 25763 31427 25877 31585
rect 25913 31460 26006 31526
tri 25913 31444 25929 31460 ne
rect 25929 31444 26006 31460
rect 25746 31345 25894 31427
rect 25634 31312 25711 31328
tri 25711 31312 25727 31328 sw
rect 25634 31246 25727 31312
rect 25634 31144 25727 31210
rect 25634 31128 25711 31144
tri 25711 31128 25727 31144 nw
rect 25763 31111 25877 31345
tri 25913 31312 25929 31328 se
rect 25929 31312 26006 31328
rect 25913 31246 26006 31312
rect 25913 31144 26006 31210
tri 25913 31128 25929 31144 ne
rect 25929 31128 26006 31144
rect 25746 31029 25894 31111
rect 25634 30996 25711 31012
tri 25711 30996 25727 31012 sw
rect 25634 30930 25727 30996
rect 25763 30871 25877 31029
tri 25913 30996 25929 31012 se
rect 25929 30996 26006 31012
rect 25913 30930 26006 30996
rect 25634 30795 26006 30871
rect 25634 30670 25727 30736
rect 25634 30654 25711 30670
tri 25711 30654 25727 30670 nw
rect 25763 30637 25877 30795
rect 25913 30670 26006 30736
tri 25913 30654 25929 30670 ne
rect 25929 30654 26006 30670
rect 25746 30555 25894 30637
rect 25634 30522 25711 30538
tri 25711 30522 25727 30538 sw
rect 25634 30456 25727 30522
rect 25634 30354 25727 30420
rect 25634 30338 25711 30354
tri 25711 30338 25727 30354 nw
rect 25763 30321 25877 30555
tri 25913 30522 25929 30538 se
rect 25929 30522 26006 30538
rect 25913 30456 26006 30522
rect 25913 30354 26006 30420
tri 25913 30338 25929 30354 ne
rect 25929 30338 26006 30354
rect 25746 30239 25894 30321
rect 25634 30206 25711 30222
tri 25711 30206 25727 30222 sw
rect 25634 30140 25727 30206
rect 25763 30081 25877 30239
tri 25913 30206 25929 30222 se
rect 25929 30206 26006 30222
rect 25913 30140 26006 30206
rect 25634 30005 26006 30081
rect 25634 29880 25727 29946
rect 25634 29864 25711 29880
tri 25711 29864 25727 29880 nw
rect 25763 29847 25877 30005
rect 25913 29880 26006 29946
tri 25913 29864 25929 29880 ne
rect 25929 29864 26006 29880
rect 25746 29765 25894 29847
rect 25634 29732 25711 29748
tri 25711 29732 25727 29748 sw
rect 25634 29666 25727 29732
rect 25634 29564 25727 29630
rect 25634 29548 25711 29564
tri 25711 29548 25727 29564 nw
rect 25763 29531 25877 29765
tri 25913 29732 25929 29748 se
rect 25929 29732 26006 29748
rect 25913 29666 26006 29732
rect 25913 29564 26006 29630
tri 25913 29548 25929 29564 ne
rect 25929 29548 26006 29564
rect 25746 29449 25894 29531
rect 25634 29416 25711 29432
tri 25711 29416 25727 29432 sw
rect 25634 29350 25727 29416
rect 25763 29291 25877 29449
tri 25913 29416 25929 29432 se
rect 25929 29416 26006 29432
rect 25913 29350 26006 29416
rect 25634 29215 26006 29291
rect 25634 29090 25727 29156
rect 25634 29074 25711 29090
tri 25711 29074 25727 29090 nw
rect 25763 29057 25877 29215
rect 25913 29090 26006 29156
tri 25913 29074 25929 29090 ne
rect 25929 29074 26006 29090
rect 25746 28975 25894 29057
rect 25634 28942 25711 28958
tri 25711 28942 25727 28958 sw
rect 25634 28876 25727 28942
rect 25763 28833 25877 28975
tri 25913 28942 25929 28958 se
rect 25929 28942 26006 28958
rect 25913 28876 26006 28942
rect 26042 28463 26078 80603
rect 26114 28463 26150 80603
rect 26186 80445 26222 80603
rect 26178 80303 26230 80445
rect 26186 28763 26222 80303
rect 26178 28621 26230 28763
rect 26186 28463 26222 28621
rect 26258 28463 26294 80603
rect 26330 28463 26366 80603
rect 26402 28833 26486 80233
rect 26522 28463 26558 80603
rect 26594 28463 26630 80603
rect 26666 80445 26702 80603
rect 26658 80303 26710 80445
rect 26666 28763 26702 80303
rect 26658 28621 26710 28763
rect 26666 28463 26702 28621
rect 26738 28463 26774 80603
rect 26810 28463 26846 80603
rect 26882 80124 26975 80190
rect 26882 80108 26959 80124
tri 26959 80108 26975 80124 nw
rect 27011 80091 27125 80233
rect 27161 80124 27254 80190
tri 27161 80108 27177 80124 ne
rect 27177 80108 27254 80124
rect 26994 80009 27142 80091
rect 26882 79976 26959 79992
tri 26959 79976 26975 79992 sw
rect 26882 79910 26975 79976
rect 27011 79851 27125 80009
tri 27161 79976 27177 79992 se
rect 27177 79976 27254 79992
rect 27161 79910 27254 79976
rect 26882 79775 27254 79851
rect 26882 79650 26975 79716
rect 26882 79634 26959 79650
tri 26959 79634 26975 79650 nw
rect 27011 79617 27125 79775
rect 27161 79650 27254 79716
tri 27161 79634 27177 79650 ne
rect 27177 79634 27254 79650
rect 26994 79535 27142 79617
rect 26882 79502 26959 79518
tri 26959 79502 26975 79518 sw
rect 26882 79436 26975 79502
rect 26882 79334 26975 79400
rect 26882 79318 26959 79334
tri 26959 79318 26975 79334 nw
rect 27011 79301 27125 79535
tri 27161 79502 27177 79518 se
rect 27177 79502 27254 79518
rect 27161 79436 27254 79502
rect 27161 79334 27254 79400
tri 27161 79318 27177 79334 ne
rect 27177 79318 27254 79334
rect 26994 79219 27142 79301
rect 26882 79186 26959 79202
tri 26959 79186 26975 79202 sw
rect 26882 79120 26975 79186
rect 27011 79061 27125 79219
tri 27161 79186 27177 79202 se
rect 27177 79186 27254 79202
rect 27161 79120 27254 79186
rect 26882 78985 27254 79061
rect 26882 78860 26975 78926
rect 26882 78844 26959 78860
tri 26959 78844 26975 78860 nw
rect 27011 78827 27125 78985
rect 27161 78860 27254 78926
tri 27161 78844 27177 78860 ne
rect 27177 78844 27254 78860
rect 26994 78745 27142 78827
rect 26882 78712 26959 78728
tri 26959 78712 26975 78728 sw
rect 26882 78646 26975 78712
rect 26882 78544 26975 78610
rect 26882 78528 26959 78544
tri 26959 78528 26975 78544 nw
rect 27011 78511 27125 78745
tri 27161 78712 27177 78728 se
rect 27177 78712 27254 78728
rect 27161 78646 27254 78712
rect 27161 78544 27254 78610
tri 27161 78528 27177 78544 ne
rect 27177 78528 27254 78544
rect 26994 78429 27142 78511
rect 26882 78396 26959 78412
tri 26959 78396 26975 78412 sw
rect 26882 78330 26975 78396
rect 27011 78271 27125 78429
tri 27161 78396 27177 78412 se
rect 27177 78396 27254 78412
rect 27161 78330 27254 78396
rect 26882 78195 27254 78271
rect 26882 78070 26975 78136
rect 26882 78054 26959 78070
tri 26959 78054 26975 78070 nw
rect 27011 78037 27125 78195
rect 27161 78070 27254 78136
tri 27161 78054 27177 78070 ne
rect 27177 78054 27254 78070
rect 26994 77955 27142 78037
rect 26882 77922 26959 77938
tri 26959 77922 26975 77938 sw
rect 26882 77856 26975 77922
rect 26882 77754 26975 77820
rect 26882 77738 26959 77754
tri 26959 77738 26975 77754 nw
rect 27011 77721 27125 77955
tri 27161 77922 27177 77938 se
rect 27177 77922 27254 77938
rect 27161 77856 27254 77922
rect 27161 77754 27254 77820
tri 27161 77738 27177 77754 ne
rect 27177 77738 27254 77754
rect 26994 77639 27142 77721
rect 26882 77606 26959 77622
tri 26959 77606 26975 77622 sw
rect 26882 77540 26975 77606
rect 27011 77481 27125 77639
tri 27161 77606 27177 77622 se
rect 27177 77606 27254 77622
rect 27161 77540 27254 77606
rect 26882 77405 27254 77481
rect 26882 77280 26975 77346
rect 26882 77264 26959 77280
tri 26959 77264 26975 77280 nw
rect 27011 77247 27125 77405
rect 27161 77280 27254 77346
tri 27161 77264 27177 77280 ne
rect 27177 77264 27254 77280
rect 26994 77165 27142 77247
rect 26882 77132 26959 77148
tri 26959 77132 26975 77148 sw
rect 26882 77066 26975 77132
rect 26882 76964 26975 77030
rect 26882 76948 26959 76964
tri 26959 76948 26975 76964 nw
rect 27011 76931 27125 77165
tri 27161 77132 27177 77148 se
rect 27177 77132 27254 77148
rect 27161 77066 27254 77132
rect 27161 76964 27254 77030
tri 27161 76948 27177 76964 ne
rect 27177 76948 27254 76964
rect 26994 76849 27142 76931
rect 26882 76816 26959 76832
tri 26959 76816 26975 76832 sw
rect 26882 76750 26975 76816
rect 27011 76691 27125 76849
tri 27161 76816 27177 76832 se
rect 27177 76816 27254 76832
rect 27161 76750 27254 76816
rect 26882 76615 27254 76691
rect 26882 76490 26975 76556
rect 26882 76474 26959 76490
tri 26959 76474 26975 76490 nw
rect 27011 76457 27125 76615
rect 27161 76490 27254 76556
tri 27161 76474 27177 76490 ne
rect 27177 76474 27254 76490
rect 26994 76375 27142 76457
rect 26882 76342 26959 76358
tri 26959 76342 26975 76358 sw
rect 26882 76276 26975 76342
rect 26882 76174 26975 76240
rect 26882 76158 26959 76174
tri 26959 76158 26975 76174 nw
rect 27011 76141 27125 76375
tri 27161 76342 27177 76358 se
rect 27177 76342 27254 76358
rect 27161 76276 27254 76342
rect 27161 76174 27254 76240
tri 27161 76158 27177 76174 ne
rect 27177 76158 27254 76174
rect 26994 76059 27142 76141
rect 26882 76026 26959 76042
tri 26959 76026 26975 76042 sw
rect 26882 75960 26975 76026
rect 27011 75901 27125 76059
tri 27161 76026 27177 76042 se
rect 27177 76026 27254 76042
rect 27161 75960 27254 76026
rect 26882 75825 27254 75901
rect 26882 75700 26975 75766
rect 26882 75684 26959 75700
tri 26959 75684 26975 75700 nw
rect 27011 75667 27125 75825
rect 27161 75700 27254 75766
tri 27161 75684 27177 75700 ne
rect 27177 75684 27254 75700
rect 26994 75585 27142 75667
rect 26882 75552 26959 75568
tri 26959 75552 26975 75568 sw
rect 26882 75486 26975 75552
rect 26882 75384 26975 75450
rect 26882 75368 26959 75384
tri 26959 75368 26975 75384 nw
rect 27011 75351 27125 75585
tri 27161 75552 27177 75568 se
rect 27177 75552 27254 75568
rect 27161 75486 27254 75552
rect 27161 75384 27254 75450
tri 27161 75368 27177 75384 ne
rect 27177 75368 27254 75384
rect 26994 75269 27142 75351
rect 26882 75236 26959 75252
tri 26959 75236 26975 75252 sw
rect 26882 75170 26975 75236
rect 27011 75111 27125 75269
tri 27161 75236 27177 75252 se
rect 27177 75236 27254 75252
rect 27161 75170 27254 75236
rect 26882 75035 27254 75111
rect 26882 74910 26975 74976
rect 26882 74894 26959 74910
tri 26959 74894 26975 74910 nw
rect 27011 74877 27125 75035
rect 27161 74910 27254 74976
tri 27161 74894 27177 74910 ne
rect 27177 74894 27254 74910
rect 26994 74795 27142 74877
rect 26882 74762 26959 74778
tri 26959 74762 26975 74778 sw
rect 26882 74696 26975 74762
rect 26882 74594 26975 74660
rect 26882 74578 26959 74594
tri 26959 74578 26975 74594 nw
rect 27011 74561 27125 74795
tri 27161 74762 27177 74778 se
rect 27177 74762 27254 74778
rect 27161 74696 27254 74762
rect 27161 74594 27254 74660
tri 27161 74578 27177 74594 ne
rect 27177 74578 27254 74594
rect 26994 74479 27142 74561
rect 26882 74446 26959 74462
tri 26959 74446 26975 74462 sw
rect 26882 74380 26975 74446
rect 27011 74321 27125 74479
tri 27161 74446 27177 74462 se
rect 27177 74446 27254 74462
rect 27161 74380 27254 74446
rect 26882 74245 27254 74321
rect 26882 74120 26975 74186
rect 26882 74104 26959 74120
tri 26959 74104 26975 74120 nw
rect 27011 74087 27125 74245
rect 27161 74120 27254 74186
tri 27161 74104 27177 74120 ne
rect 27177 74104 27254 74120
rect 26994 74005 27142 74087
rect 26882 73972 26959 73988
tri 26959 73972 26975 73988 sw
rect 26882 73906 26975 73972
rect 26882 73804 26975 73870
rect 26882 73788 26959 73804
tri 26959 73788 26975 73804 nw
rect 27011 73771 27125 74005
tri 27161 73972 27177 73988 se
rect 27177 73972 27254 73988
rect 27161 73906 27254 73972
rect 27161 73804 27254 73870
tri 27161 73788 27177 73804 ne
rect 27177 73788 27254 73804
rect 26994 73689 27142 73771
rect 26882 73656 26959 73672
tri 26959 73656 26975 73672 sw
rect 26882 73590 26975 73656
rect 27011 73531 27125 73689
tri 27161 73656 27177 73672 se
rect 27177 73656 27254 73672
rect 27161 73590 27254 73656
rect 26882 73455 27254 73531
rect 26882 73330 26975 73396
rect 26882 73314 26959 73330
tri 26959 73314 26975 73330 nw
rect 27011 73297 27125 73455
rect 27161 73330 27254 73396
tri 27161 73314 27177 73330 ne
rect 27177 73314 27254 73330
rect 26994 73215 27142 73297
rect 26882 73182 26959 73198
tri 26959 73182 26975 73198 sw
rect 26882 73116 26975 73182
rect 26882 73014 26975 73080
rect 26882 72998 26959 73014
tri 26959 72998 26975 73014 nw
rect 27011 72981 27125 73215
tri 27161 73182 27177 73198 se
rect 27177 73182 27254 73198
rect 27161 73116 27254 73182
rect 27161 73014 27254 73080
tri 27161 72998 27177 73014 ne
rect 27177 72998 27254 73014
rect 26994 72899 27142 72981
rect 26882 72866 26959 72882
tri 26959 72866 26975 72882 sw
rect 26882 72800 26975 72866
rect 27011 72741 27125 72899
tri 27161 72866 27177 72882 se
rect 27177 72866 27254 72882
rect 27161 72800 27254 72866
rect 26882 72665 27254 72741
rect 26882 72540 26975 72606
rect 26882 72524 26959 72540
tri 26959 72524 26975 72540 nw
rect 27011 72507 27125 72665
rect 27161 72540 27254 72606
tri 27161 72524 27177 72540 ne
rect 27177 72524 27254 72540
rect 26994 72425 27142 72507
rect 26882 72392 26959 72408
tri 26959 72392 26975 72408 sw
rect 26882 72326 26975 72392
rect 26882 72224 26975 72290
rect 26882 72208 26959 72224
tri 26959 72208 26975 72224 nw
rect 27011 72191 27125 72425
tri 27161 72392 27177 72408 se
rect 27177 72392 27254 72408
rect 27161 72326 27254 72392
rect 27161 72224 27254 72290
tri 27161 72208 27177 72224 ne
rect 27177 72208 27254 72224
rect 26994 72109 27142 72191
rect 26882 72076 26959 72092
tri 26959 72076 26975 72092 sw
rect 26882 72010 26975 72076
rect 27011 71951 27125 72109
tri 27161 72076 27177 72092 se
rect 27177 72076 27254 72092
rect 27161 72010 27254 72076
rect 26882 71875 27254 71951
rect 26882 71750 26975 71816
rect 26882 71734 26959 71750
tri 26959 71734 26975 71750 nw
rect 27011 71717 27125 71875
rect 27161 71750 27254 71816
tri 27161 71734 27177 71750 ne
rect 27177 71734 27254 71750
rect 26994 71635 27142 71717
rect 26882 71602 26959 71618
tri 26959 71602 26975 71618 sw
rect 26882 71536 26975 71602
rect 26882 71434 26975 71500
rect 26882 71418 26959 71434
tri 26959 71418 26975 71434 nw
rect 27011 71401 27125 71635
tri 27161 71602 27177 71618 se
rect 27177 71602 27254 71618
rect 27161 71536 27254 71602
rect 27161 71434 27254 71500
tri 27161 71418 27177 71434 ne
rect 27177 71418 27254 71434
rect 26994 71319 27142 71401
rect 26882 71286 26959 71302
tri 26959 71286 26975 71302 sw
rect 26882 71220 26975 71286
rect 27011 71161 27125 71319
tri 27161 71286 27177 71302 se
rect 27177 71286 27254 71302
rect 27161 71220 27254 71286
rect 26882 71085 27254 71161
rect 26882 70960 26975 71026
rect 26882 70944 26959 70960
tri 26959 70944 26975 70960 nw
rect 27011 70927 27125 71085
rect 27161 70960 27254 71026
tri 27161 70944 27177 70960 ne
rect 27177 70944 27254 70960
rect 26994 70845 27142 70927
rect 26882 70812 26959 70828
tri 26959 70812 26975 70828 sw
rect 26882 70746 26975 70812
rect 26882 70644 26975 70710
rect 26882 70628 26959 70644
tri 26959 70628 26975 70644 nw
rect 27011 70611 27125 70845
tri 27161 70812 27177 70828 se
rect 27177 70812 27254 70828
rect 27161 70746 27254 70812
rect 27161 70644 27254 70710
tri 27161 70628 27177 70644 ne
rect 27177 70628 27254 70644
rect 26994 70529 27142 70611
rect 26882 70496 26959 70512
tri 26959 70496 26975 70512 sw
rect 26882 70430 26975 70496
rect 27011 70371 27125 70529
tri 27161 70496 27177 70512 se
rect 27177 70496 27254 70512
rect 27161 70430 27254 70496
rect 26882 70295 27254 70371
rect 26882 70170 26975 70236
rect 26882 70154 26959 70170
tri 26959 70154 26975 70170 nw
rect 27011 70137 27125 70295
rect 27161 70170 27254 70236
tri 27161 70154 27177 70170 ne
rect 27177 70154 27254 70170
rect 26994 70055 27142 70137
rect 26882 70022 26959 70038
tri 26959 70022 26975 70038 sw
rect 26882 69956 26975 70022
rect 26882 69854 26975 69920
rect 26882 69838 26959 69854
tri 26959 69838 26975 69854 nw
rect 27011 69821 27125 70055
tri 27161 70022 27177 70038 se
rect 27177 70022 27254 70038
rect 27161 69956 27254 70022
rect 27161 69854 27254 69920
tri 27161 69838 27177 69854 ne
rect 27177 69838 27254 69854
rect 26994 69739 27142 69821
rect 26882 69706 26959 69722
tri 26959 69706 26975 69722 sw
rect 26882 69640 26975 69706
rect 27011 69581 27125 69739
tri 27161 69706 27177 69722 se
rect 27177 69706 27254 69722
rect 27161 69640 27254 69706
rect 26882 69505 27254 69581
rect 26882 69380 26975 69446
rect 26882 69364 26959 69380
tri 26959 69364 26975 69380 nw
rect 27011 69347 27125 69505
rect 27161 69380 27254 69446
tri 27161 69364 27177 69380 ne
rect 27177 69364 27254 69380
rect 26994 69265 27142 69347
rect 26882 69232 26959 69248
tri 26959 69232 26975 69248 sw
rect 26882 69166 26975 69232
rect 26882 69064 26975 69130
rect 26882 69048 26959 69064
tri 26959 69048 26975 69064 nw
rect 27011 69031 27125 69265
tri 27161 69232 27177 69248 se
rect 27177 69232 27254 69248
rect 27161 69166 27254 69232
rect 27161 69064 27254 69130
tri 27161 69048 27177 69064 ne
rect 27177 69048 27254 69064
rect 26994 68949 27142 69031
rect 26882 68916 26959 68932
tri 26959 68916 26975 68932 sw
rect 26882 68850 26975 68916
rect 27011 68791 27125 68949
tri 27161 68916 27177 68932 se
rect 27177 68916 27254 68932
rect 27161 68850 27254 68916
rect 26882 68715 27254 68791
rect 26882 68590 26975 68656
rect 26882 68574 26959 68590
tri 26959 68574 26975 68590 nw
rect 27011 68557 27125 68715
rect 27161 68590 27254 68656
tri 27161 68574 27177 68590 ne
rect 27177 68574 27254 68590
rect 26994 68475 27142 68557
rect 26882 68442 26959 68458
tri 26959 68442 26975 68458 sw
rect 26882 68376 26975 68442
rect 26882 68274 26975 68340
rect 26882 68258 26959 68274
tri 26959 68258 26975 68274 nw
rect 27011 68241 27125 68475
tri 27161 68442 27177 68458 se
rect 27177 68442 27254 68458
rect 27161 68376 27254 68442
rect 27161 68274 27254 68340
tri 27161 68258 27177 68274 ne
rect 27177 68258 27254 68274
rect 26994 68159 27142 68241
rect 26882 68126 26959 68142
tri 26959 68126 26975 68142 sw
rect 26882 68060 26975 68126
rect 27011 68001 27125 68159
tri 27161 68126 27177 68142 se
rect 27177 68126 27254 68142
rect 27161 68060 27254 68126
rect 26882 67925 27254 68001
rect 26882 67800 26975 67866
rect 26882 67784 26959 67800
tri 26959 67784 26975 67800 nw
rect 27011 67767 27125 67925
rect 27161 67800 27254 67866
tri 27161 67784 27177 67800 ne
rect 27177 67784 27254 67800
rect 26994 67685 27142 67767
rect 26882 67652 26959 67668
tri 26959 67652 26975 67668 sw
rect 26882 67586 26975 67652
rect 26882 67484 26975 67550
rect 26882 67468 26959 67484
tri 26959 67468 26975 67484 nw
rect 27011 67451 27125 67685
tri 27161 67652 27177 67668 se
rect 27177 67652 27254 67668
rect 27161 67586 27254 67652
rect 27161 67484 27254 67550
tri 27161 67468 27177 67484 ne
rect 27177 67468 27254 67484
rect 26994 67369 27142 67451
rect 26882 67336 26959 67352
tri 26959 67336 26975 67352 sw
rect 26882 67270 26975 67336
rect 27011 67211 27125 67369
tri 27161 67336 27177 67352 se
rect 27177 67336 27254 67352
rect 27161 67270 27254 67336
rect 26882 67135 27254 67211
rect 26882 67010 26975 67076
rect 26882 66994 26959 67010
tri 26959 66994 26975 67010 nw
rect 27011 66977 27125 67135
rect 27161 67010 27254 67076
tri 27161 66994 27177 67010 ne
rect 27177 66994 27254 67010
rect 26994 66895 27142 66977
rect 26882 66862 26959 66878
tri 26959 66862 26975 66878 sw
rect 26882 66796 26975 66862
rect 26882 66694 26975 66760
rect 26882 66678 26959 66694
tri 26959 66678 26975 66694 nw
rect 27011 66661 27125 66895
tri 27161 66862 27177 66878 se
rect 27177 66862 27254 66878
rect 27161 66796 27254 66862
rect 27161 66694 27254 66760
tri 27161 66678 27177 66694 ne
rect 27177 66678 27254 66694
rect 26994 66579 27142 66661
rect 26882 66546 26959 66562
tri 26959 66546 26975 66562 sw
rect 26882 66480 26975 66546
rect 27011 66421 27125 66579
tri 27161 66546 27177 66562 se
rect 27177 66546 27254 66562
rect 27161 66480 27254 66546
rect 26882 66345 27254 66421
rect 26882 66220 26975 66286
rect 26882 66204 26959 66220
tri 26959 66204 26975 66220 nw
rect 27011 66187 27125 66345
rect 27161 66220 27254 66286
tri 27161 66204 27177 66220 ne
rect 27177 66204 27254 66220
rect 26994 66105 27142 66187
rect 26882 66072 26959 66088
tri 26959 66072 26975 66088 sw
rect 26882 66006 26975 66072
rect 26882 65904 26975 65970
rect 26882 65888 26959 65904
tri 26959 65888 26975 65904 nw
rect 27011 65871 27125 66105
tri 27161 66072 27177 66088 se
rect 27177 66072 27254 66088
rect 27161 66006 27254 66072
rect 27161 65904 27254 65970
tri 27161 65888 27177 65904 ne
rect 27177 65888 27254 65904
rect 26994 65789 27142 65871
rect 26882 65756 26959 65772
tri 26959 65756 26975 65772 sw
rect 26882 65690 26975 65756
rect 27011 65631 27125 65789
tri 27161 65756 27177 65772 se
rect 27177 65756 27254 65772
rect 27161 65690 27254 65756
rect 26882 65555 27254 65631
rect 26882 65430 26975 65496
rect 26882 65414 26959 65430
tri 26959 65414 26975 65430 nw
rect 27011 65397 27125 65555
rect 27161 65430 27254 65496
tri 27161 65414 27177 65430 ne
rect 27177 65414 27254 65430
rect 26994 65315 27142 65397
rect 26882 65282 26959 65298
tri 26959 65282 26975 65298 sw
rect 26882 65216 26975 65282
rect 26882 65114 26975 65180
rect 26882 65098 26959 65114
tri 26959 65098 26975 65114 nw
rect 27011 65081 27125 65315
tri 27161 65282 27177 65298 se
rect 27177 65282 27254 65298
rect 27161 65216 27254 65282
rect 27161 65114 27254 65180
tri 27161 65098 27177 65114 ne
rect 27177 65098 27254 65114
rect 26994 64999 27142 65081
rect 26882 64966 26959 64982
tri 26959 64966 26975 64982 sw
rect 26882 64900 26975 64966
rect 27011 64841 27125 64999
tri 27161 64966 27177 64982 se
rect 27177 64966 27254 64982
rect 27161 64900 27254 64966
rect 26882 64765 27254 64841
rect 26882 64640 26975 64706
rect 26882 64624 26959 64640
tri 26959 64624 26975 64640 nw
rect 27011 64607 27125 64765
rect 27161 64640 27254 64706
tri 27161 64624 27177 64640 ne
rect 27177 64624 27254 64640
rect 26994 64525 27142 64607
rect 26882 64492 26959 64508
tri 26959 64492 26975 64508 sw
rect 26882 64426 26975 64492
rect 26882 64324 26975 64390
rect 26882 64308 26959 64324
tri 26959 64308 26975 64324 nw
rect 27011 64291 27125 64525
tri 27161 64492 27177 64508 se
rect 27177 64492 27254 64508
rect 27161 64426 27254 64492
rect 27161 64324 27254 64390
tri 27161 64308 27177 64324 ne
rect 27177 64308 27254 64324
rect 26994 64209 27142 64291
rect 26882 64176 26959 64192
tri 26959 64176 26975 64192 sw
rect 26882 64110 26975 64176
rect 27011 64051 27125 64209
tri 27161 64176 27177 64192 se
rect 27177 64176 27254 64192
rect 27161 64110 27254 64176
rect 26882 63975 27254 64051
rect 26882 63850 26975 63916
rect 26882 63834 26959 63850
tri 26959 63834 26975 63850 nw
rect 27011 63817 27125 63975
rect 27161 63850 27254 63916
tri 27161 63834 27177 63850 ne
rect 27177 63834 27254 63850
rect 26994 63735 27142 63817
rect 26882 63702 26959 63718
tri 26959 63702 26975 63718 sw
rect 26882 63636 26975 63702
rect 26882 63534 26975 63600
rect 26882 63518 26959 63534
tri 26959 63518 26975 63534 nw
rect 27011 63501 27125 63735
tri 27161 63702 27177 63718 se
rect 27177 63702 27254 63718
rect 27161 63636 27254 63702
rect 27161 63534 27254 63600
tri 27161 63518 27177 63534 ne
rect 27177 63518 27254 63534
rect 26994 63419 27142 63501
rect 26882 63386 26959 63402
tri 26959 63386 26975 63402 sw
rect 26882 63320 26975 63386
rect 27011 63261 27125 63419
tri 27161 63386 27177 63402 se
rect 27177 63386 27254 63402
rect 27161 63320 27254 63386
rect 26882 63185 27254 63261
rect 26882 63060 26975 63126
rect 26882 63044 26959 63060
tri 26959 63044 26975 63060 nw
rect 27011 63027 27125 63185
rect 27161 63060 27254 63126
tri 27161 63044 27177 63060 ne
rect 27177 63044 27254 63060
rect 26994 62945 27142 63027
rect 26882 62912 26959 62928
tri 26959 62912 26975 62928 sw
rect 26882 62846 26975 62912
rect 26882 62744 26975 62810
rect 26882 62728 26959 62744
tri 26959 62728 26975 62744 nw
rect 27011 62711 27125 62945
tri 27161 62912 27177 62928 se
rect 27177 62912 27254 62928
rect 27161 62846 27254 62912
rect 27161 62744 27254 62810
tri 27161 62728 27177 62744 ne
rect 27177 62728 27254 62744
rect 26994 62629 27142 62711
rect 26882 62596 26959 62612
tri 26959 62596 26975 62612 sw
rect 26882 62530 26975 62596
rect 27011 62471 27125 62629
tri 27161 62596 27177 62612 se
rect 27177 62596 27254 62612
rect 27161 62530 27254 62596
rect 26882 62395 27254 62471
rect 26882 62270 26975 62336
rect 26882 62254 26959 62270
tri 26959 62254 26975 62270 nw
rect 27011 62237 27125 62395
rect 27161 62270 27254 62336
tri 27161 62254 27177 62270 ne
rect 27177 62254 27254 62270
rect 26994 62155 27142 62237
rect 26882 62122 26959 62138
tri 26959 62122 26975 62138 sw
rect 26882 62056 26975 62122
rect 26882 61954 26975 62020
rect 26882 61938 26959 61954
tri 26959 61938 26975 61954 nw
rect 27011 61921 27125 62155
tri 27161 62122 27177 62138 se
rect 27177 62122 27254 62138
rect 27161 62056 27254 62122
rect 27161 61954 27254 62020
tri 27161 61938 27177 61954 ne
rect 27177 61938 27254 61954
rect 26994 61839 27142 61921
rect 26882 61806 26959 61822
tri 26959 61806 26975 61822 sw
rect 26882 61740 26975 61806
rect 27011 61681 27125 61839
tri 27161 61806 27177 61822 se
rect 27177 61806 27254 61822
rect 27161 61740 27254 61806
rect 26882 61605 27254 61681
rect 26882 61480 26975 61546
rect 26882 61464 26959 61480
tri 26959 61464 26975 61480 nw
rect 27011 61447 27125 61605
rect 27161 61480 27254 61546
tri 27161 61464 27177 61480 ne
rect 27177 61464 27254 61480
rect 26994 61365 27142 61447
rect 26882 61332 26959 61348
tri 26959 61332 26975 61348 sw
rect 26882 61266 26975 61332
rect 26882 61164 26975 61230
rect 26882 61148 26959 61164
tri 26959 61148 26975 61164 nw
rect 27011 61131 27125 61365
tri 27161 61332 27177 61348 se
rect 27177 61332 27254 61348
rect 27161 61266 27254 61332
rect 27161 61164 27254 61230
tri 27161 61148 27177 61164 ne
rect 27177 61148 27254 61164
rect 26994 61049 27142 61131
rect 26882 61016 26959 61032
tri 26959 61016 26975 61032 sw
rect 26882 60950 26975 61016
rect 27011 60891 27125 61049
tri 27161 61016 27177 61032 se
rect 27177 61016 27254 61032
rect 27161 60950 27254 61016
rect 26882 60815 27254 60891
rect 26882 60690 26975 60756
rect 26882 60674 26959 60690
tri 26959 60674 26975 60690 nw
rect 27011 60657 27125 60815
rect 27161 60690 27254 60756
tri 27161 60674 27177 60690 ne
rect 27177 60674 27254 60690
rect 26994 60575 27142 60657
rect 26882 60542 26959 60558
tri 26959 60542 26975 60558 sw
rect 26882 60476 26975 60542
rect 26882 60374 26975 60440
rect 26882 60358 26959 60374
tri 26959 60358 26975 60374 nw
rect 27011 60341 27125 60575
tri 27161 60542 27177 60558 se
rect 27177 60542 27254 60558
rect 27161 60476 27254 60542
rect 27161 60374 27254 60440
tri 27161 60358 27177 60374 ne
rect 27177 60358 27254 60374
rect 26994 60259 27142 60341
rect 26882 60226 26959 60242
tri 26959 60226 26975 60242 sw
rect 26882 60160 26975 60226
rect 27011 60101 27125 60259
tri 27161 60226 27177 60242 se
rect 27177 60226 27254 60242
rect 27161 60160 27254 60226
rect 26882 60025 27254 60101
rect 26882 59900 26975 59966
rect 26882 59884 26959 59900
tri 26959 59884 26975 59900 nw
rect 27011 59867 27125 60025
rect 27161 59900 27254 59966
tri 27161 59884 27177 59900 ne
rect 27177 59884 27254 59900
rect 26994 59785 27142 59867
rect 26882 59752 26959 59768
tri 26959 59752 26975 59768 sw
rect 26882 59686 26975 59752
rect 26882 59584 26975 59650
rect 26882 59568 26959 59584
tri 26959 59568 26975 59584 nw
rect 27011 59551 27125 59785
tri 27161 59752 27177 59768 se
rect 27177 59752 27254 59768
rect 27161 59686 27254 59752
rect 27161 59584 27254 59650
tri 27161 59568 27177 59584 ne
rect 27177 59568 27254 59584
rect 26994 59469 27142 59551
rect 26882 59436 26959 59452
tri 26959 59436 26975 59452 sw
rect 26882 59370 26975 59436
rect 27011 59311 27125 59469
tri 27161 59436 27177 59452 se
rect 27177 59436 27254 59452
rect 27161 59370 27254 59436
rect 26882 59235 27254 59311
rect 26882 59110 26975 59176
rect 26882 59094 26959 59110
tri 26959 59094 26975 59110 nw
rect 27011 59077 27125 59235
rect 27161 59110 27254 59176
tri 27161 59094 27177 59110 ne
rect 27177 59094 27254 59110
rect 26994 58995 27142 59077
rect 26882 58962 26959 58978
tri 26959 58962 26975 58978 sw
rect 26882 58896 26975 58962
rect 26882 58794 26975 58860
rect 26882 58778 26959 58794
tri 26959 58778 26975 58794 nw
rect 27011 58761 27125 58995
tri 27161 58962 27177 58978 se
rect 27177 58962 27254 58978
rect 27161 58896 27254 58962
rect 27161 58794 27254 58860
tri 27161 58778 27177 58794 ne
rect 27177 58778 27254 58794
rect 26994 58679 27142 58761
rect 26882 58646 26959 58662
tri 26959 58646 26975 58662 sw
rect 26882 58580 26975 58646
rect 27011 58521 27125 58679
tri 27161 58646 27177 58662 se
rect 27177 58646 27254 58662
rect 27161 58580 27254 58646
rect 26882 58445 27254 58521
rect 26882 58320 26975 58386
rect 26882 58304 26959 58320
tri 26959 58304 26975 58320 nw
rect 27011 58287 27125 58445
rect 27161 58320 27254 58386
tri 27161 58304 27177 58320 ne
rect 27177 58304 27254 58320
rect 26994 58205 27142 58287
rect 26882 58172 26959 58188
tri 26959 58172 26975 58188 sw
rect 26882 58106 26975 58172
rect 26882 58004 26975 58070
rect 26882 57988 26959 58004
tri 26959 57988 26975 58004 nw
rect 27011 57971 27125 58205
tri 27161 58172 27177 58188 se
rect 27177 58172 27254 58188
rect 27161 58106 27254 58172
rect 27161 58004 27254 58070
tri 27161 57988 27177 58004 ne
rect 27177 57988 27254 58004
rect 26994 57889 27142 57971
rect 26882 57856 26959 57872
tri 26959 57856 26975 57872 sw
rect 26882 57790 26975 57856
rect 27011 57731 27125 57889
tri 27161 57856 27177 57872 se
rect 27177 57856 27254 57872
rect 27161 57790 27254 57856
rect 26882 57655 27254 57731
rect 26882 57530 26975 57596
rect 26882 57514 26959 57530
tri 26959 57514 26975 57530 nw
rect 27011 57497 27125 57655
rect 27161 57530 27254 57596
tri 27161 57514 27177 57530 ne
rect 27177 57514 27254 57530
rect 26994 57415 27142 57497
rect 26882 57382 26959 57398
tri 26959 57382 26975 57398 sw
rect 26882 57316 26975 57382
rect 26882 57214 26975 57280
rect 26882 57198 26959 57214
tri 26959 57198 26975 57214 nw
rect 27011 57181 27125 57415
tri 27161 57382 27177 57398 se
rect 27177 57382 27254 57398
rect 27161 57316 27254 57382
rect 27161 57214 27254 57280
tri 27161 57198 27177 57214 ne
rect 27177 57198 27254 57214
rect 26994 57099 27142 57181
rect 26882 57066 26959 57082
tri 26959 57066 26975 57082 sw
rect 26882 57000 26975 57066
rect 27011 56941 27125 57099
tri 27161 57066 27177 57082 se
rect 27177 57066 27254 57082
rect 27161 57000 27254 57066
rect 26882 56865 27254 56941
rect 26882 56740 26975 56806
rect 26882 56724 26959 56740
tri 26959 56724 26975 56740 nw
rect 27011 56707 27125 56865
rect 27161 56740 27254 56806
tri 27161 56724 27177 56740 ne
rect 27177 56724 27254 56740
rect 26994 56625 27142 56707
rect 26882 56592 26959 56608
tri 26959 56592 26975 56608 sw
rect 26882 56526 26975 56592
rect 26882 56424 26975 56490
rect 26882 56408 26959 56424
tri 26959 56408 26975 56424 nw
rect 27011 56391 27125 56625
tri 27161 56592 27177 56608 se
rect 27177 56592 27254 56608
rect 27161 56526 27254 56592
rect 27161 56424 27254 56490
tri 27161 56408 27177 56424 ne
rect 27177 56408 27254 56424
rect 26994 56309 27142 56391
rect 26882 56276 26959 56292
tri 26959 56276 26975 56292 sw
rect 26882 56210 26975 56276
rect 27011 56151 27125 56309
tri 27161 56276 27177 56292 se
rect 27177 56276 27254 56292
rect 27161 56210 27254 56276
rect 26882 56075 27254 56151
rect 26882 55950 26975 56016
rect 26882 55934 26959 55950
tri 26959 55934 26975 55950 nw
rect 27011 55917 27125 56075
rect 27161 55950 27254 56016
tri 27161 55934 27177 55950 ne
rect 27177 55934 27254 55950
rect 26994 55835 27142 55917
rect 26882 55802 26959 55818
tri 26959 55802 26975 55818 sw
rect 26882 55736 26975 55802
rect 26882 55634 26975 55700
rect 26882 55618 26959 55634
tri 26959 55618 26975 55634 nw
rect 27011 55601 27125 55835
tri 27161 55802 27177 55818 se
rect 27177 55802 27254 55818
rect 27161 55736 27254 55802
rect 27161 55634 27254 55700
tri 27161 55618 27177 55634 ne
rect 27177 55618 27254 55634
rect 26994 55519 27142 55601
rect 26882 55486 26959 55502
tri 26959 55486 26975 55502 sw
rect 26882 55420 26975 55486
rect 27011 55361 27125 55519
tri 27161 55486 27177 55502 se
rect 27177 55486 27254 55502
rect 27161 55420 27254 55486
rect 26882 55285 27254 55361
rect 26882 55160 26975 55226
rect 26882 55144 26959 55160
tri 26959 55144 26975 55160 nw
rect 27011 55127 27125 55285
rect 27161 55160 27254 55226
tri 27161 55144 27177 55160 ne
rect 27177 55144 27254 55160
rect 26994 55045 27142 55127
rect 26882 55012 26959 55028
tri 26959 55012 26975 55028 sw
rect 26882 54946 26975 55012
rect 26882 54844 26975 54910
rect 26882 54828 26959 54844
tri 26959 54828 26975 54844 nw
rect 27011 54811 27125 55045
tri 27161 55012 27177 55028 se
rect 27177 55012 27254 55028
rect 27161 54946 27254 55012
rect 27161 54844 27254 54910
tri 27161 54828 27177 54844 ne
rect 27177 54828 27254 54844
rect 26994 54729 27142 54811
rect 26882 54696 26959 54712
tri 26959 54696 26975 54712 sw
rect 26882 54630 26975 54696
rect 27011 54571 27125 54729
tri 27161 54696 27177 54712 se
rect 27177 54696 27254 54712
rect 27161 54630 27254 54696
rect 26882 54495 27254 54571
rect 26882 54370 26975 54436
rect 26882 54354 26959 54370
tri 26959 54354 26975 54370 nw
rect 27011 54337 27125 54495
rect 27161 54370 27254 54436
tri 27161 54354 27177 54370 ne
rect 27177 54354 27254 54370
rect 26994 54255 27142 54337
rect 26882 54222 26959 54238
tri 26959 54222 26975 54238 sw
rect 26882 54156 26975 54222
rect 26882 54054 26975 54120
rect 26882 54038 26959 54054
tri 26959 54038 26975 54054 nw
rect 27011 54021 27125 54255
tri 27161 54222 27177 54238 se
rect 27177 54222 27254 54238
rect 27161 54156 27254 54222
rect 27161 54054 27254 54120
tri 27161 54038 27177 54054 ne
rect 27177 54038 27254 54054
rect 26994 53939 27142 54021
rect 26882 53906 26959 53922
tri 26959 53906 26975 53922 sw
rect 26882 53840 26975 53906
rect 27011 53781 27125 53939
tri 27161 53906 27177 53922 se
rect 27177 53906 27254 53922
rect 27161 53840 27254 53906
rect 26882 53705 27254 53781
rect 26882 53580 26975 53646
rect 26882 53564 26959 53580
tri 26959 53564 26975 53580 nw
rect 27011 53547 27125 53705
rect 27161 53580 27254 53646
tri 27161 53564 27177 53580 ne
rect 27177 53564 27254 53580
rect 26994 53465 27142 53547
rect 26882 53432 26959 53448
tri 26959 53432 26975 53448 sw
rect 26882 53366 26975 53432
rect 26882 53264 26975 53330
rect 26882 53248 26959 53264
tri 26959 53248 26975 53264 nw
rect 27011 53231 27125 53465
tri 27161 53432 27177 53448 se
rect 27177 53432 27254 53448
rect 27161 53366 27254 53432
rect 27161 53264 27254 53330
tri 27161 53248 27177 53264 ne
rect 27177 53248 27254 53264
rect 26994 53149 27142 53231
rect 26882 53116 26959 53132
tri 26959 53116 26975 53132 sw
rect 26882 53050 26975 53116
rect 27011 52991 27125 53149
tri 27161 53116 27177 53132 se
rect 27177 53116 27254 53132
rect 27161 53050 27254 53116
rect 26882 52915 27254 52991
rect 26882 52790 26975 52856
rect 26882 52774 26959 52790
tri 26959 52774 26975 52790 nw
rect 27011 52757 27125 52915
rect 27161 52790 27254 52856
tri 27161 52774 27177 52790 ne
rect 27177 52774 27254 52790
rect 26994 52675 27142 52757
rect 26882 52642 26959 52658
tri 26959 52642 26975 52658 sw
rect 26882 52576 26975 52642
rect 26882 52474 26975 52540
rect 26882 52458 26959 52474
tri 26959 52458 26975 52474 nw
rect 27011 52441 27125 52675
tri 27161 52642 27177 52658 se
rect 27177 52642 27254 52658
rect 27161 52576 27254 52642
rect 27161 52474 27254 52540
tri 27161 52458 27177 52474 ne
rect 27177 52458 27254 52474
rect 26994 52359 27142 52441
rect 26882 52326 26959 52342
tri 26959 52326 26975 52342 sw
rect 26882 52260 26975 52326
rect 27011 52201 27125 52359
tri 27161 52326 27177 52342 se
rect 27177 52326 27254 52342
rect 27161 52260 27254 52326
rect 26882 52125 27254 52201
rect 26882 52000 26975 52066
rect 26882 51984 26959 52000
tri 26959 51984 26975 52000 nw
rect 27011 51967 27125 52125
rect 27161 52000 27254 52066
tri 27161 51984 27177 52000 ne
rect 27177 51984 27254 52000
rect 26994 51885 27142 51967
rect 26882 51852 26959 51868
tri 26959 51852 26975 51868 sw
rect 26882 51786 26975 51852
rect 26882 51684 26975 51750
rect 26882 51668 26959 51684
tri 26959 51668 26975 51684 nw
rect 27011 51651 27125 51885
tri 27161 51852 27177 51868 se
rect 27177 51852 27254 51868
rect 27161 51786 27254 51852
rect 27161 51684 27254 51750
tri 27161 51668 27177 51684 ne
rect 27177 51668 27254 51684
rect 26994 51569 27142 51651
rect 26882 51536 26959 51552
tri 26959 51536 26975 51552 sw
rect 26882 51470 26975 51536
rect 27011 51411 27125 51569
tri 27161 51536 27177 51552 se
rect 27177 51536 27254 51552
rect 27161 51470 27254 51536
rect 26882 51335 27254 51411
rect 26882 51210 26975 51276
rect 26882 51194 26959 51210
tri 26959 51194 26975 51210 nw
rect 27011 51177 27125 51335
rect 27161 51210 27254 51276
tri 27161 51194 27177 51210 ne
rect 27177 51194 27254 51210
rect 26994 51095 27142 51177
rect 26882 51062 26959 51078
tri 26959 51062 26975 51078 sw
rect 26882 50996 26975 51062
rect 26882 50894 26975 50960
rect 26882 50878 26959 50894
tri 26959 50878 26975 50894 nw
rect 27011 50861 27125 51095
tri 27161 51062 27177 51078 se
rect 27177 51062 27254 51078
rect 27161 50996 27254 51062
rect 27161 50894 27254 50960
tri 27161 50878 27177 50894 ne
rect 27177 50878 27254 50894
rect 26994 50779 27142 50861
rect 26882 50746 26959 50762
tri 26959 50746 26975 50762 sw
rect 26882 50680 26975 50746
rect 27011 50621 27125 50779
tri 27161 50746 27177 50762 se
rect 27177 50746 27254 50762
rect 27161 50680 27254 50746
rect 26882 50545 27254 50621
rect 26882 50420 26975 50486
rect 26882 50404 26959 50420
tri 26959 50404 26975 50420 nw
rect 27011 50387 27125 50545
rect 27161 50420 27254 50486
tri 27161 50404 27177 50420 ne
rect 27177 50404 27254 50420
rect 26994 50305 27142 50387
rect 26882 50272 26959 50288
tri 26959 50272 26975 50288 sw
rect 26882 50206 26975 50272
rect 26882 50104 26975 50170
rect 26882 50088 26959 50104
tri 26959 50088 26975 50104 nw
rect 27011 50071 27125 50305
tri 27161 50272 27177 50288 se
rect 27177 50272 27254 50288
rect 27161 50206 27254 50272
rect 27161 50104 27254 50170
tri 27161 50088 27177 50104 ne
rect 27177 50088 27254 50104
rect 26994 49989 27142 50071
rect 26882 49956 26959 49972
tri 26959 49956 26975 49972 sw
rect 26882 49890 26975 49956
rect 27011 49831 27125 49989
tri 27161 49956 27177 49972 se
rect 27177 49956 27254 49972
rect 27161 49890 27254 49956
rect 26882 49755 27254 49831
rect 26882 49630 26975 49696
rect 26882 49614 26959 49630
tri 26959 49614 26975 49630 nw
rect 27011 49597 27125 49755
rect 27161 49630 27254 49696
tri 27161 49614 27177 49630 ne
rect 27177 49614 27254 49630
rect 26994 49515 27142 49597
rect 26882 49482 26959 49498
tri 26959 49482 26975 49498 sw
rect 26882 49416 26975 49482
rect 26882 49314 26975 49380
rect 26882 49298 26959 49314
tri 26959 49298 26975 49314 nw
rect 27011 49281 27125 49515
tri 27161 49482 27177 49498 se
rect 27177 49482 27254 49498
rect 27161 49416 27254 49482
rect 27161 49314 27254 49380
tri 27161 49298 27177 49314 ne
rect 27177 49298 27254 49314
rect 26994 49199 27142 49281
rect 26882 49166 26959 49182
tri 26959 49166 26975 49182 sw
rect 26882 49100 26975 49166
rect 27011 49041 27125 49199
tri 27161 49166 27177 49182 se
rect 27177 49166 27254 49182
rect 27161 49100 27254 49166
rect 26882 48965 27254 49041
rect 26882 48840 26975 48906
rect 26882 48824 26959 48840
tri 26959 48824 26975 48840 nw
rect 27011 48807 27125 48965
rect 27161 48840 27254 48906
tri 27161 48824 27177 48840 ne
rect 27177 48824 27254 48840
rect 26994 48725 27142 48807
rect 26882 48692 26959 48708
tri 26959 48692 26975 48708 sw
rect 26882 48626 26975 48692
rect 26882 48524 26975 48590
rect 26882 48508 26959 48524
tri 26959 48508 26975 48524 nw
rect 27011 48491 27125 48725
tri 27161 48692 27177 48708 se
rect 27177 48692 27254 48708
rect 27161 48626 27254 48692
rect 27161 48524 27254 48590
tri 27161 48508 27177 48524 ne
rect 27177 48508 27254 48524
rect 26994 48409 27142 48491
rect 26882 48376 26959 48392
tri 26959 48376 26975 48392 sw
rect 26882 48310 26975 48376
rect 27011 48251 27125 48409
tri 27161 48376 27177 48392 se
rect 27177 48376 27254 48392
rect 27161 48310 27254 48376
rect 26882 48175 27254 48251
rect 26882 48050 26975 48116
rect 26882 48034 26959 48050
tri 26959 48034 26975 48050 nw
rect 27011 48017 27125 48175
rect 27161 48050 27254 48116
tri 27161 48034 27177 48050 ne
rect 27177 48034 27254 48050
rect 26994 47935 27142 48017
rect 26882 47902 26959 47918
tri 26959 47902 26975 47918 sw
rect 26882 47836 26975 47902
rect 26882 47734 26975 47800
rect 26882 47718 26959 47734
tri 26959 47718 26975 47734 nw
rect 27011 47701 27125 47935
tri 27161 47902 27177 47918 se
rect 27177 47902 27254 47918
rect 27161 47836 27254 47902
rect 27161 47734 27254 47800
tri 27161 47718 27177 47734 ne
rect 27177 47718 27254 47734
rect 26994 47619 27142 47701
rect 26882 47586 26959 47602
tri 26959 47586 26975 47602 sw
rect 26882 47520 26975 47586
rect 27011 47461 27125 47619
tri 27161 47586 27177 47602 se
rect 27177 47586 27254 47602
rect 27161 47520 27254 47586
rect 26882 47385 27254 47461
rect 26882 47260 26975 47326
rect 26882 47244 26959 47260
tri 26959 47244 26975 47260 nw
rect 27011 47227 27125 47385
rect 27161 47260 27254 47326
tri 27161 47244 27177 47260 ne
rect 27177 47244 27254 47260
rect 26994 47145 27142 47227
rect 26882 47112 26959 47128
tri 26959 47112 26975 47128 sw
rect 26882 47046 26975 47112
rect 26882 46944 26975 47010
rect 26882 46928 26959 46944
tri 26959 46928 26975 46944 nw
rect 27011 46911 27125 47145
tri 27161 47112 27177 47128 se
rect 27177 47112 27254 47128
rect 27161 47046 27254 47112
rect 27161 46944 27254 47010
tri 27161 46928 27177 46944 ne
rect 27177 46928 27254 46944
rect 26994 46829 27142 46911
rect 26882 46796 26959 46812
tri 26959 46796 26975 46812 sw
rect 26882 46730 26975 46796
rect 27011 46671 27125 46829
tri 27161 46796 27177 46812 se
rect 27177 46796 27254 46812
rect 27161 46730 27254 46796
rect 26882 46595 27254 46671
rect 26882 46470 26975 46536
rect 26882 46454 26959 46470
tri 26959 46454 26975 46470 nw
rect 27011 46437 27125 46595
rect 27161 46470 27254 46536
tri 27161 46454 27177 46470 ne
rect 27177 46454 27254 46470
rect 26994 46355 27142 46437
rect 26882 46322 26959 46338
tri 26959 46322 26975 46338 sw
rect 26882 46256 26975 46322
rect 26882 46154 26975 46220
rect 26882 46138 26959 46154
tri 26959 46138 26975 46154 nw
rect 27011 46121 27125 46355
tri 27161 46322 27177 46338 se
rect 27177 46322 27254 46338
rect 27161 46256 27254 46322
rect 27161 46154 27254 46220
tri 27161 46138 27177 46154 ne
rect 27177 46138 27254 46154
rect 26994 46039 27142 46121
rect 26882 46006 26959 46022
tri 26959 46006 26975 46022 sw
rect 26882 45940 26975 46006
rect 27011 45881 27125 46039
tri 27161 46006 27177 46022 se
rect 27177 46006 27254 46022
rect 27161 45940 27254 46006
rect 26882 45805 27254 45881
rect 26882 45680 26975 45746
rect 26882 45664 26959 45680
tri 26959 45664 26975 45680 nw
rect 27011 45647 27125 45805
rect 27161 45680 27254 45746
tri 27161 45664 27177 45680 ne
rect 27177 45664 27254 45680
rect 26994 45565 27142 45647
rect 26882 45532 26959 45548
tri 26959 45532 26975 45548 sw
rect 26882 45466 26975 45532
rect 26882 45364 26975 45430
rect 26882 45348 26959 45364
tri 26959 45348 26975 45364 nw
rect 27011 45331 27125 45565
tri 27161 45532 27177 45548 se
rect 27177 45532 27254 45548
rect 27161 45466 27254 45532
rect 27161 45364 27254 45430
tri 27161 45348 27177 45364 ne
rect 27177 45348 27254 45364
rect 26994 45249 27142 45331
rect 26882 45216 26959 45232
tri 26959 45216 26975 45232 sw
rect 26882 45150 26975 45216
rect 27011 45091 27125 45249
tri 27161 45216 27177 45232 se
rect 27177 45216 27254 45232
rect 27161 45150 27254 45216
rect 26882 45015 27254 45091
rect 26882 44890 26975 44956
rect 26882 44874 26959 44890
tri 26959 44874 26975 44890 nw
rect 27011 44857 27125 45015
rect 27161 44890 27254 44956
tri 27161 44874 27177 44890 ne
rect 27177 44874 27254 44890
rect 26994 44775 27142 44857
rect 26882 44742 26959 44758
tri 26959 44742 26975 44758 sw
rect 26882 44676 26975 44742
rect 26882 44574 26975 44640
rect 26882 44558 26959 44574
tri 26959 44558 26975 44574 nw
rect 27011 44541 27125 44775
tri 27161 44742 27177 44758 se
rect 27177 44742 27254 44758
rect 27161 44676 27254 44742
rect 27161 44574 27254 44640
tri 27161 44558 27177 44574 ne
rect 27177 44558 27254 44574
rect 26994 44459 27142 44541
rect 26882 44426 26959 44442
tri 26959 44426 26975 44442 sw
rect 26882 44360 26975 44426
rect 27011 44301 27125 44459
tri 27161 44426 27177 44442 se
rect 27177 44426 27254 44442
rect 27161 44360 27254 44426
rect 26882 44225 27254 44301
rect 26882 44100 26975 44166
rect 26882 44084 26959 44100
tri 26959 44084 26975 44100 nw
rect 27011 44067 27125 44225
rect 27161 44100 27254 44166
tri 27161 44084 27177 44100 ne
rect 27177 44084 27254 44100
rect 26994 43985 27142 44067
rect 26882 43952 26959 43968
tri 26959 43952 26975 43968 sw
rect 26882 43886 26975 43952
rect 26882 43784 26975 43850
rect 26882 43768 26959 43784
tri 26959 43768 26975 43784 nw
rect 27011 43751 27125 43985
tri 27161 43952 27177 43968 se
rect 27177 43952 27254 43968
rect 27161 43886 27254 43952
rect 27161 43784 27254 43850
tri 27161 43768 27177 43784 ne
rect 27177 43768 27254 43784
rect 26994 43669 27142 43751
rect 26882 43636 26959 43652
tri 26959 43636 26975 43652 sw
rect 26882 43570 26975 43636
rect 27011 43511 27125 43669
tri 27161 43636 27177 43652 se
rect 27177 43636 27254 43652
rect 27161 43570 27254 43636
rect 26882 43435 27254 43511
rect 26882 43310 26975 43376
rect 26882 43294 26959 43310
tri 26959 43294 26975 43310 nw
rect 27011 43277 27125 43435
rect 27161 43310 27254 43376
tri 27161 43294 27177 43310 ne
rect 27177 43294 27254 43310
rect 26994 43195 27142 43277
rect 26882 43162 26959 43178
tri 26959 43162 26975 43178 sw
rect 26882 43096 26975 43162
rect 26882 42994 26975 43060
rect 26882 42978 26959 42994
tri 26959 42978 26975 42994 nw
rect 27011 42961 27125 43195
tri 27161 43162 27177 43178 se
rect 27177 43162 27254 43178
rect 27161 43096 27254 43162
rect 27161 42994 27254 43060
tri 27161 42978 27177 42994 ne
rect 27177 42978 27254 42994
rect 26994 42879 27142 42961
rect 26882 42846 26959 42862
tri 26959 42846 26975 42862 sw
rect 26882 42780 26975 42846
rect 27011 42721 27125 42879
tri 27161 42846 27177 42862 se
rect 27177 42846 27254 42862
rect 27161 42780 27254 42846
rect 26882 42645 27254 42721
rect 26882 42520 26975 42586
rect 26882 42504 26959 42520
tri 26959 42504 26975 42520 nw
rect 27011 42487 27125 42645
rect 27161 42520 27254 42586
tri 27161 42504 27177 42520 ne
rect 27177 42504 27254 42520
rect 26994 42405 27142 42487
rect 26882 42372 26959 42388
tri 26959 42372 26975 42388 sw
rect 26882 42306 26975 42372
rect 26882 42204 26975 42270
rect 26882 42188 26959 42204
tri 26959 42188 26975 42204 nw
rect 27011 42171 27125 42405
tri 27161 42372 27177 42388 se
rect 27177 42372 27254 42388
rect 27161 42306 27254 42372
rect 27161 42204 27254 42270
tri 27161 42188 27177 42204 ne
rect 27177 42188 27254 42204
rect 26994 42089 27142 42171
rect 26882 42056 26959 42072
tri 26959 42056 26975 42072 sw
rect 26882 41990 26975 42056
rect 27011 41931 27125 42089
tri 27161 42056 27177 42072 se
rect 27177 42056 27254 42072
rect 27161 41990 27254 42056
rect 26882 41855 27254 41931
rect 26882 41730 26975 41796
rect 26882 41714 26959 41730
tri 26959 41714 26975 41730 nw
rect 27011 41697 27125 41855
rect 27161 41730 27254 41796
tri 27161 41714 27177 41730 ne
rect 27177 41714 27254 41730
rect 26994 41615 27142 41697
rect 26882 41582 26959 41598
tri 26959 41582 26975 41598 sw
rect 26882 41516 26975 41582
rect 26882 41414 26975 41480
rect 26882 41398 26959 41414
tri 26959 41398 26975 41414 nw
rect 27011 41381 27125 41615
tri 27161 41582 27177 41598 se
rect 27177 41582 27254 41598
rect 27161 41516 27254 41582
rect 27161 41414 27254 41480
tri 27161 41398 27177 41414 ne
rect 27177 41398 27254 41414
rect 26994 41299 27142 41381
rect 26882 41266 26959 41282
tri 26959 41266 26975 41282 sw
rect 26882 41200 26975 41266
rect 27011 41141 27125 41299
tri 27161 41266 27177 41282 se
rect 27177 41266 27254 41282
rect 27161 41200 27254 41266
rect 26882 41065 27254 41141
rect 26882 40940 26975 41006
rect 26882 40924 26959 40940
tri 26959 40924 26975 40940 nw
rect 27011 40907 27125 41065
rect 27161 40940 27254 41006
tri 27161 40924 27177 40940 ne
rect 27177 40924 27254 40940
rect 26994 40825 27142 40907
rect 26882 40792 26959 40808
tri 26959 40792 26975 40808 sw
rect 26882 40726 26975 40792
rect 26882 40624 26975 40690
rect 26882 40608 26959 40624
tri 26959 40608 26975 40624 nw
rect 27011 40591 27125 40825
tri 27161 40792 27177 40808 se
rect 27177 40792 27254 40808
rect 27161 40726 27254 40792
rect 27161 40624 27254 40690
tri 27161 40608 27177 40624 ne
rect 27177 40608 27254 40624
rect 26994 40509 27142 40591
rect 26882 40476 26959 40492
tri 26959 40476 26975 40492 sw
rect 26882 40410 26975 40476
rect 27011 40351 27125 40509
tri 27161 40476 27177 40492 se
rect 27177 40476 27254 40492
rect 27161 40410 27254 40476
rect 26882 40275 27254 40351
rect 26882 40150 26975 40216
rect 26882 40134 26959 40150
tri 26959 40134 26975 40150 nw
rect 27011 40117 27125 40275
rect 27161 40150 27254 40216
tri 27161 40134 27177 40150 ne
rect 27177 40134 27254 40150
rect 26994 40035 27142 40117
rect 26882 40002 26959 40018
tri 26959 40002 26975 40018 sw
rect 26882 39936 26975 40002
rect 26882 39834 26975 39900
rect 26882 39818 26959 39834
tri 26959 39818 26975 39834 nw
rect 27011 39801 27125 40035
tri 27161 40002 27177 40018 se
rect 27177 40002 27254 40018
rect 27161 39936 27254 40002
rect 27161 39834 27254 39900
tri 27161 39818 27177 39834 ne
rect 27177 39818 27254 39834
rect 26994 39719 27142 39801
rect 26882 39686 26959 39702
tri 26959 39686 26975 39702 sw
rect 26882 39620 26975 39686
rect 27011 39561 27125 39719
tri 27161 39686 27177 39702 se
rect 27177 39686 27254 39702
rect 27161 39620 27254 39686
rect 26882 39485 27254 39561
rect 26882 39360 26975 39426
rect 26882 39344 26959 39360
tri 26959 39344 26975 39360 nw
rect 27011 39327 27125 39485
rect 27161 39360 27254 39426
tri 27161 39344 27177 39360 ne
rect 27177 39344 27254 39360
rect 26994 39245 27142 39327
rect 26882 39212 26959 39228
tri 26959 39212 26975 39228 sw
rect 26882 39146 26975 39212
rect 26882 39044 26975 39110
rect 26882 39028 26959 39044
tri 26959 39028 26975 39044 nw
rect 27011 39011 27125 39245
tri 27161 39212 27177 39228 se
rect 27177 39212 27254 39228
rect 27161 39146 27254 39212
rect 27161 39044 27254 39110
tri 27161 39028 27177 39044 ne
rect 27177 39028 27254 39044
rect 26994 38929 27142 39011
rect 26882 38896 26959 38912
tri 26959 38896 26975 38912 sw
rect 26882 38830 26975 38896
rect 27011 38771 27125 38929
tri 27161 38896 27177 38912 se
rect 27177 38896 27254 38912
rect 27161 38830 27254 38896
rect 26882 38695 27254 38771
rect 26882 38570 26975 38636
rect 26882 38554 26959 38570
tri 26959 38554 26975 38570 nw
rect 27011 38537 27125 38695
rect 27161 38570 27254 38636
tri 27161 38554 27177 38570 ne
rect 27177 38554 27254 38570
rect 26994 38455 27142 38537
rect 26882 38422 26959 38438
tri 26959 38422 26975 38438 sw
rect 26882 38356 26975 38422
rect 26882 38254 26975 38320
rect 26882 38238 26959 38254
tri 26959 38238 26975 38254 nw
rect 27011 38221 27125 38455
tri 27161 38422 27177 38438 se
rect 27177 38422 27254 38438
rect 27161 38356 27254 38422
rect 27161 38254 27254 38320
tri 27161 38238 27177 38254 ne
rect 27177 38238 27254 38254
rect 26994 38139 27142 38221
rect 26882 38106 26959 38122
tri 26959 38106 26975 38122 sw
rect 26882 38040 26975 38106
rect 27011 37981 27125 38139
tri 27161 38106 27177 38122 se
rect 27177 38106 27254 38122
rect 27161 38040 27254 38106
rect 26882 37905 27254 37981
rect 26882 37780 26975 37846
rect 26882 37764 26959 37780
tri 26959 37764 26975 37780 nw
rect 27011 37747 27125 37905
rect 27161 37780 27254 37846
tri 27161 37764 27177 37780 ne
rect 27177 37764 27254 37780
rect 26994 37665 27142 37747
rect 26882 37632 26959 37648
tri 26959 37632 26975 37648 sw
rect 26882 37566 26975 37632
rect 26882 37464 26975 37530
rect 26882 37448 26959 37464
tri 26959 37448 26975 37464 nw
rect 27011 37431 27125 37665
tri 27161 37632 27177 37648 se
rect 27177 37632 27254 37648
rect 27161 37566 27254 37632
rect 27161 37464 27254 37530
tri 27161 37448 27177 37464 ne
rect 27177 37448 27254 37464
rect 26994 37349 27142 37431
rect 26882 37316 26959 37332
tri 26959 37316 26975 37332 sw
rect 26882 37250 26975 37316
rect 27011 37191 27125 37349
tri 27161 37316 27177 37332 se
rect 27177 37316 27254 37332
rect 27161 37250 27254 37316
rect 26882 37115 27254 37191
rect 26882 36990 26975 37056
rect 26882 36974 26959 36990
tri 26959 36974 26975 36990 nw
rect 27011 36957 27125 37115
rect 27161 36990 27254 37056
tri 27161 36974 27177 36990 ne
rect 27177 36974 27254 36990
rect 26994 36875 27142 36957
rect 26882 36842 26959 36858
tri 26959 36842 26975 36858 sw
rect 26882 36776 26975 36842
rect 26882 36674 26975 36740
rect 26882 36658 26959 36674
tri 26959 36658 26975 36674 nw
rect 27011 36641 27125 36875
tri 27161 36842 27177 36858 se
rect 27177 36842 27254 36858
rect 27161 36776 27254 36842
rect 27161 36674 27254 36740
tri 27161 36658 27177 36674 ne
rect 27177 36658 27254 36674
rect 26994 36559 27142 36641
rect 26882 36526 26959 36542
tri 26959 36526 26975 36542 sw
rect 26882 36460 26975 36526
rect 27011 36401 27125 36559
tri 27161 36526 27177 36542 se
rect 27177 36526 27254 36542
rect 27161 36460 27254 36526
rect 26882 36325 27254 36401
rect 26882 36200 26975 36266
rect 26882 36184 26959 36200
tri 26959 36184 26975 36200 nw
rect 27011 36167 27125 36325
rect 27161 36200 27254 36266
tri 27161 36184 27177 36200 ne
rect 27177 36184 27254 36200
rect 26994 36085 27142 36167
rect 26882 36052 26959 36068
tri 26959 36052 26975 36068 sw
rect 26882 35986 26975 36052
rect 26882 35884 26975 35950
rect 26882 35868 26959 35884
tri 26959 35868 26975 35884 nw
rect 27011 35851 27125 36085
tri 27161 36052 27177 36068 se
rect 27177 36052 27254 36068
rect 27161 35986 27254 36052
rect 27161 35884 27254 35950
tri 27161 35868 27177 35884 ne
rect 27177 35868 27254 35884
rect 26994 35769 27142 35851
rect 26882 35736 26959 35752
tri 26959 35736 26975 35752 sw
rect 26882 35670 26975 35736
rect 27011 35611 27125 35769
tri 27161 35736 27177 35752 se
rect 27177 35736 27254 35752
rect 27161 35670 27254 35736
rect 26882 35535 27254 35611
rect 26882 35410 26975 35476
rect 26882 35394 26959 35410
tri 26959 35394 26975 35410 nw
rect 27011 35377 27125 35535
rect 27161 35410 27254 35476
tri 27161 35394 27177 35410 ne
rect 27177 35394 27254 35410
rect 26994 35295 27142 35377
rect 26882 35262 26959 35278
tri 26959 35262 26975 35278 sw
rect 26882 35196 26975 35262
rect 26882 35094 26975 35160
rect 26882 35078 26959 35094
tri 26959 35078 26975 35094 nw
rect 27011 35061 27125 35295
tri 27161 35262 27177 35278 se
rect 27177 35262 27254 35278
rect 27161 35196 27254 35262
rect 27161 35094 27254 35160
tri 27161 35078 27177 35094 ne
rect 27177 35078 27254 35094
rect 26994 34979 27142 35061
rect 26882 34946 26959 34962
tri 26959 34946 26975 34962 sw
rect 26882 34880 26975 34946
rect 27011 34821 27125 34979
tri 27161 34946 27177 34962 se
rect 27177 34946 27254 34962
rect 27161 34880 27254 34946
rect 26882 34745 27254 34821
rect 26882 34620 26975 34686
rect 26882 34604 26959 34620
tri 26959 34604 26975 34620 nw
rect 27011 34587 27125 34745
rect 27161 34620 27254 34686
tri 27161 34604 27177 34620 ne
rect 27177 34604 27254 34620
rect 26994 34505 27142 34587
rect 26882 34472 26959 34488
tri 26959 34472 26975 34488 sw
rect 26882 34406 26975 34472
rect 26882 34304 26975 34370
rect 26882 34288 26959 34304
tri 26959 34288 26975 34304 nw
rect 27011 34271 27125 34505
tri 27161 34472 27177 34488 se
rect 27177 34472 27254 34488
rect 27161 34406 27254 34472
rect 27161 34304 27254 34370
tri 27161 34288 27177 34304 ne
rect 27177 34288 27254 34304
rect 26994 34189 27142 34271
rect 26882 34156 26959 34172
tri 26959 34156 26975 34172 sw
rect 26882 34090 26975 34156
rect 27011 34031 27125 34189
tri 27161 34156 27177 34172 se
rect 27177 34156 27254 34172
rect 27161 34090 27254 34156
rect 26882 33955 27254 34031
rect 26882 33830 26975 33896
rect 26882 33814 26959 33830
tri 26959 33814 26975 33830 nw
rect 27011 33797 27125 33955
rect 27161 33830 27254 33896
tri 27161 33814 27177 33830 ne
rect 27177 33814 27254 33830
rect 26994 33715 27142 33797
rect 26882 33682 26959 33698
tri 26959 33682 26975 33698 sw
rect 26882 33616 26975 33682
rect 26882 33514 26975 33580
rect 26882 33498 26959 33514
tri 26959 33498 26975 33514 nw
rect 27011 33481 27125 33715
tri 27161 33682 27177 33698 se
rect 27177 33682 27254 33698
rect 27161 33616 27254 33682
rect 27161 33514 27254 33580
tri 27161 33498 27177 33514 ne
rect 27177 33498 27254 33514
rect 26994 33399 27142 33481
rect 26882 33366 26959 33382
tri 26959 33366 26975 33382 sw
rect 26882 33300 26975 33366
rect 27011 33241 27125 33399
tri 27161 33366 27177 33382 se
rect 27177 33366 27254 33382
rect 27161 33300 27254 33366
rect 26882 33165 27254 33241
rect 26882 33040 26975 33106
rect 26882 33024 26959 33040
tri 26959 33024 26975 33040 nw
rect 27011 33007 27125 33165
rect 27161 33040 27254 33106
tri 27161 33024 27177 33040 ne
rect 27177 33024 27254 33040
rect 26994 32925 27142 33007
rect 26882 32892 26959 32908
tri 26959 32892 26975 32908 sw
rect 26882 32826 26975 32892
rect 26882 32724 26975 32790
rect 26882 32708 26959 32724
tri 26959 32708 26975 32724 nw
rect 27011 32691 27125 32925
tri 27161 32892 27177 32908 se
rect 27177 32892 27254 32908
rect 27161 32826 27254 32892
rect 27161 32724 27254 32790
tri 27161 32708 27177 32724 ne
rect 27177 32708 27254 32724
rect 26994 32609 27142 32691
rect 26882 32576 26959 32592
tri 26959 32576 26975 32592 sw
rect 26882 32510 26975 32576
rect 27011 32451 27125 32609
tri 27161 32576 27177 32592 se
rect 27177 32576 27254 32592
rect 27161 32510 27254 32576
rect 26882 32375 27254 32451
rect 26882 32250 26975 32316
rect 26882 32234 26959 32250
tri 26959 32234 26975 32250 nw
rect 27011 32217 27125 32375
rect 27161 32250 27254 32316
tri 27161 32234 27177 32250 ne
rect 27177 32234 27254 32250
rect 26994 32135 27142 32217
rect 26882 32102 26959 32118
tri 26959 32102 26975 32118 sw
rect 26882 32036 26975 32102
rect 26882 31934 26975 32000
rect 26882 31918 26959 31934
tri 26959 31918 26975 31934 nw
rect 27011 31901 27125 32135
tri 27161 32102 27177 32118 se
rect 27177 32102 27254 32118
rect 27161 32036 27254 32102
rect 27161 31934 27254 32000
tri 27161 31918 27177 31934 ne
rect 27177 31918 27254 31934
rect 26994 31819 27142 31901
rect 26882 31786 26959 31802
tri 26959 31786 26975 31802 sw
rect 26882 31720 26975 31786
rect 27011 31661 27125 31819
tri 27161 31786 27177 31802 se
rect 27177 31786 27254 31802
rect 27161 31720 27254 31786
rect 26882 31585 27254 31661
rect 26882 31460 26975 31526
rect 26882 31444 26959 31460
tri 26959 31444 26975 31460 nw
rect 27011 31427 27125 31585
rect 27161 31460 27254 31526
tri 27161 31444 27177 31460 ne
rect 27177 31444 27254 31460
rect 26994 31345 27142 31427
rect 26882 31312 26959 31328
tri 26959 31312 26975 31328 sw
rect 26882 31246 26975 31312
rect 26882 31144 26975 31210
rect 26882 31128 26959 31144
tri 26959 31128 26975 31144 nw
rect 27011 31111 27125 31345
tri 27161 31312 27177 31328 se
rect 27177 31312 27254 31328
rect 27161 31246 27254 31312
rect 27161 31144 27254 31210
tri 27161 31128 27177 31144 ne
rect 27177 31128 27254 31144
rect 26994 31029 27142 31111
rect 26882 30996 26959 31012
tri 26959 30996 26975 31012 sw
rect 26882 30930 26975 30996
rect 27011 30871 27125 31029
tri 27161 30996 27177 31012 se
rect 27177 30996 27254 31012
rect 27161 30930 27254 30996
rect 26882 30795 27254 30871
rect 26882 30670 26975 30736
rect 26882 30654 26959 30670
tri 26959 30654 26975 30670 nw
rect 27011 30637 27125 30795
rect 27161 30670 27254 30736
tri 27161 30654 27177 30670 ne
rect 27177 30654 27254 30670
rect 26994 30555 27142 30637
rect 26882 30522 26959 30538
tri 26959 30522 26975 30538 sw
rect 26882 30456 26975 30522
rect 26882 30354 26975 30420
rect 26882 30338 26959 30354
tri 26959 30338 26975 30354 nw
rect 27011 30321 27125 30555
tri 27161 30522 27177 30538 se
rect 27177 30522 27254 30538
rect 27161 30456 27254 30522
rect 27161 30354 27254 30420
tri 27161 30338 27177 30354 ne
rect 27177 30338 27254 30354
rect 26994 30239 27142 30321
rect 26882 30206 26959 30222
tri 26959 30206 26975 30222 sw
rect 26882 30140 26975 30206
rect 27011 30081 27125 30239
tri 27161 30206 27177 30222 se
rect 27177 30206 27254 30222
rect 27161 30140 27254 30206
rect 26882 30005 27254 30081
rect 26882 29880 26975 29946
rect 26882 29864 26959 29880
tri 26959 29864 26975 29880 nw
rect 27011 29847 27125 30005
rect 27161 29880 27254 29946
tri 27161 29864 27177 29880 ne
rect 27177 29864 27254 29880
rect 26994 29765 27142 29847
rect 26882 29732 26959 29748
tri 26959 29732 26975 29748 sw
rect 26882 29666 26975 29732
rect 26882 29564 26975 29630
rect 26882 29548 26959 29564
tri 26959 29548 26975 29564 nw
rect 27011 29531 27125 29765
tri 27161 29732 27177 29748 se
rect 27177 29732 27254 29748
rect 27161 29666 27254 29732
rect 27161 29564 27254 29630
tri 27161 29548 27177 29564 ne
rect 27177 29548 27254 29564
rect 26994 29449 27142 29531
rect 26882 29416 26959 29432
tri 26959 29416 26975 29432 sw
rect 26882 29350 26975 29416
rect 27011 29291 27125 29449
tri 27161 29416 27177 29432 se
rect 27177 29416 27254 29432
rect 27161 29350 27254 29416
rect 26882 29215 27254 29291
rect 26882 29090 26975 29156
rect 26882 29074 26959 29090
tri 26959 29074 26975 29090 nw
rect 27011 29057 27125 29215
rect 27161 29090 27254 29156
tri 27161 29074 27177 29090 ne
rect 27177 29074 27254 29090
rect 26994 28975 27142 29057
rect 26882 28942 26959 28958
tri 26959 28942 26975 28958 sw
rect 26882 28876 26975 28942
rect 27011 28833 27125 28975
tri 27161 28942 27177 28958 se
rect 27177 28942 27254 28958
rect 27161 28876 27254 28942
rect 27290 28463 27326 80603
rect 27362 28463 27398 80603
rect 27434 80445 27470 80603
rect 27426 80303 27478 80445
rect 27434 28763 27470 80303
rect 27426 28621 27478 28763
rect 27434 28463 27470 28621
rect 27506 28463 27542 80603
rect 27578 28463 27614 80603
rect 27650 28833 27734 80233
rect 27770 28463 27806 80603
rect 27842 28463 27878 80603
rect 27914 80445 27950 80603
rect 27906 80303 27958 80445
rect 27914 28763 27950 80303
rect 27906 28621 27958 28763
rect 27914 28463 27950 28621
rect 27986 28463 28022 80603
rect 28058 28463 28094 80603
rect 28130 80124 28223 80190
rect 28130 80108 28207 80124
tri 28207 80108 28223 80124 nw
rect 28259 80091 28373 80233
rect 28409 80124 28502 80190
tri 28409 80108 28425 80124 ne
rect 28425 80108 28502 80124
rect 28242 80009 28390 80091
rect 28130 79976 28207 79992
tri 28207 79976 28223 79992 sw
rect 28130 79910 28223 79976
rect 28259 79851 28373 80009
tri 28409 79976 28425 79992 se
rect 28425 79976 28502 79992
rect 28409 79910 28502 79976
rect 28130 79775 28502 79851
rect 28130 79650 28223 79716
rect 28130 79634 28207 79650
tri 28207 79634 28223 79650 nw
rect 28259 79617 28373 79775
rect 28409 79650 28502 79716
tri 28409 79634 28425 79650 ne
rect 28425 79634 28502 79650
rect 28242 79535 28390 79617
rect 28130 79502 28207 79518
tri 28207 79502 28223 79518 sw
rect 28130 79436 28223 79502
rect 28130 79334 28223 79400
rect 28130 79318 28207 79334
tri 28207 79318 28223 79334 nw
rect 28259 79301 28373 79535
tri 28409 79502 28425 79518 se
rect 28425 79502 28502 79518
rect 28409 79436 28502 79502
rect 28409 79334 28502 79400
tri 28409 79318 28425 79334 ne
rect 28425 79318 28502 79334
rect 28242 79219 28390 79301
rect 28130 79186 28207 79202
tri 28207 79186 28223 79202 sw
rect 28130 79120 28223 79186
rect 28259 79061 28373 79219
tri 28409 79186 28425 79202 se
rect 28425 79186 28502 79202
rect 28409 79120 28502 79186
rect 28130 78985 28502 79061
rect 28130 78860 28223 78926
rect 28130 78844 28207 78860
tri 28207 78844 28223 78860 nw
rect 28259 78827 28373 78985
rect 28409 78860 28502 78926
tri 28409 78844 28425 78860 ne
rect 28425 78844 28502 78860
rect 28242 78745 28390 78827
rect 28130 78712 28207 78728
tri 28207 78712 28223 78728 sw
rect 28130 78646 28223 78712
rect 28130 78544 28223 78610
rect 28130 78528 28207 78544
tri 28207 78528 28223 78544 nw
rect 28259 78511 28373 78745
tri 28409 78712 28425 78728 se
rect 28425 78712 28502 78728
rect 28409 78646 28502 78712
rect 28409 78544 28502 78610
tri 28409 78528 28425 78544 ne
rect 28425 78528 28502 78544
rect 28242 78429 28390 78511
rect 28130 78396 28207 78412
tri 28207 78396 28223 78412 sw
rect 28130 78330 28223 78396
rect 28259 78271 28373 78429
tri 28409 78396 28425 78412 se
rect 28425 78396 28502 78412
rect 28409 78330 28502 78396
rect 28130 78195 28502 78271
rect 28130 78070 28223 78136
rect 28130 78054 28207 78070
tri 28207 78054 28223 78070 nw
rect 28259 78037 28373 78195
rect 28409 78070 28502 78136
tri 28409 78054 28425 78070 ne
rect 28425 78054 28502 78070
rect 28242 77955 28390 78037
rect 28130 77922 28207 77938
tri 28207 77922 28223 77938 sw
rect 28130 77856 28223 77922
rect 28130 77754 28223 77820
rect 28130 77738 28207 77754
tri 28207 77738 28223 77754 nw
rect 28259 77721 28373 77955
tri 28409 77922 28425 77938 se
rect 28425 77922 28502 77938
rect 28409 77856 28502 77922
rect 28409 77754 28502 77820
tri 28409 77738 28425 77754 ne
rect 28425 77738 28502 77754
rect 28242 77639 28390 77721
rect 28130 77606 28207 77622
tri 28207 77606 28223 77622 sw
rect 28130 77540 28223 77606
rect 28259 77481 28373 77639
tri 28409 77606 28425 77622 se
rect 28425 77606 28502 77622
rect 28409 77540 28502 77606
rect 28130 77405 28502 77481
rect 28130 77280 28223 77346
rect 28130 77264 28207 77280
tri 28207 77264 28223 77280 nw
rect 28259 77247 28373 77405
rect 28409 77280 28502 77346
tri 28409 77264 28425 77280 ne
rect 28425 77264 28502 77280
rect 28242 77165 28390 77247
rect 28130 77132 28207 77148
tri 28207 77132 28223 77148 sw
rect 28130 77066 28223 77132
rect 28130 76964 28223 77030
rect 28130 76948 28207 76964
tri 28207 76948 28223 76964 nw
rect 28259 76931 28373 77165
tri 28409 77132 28425 77148 se
rect 28425 77132 28502 77148
rect 28409 77066 28502 77132
rect 28409 76964 28502 77030
tri 28409 76948 28425 76964 ne
rect 28425 76948 28502 76964
rect 28242 76849 28390 76931
rect 28130 76816 28207 76832
tri 28207 76816 28223 76832 sw
rect 28130 76750 28223 76816
rect 28259 76691 28373 76849
tri 28409 76816 28425 76832 se
rect 28425 76816 28502 76832
rect 28409 76750 28502 76816
rect 28130 76615 28502 76691
rect 28130 76490 28223 76556
rect 28130 76474 28207 76490
tri 28207 76474 28223 76490 nw
rect 28259 76457 28373 76615
rect 28409 76490 28502 76556
tri 28409 76474 28425 76490 ne
rect 28425 76474 28502 76490
rect 28242 76375 28390 76457
rect 28130 76342 28207 76358
tri 28207 76342 28223 76358 sw
rect 28130 76276 28223 76342
rect 28130 76174 28223 76240
rect 28130 76158 28207 76174
tri 28207 76158 28223 76174 nw
rect 28259 76141 28373 76375
tri 28409 76342 28425 76358 se
rect 28425 76342 28502 76358
rect 28409 76276 28502 76342
rect 28409 76174 28502 76240
tri 28409 76158 28425 76174 ne
rect 28425 76158 28502 76174
rect 28242 76059 28390 76141
rect 28130 76026 28207 76042
tri 28207 76026 28223 76042 sw
rect 28130 75960 28223 76026
rect 28259 75901 28373 76059
tri 28409 76026 28425 76042 se
rect 28425 76026 28502 76042
rect 28409 75960 28502 76026
rect 28130 75825 28502 75901
rect 28130 75700 28223 75766
rect 28130 75684 28207 75700
tri 28207 75684 28223 75700 nw
rect 28259 75667 28373 75825
rect 28409 75700 28502 75766
tri 28409 75684 28425 75700 ne
rect 28425 75684 28502 75700
rect 28242 75585 28390 75667
rect 28130 75552 28207 75568
tri 28207 75552 28223 75568 sw
rect 28130 75486 28223 75552
rect 28130 75384 28223 75450
rect 28130 75368 28207 75384
tri 28207 75368 28223 75384 nw
rect 28259 75351 28373 75585
tri 28409 75552 28425 75568 se
rect 28425 75552 28502 75568
rect 28409 75486 28502 75552
rect 28409 75384 28502 75450
tri 28409 75368 28425 75384 ne
rect 28425 75368 28502 75384
rect 28242 75269 28390 75351
rect 28130 75236 28207 75252
tri 28207 75236 28223 75252 sw
rect 28130 75170 28223 75236
rect 28259 75111 28373 75269
tri 28409 75236 28425 75252 se
rect 28425 75236 28502 75252
rect 28409 75170 28502 75236
rect 28130 75035 28502 75111
rect 28130 74910 28223 74976
rect 28130 74894 28207 74910
tri 28207 74894 28223 74910 nw
rect 28259 74877 28373 75035
rect 28409 74910 28502 74976
tri 28409 74894 28425 74910 ne
rect 28425 74894 28502 74910
rect 28242 74795 28390 74877
rect 28130 74762 28207 74778
tri 28207 74762 28223 74778 sw
rect 28130 74696 28223 74762
rect 28130 74594 28223 74660
rect 28130 74578 28207 74594
tri 28207 74578 28223 74594 nw
rect 28259 74561 28373 74795
tri 28409 74762 28425 74778 se
rect 28425 74762 28502 74778
rect 28409 74696 28502 74762
rect 28409 74594 28502 74660
tri 28409 74578 28425 74594 ne
rect 28425 74578 28502 74594
rect 28242 74479 28390 74561
rect 28130 74446 28207 74462
tri 28207 74446 28223 74462 sw
rect 28130 74380 28223 74446
rect 28259 74321 28373 74479
tri 28409 74446 28425 74462 se
rect 28425 74446 28502 74462
rect 28409 74380 28502 74446
rect 28130 74245 28502 74321
rect 28130 74120 28223 74186
rect 28130 74104 28207 74120
tri 28207 74104 28223 74120 nw
rect 28259 74087 28373 74245
rect 28409 74120 28502 74186
tri 28409 74104 28425 74120 ne
rect 28425 74104 28502 74120
rect 28242 74005 28390 74087
rect 28130 73972 28207 73988
tri 28207 73972 28223 73988 sw
rect 28130 73906 28223 73972
rect 28130 73804 28223 73870
rect 28130 73788 28207 73804
tri 28207 73788 28223 73804 nw
rect 28259 73771 28373 74005
tri 28409 73972 28425 73988 se
rect 28425 73972 28502 73988
rect 28409 73906 28502 73972
rect 28409 73804 28502 73870
tri 28409 73788 28425 73804 ne
rect 28425 73788 28502 73804
rect 28242 73689 28390 73771
rect 28130 73656 28207 73672
tri 28207 73656 28223 73672 sw
rect 28130 73590 28223 73656
rect 28259 73531 28373 73689
tri 28409 73656 28425 73672 se
rect 28425 73656 28502 73672
rect 28409 73590 28502 73656
rect 28130 73455 28502 73531
rect 28130 73330 28223 73396
rect 28130 73314 28207 73330
tri 28207 73314 28223 73330 nw
rect 28259 73297 28373 73455
rect 28409 73330 28502 73396
tri 28409 73314 28425 73330 ne
rect 28425 73314 28502 73330
rect 28242 73215 28390 73297
rect 28130 73182 28207 73198
tri 28207 73182 28223 73198 sw
rect 28130 73116 28223 73182
rect 28130 73014 28223 73080
rect 28130 72998 28207 73014
tri 28207 72998 28223 73014 nw
rect 28259 72981 28373 73215
tri 28409 73182 28425 73198 se
rect 28425 73182 28502 73198
rect 28409 73116 28502 73182
rect 28409 73014 28502 73080
tri 28409 72998 28425 73014 ne
rect 28425 72998 28502 73014
rect 28242 72899 28390 72981
rect 28130 72866 28207 72882
tri 28207 72866 28223 72882 sw
rect 28130 72800 28223 72866
rect 28259 72741 28373 72899
tri 28409 72866 28425 72882 se
rect 28425 72866 28502 72882
rect 28409 72800 28502 72866
rect 28130 72665 28502 72741
rect 28130 72540 28223 72606
rect 28130 72524 28207 72540
tri 28207 72524 28223 72540 nw
rect 28259 72507 28373 72665
rect 28409 72540 28502 72606
tri 28409 72524 28425 72540 ne
rect 28425 72524 28502 72540
rect 28242 72425 28390 72507
rect 28130 72392 28207 72408
tri 28207 72392 28223 72408 sw
rect 28130 72326 28223 72392
rect 28130 72224 28223 72290
rect 28130 72208 28207 72224
tri 28207 72208 28223 72224 nw
rect 28259 72191 28373 72425
tri 28409 72392 28425 72408 se
rect 28425 72392 28502 72408
rect 28409 72326 28502 72392
rect 28409 72224 28502 72290
tri 28409 72208 28425 72224 ne
rect 28425 72208 28502 72224
rect 28242 72109 28390 72191
rect 28130 72076 28207 72092
tri 28207 72076 28223 72092 sw
rect 28130 72010 28223 72076
rect 28259 71951 28373 72109
tri 28409 72076 28425 72092 se
rect 28425 72076 28502 72092
rect 28409 72010 28502 72076
rect 28130 71875 28502 71951
rect 28130 71750 28223 71816
rect 28130 71734 28207 71750
tri 28207 71734 28223 71750 nw
rect 28259 71717 28373 71875
rect 28409 71750 28502 71816
tri 28409 71734 28425 71750 ne
rect 28425 71734 28502 71750
rect 28242 71635 28390 71717
rect 28130 71602 28207 71618
tri 28207 71602 28223 71618 sw
rect 28130 71536 28223 71602
rect 28130 71434 28223 71500
rect 28130 71418 28207 71434
tri 28207 71418 28223 71434 nw
rect 28259 71401 28373 71635
tri 28409 71602 28425 71618 se
rect 28425 71602 28502 71618
rect 28409 71536 28502 71602
rect 28409 71434 28502 71500
tri 28409 71418 28425 71434 ne
rect 28425 71418 28502 71434
rect 28242 71319 28390 71401
rect 28130 71286 28207 71302
tri 28207 71286 28223 71302 sw
rect 28130 71220 28223 71286
rect 28259 71161 28373 71319
tri 28409 71286 28425 71302 se
rect 28425 71286 28502 71302
rect 28409 71220 28502 71286
rect 28130 71085 28502 71161
rect 28130 70960 28223 71026
rect 28130 70944 28207 70960
tri 28207 70944 28223 70960 nw
rect 28259 70927 28373 71085
rect 28409 70960 28502 71026
tri 28409 70944 28425 70960 ne
rect 28425 70944 28502 70960
rect 28242 70845 28390 70927
rect 28130 70812 28207 70828
tri 28207 70812 28223 70828 sw
rect 28130 70746 28223 70812
rect 28130 70644 28223 70710
rect 28130 70628 28207 70644
tri 28207 70628 28223 70644 nw
rect 28259 70611 28373 70845
tri 28409 70812 28425 70828 se
rect 28425 70812 28502 70828
rect 28409 70746 28502 70812
rect 28409 70644 28502 70710
tri 28409 70628 28425 70644 ne
rect 28425 70628 28502 70644
rect 28242 70529 28390 70611
rect 28130 70496 28207 70512
tri 28207 70496 28223 70512 sw
rect 28130 70430 28223 70496
rect 28259 70371 28373 70529
tri 28409 70496 28425 70512 se
rect 28425 70496 28502 70512
rect 28409 70430 28502 70496
rect 28130 70295 28502 70371
rect 28130 70170 28223 70236
rect 28130 70154 28207 70170
tri 28207 70154 28223 70170 nw
rect 28259 70137 28373 70295
rect 28409 70170 28502 70236
tri 28409 70154 28425 70170 ne
rect 28425 70154 28502 70170
rect 28242 70055 28390 70137
rect 28130 70022 28207 70038
tri 28207 70022 28223 70038 sw
rect 28130 69956 28223 70022
rect 28130 69854 28223 69920
rect 28130 69838 28207 69854
tri 28207 69838 28223 69854 nw
rect 28259 69821 28373 70055
tri 28409 70022 28425 70038 se
rect 28425 70022 28502 70038
rect 28409 69956 28502 70022
rect 28409 69854 28502 69920
tri 28409 69838 28425 69854 ne
rect 28425 69838 28502 69854
rect 28242 69739 28390 69821
rect 28130 69706 28207 69722
tri 28207 69706 28223 69722 sw
rect 28130 69640 28223 69706
rect 28259 69581 28373 69739
tri 28409 69706 28425 69722 se
rect 28425 69706 28502 69722
rect 28409 69640 28502 69706
rect 28130 69505 28502 69581
rect 28130 69380 28223 69446
rect 28130 69364 28207 69380
tri 28207 69364 28223 69380 nw
rect 28259 69347 28373 69505
rect 28409 69380 28502 69446
tri 28409 69364 28425 69380 ne
rect 28425 69364 28502 69380
rect 28242 69265 28390 69347
rect 28130 69232 28207 69248
tri 28207 69232 28223 69248 sw
rect 28130 69166 28223 69232
rect 28130 69064 28223 69130
rect 28130 69048 28207 69064
tri 28207 69048 28223 69064 nw
rect 28259 69031 28373 69265
tri 28409 69232 28425 69248 se
rect 28425 69232 28502 69248
rect 28409 69166 28502 69232
rect 28409 69064 28502 69130
tri 28409 69048 28425 69064 ne
rect 28425 69048 28502 69064
rect 28242 68949 28390 69031
rect 28130 68916 28207 68932
tri 28207 68916 28223 68932 sw
rect 28130 68850 28223 68916
rect 28259 68791 28373 68949
tri 28409 68916 28425 68932 se
rect 28425 68916 28502 68932
rect 28409 68850 28502 68916
rect 28130 68715 28502 68791
rect 28130 68590 28223 68656
rect 28130 68574 28207 68590
tri 28207 68574 28223 68590 nw
rect 28259 68557 28373 68715
rect 28409 68590 28502 68656
tri 28409 68574 28425 68590 ne
rect 28425 68574 28502 68590
rect 28242 68475 28390 68557
rect 28130 68442 28207 68458
tri 28207 68442 28223 68458 sw
rect 28130 68376 28223 68442
rect 28130 68274 28223 68340
rect 28130 68258 28207 68274
tri 28207 68258 28223 68274 nw
rect 28259 68241 28373 68475
tri 28409 68442 28425 68458 se
rect 28425 68442 28502 68458
rect 28409 68376 28502 68442
rect 28409 68274 28502 68340
tri 28409 68258 28425 68274 ne
rect 28425 68258 28502 68274
rect 28242 68159 28390 68241
rect 28130 68126 28207 68142
tri 28207 68126 28223 68142 sw
rect 28130 68060 28223 68126
rect 28259 68001 28373 68159
tri 28409 68126 28425 68142 se
rect 28425 68126 28502 68142
rect 28409 68060 28502 68126
rect 28130 67925 28502 68001
rect 28130 67800 28223 67866
rect 28130 67784 28207 67800
tri 28207 67784 28223 67800 nw
rect 28259 67767 28373 67925
rect 28409 67800 28502 67866
tri 28409 67784 28425 67800 ne
rect 28425 67784 28502 67800
rect 28242 67685 28390 67767
rect 28130 67652 28207 67668
tri 28207 67652 28223 67668 sw
rect 28130 67586 28223 67652
rect 28130 67484 28223 67550
rect 28130 67468 28207 67484
tri 28207 67468 28223 67484 nw
rect 28259 67451 28373 67685
tri 28409 67652 28425 67668 se
rect 28425 67652 28502 67668
rect 28409 67586 28502 67652
rect 28409 67484 28502 67550
tri 28409 67468 28425 67484 ne
rect 28425 67468 28502 67484
rect 28242 67369 28390 67451
rect 28130 67336 28207 67352
tri 28207 67336 28223 67352 sw
rect 28130 67270 28223 67336
rect 28259 67211 28373 67369
tri 28409 67336 28425 67352 se
rect 28425 67336 28502 67352
rect 28409 67270 28502 67336
rect 28130 67135 28502 67211
rect 28130 67010 28223 67076
rect 28130 66994 28207 67010
tri 28207 66994 28223 67010 nw
rect 28259 66977 28373 67135
rect 28409 67010 28502 67076
tri 28409 66994 28425 67010 ne
rect 28425 66994 28502 67010
rect 28242 66895 28390 66977
rect 28130 66862 28207 66878
tri 28207 66862 28223 66878 sw
rect 28130 66796 28223 66862
rect 28130 66694 28223 66760
rect 28130 66678 28207 66694
tri 28207 66678 28223 66694 nw
rect 28259 66661 28373 66895
tri 28409 66862 28425 66878 se
rect 28425 66862 28502 66878
rect 28409 66796 28502 66862
rect 28409 66694 28502 66760
tri 28409 66678 28425 66694 ne
rect 28425 66678 28502 66694
rect 28242 66579 28390 66661
rect 28130 66546 28207 66562
tri 28207 66546 28223 66562 sw
rect 28130 66480 28223 66546
rect 28259 66421 28373 66579
tri 28409 66546 28425 66562 se
rect 28425 66546 28502 66562
rect 28409 66480 28502 66546
rect 28130 66345 28502 66421
rect 28130 66220 28223 66286
rect 28130 66204 28207 66220
tri 28207 66204 28223 66220 nw
rect 28259 66187 28373 66345
rect 28409 66220 28502 66286
tri 28409 66204 28425 66220 ne
rect 28425 66204 28502 66220
rect 28242 66105 28390 66187
rect 28130 66072 28207 66088
tri 28207 66072 28223 66088 sw
rect 28130 66006 28223 66072
rect 28130 65904 28223 65970
rect 28130 65888 28207 65904
tri 28207 65888 28223 65904 nw
rect 28259 65871 28373 66105
tri 28409 66072 28425 66088 se
rect 28425 66072 28502 66088
rect 28409 66006 28502 66072
rect 28409 65904 28502 65970
tri 28409 65888 28425 65904 ne
rect 28425 65888 28502 65904
rect 28242 65789 28390 65871
rect 28130 65756 28207 65772
tri 28207 65756 28223 65772 sw
rect 28130 65690 28223 65756
rect 28259 65631 28373 65789
tri 28409 65756 28425 65772 se
rect 28425 65756 28502 65772
rect 28409 65690 28502 65756
rect 28130 65555 28502 65631
rect 28130 65430 28223 65496
rect 28130 65414 28207 65430
tri 28207 65414 28223 65430 nw
rect 28259 65397 28373 65555
rect 28409 65430 28502 65496
tri 28409 65414 28425 65430 ne
rect 28425 65414 28502 65430
rect 28242 65315 28390 65397
rect 28130 65282 28207 65298
tri 28207 65282 28223 65298 sw
rect 28130 65216 28223 65282
rect 28130 65114 28223 65180
rect 28130 65098 28207 65114
tri 28207 65098 28223 65114 nw
rect 28259 65081 28373 65315
tri 28409 65282 28425 65298 se
rect 28425 65282 28502 65298
rect 28409 65216 28502 65282
rect 28409 65114 28502 65180
tri 28409 65098 28425 65114 ne
rect 28425 65098 28502 65114
rect 28242 64999 28390 65081
rect 28130 64966 28207 64982
tri 28207 64966 28223 64982 sw
rect 28130 64900 28223 64966
rect 28259 64841 28373 64999
tri 28409 64966 28425 64982 se
rect 28425 64966 28502 64982
rect 28409 64900 28502 64966
rect 28130 64765 28502 64841
rect 28130 64640 28223 64706
rect 28130 64624 28207 64640
tri 28207 64624 28223 64640 nw
rect 28259 64607 28373 64765
rect 28409 64640 28502 64706
tri 28409 64624 28425 64640 ne
rect 28425 64624 28502 64640
rect 28242 64525 28390 64607
rect 28130 64492 28207 64508
tri 28207 64492 28223 64508 sw
rect 28130 64426 28223 64492
rect 28130 64324 28223 64390
rect 28130 64308 28207 64324
tri 28207 64308 28223 64324 nw
rect 28259 64291 28373 64525
tri 28409 64492 28425 64508 se
rect 28425 64492 28502 64508
rect 28409 64426 28502 64492
rect 28409 64324 28502 64390
tri 28409 64308 28425 64324 ne
rect 28425 64308 28502 64324
rect 28242 64209 28390 64291
rect 28130 64176 28207 64192
tri 28207 64176 28223 64192 sw
rect 28130 64110 28223 64176
rect 28259 64051 28373 64209
tri 28409 64176 28425 64192 se
rect 28425 64176 28502 64192
rect 28409 64110 28502 64176
rect 28130 63975 28502 64051
rect 28130 63850 28223 63916
rect 28130 63834 28207 63850
tri 28207 63834 28223 63850 nw
rect 28259 63817 28373 63975
rect 28409 63850 28502 63916
tri 28409 63834 28425 63850 ne
rect 28425 63834 28502 63850
rect 28242 63735 28390 63817
rect 28130 63702 28207 63718
tri 28207 63702 28223 63718 sw
rect 28130 63636 28223 63702
rect 28130 63534 28223 63600
rect 28130 63518 28207 63534
tri 28207 63518 28223 63534 nw
rect 28259 63501 28373 63735
tri 28409 63702 28425 63718 se
rect 28425 63702 28502 63718
rect 28409 63636 28502 63702
rect 28409 63534 28502 63600
tri 28409 63518 28425 63534 ne
rect 28425 63518 28502 63534
rect 28242 63419 28390 63501
rect 28130 63386 28207 63402
tri 28207 63386 28223 63402 sw
rect 28130 63320 28223 63386
rect 28259 63261 28373 63419
tri 28409 63386 28425 63402 se
rect 28425 63386 28502 63402
rect 28409 63320 28502 63386
rect 28130 63185 28502 63261
rect 28130 63060 28223 63126
rect 28130 63044 28207 63060
tri 28207 63044 28223 63060 nw
rect 28259 63027 28373 63185
rect 28409 63060 28502 63126
tri 28409 63044 28425 63060 ne
rect 28425 63044 28502 63060
rect 28242 62945 28390 63027
rect 28130 62912 28207 62928
tri 28207 62912 28223 62928 sw
rect 28130 62846 28223 62912
rect 28130 62744 28223 62810
rect 28130 62728 28207 62744
tri 28207 62728 28223 62744 nw
rect 28259 62711 28373 62945
tri 28409 62912 28425 62928 se
rect 28425 62912 28502 62928
rect 28409 62846 28502 62912
rect 28409 62744 28502 62810
tri 28409 62728 28425 62744 ne
rect 28425 62728 28502 62744
rect 28242 62629 28390 62711
rect 28130 62596 28207 62612
tri 28207 62596 28223 62612 sw
rect 28130 62530 28223 62596
rect 28259 62471 28373 62629
tri 28409 62596 28425 62612 se
rect 28425 62596 28502 62612
rect 28409 62530 28502 62596
rect 28130 62395 28502 62471
rect 28130 62270 28223 62336
rect 28130 62254 28207 62270
tri 28207 62254 28223 62270 nw
rect 28259 62237 28373 62395
rect 28409 62270 28502 62336
tri 28409 62254 28425 62270 ne
rect 28425 62254 28502 62270
rect 28242 62155 28390 62237
rect 28130 62122 28207 62138
tri 28207 62122 28223 62138 sw
rect 28130 62056 28223 62122
rect 28130 61954 28223 62020
rect 28130 61938 28207 61954
tri 28207 61938 28223 61954 nw
rect 28259 61921 28373 62155
tri 28409 62122 28425 62138 se
rect 28425 62122 28502 62138
rect 28409 62056 28502 62122
rect 28409 61954 28502 62020
tri 28409 61938 28425 61954 ne
rect 28425 61938 28502 61954
rect 28242 61839 28390 61921
rect 28130 61806 28207 61822
tri 28207 61806 28223 61822 sw
rect 28130 61740 28223 61806
rect 28259 61681 28373 61839
tri 28409 61806 28425 61822 se
rect 28425 61806 28502 61822
rect 28409 61740 28502 61806
rect 28130 61605 28502 61681
rect 28130 61480 28223 61546
rect 28130 61464 28207 61480
tri 28207 61464 28223 61480 nw
rect 28259 61447 28373 61605
rect 28409 61480 28502 61546
tri 28409 61464 28425 61480 ne
rect 28425 61464 28502 61480
rect 28242 61365 28390 61447
rect 28130 61332 28207 61348
tri 28207 61332 28223 61348 sw
rect 28130 61266 28223 61332
rect 28130 61164 28223 61230
rect 28130 61148 28207 61164
tri 28207 61148 28223 61164 nw
rect 28259 61131 28373 61365
tri 28409 61332 28425 61348 se
rect 28425 61332 28502 61348
rect 28409 61266 28502 61332
rect 28409 61164 28502 61230
tri 28409 61148 28425 61164 ne
rect 28425 61148 28502 61164
rect 28242 61049 28390 61131
rect 28130 61016 28207 61032
tri 28207 61016 28223 61032 sw
rect 28130 60950 28223 61016
rect 28259 60891 28373 61049
tri 28409 61016 28425 61032 se
rect 28425 61016 28502 61032
rect 28409 60950 28502 61016
rect 28130 60815 28502 60891
rect 28130 60690 28223 60756
rect 28130 60674 28207 60690
tri 28207 60674 28223 60690 nw
rect 28259 60657 28373 60815
rect 28409 60690 28502 60756
tri 28409 60674 28425 60690 ne
rect 28425 60674 28502 60690
rect 28242 60575 28390 60657
rect 28130 60542 28207 60558
tri 28207 60542 28223 60558 sw
rect 28130 60476 28223 60542
rect 28130 60374 28223 60440
rect 28130 60358 28207 60374
tri 28207 60358 28223 60374 nw
rect 28259 60341 28373 60575
tri 28409 60542 28425 60558 se
rect 28425 60542 28502 60558
rect 28409 60476 28502 60542
rect 28409 60374 28502 60440
tri 28409 60358 28425 60374 ne
rect 28425 60358 28502 60374
rect 28242 60259 28390 60341
rect 28130 60226 28207 60242
tri 28207 60226 28223 60242 sw
rect 28130 60160 28223 60226
rect 28259 60101 28373 60259
tri 28409 60226 28425 60242 se
rect 28425 60226 28502 60242
rect 28409 60160 28502 60226
rect 28130 60025 28502 60101
rect 28130 59900 28223 59966
rect 28130 59884 28207 59900
tri 28207 59884 28223 59900 nw
rect 28259 59867 28373 60025
rect 28409 59900 28502 59966
tri 28409 59884 28425 59900 ne
rect 28425 59884 28502 59900
rect 28242 59785 28390 59867
rect 28130 59752 28207 59768
tri 28207 59752 28223 59768 sw
rect 28130 59686 28223 59752
rect 28130 59584 28223 59650
rect 28130 59568 28207 59584
tri 28207 59568 28223 59584 nw
rect 28259 59551 28373 59785
tri 28409 59752 28425 59768 se
rect 28425 59752 28502 59768
rect 28409 59686 28502 59752
rect 28409 59584 28502 59650
tri 28409 59568 28425 59584 ne
rect 28425 59568 28502 59584
rect 28242 59469 28390 59551
rect 28130 59436 28207 59452
tri 28207 59436 28223 59452 sw
rect 28130 59370 28223 59436
rect 28259 59311 28373 59469
tri 28409 59436 28425 59452 se
rect 28425 59436 28502 59452
rect 28409 59370 28502 59436
rect 28130 59235 28502 59311
rect 28130 59110 28223 59176
rect 28130 59094 28207 59110
tri 28207 59094 28223 59110 nw
rect 28259 59077 28373 59235
rect 28409 59110 28502 59176
tri 28409 59094 28425 59110 ne
rect 28425 59094 28502 59110
rect 28242 58995 28390 59077
rect 28130 58962 28207 58978
tri 28207 58962 28223 58978 sw
rect 28130 58896 28223 58962
rect 28130 58794 28223 58860
rect 28130 58778 28207 58794
tri 28207 58778 28223 58794 nw
rect 28259 58761 28373 58995
tri 28409 58962 28425 58978 se
rect 28425 58962 28502 58978
rect 28409 58896 28502 58962
rect 28409 58794 28502 58860
tri 28409 58778 28425 58794 ne
rect 28425 58778 28502 58794
rect 28242 58679 28390 58761
rect 28130 58646 28207 58662
tri 28207 58646 28223 58662 sw
rect 28130 58580 28223 58646
rect 28259 58521 28373 58679
tri 28409 58646 28425 58662 se
rect 28425 58646 28502 58662
rect 28409 58580 28502 58646
rect 28130 58445 28502 58521
rect 28130 58320 28223 58386
rect 28130 58304 28207 58320
tri 28207 58304 28223 58320 nw
rect 28259 58287 28373 58445
rect 28409 58320 28502 58386
tri 28409 58304 28425 58320 ne
rect 28425 58304 28502 58320
rect 28242 58205 28390 58287
rect 28130 58172 28207 58188
tri 28207 58172 28223 58188 sw
rect 28130 58106 28223 58172
rect 28130 58004 28223 58070
rect 28130 57988 28207 58004
tri 28207 57988 28223 58004 nw
rect 28259 57971 28373 58205
tri 28409 58172 28425 58188 se
rect 28425 58172 28502 58188
rect 28409 58106 28502 58172
rect 28409 58004 28502 58070
tri 28409 57988 28425 58004 ne
rect 28425 57988 28502 58004
rect 28242 57889 28390 57971
rect 28130 57856 28207 57872
tri 28207 57856 28223 57872 sw
rect 28130 57790 28223 57856
rect 28259 57731 28373 57889
tri 28409 57856 28425 57872 se
rect 28425 57856 28502 57872
rect 28409 57790 28502 57856
rect 28130 57655 28502 57731
rect 28130 57530 28223 57596
rect 28130 57514 28207 57530
tri 28207 57514 28223 57530 nw
rect 28259 57497 28373 57655
rect 28409 57530 28502 57596
tri 28409 57514 28425 57530 ne
rect 28425 57514 28502 57530
rect 28242 57415 28390 57497
rect 28130 57382 28207 57398
tri 28207 57382 28223 57398 sw
rect 28130 57316 28223 57382
rect 28130 57214 28223 57280
rect 28130 57198 28207 57214
tri 28207 57198 28223 57214 nw
rect 28259 57181 28373 57415
tri 28409 57382 28425 57398 se
rect 28425 57382 28502 57398
rect 28409 57316 28502 57382
rect 28409 57214 28502 57280
tri 28409 57198 28425 57214 ne
rect 28425 57198 28502 57214
rect 28242 57099 28390 57181
rect 28130 57066 28207 57082
tri 28207 57066 28223 57082 sw
rect 28130 57000 28223 57066
rect 28259 56941 28373 57099
tri 28409 57066 28425 57082 se
rect 28425 57066 28502 57082
rect 28409 57000 28502 57066
rect 28130 56865 28502 56941
rect 28130 56740 28223 56806
rect 28130 56724 28207 56740
tri 28207 56724 28223 56740 nw
rect 28259 56707 28373 56865
rect 28409 56740 28502 56806
tri 28409 56724 28425 56740 ne
rect 28425 56724 28502 56740
rect 28242 56625 28390 56707
rect 28130 56592 28207 56608
tri 28207 56592 28223 56608 sw
rect 28130 56526 28223 56592
rect 28130 56424 28223 56490
rect 28130 56408 28207 56424
tri 28207 56408 28223 56424 nw
rect 28259 56391 28373 56625
tri 28409 56592 28425 56608 se
rect 28425 56592 28502 56608
rect 28409 56526 28502 56592
rect 28409 56424 28502 56490
tri 28409 56408 28425 56424 ne
rect 28425 56408 28502 56424
rect 28242 56309 28390 56391
rect 28130 56276 28207 56292
tri 28207 56276 28223 56292 sw
rect 28130 56210 28223 56276
rect 28259 56151 28373 56309
tri 28409 56276 28425 56292 se
rect 28425 56276 28502 56292
rect 28409 56210 28502 56276
rect 28130 56075 28502 56151
rect 28130 55950 28223 56016
rect 28130 55934 28207 55950
tri 28207 55934 28223 55950 nw
rect 28259 55917 28373 56075
rect 28409 55950 28502 56016
tri 28409 55934 28425 55950 ne
rect 28425 55934 28502 55950
rect 28242 55835 28390 55917
rect 28130 55802 28207 55818
tri 28207 55802 28223 55818 sw
rect 28130 55736 28223 55802
rect 28130 55634 28223 55700
rect 28130 55618 28207 55634
tri 28207 55618 28223 55634 nw
rect 28259 55601 28373 55835
tri 28409 55802 28425 55818 se
rect 28425 55802 28502 55818
rect 28409 55736 28502 55802
rect 28409 55634 28502 55700
tri 28409 55618 28425 55634 ne
rect 28425 55618 28502 55634
rect 28242 55519 28390 55601
rect 28130 55486 28207 55502
tri 28207 55486 28223 55502 sw
rect 28130 55420 28223 55486
rect 28259 55361 28373 55519
tri 28409 55486 28425 55502 se
rect 28425 55486 28502 55502
rect 28409 55420 28502 55486
rect 28130 55285 28502 55361
rect 28130 55160 28223 55226
rect 28130 55144 28207 55160
tri 28207 55144 28223 55160 nw
rect 28259 55127 28373 55285
rect 28409 55160 28502 55226
tri 28409 55144 28425 55160 ne
rect 28425 55144 28502 55160
rect 28242 55045 28390 55127
rect 28130 55012 28207 55028
tri 28207 55012 28223 55028 sw
rect 28130 54946 28223 55012
rect 28130 54844 28223 54910
rect 28130 54828 28207 54844
tri 28207 54828 28223 54844 nw
rect 28259 54811 28373 55045
tri 28409 55012 28425 55028 se
rect 28425 55012 28502 55028
rect 28409 54946 28502 55012
rect 28409 54844 28502 54910
tri 28409 54828 28425 54844 ne
rect 28425 54828 28502 54844
rect 28242 54729 28390 54811
rect 28130 54696 28207 54712
tri 28207 54696 28223 54712 sw
rect 28130 54630 28223 54696
rect 28259 54571 28373 54729
tri 28409 54696 28425 54712 se
rect 28425 54696 28502 54712
rect 28409 54630 28502 54696
rect 28130 54495 28502 54571
rect 28130 54370 28223 54436
rect 28130 54354 28207 54370
tri 28207 54354 28223 54370 nw
rect 28259 54337 28373 54495
rect 28409 54370 28502 54436
tri 28409 54354 28425 54370 ne
rect 28425 54354 28502 54370
rect 28242 54255 28390 54337
rect 28130 54222 28207 54238
tri 28207 54222 28223 54238 sw
rect 28130 54156 28223 54222
rect 28130 54054 28223 54120
rect 28130 54038 28207 54054
tri 28207 54038 28223 54054 nw
rect 28259 54021 28373 54255
tri 28409 54222 28425 54238 se
rect 28425 54222 28502 54238
rect 28409 54156 28502 54222
rect 28409 54054 28502 54120
tri 28409 54038 28425 54054 ne
rect 28425 54038 28502 54054
rect 28242 53939 28390 54021
rect 28130 53906 28207 53922
tri 28207 53906 28223 53922 sw
rect 28130 53840 28223 53906
rect 28259 53781 28373 53939
tri 28409 53906 28425 53922 se
rect 28425 53906 28502 53922
rect 28409 53840 28502 53906
rect 28130 53705 28502 53781
rect 28130 53580 28223 53646
rect 28130 53564 28207 53580
tri 28207 53564 28223 53580 nw
rect 28259 53547 28373 53705
rect 28409 53580 28502 53646
tri 28409 53564 28425 53580 ne
rect 28425 53564 28502 53580
rect 28242 53465 28390 53547
rect 28130 53432 28207 53448
tri 28207 53432 28223 53448 sw
rect 28130 53366 28223 53432
rect 28130 53264 28223 53330
rect 28130 53248 28207 53264
tri 28207 53248 28223 53264 nw
rect 28259 53231 28373 53465
tri 28409 53432 28425 53448 se
rect 28425 53432 28502 53448
rect 28409 53366 28502 53432
rect 28409 53264 28502 53330
tri 28409 53248 28425 53264 ne
rect 28425 53248 28502 53264
rect 28242 53149 28390 53231
rect 28130 53116 28207 53132
tri 28207 53116 28223 53132 sw
rect 28130 53050 28223 53116
rect 28259 52991 28373 53149
tri 28409 53116 28425 53132 se
rect 28425 53116 28502 53132
rect 28409 53050 28502 53116
rect 28130 52915 28502 52991
rect 28130 52790 28223 52856
rect 28130 52774 28207 52790
tri 28207 52774 28223 52790 nw
rect 28259 52757 28373 52915
rect 28409 52790 28502 52856
tri 28409 52774 28425 52790 ne
rect 28425 52774 28502 52790
rect 28242 52675 28390 52757
rect 28130 52642 28207 52658
tri 28207 52642 28223 52658 sw
rect 28130 52576 28223 52642
rect 28130 52474 28223 52540
rect 28130 52458 28207 52474
tri 28207 52458 28223 52474 nw
rect 28259 52441 28373 52675
tri 28409 52642 28425 52658 se
rect 28425 52642 28502 52658
rect 28409 52576 28502 52642
rect 28409 52474 28502 52540
tri 28409 52458 28425 52474 ne
rect 28425 52458 28502 52474
rect 28242 52359 28390 52441
rect 28130 52326 28207 52342
tri 28207 52326 28223 52342 sw
rect 28130 52260 28223 52326
rect 28259 52201 28373 52359
tri 28409 52326 28425 52342 se
rect 28425 52326 28502 52342
rect 28409 52260 28502 52326
rect 28130 52125 28502 52201
rect 28130 52000 28223 52066
rect 28130 51984 28207 52000
tri 28207 51984 28223 52000 nw
rect 28259 51967 28373 52125
rect 28409 52000 28502 52066
tri 28409 51984 28425 52000 ne
rect 28425 51984 28502 52000
rect 28242 51885 28390 51967
rect 28130 51852 28207 51868
tri 28207 51852 28223 51868 sw
rect 28130 51786 28223 51852
rect 28130 51684 28223 51750
rect 28130 51668 28207 51684
tri 28207 51668 28223 51684 nw
rect 28259 51651 28373 51885
tri 28409 51852 28425 51868 se
rect 28425 51852 28502 51868
rect 28409 51786 28502 51852
rect 28409 51684 28502 51750
tri 28409 51668 28425 51684 ne
rect 28425 51668 28502 51684
rect 28242 51569 28390 51651
rect 28130 51536 28207 51552
tri 28207 51536 28223 51552 sw
rect 28130 51470 28223 51536
rect 28259 51411 28373 51569
tri 28409 51536 28425 51552 se
rect 28425 51536 28502 51552
rect 28409 51470 28502 51536
rect 28130 51335 28502 51411
rect 28130 51210 28223 51276
rect 28130 51194 28207 51210
tri 28207 51194 28223 51210 nw
rect 28259 51177 28373 51335
rect 28409 51210 28502 51276
tri 28409 51194 28425 51210 ne
rect 28425 51194 28502 51210
rect 28242 51095 28390 51177
rect 28130 51062 28207 51078
tri 28207 51062 28223 51078 sw
rect 28130 50996 28223 51062
rect 28130 50894 28223 50960
rect 28130 50878 28207 50894
tri 28207 50878 28223 50894 nw
rect 28259 50861 28373 51095
tri 28409 51062 28425 51078 se
rect 28425 51062 28502 51078
rect 28409 50996 28502 51062
rect 28409 50894 28502 50960
tri 28409 50878 28425 50894 ne
rect 28425 50878 28502 50894
rect 28242 50779 28390 50861
rect 28130 50746 28207 50762
tri 28207 50746 28223 50762 sw
rect 28130 50680 28223 50746
rect 28259 50621 28373 50779
tri 28409 50746 28425 50762 se
rect 28425 50746 28502 50762
rect 28409 50680 28502 50746
rect 28130 50545 28502 50621
rect 28130 50420 28223 50486
rect 28130 50404 28207 50420
tri 28207 50404 28223 50420 nw
rect 28259 50387 28373 50545
rect 28409 50420 28502 50486
tri 28409 50404 28425 50420 ne
rect 28425 50404 28502 50420
rect 28242 50305 28390 50387
rect 28130 50272 28207 50288
tri 28207 50272 28223 50288 sw
rect 28130 50206 28223 50272
rect 28130 50104 28223 50170
rect 28130 50088 28207 50104
tri 28207 50088 28223 50104 nw
rect 28259 50071 28373 50305
tri 28409 50272 28425 50288 se
rect 28425 50272 28502 50288
rect 28409 50206 28502 50272
rect 28409 50104 28502 50170
tri 28409 50088 28425 50104 ne
rect 28425 50088 28502 50104
rect 28242 49989 28390 50071
rect 28130 49956 28207 49972
tri 28207 49956 28223 49972 sw
rect 28130 49890 28223 49956
rect 28259 49831 28373 49989
tri 28409 49956 28425 49972 se
rect 28425 49956 28502 49972
rect 28409 49890 28502 49956
rect 28130 49755 28502 49831
rect 28130 49630 28223 49696
rect 28130 49614 28207 49630
tri 28207 49614 28223 49630 nw
rect 28259 49597 28373 49755
rect 28409 49630 28502 49696
tri 28409 49614 28425 49630 ne
rect 28425 49614 28502 49630
rect 28242 49515 28390 49597
rect 28130 49482 28207 49498
tri 28207 49482 28223 49498 sw
rect 28130 49416 28223 49482
rect 28130 49314 28223 49380
rect 28130 49298 28207 49314
tri 28207 49298 28223 49314 nw
rect 28259 49281 28373 49515
tri 28409 49482 28425 49498 se
rect 28425 49482 28502 49498
rect 28409 49416 28502 49482
rect 28409 49314 28502 49380
tri 28409 49298 28425 49314 ne
rect 28425 49298 28502 49314
rect 28242 49199 28390 49281
rect 28130 49166 28207 49182
tri 28207 49166 28223 49182 sw
rect 28130 49100 28223 49166
rect 28259 49041 28373 49199
tri 28409 49166 28425 49182 se
rect 28425 49166 28502 49182
rect 28409 49100 28502 49166
rect 28130 48965 28502 49041
rect 28130 48840 28223 48906
rect 28130 48824 28207 48840
tri 28207 48824 28223 48840 nw
rect 28259 48807 28373 48965
rect 28409 48840 28502 48906
tri 28409 48824 28425 48840 ne
rect 28425 48824 28502 48840
rect 28242 48725 28390 48807
rect 28130 48692 28207 48708
tri 28207 48692 28223 48708 sw
rect 28130 48626 28223 48692
rect 28130 48524 28223 48590
rect 28130 48508 28207 48524
tri 28207 48508 28223 48524 nw
rect 28259 48491 28373 48725
tri 28409 48692 28425 48708 se
rect 28425 48692 28502 48708
rect 28409 48626 28502 48692
rect 28409 48524 28502 48590
tri 28409 48508 28425 48524 ne
rect 28425 48508 28502 48524
rect 28242 48409 28390 48491
rect 28130 48376 28207 48392
tri 28207 48376 28223 48392 sw
rect 28130 48310 28223 48376
rect 28259 48251 28373 48409
tri 28409 48376 28425 48392 se
rect 28425 48376 28502 48392
rect 28409 48310 28502 48376
rect 28130 48175 28502 48251
rect 28130 48050 28223 48116
rect 28130 48034 28207 48050
tri 28207 48034 28223 48050 nw
rect 28259 48017 28373 48175
rect 28409 48050 28502 48116
tri 28409 48034 28425 48050 ne
rect 28425 48034 28502 48050
rect 28242 47935 28390 48017
rect 28130 47902 28207 47918
tri 28207 47902 28223 47918 sw
rect 28130 47836 28223 47902
rect 28130 47734 28223 47800
rect 28130 47718 28207 47734
tri 28207 47718 28223 47734 nw
rect 28259 47701 28373 47935
tri 28409 47902 28425 47918 se
rect 28425 47902 28502 47918
rect 28409 47836 28502 47902
rect 28409 47734 28502 47800
tri 28409 47718 28425 47734 ne
rect 28425 47718 28502 47734
rect 28242 47619 28390 47701
rect 28130 47586 28207 47602
tri 28207 47586 28223 47602 sw
rect 28130 47520 28223 47586
rect 28259 47461 28373 47619
tri 28409 47586 28425 47602 se
rect 28425 47586 28502 47602
rect 28409 47520 28502 47586
rect 28130 47385 28502 47461
rect 28130 47260 28223 47326
rect 28130 47244 28207 47260
tri 28207 47244 28223 47260 nw
rect 28259 47227 28373 47385
rect 28409 47260 28502 47326
tri 28409 47244 28425 47260 ne
rect 28425 47244 28502 47260
rect 28242 47145 28390 47227
rect 28130 47112 28207 47128
tri 28207 47112 28223 47128 sw
rect 28130 47046 28223 47112
rect 28130 46944 28223 47010
rect 28130 46928 28207 46944
tri 28207 46928 28223 46944 nw
rect 28259 46911 28373 47145
tri 28409 47112 28425 47128 se
rect 28425 47112 28502 47128
rect 28409 47046 28502 47112
rect 28409 46944 28502 47010
tri 28409 46928 28425 46944 ne
rect 28425 46928 28502 46944
rect 28242 46829 28390 46911
rect 28130 46796 28207 46812
tri 28207 46796 28223 46812 sw
rect 28130 46730 28223 46796
rect 28259 46671 28373 46829
tri 28409 46796 28425 46812 se
rect 28425 46796 28502 46812
rect 28409 46730 28502 46796
rect 28130 46595 28502 46671
rect 28130 46470 28223 46536
rect 28130 46454 28207 46470
tri 28207 46454 28223 46470 nw
rect 28259 46437 28373 46595
rect 28409 46470 28502 46536
tri 28409 46454 28425 46470 ne
rect 28425 46454 28502 46470
rect 28242 46355 28390 46437
rect 28130 46322 28207 46338
tri 28207 46322 28223 46338 sw
rect 28130 46256 28223 46322
rect 28130 46154 28223 46220
rect 28130 46138 28207 46154
tri 28207 46138 28223 46154 nw
rect 28259 46121 28373 46355
tri 28409 46322 28425 46338 se
rect 28425 46322 28502 46338
rect 28409 46256 28502 46322
rect 28409 46154 28502 46220
tri 28409 46138 28425 46154 ne
rect 28425 46138 28502 46154
rect 28242 46039 28390 46121
rect 28130 46006 28207 46022
tri 28207 46006 28223 46022 sw
rect 28130 45940 28223 46006
rect 28259 45881 28373 46039
tri 28409 46006 28425 46022 se
rect 28425 46006 28502 46022
rect 28409 45940 28502 46006
rect 28130 45805 28502 45881
rect 28130 45680 28223 45746
rect 28130 45664 28207 45680
tri 28207 45664 28223 45680 nw
rect 28259 45647 28373 45805
rect 28409 45680 28502 45746
tri 28409 45664 28425 45680 ne
rect 28425 45664 28502 45680
rect 28242 45565 28390 45647
rect 28130 45532 28207 45548
tri 28207 45532 28223 45548 sw
rect 28130 45466 28223 45532
rect 28130 45364 28223 45430
rect 28130 45348 28207 45364
tri 28207 45348 28223 45364 nw
rect 28259 45331 28373 45565
tri 28409 45532 28425 45548 se
rect 28425 45532 28502 45548
rect 28409 45466 28502 45532
rect 28409 45364 28502 45430
tri 28409 45348 28425 45364 ne
rect 28425 45348 28502 45364
rect 28242 45249 28390 45331
rect 28130 45216 28207 45232
tri 28207 45216 28223 45232 sw
rect 28130 45150 28223 45216
rect 28259 45091 28373 45249
tri 28409 45216 28425 45232 se
rect 28425 45216 28502 45232
rect 28409 45150 28502 45216
rect 28130 45015 28502 45091
rect 28130 44890 28223 44956
rect 28130 44874 28207 44890
tri 28207 44874 28223 44890 nw
rect 28259 44857 28373 45015
rect 28409 44890 28502 44956
tri 28409 44874 28425 44890 ne
rect 28425 44874 28502 44890
rect 28242 44775 28390 44857
rect 28130 44742 28207 44758
tri 28207 44742 28223 44758 sw
rect 28130 44676 28223 44742
rect 28130 44574 28223 44640
rect 28130 44558 28207 44574
tri 28207 44558 28223 44574 nw
rect 28259 44541 28373 44775
tri 28409 44742 28425 44758 se
rect 28425 44742 28502 44758
rect 28409 44676 28502 44742
rect 28409 44574 28502 44640
tri 28409 44558 28425 44574 ne
rect 28425 44558 28502 44574
rect 28242 44459 28390 44541
rect 28130 44426 28207 44442
tri 28207 44426 28223 44442 sw
rect 28130 44360 28223 44426
rect 28259 44301 28373 44459
tri 28409 44426 28425 44442 se
rect 28425 44426 28502 44442
rect 28409 44360 28502 44426
rect 28130 44225 28502 44301
rect 28130 44100 28223 44166
rect 28130 44084 28207 44100
tri 28207 44084 28223 44100 nw
rect 28259 44067 28373 44225
rect 28409 44100 28502 44166
tri 28409 44084 28425 44100 ne
rect 28425 44084 28502 44100
rect 28242 43985 28390 44067
rect 28130 43952 28207 43968
tri 28207 43952 28223 43968 sw
rect 28130 43886 28223 43952
rect 28130 43784 28223 43850
rect 28130 43768 28207 43784
tri 28207 43768 28223 43784 nw
rect 28259 43751 28373 43985
tri 28409 43952 28425 43968 se
rect 28425 43952 28502 43968
rect 28409 43886 28502 43952
rect 28409 43784 28502 43850
tri 28409 43768 28425 43784 ne
rect 28425 43768 28502 43784
rect 28242 43669 28390 43751
rect 28130 43636 28207 43652
tri 28207 43636 28223 43652 sw
rect 28130 43570 28223 43636
rect 28259 43511 28373 43669
tri 28409 43636 28425 43652 se
rect 28425 43636 28502 43652
rect 28409 43570 28502 43636
rect 28130 43435 28502 43511
rect 28130 43310 28223 43376
rect 28130 43294 28207 43310
tri 28207 43294 28223 43310 nw
rect 28259 43277 28373 43435
rect 28409 43310 28502 43376
tri 28409 43294 28425 43310 ne
rect 28425 43294 28502 43310
rect 28242 43195 28390 43277
rect 28130 43162 28207 43178
tri 28207 43162 28223 43178 sw
rect 28130 43096 28223 43162
rect 28130 42994 28223 43060
rect 28130 42978 28207 42994
tri 28207 42978 28223 42994 nw
rect 28259 42961 28373 43195
tri 28409 43162 28425 43178 se
rect 28425 43162 28502 43178
rect 28409 43096 28502 43162
rect 28409 42994 28502 43060
tri 28409 42978 28425 42994 ne
rect 28425 42978 28502 42994
rect 28242 42879 28390 42961
rect 28130 42846 28207 42862
tri 28207 42846 28223 42862 sw
rect 28130 42780 28223 42846
rect 28259 42721 28373 42879
tri 28409 42846 28425 42862 se
rect 28425 42846 28502 42862
rect 28409 42780 28502 42846
rect 28130 42645 28502 42721
rect 28130 42520 28223 42586
rect 28130 42504 28207 42520
tri 28207 42504 28223 42520 nw
rect 28259 42487 28373 42645
rect 28409 42520 28502 42586
tri 28409 42504 28425 42520 ne
rect 28425 42504 28502 42520
rect 28242 42405 28390 42487
rect 28130 42372 28207 42388
tri 28207 42372 28223 42388 sw
rect 28130 42306 28223 42372
rect 28130 42204 28223 42270
rect 28130 42188 28207 42204
tri 28207 42188 28223 42204 nw
rect 28259 42171 28373 42405
tri 28409 42372 28425 42388 se
rect 28425 42372 28502 42388
rect 28409 42306 28502 42372
rect 28409 42204 28502 42270
tri 28409 42188 28425 42204 ne
rect 28425 42188 28502 42204
rect 28242 42089 28390 42171
rect 28130 42056 28207 42072
tri 28207 42056 28223 42072 sw
rect 28130 41990 28223 42056
rect 28259 41931 28373 42089
tri 28409 42056 28425 42072 se
rect 28425 42056 28502 42072
rect 28409 41990 28502 42056
rect 28130 41855 28502 41931
rect 28130 41730 28223 41796
rect 28130 41714 28207 41730
tri 28207 41714 28223 41730 nw
rect 28259 41697 28373 41855
rect 28409 41730 28502 41796
tri 28409 41714 28425 41730 ne
rect 28425 41714 28502 41730
rect 28242 41615 28390 41697
rect 28130 41582 28207 41598
tri 28207 41582 28223 41598 sw
rect 28130 41516 28223 41582
rect 28130 41414 28223 41480
rect 28130 41398 28207 41414
tri 28207 41398 28223 41414 nw
rect 28259 41381 28373 41615
tri 28409 41582 28425 41598 se
rect 28425 41582 28502 41598
rect 28409 41516 28502 41582
rect 28409 41414 28502 41480
tri 28409 41398 28425 41414 ne
rect 28425 41398 28502 41414
rect 28242 41299 28390 41381
rect 28130 41266 28207 41282
tri 28207 41266 28223 41282 sw
rect 28130 41200 28223 41266
rect 28259 41141 28373 41299
tri 28409 41266 28425 41282 se
rect 28425 41266 28502 41282
rect 28409 41200 28502 41266
rect 28130 41065 28502 41141
rect 28130 40940 28223 41006
rect 28130 40924 28207 40940
tri 28207 40924 28223 40940 nw
rect 28259 40907 28373 41065
rect 28409 40940 28502 41006
tri 28409 40924 28425 40940 ne
rect 28425 40924 28502 40940
rect 28242 40825 28390 40907
rect 28130 40792 28207 40808
tri 28207 40792 28223 40808 sw
rect 28130 40726 28223 40792
rect 28130 40624 28223 40690
rect 28130 40608 28207 40624
tri 28207 40608 28223 40624 nw
rect 28259 40591 28373 40825
tri 28409 40792 28425 40808 se
rect 28425 40792 28502 40808
rect 28409 40726 28502 40792
rect 28409 40624 28502 40690
tri 28409 40608 28425 40624 ne
rect 28425 40608 28502 40624
rect 28242 40509 28390 40591
rect 28130 40476 28207 40492
tri 28207 40476 28223 40492 sw
rect 28130 40410 28223 40476
rect 28259 40351 28373 40509
tri 28409 40476 28425 40492 se
rect 28425 40476 28502 40492
rect 28409 40410 28502 40476
rect 28130 40275 28502 40351
rect 28130 40150 28223 40216
rect 28130 40134 28207 40150
tri 28207 40134 28223 40150 nw
rect 28259 40117 28373 40275
rect 28409 40150 28502 40216
tri 28409 40134 28425 40150 ne
rect 28425 40134 28502 40150
rect 28242 40035 28390 40117
rect 28130 40002 28207 40018
tri 28207 40002 28223 40018 sw
rect 28130 39936 28223 40002
rect 28130 39834 28223 39900
rect 28130 39818 28207 39834
tri 28207 39818 28223 39834 nw
rect 28259 39801 28373 40035
tri 28409 40002 28425 40018 se
rect 28425 40002 28502 40018
rect 28409 39936 28502 40002
rect 28409 39834 28502 39900
tri 28409 39818 28425 39834 ne
rect 28425 39818 28502 39834
rect 28242 39719 28390 39801
rect 28130 39686 28207 39702
tri 28207 39686 28223 39702 sw
rect 28130 39620 28223 39686
rect 28259 39561 28373 39719
tri 28409 39686 28425 39702 se
rect 28425 39686 28502 39702
rect 28409 39620 28502 39686
rect 28130 39485 28502 39561
rect 28130 39360 28223 39426
rect 28130 39344 28207 39360
tri 28207 39344 28223 39360 nw
rect 28259 39327 28373 39485
rect 28409 39360 28502 39426
tri 28409 39344 28425 39360 ne
rect 28425 39344 28502 39360
rect 28242 39245 28390 39327
rect 28130 39212 28207 39228
tri 28207 39212 28223 39228 sw
rect 28130 39146 28223 39212
rect 28130 39044 28223 39110
rect 28130 39028 28207 39044
tri 28207 39028 28223 39044 nw
rect 28259 39011 28373 39245
tri 28409 39212 28425 39228 se
rect 28425 39212 28502 39228
rect 28409 39146 28502 39212
rect 28409 39044 28502 39110
tri 28409 39028 28425 39044 ne
rect 28425 39028 28502 39044
rect 28242 38929 28390 39011
rect 28130 38896 28207 38912
tri 28207 38896 28223 38912 sw
rect 28130 38830 28223 38896
rect 28259 38771 28373 38929
tri 28409 38896 28425 38912 se
rect 28425 38896 28502 38912
rect 28409 38830 28502 38896
rect 28130 38695 28502 38771
rect 28130 38570 28223 38636
rect 28130 38554 28207 38570
tri 28207 38554 28223 38570 nw
rect 28259 38537 28373 38695
rect 28409 38570 28502 38636
tri 28409 38554 28425 38570 ne
rect 28425 38554 28502 38570
rect 28242 38455 28390 38537
rect 28130 38422 28207 38438
tri 28207 38422 28223 38438 sw
rect 28130 38356 28223 38422
rect 28130 38254 28223 38320
rect 28130 38238 28207 38254
tri 28207 38238 28223 38254 nw
rect 28259 38221 28373 38455
tri 28409 38422 28425 38438 se
rect 28425 38422 28502 38438
rect 28409 38356 28502 38422
rect 28409 38254 28502 38320
tri 28409 38238 28425 38254 ne
rect 28425 38238 28502 38254
rect 28242 38139 28390 38221
rect 28130 38106 28207 38122
tri 28207 38106 28223 38122 sw
rect 28130 38040 28223 38106
rect 28259 37981 28373 38139
tri 28409 38106 28425 38122 se
rect 28425 38106 28502 38122
rect 28409 38040 28502 38106
rect 28130 37905 28502 37981
rect 28130 37780 28223 37846
rect 28130 37764 28207 37780
tri 28207 37764 28223 37780 nw
rect 28259 37747 28373 37905
rect 28409 37780 28502 37846
tri 28409 37764 28425 37780 ne
rect 28425 37764 28502 37780
rect 28242 37665 28390 37747
rect 28130 37632 28207 37648
tri 28207 37632 28223 37648 sw
rect 28130 37566 28223 37632
rect 28130 37464 28223 37530
rect 28130 37448 28207 37464
tri 28207 37448 28223 37464 nw
rect 28259 37431 28373 37665
tri 28409 37632 28425 37648 se
rect 28425 37632 28502 37648
rect 28409 37566 28502 37632
rect 28409 37464 28502 37530
tri 28409 37448 28425 37464 ne
rect 28425 37448 28502 37464
rect 28242 37349 28390 37431
rect 28130 37316 28207 37332
tri 28207 37316 28223 37332 sw
rect 28130 37250 28223 37316
rect 28259 37191 28373 37349
tri 28409 37316 28425 37332 se
rect 28425 37316 28502 37332
rect 28409 37250 28502 37316
rect 28130 37115 28502 37191
rect 28130 36990 28223 37056
rect 28130 36974 28207 36990
tri 28207 36974 28223 36990 nw
rect 28259 36957 28373 37115
rect 28409 36990 28502 37056
tri 28409 36974 28425 36990 ne
rect 28425 36974 28502 36990
rect 28242 36875 28390 36957
rect 28130 36842 28207 36858
tri 28207 36842 28223 36858 sw
rect 28130 36776 28223 36842
rect 28130 36674 28223 36740
rect 28130 36658 28207 36674
tri 28207 36658 28223 36674 nw
rect 28259 36641 28373 36875
tri 28409 36842 28425 36858 se
rect 28425 36842 28502 36858
rect 28409 36776 28502 36842
rect 28409 36674 28502 36740
tri 28409 36658 28425 36674 ne
rect 28425 36658 28502 36674
rect 28242 36559 28390 36641
rect 28130 36526 28207 36542
tri 28207 36526 28223 36542 sw
rect 28130 36460 28223 36526
rect 28259 36401 28373 36559
tri 28409 36526 28425 36542 se
rect 28425 36526 28502 36542
rect 28409 36460 28502 36526
rect 28130 36325 28502 36401
rect 28130 36200 28223 36266
rect 28130 36184 28207 36200
tri 28207 36184 28223 36200 nw
rect 28259 36167 28373 36325
rect 28409 36200 28502 36266
tri 28409 36184 28425 36200 ne
rect 28425 36184 28502 36200
rect 28242 36085 28390 36167
rect 28130 36052 28207 36068
tri 28207 36052 28223 36068 sw
rect 28130 35986 28223 36052
rect 28130 35884 28223 35950
rect 28130 35868 28207 35884
tri 28207 35868 28223 35884 nw
rect 28259 35851 28373 36085
tri 28409 36052 28425 36068 se
rect 28425 36052 28502 36068
rect 28409 35986 28502 36052
rect 28409 35884 28502 35950
tri 28409 35868 28425 35884 ne
rect 28425 35868 28502 35884
rect 28242 35769 28390 35851
rect 28130 35736 28207 35752
tri 28207 35736 28223 35752 sw
rect 28130 35670 28223 35736
rect 28259 35611 28373 35769
tri 28409 35736 28425 35752 se
rect 28425 35736 28502 35752
rect 28409 35670 28502 35736
rect 28130 35535 28502 35611
rect 28130 35410 28223 35476
rect 28130 35394 28207 35410
tri 28207 35394 28223 35410 nw
rect 28259 35377 28373 35535
rect 28409 35410 28502 35476
tri 28409 35394 28425 35410 ne
rect 28425 35394 28502 35410
rect 28242 35295 28390 35377
rect 28130 35262 28207 35278
tri 28207 35262 28223 35278 sw
rect 28130 35196 28223 35262
rect 28130 35094 28223 35160
rect 28130 35078 28207 35094
tri 28207 35078 28223 35094 nw
rect 28259 35061 28373 35295
tri 28409 35262 28425 35278 se
rect 28425 35262 28502 35278
rect 28409 35196 28502 35262
rect 28409 35094 28502 35160
tri 28409 35078 28425 35094 ne
rect 28425 35078 28502 35094
rect 28242 34979 28390 35061
rect 28130 34946 28207 34962
tri 28207 34946 28223 34962 sw
rect 28130 34880 28223 34946
rect 28259 34821 28373 34979
tri 28409 34946 28425 34962 se
rect 28425 34946 28502 34962
rect 28409 34880 28502 34946
rect 28130 34745 28502 34821
rect 28130 34620 28223 34686
rect 28130 34604 28207 34620
tri 28207 34604 28223 34620 nw
rect 28259 34587 28373 34745
rect 28409 34620 28502 34686
tri 28409 34604 28425 34620 ne
rect 28425 34604 28502 34620
rect 28242 34505 28390 34587
rect 28130 34472 28207 34488
tri 28207 34472 28223 34488 sw
rect 28130 34406 28223 34472
rect 28130 34304 28223 34370
rect 28130 34288 28207 34304
tri 28207 34288 28223 34304 nw
rect 28259 34271 28373 34505
tri 28409 34472 28425 34488 se
rect 28425 34472 28502 34488
rect 28409 34406 28502 34472
rect 28409 34304 28502 34370
tri 28409 34288 28425 34304 ne
rect 28425 34288 28502 34304
rect 28242 34189 28390 34271
rect 28130 34156 28207 34172
tri 28207 34156 28223 34172 sw
rect 28130 34090 28223 34156
rect 28259 34031 28373 34189
tri 28409 34156 28425 34172 se
rect 28425 34156 28502 34172
rect 28409 34090 28502 34156
rect 28130 33955 28502 34031
rect 28130 33830 28223 33896
rect 28130 33814 28207 33830
tri 28207 33814 28223 33830 nw
rect 28259 33797 28373 33955
rect 28409 33830 28502 33896
tri 28409 33814 28425 33830 ne
rect 28425 33814 28502 33830
rect 28242 33715 28390 33797
rect 28130 33682 28207 33698
tri 28207 33682 28223 33698 sw
rect 28130 33616 28223 33682
rect 28130 33514 28223 33580
rect 28130 33498 28207 33514
tri 28207 33498 28223 33514 nw
rect 28259 33481 28373 33715
tri 28409 33682 28425 33698 se
rect 28425 33682 28502 33698
rect 28409 33616 28502 33682
rect 28409 33514 28502 33580
tri 28409 33498 28425 33514 ne
rect 28425 33498 28502 33514
rect 28242 33399 28390 33481
rect 28130 33366 28207 33382
tri 28207 33366 28223 33382 sw
rect 28130 33300 28223 33366
rect 28259 33241 28373 33399
tri 28409 33366 28425 33382 se
rect 28425 33366 28502 33382
rect 28409 33300 28502 33366
rect 28130 33165 28502 33241
rect 28130 33040 28223 33106
rect 28130 33024 28207 33040
tri 28207 33024 28223 33040 nw
rect 28259 33007 28373 33165
rect 28409 33040 28502 33106
tri 28409 33024 28425 33040 ne
rect 28425 33024 28502 33040
rect 28242 32925 28390 33007
rect 28130 32892 28207 32908
tri 28207 32892 28223 32908 sw
rect 28130 32826 28223 32892
rect 28130 32724 28223 32790
rect 28130 32708 28207 32724
tri 28207 32708 28223 32724 nw
rect 28259 32691 28373 32925
tri 28409 32892 28425 32908 se
rect 28425 32892 28502 32908
rect 28409 32826 28502 32892
rect 28409 32724 28502 32790
tri 28409 32708 28425 32724 ne
rect 28425 32708 28502 32724
rect 28242 32609 28390 32691
rect 28130 32576 28207 32592
tri 28207 32576 28223 32592 sw
rect 28130 32510 28223 32576
rect 28259 32451 28373 32609
tri 28409 32576 28425 32592 se
rect 28425 32576 28502 32592
rect 28409 32510 28502 32576
rect 28130 32375 28502 32451
rect 28130 32250 28223 32316
rect 28130 32234 28207 32250
tri 28207 32234 28223 32250 nw
rect 28259 32217 28373 32375
rect 28409 32250 28502 32316
tri 28409 32234 28425 32250 ne
rect 28425 32234 28502 32250
rect 28242 32135 28390 32217
rect 28130 32102 28207 32118
tri 28207 32102 28223 32118 sw
rect 28130 32036 28223 32102
rect 28130 31934 28223 32000
rect 28130 31918 28207 31934
tri 28207 31918 28223 31934 nw
rect 28259 31901 28373 32135
tri 28409 32102 28425 32118 se
rect 28425 32102 28502 32118
rect 28409 32036 28502 32102
rect 28409 31934 28502 32000
tri 28409 31918 28425 31934 ne
rect 28425 31918 28502 31934
rect 28242 31819 28390 31901
rect 28130 31786 28207 31802
tri 28207 31786 28223 31802 sw
rect 28130 31720 28223 31786
rect 28259 31661 28373 31819
tri 28409 31786 28425 31802 se
rect 28425 31786 28502 31802
rect 28409 31720 28502 31786
rect 28130 31585 28502 31661
rect 28130 31460 28223 31526
rect 28130 31444 28207 31460
tri 28207 31444 28223 31460 nw
rect 28259 31427 28373 31585
rect 28409 31460 28502 31526
tri 28409 31444 28425 31460 ne
rect 28425 31444 28502 31460
rect 28242 31345 28390 31427
rect 28130 31312 28207 31328
tri 28207 31312 28223 31328 sw
rect 28130 31246 28223 31312
rect 28130 31144 28223 31210
rect 28130 31128 28207 31144
tri 28207 31128 28223 31144 nw
rect 28259 31111 28373 31345
tri 28409 31312 28425 31328 se
rect 28425 31312 28502 31328
rect 28409 31246 28502 31312
rect 28409 31144 28502 31210
tri 28409 31128 28425 31144 ne
rect 28425 31128 28502 31144
rect 28242 31029 28390 31111
rect 28130 30996 28207 31012
tri 28207 30996 28223 31012 sw
rect 28130 30930 28223 30996
rect 28259 30871 28373 31029
tri 28409 30996 28425 31012 se
rect 28425 30996 28502 31012
rect 28409 30930 28502 30996
rect 28130 30795 28502 30871
rect 28130 30670 28223 30736
rect 28130 30654 28207 30670
tri 28207 30654 28223 30670 nw
rect 28259 30637 28373 30795
rect 28409 30670 28502 30736
tri 28409 30654 28425 30670 ne
rect 28425 30654 28502 30670
rect 28242 30555 28390 30637
rect 28130 30522 28207 30538
tri 28207 30522 28223 30538 sw
rect 28130 30456 28223 30522
rect 28130 30354 28223 30420
rect 28130 30338 28207 30354
tri 28207 30338 28223 30354 nw
rect 28259 30321 28373 30555
tri 28409 30522 28425 30538 se
rect 28425 30522 28502 30538
rect 28409 30456 28502 30522
rect 28409 30354 28502 30420
tri 28409 30338 28425 30354 ne
rect 28425 30338 28502 30354
rect 28242 30239 28390 30321
rect 28130 30206 28207 30222
tri 28207 30206 28223 30222 sw
rect 28130 30140 28223 30206
rect 28259 30081 28373 30239
tri 28409 30206 28425 30222 se
rect 28425 30206 28502 30222
rect 28409 30140 28502 30206
rect 28130 30005 28502 30081
rect 28130 29880 28223 29946
rect 28130 29864 28207 29880
tri 28207 29864 28223 29880 nw
rect 28259 29847 28373 30005
rect 28409 29880 28502 29946
tri 28409 29864 28425 29880 ne
rect 28425 29864 28502 29880
rect 28242 29765 28390 29847
rect 28130 29732 28207 29748
tri 28207 29732 28223 29748 sw
rect 28130 29666 28223 29732
rect 28130 29564 28223 29630
rect 28130 29548 28207 29564
tri 28207 29548 28223 29564 nw
rect 28259 29531 28373 29765
tri 28409 29732 28425 29748 se
rect 28425 29732 28502 29748
rect 28409 29666 28502 29732
rect 28409 29564 28502 29630
tri 28409 29548 28425 29564 ne
rect 28425 29548 28502 29564
rect 28242 29449 28390 29531
rect 28130 29416 28207 29432
tri 28207 29416 28223 29432 sw
rect 28130 29350 28223 29416
rect 28259 29291 28373 29449
tri 28409 29416 28425 29432 se
rect 28425 29416 28502 29432
rect 28409 29350 28502 29416
rect 28130 29215 28502 29291
rect 28130 29090 28223 29156
rect 28130 29074 28207 29090
tri 28207 29074 28223 29090 nw
rect 28259 29057 28373 29215
rect 28409 29090 28502 29156
tri 28409 29074 28425 29090 ne
rect 28425 29074 28502 29090
rect 28242 28975 28390 29057
rect 28130 28942 28207 28958
tri 28207 28942 28223 28958 sw
rect 28130 28876 28223 28942
rect 28259 28833 28373 28975
tri 28409 28942 28425 28958 se
rect 28425 28942 28502 28958
rect 28409 28876 28502 28942
rect 28538 28463 28574 80603
rect 28610 28463 28646 80603
rect 28682 80445 28718 80603
rect 28674 80303 28726 80445
rect 28682 28763 28718 80303
rect 28674 28621 28726 28763
rect 28682 28463 28718 28621
rect 28754 28463 28790 80603
rect 28826 28463 28862 80603
rect 28898 28833 28982 80233
rect 29018 28463 29054 80603
rect 29090 28463 29126 80603
rect 29162 80445 29198 80603
rect 29154 80303 29206 80445
rect 29162 28763 29198 80303
rect 29154 28621 29206 28763
rect 29162 28463 29198 28621
rect 29234 28463 29270 80603
rect 29306 28463 29342 80603
rect 29378 80124 29471 80190
rect 29378 80108 29455 80124
tri 29455 80108 29471 80124 nw
rect 29507 80091 29621 80233
rect 29657 80124 29750 80190
tri 29657 80108 29673 80124 ne
rect 29673 80108 29750 80124
rect 29490 80009 29638 80091
rect 29378 79976 29455 79992
tri 29455 79976 29471 79992 sw
rect 29378 79910 29471 79976
rect 29507 79851 29621 80009
tri 29657 79976 29673 79992 se
rect 29673 79976 29750 79992
rect 29657 79910 29750 79976
rect 29378 79775 29750 79851
rect 29378 79650 29471 79716
rect 29378 79634 29455 79650
tri 29455 79634 29471 79650 nw
rect 29507 79617 29621 79775
rect 29657 79650 29750 79716
tri 29657 79634 29673 79650 ne
rect 29673 79634 29750 79650
rect 29490 79535 29638 79617
rect 29378 79502 29455 79518
tri 29455 79502 29471 79518 sw
rect 29378 79436 29471 79502
rect 29378 79334 29471 79400
rect 29378 79318 29455 79334
tri 29455 79318 29471 79334 nw
rect 29507 79301 29621 79535
tri 29657 79502 29673 79518 se
rect 29673 79502 29750 79518
rect 29657 79436 29750 79502
rect 29657 79334 29750 79400
tri 29657 79318 29673 79334 ne
rect 29673 79318 29750 79334
rect 29490 79219 29638 79301
rect 29378 79186 29455 79202
tri 29455 79186 29471 79202 sw
rect 29378 79120 29471 79186
rect 29507 79061 29621 79219
tri 29657 79186 29673 79202 se
rect 29673 79186 29750 79202
rect 29657 79120 29750 79186
rect 29378 78985 29750 79061
rect 29378 78860 29471 78926
rect 29378 78844 29455 78860
tri 29455 78844 29471 78860 nw
rect 29507 78827 29621 78985
rect 29657 78860 29750 78926
tri 29657 78844 29673 78860 ne
rect 29673 78844 29750 78860
rect 29490 78745 29638 78827
rect 29378 78712 29455 78728
tri 29455 78712 29471 78728 sw
rect 29378 78646 29471 78712
rect 29378 78544 29471 78610
rect 29378 78528 29455 78544
tri 29455 78528 29471 78544 nw
rect 29507 78511 29621 78745
tri 29657 78712 29673 78728 se
rect 29673 78712 29750 78728
rect 29657 78646 29750 78712
rect 29657 78544 29750 78610
tri 29657 78528 29673 78544 ne
rect 29673 78528 29750 78544
rect 29490 78429 29638 78511
rect 29378 78396 29455 78412
tri 29455 78396 29471 78412 sw
rect 29378 78330 29471 78396
rect 29507 78271 29621 78429
tri 29657 78396 29673 78412 se
rect 29673 78396 29750 78412
rect 29657 78330 29750 78396
rect 29378 78195 29750 78271
rect 29378 78070 29471 78136
rect 29378 78054 29455 78070
tri 29455 78054 29471 78070 nw
rect 29507 78037 29621 78195
rect 29657 78070 29750 78136
tri 29657 78054 29673 78070 ne
rect 29673 78054 29750 78070
rect 29490 77955 29638 78037
rect 29378 77922 29455 77938
tri 29455 77922 29471 77938 sw
rect 29378 77856 29471 77922
rect 29378 77754 29471 77820
rect 29378 77738 29455 77754
tri 29455 77738 29471 77754 nw
rect 29507 77721 29621 77955
tri 29657 77922 29673 77938 se
rect 29673 77922 29750 77938
rect 29657 77856 29750 77922
rect 29657 77754 29750 77820
tri 29657 77738 29673 77754 ne
rect 29673 77738 29750 77754
rect 29490 77639 29638 77721
rect 29378 77606 29455 77622
tri 29455 77606 29471 77622 sw
rect 29378 77540 29471 77606
rect 29507 77481 29621 77639
tri 29657 77606 29673 77622 se
rect 29673 77606 29750 77622
rect 29657 77540 29750 77606
rect 29378 77405 29750 77481
rect 29378 77280 29471 77346
rect 29378 77264 29455 77280
tri 29455 77264 29471 77280 nw
rect 29507 77247 29621 77405
rect 29657 77280 29750 77346
tri 29657 77264 29673 77280 ne
rect 29673 77264 29750 77280
rect 29490 77165 29638 77247
rect 29378 77132 29455 77148
tri 29455 77132 29471 77148 sw
rect 29378 77066 29471 77132
rect 29378 76964 29471 77030
rect 29378 76948 29455 76964
tri 29455 76948 29471 76964 nw
rect 29507 76931 29621 77165
tri 29657 77132 29673 77148 se
rect 29673 77132 29750 77148
rect 29657 77066 29750 77132
rect 29657 76964 29750 77030
tri 29657 76948 29673 76964 ne
rect 29673 76948 29750 76964
rect 29490 76849 29638 76931
rect 29378 76816 29455 76832
tri 29455 76816 29471 76832 sw
rect 29378 76750 29471 76816
rect 29507 76691 29621 76849
tri 29657 76816 29673 76832 se
rect 29673 76816 29750 76832
rect 29657 76750 29750 76816
rect 29378 76615 29750 76691
rect 29378 76490 29471 76556
rect 29378 76474 29455 76490
tri 29455 76474 29471 76490 nw
rect 29507 76457 29621 76615
rect 29657 76490 29750 76556
tri 29657 76474 29673 76490 ne
rect 29673 76474 29750 76490
rect 29490 76375 29638 76457
rect 29378 76342 29455 76358
tri 29455 76342 29471 76358 sw
rect 29378 76276 29471 76342
rect 29378 76174 29471 76240
rect 29378 76158 29455 76174
tri 29455 76158 29471 76174 nw
rect 29507 76141 29621 76375
tri 29657 76342 29673 76358 se
rect 29673 76342 29750 76358
rect 29657 76276 29750 76342
rect 29657 76174 29750 76240
tri 29657 76158 29673 76174 ne
rect 29673 76158 29750 76174
rect 29490 76059 29638 76141
rect 29378 76026 29455 76042
tri 29455 76026 29471 76042 sw
rect 29378 75960 29471 76026
rect 29507 75901 29621 76059
tri 29657 76026 29673 76042 se
rect 29673 76026 29750 76042
rect 29657 75960 29750 76026
rect 29378 75825 29750 75901
rect 29378 75700 29471 75766
rect 29378 75684 29455 75700
tri 29455 75684 29471 75700 nw
rect 29507 75667 29621 75825
rect 29657 75700 29750 75766
tri 29657 75684 29673 75700 ne
rect 29673 75684 29750 75700
rect 29490 75585 29638 75667
rect 29378 75552 29455 75568
tri 29455 75552 29471 75568 sw
rect 29378 75486 29471 75552
rect 29378 75384 29471 75450
rect 29378 75368 29455 75384
tri 29455 75368 29471 75384 nw
rect 29507 75351 29621 75585
tri 29657 75552 29673 75568 se
rect 29673 75552 29750 75568
rect 29657 75486 29750 75552
rect 29657 75384 29750 75450
tri 29657 75368 29673 75384 ne
rect 29673 75368 29750 75384
rect 29490 75269 29638 75351
rect 29378 75236 29455 75252
tri 29455 75236 29471 75252 sw
rect 29378 75170 29471 75236
rect 29507 75111 29621 75269
tri 29657 75236 29673 75252 se
rect 29673 75236 29750 75252
rect 29657 75170 29750 75236
rect 29378 75035 29750 75111
rect 29378 74910 29471 74976
rect 29378 74894 29455 74910
tri 29455 74894 29471 74910 nw
rect 29507 74877 29621 75035
rect 29657 74910 29750 74976
tri 29657 74894 29673 74910 ne
rect 29673 74894 29750 74910
rect 29490 74795 29638 74877
rect 29378 74762 29455 74778
tri 29455 74762 29471 74778 sw
rect 29378 74696 29471 74762
rect 29378 74594 29471 74660
rect 29378 74578 29455 74594
tri 29455 74578 29471 74594 nw
rect 29507 74561 29621 74795
tri 29657 74762 29673 74778 se
rect 29673 74762 29750 74778
rect 29657 74696 29750 74762
rect 29657 74594 29750 74660
tri 29657 74578 29673 74594 ne
rect 29673 74578 29750 74594
rect 29490 74479 29638 74561
rect 29378 74446 29455 74462
tri 29455 74446 29471 74462 sw
rect 29378 74380 29471 74446
rect 29507 74321 29621 74479
tri 29657 74446 29673 74462 se
rect 29673 74446 29750 74462
rect 29657 74380 29750 74446
rect 29378 74245 29750 74321
rect 29378 74120 29471 74186
rect 29378 74104 29455 74120
tri 29455 74104 29471 74120 nw
rect 29507 74087 29621 74245
rect 29657 74120 29750 74186
tri 29657 74104 29673 74120 ne
rect 29673 74104 29750 74120
rect 29490 74005 29638 74087
rect 29378 73972 29455 73988
tri 29455 73972 29471 73988 sw
rect 29378 73906 29471 73972
rect 29378 73804 29471 73870
rect 29378 73788 29455 73804
tri 29455 73788 29471 73804 nw
rect 29507 73771 29621 74005
tri 29657 73972 29673 73988 se
rect 29673 73972 29750 73988
rect 29657 73906 29750 73972
rect 29657 73804 29750 73870
tri 29657 73788 29673 73804 ne
rect 29673 73788 29750 73804
rect 29490 73689 29638 73771
rect 29378 73656 29455 73672
tri 29455 73656 29471 73672 sw
rect 29378 73590 29471 73656
rect 29507 73531 29621 73689
tri 29657 73656 29673 73672 se
rect 29673 73656 29750 73672
rect 29657 73590 29750 73656
rect 29378 73455 29750 73531
rect 29378 73330 29471 73396
rect 29378 73314 29455 73330
tri 29455 73314 29471 73330 nw
rect 29507 73297 29621 73455
rect 29657 73330 29750 73396
tri 29657 73314 29673 73330 ne
rect 29673 73314 29750 73330
rect 29490 73215 29638 73297
rect 29378 73182 29455 73198
tri 29455 73182 29471 73198 sw
rect 29378 73116 29471 73182
rect 29378 73014 29471 73080
rect 29378 72998 29455 73014
tri 29455 72998 29471 73014 nw
rect 29507 72981 29621 73215
tri 29657 73182 29673 73198 se
rect 29673 73182 29750 73198
rect 29657 73116 29750 73182
rect 29657 73014 29750 73080
tri 29657 72998 29673 73014 ne
rect 29673 72998 29750 73014
rect 29490 72899 29638 72981
rect 29378 72866 29455 72882
tri 29455 72866 29471 72882 sw
rect 29378 72800 29471 72866
rect 29507 72741 29621 72899
tri 29657 72866 29673 72882 se
rect 29673 72866 29750 72882
rect 29657 72800 29750 72866
rect 29378 72665 29750 72741
rect 29378 72540 29471 72606
rect 29378 72524 29455 72540
tri 29455 72524 29471 72540 nw
rect 29507 72507 29621 72665
rect 29657 72540 29750 72606
tri 29657 72524 29673 72540 ne
rect 29673 72524 29750 72540
rect 29490 72425 29638 72507
rect 29378 72392 29455 72408
tri 29455 72392 29471 72408 sw
rect 29378 72326 29471 72392
rect 29378 72224 29471 72290
rect 29378 72208 29455 72224
tri 29455 72208 29471 72224 nw
rect 29507 72191 29621 72425
tri 29657 72392 29673 72408 se
rect 29673 72392 29750 72408
rect 29657 72326 29750 72392
rect 29657 72224 29750 72290
tri 29657 72208 29673 72224 ne
rect 29673 72208 29750 72224
rect 29490 72109 29638 72191
rect 29378 72076 29455 72092
tri 29455 72076 29471 72092 sw
rect 29378 72010 29471 72076
rect 29507 71951 29621 72109
tri 29657 72076 29673 72092 se
rect 29673 72076 29750 72092
rect 29657 72010 29750 72076
rect 29378 71875 29750 71951
rect 29378 71750 29471 71816
rect 29378 71734 29455 71750
tri 29455 71734 29471 71750 nw
rect 29507 71717 29621 71875
rect 29657 71750 29750 71816
tri 29657 71734 29673 71750 ne
rect 29673 71734 29750 71750
rect 29490 71635 29638 71717
rect 29378 71602 29455 71618
tri 29455 71602 29471 71618 sw
rect 29378 71536 29471 71602
rect 29378 71434 29471 71500
rect 29378 71418 29455 71434
tri 29455 71418 29471 71434 nw
rect 29507 71401 29621 71635
tri 29657 71602 29673 71618 se
rect 29673 71602 29750 71618
rect 29657 71536 29750 71602
rect 29657 71434 29750 71500
tri 29657 71418 29673 71434 ne
rect 29673 71418 29750 71434
rect 29490 71319 29638 71401
rect 29378 71286 29455 71302
tri 29455 71286 29471 71302 sw
rect 29378 71220 29471 71286
rect 29507 71161 29621 71319
tri 29657 71286 29673 71302 se
rect 29673 71286 29750 71302
rect 29657 71220 29750 71286
rect 29378 71085 29750 71161
rect 29378 70960 29471 71026
rect 29378 70944 29455 70960
tri 29455 70944 29471 70960 nw
rect 29507 70927 29621 71085
rect 29657 70960 29750 71026
tri 29657 70944 29673 70960 ne
rect 29673 70944 29750 70960
rect 29490 70845 29638 70927
rect 29378 70812 29455 70828
tri 29455 70812 29471 70828 sw
rect 29378 70746 29471 70812
rect 29378 70644 29471 70710
rect 29378 70628 29455 70644
tri 29455 70628 29471 70644 nw
rect 29507 70611 29621 70845
tri 29657 70812 29673 70828 se
rect 29673 70812 29750 70828
rect 29657 70746 29750 70812
rect 29657 70644 29750 70710
tri 29657 70628 29673 70644 ne
rect 29673 70628 29750 70644
rect 29490 70529 29638 70611
rect 29378 70496 29455 70512
tri 29455 70496 29471 70512 sw
rect 29378 70430 29471 70496
rect 29507 70371 29621 70529
tri 29657 70496 29673 70512 se
rect 29673 70496 29750 70512
rect 29657 70430 29750 70496
rect 29378 70295 29750 70371
rect 29378 70170 29471 70236
rect 29378 70154 29455 70170
tri 29455 70154 29471 70170 nw
rect 29507 70137 29621 70295
rect 29657 70170 29750 70236
tri 29657 70154 29673 70170 ne
rect 29673 70154 29750 70170
rect 29490 70055 29638 70137
rect 29378 70022 29455 70038
tri 29455 70022 29471 70038 sw
rect 29378 69956 29471 70022
rect 29378 69854 29471 69920
rect 29378 69838 29455 69854
tri 29455 69838 29471 69854 nw
rect 29507 69821 29621 70055
tri 29657 70022 29673 70038 se
rect 29673 70022 29750 70038
rect 29657 69956 29750 70022
rect 29657 69854 29750 69920
tri 29657 69838 29673 69854 ne
rect 29673 69838 29750 69854
rect 29490 69739 29638 69821
rect 29378 69706 29455 69722
tri 29455 69706 29471 69722 sw
rect 29378 69640 29471 69706
rect 29507 69581 29621 69739
tri 29657 69706 29673 69722 se
rect 29673 69706 29750 69722
rect 29657 69640 29750 69706
rect 29378 69505 29750 69581
rect 29378 69380 29471 69446
rect 29378 69364 29455 69380
tri 29455 69364 29471 69380 nw
rect 29507 69347 29621 69505
rect 29657 69380 29750 69446
tri 29657 69364 29673 69380 ne
rect 29673 69364 29750 69380
rect 29490 69265 29638 69347
rect 29378 69232 29455 69248
tri 29455 69232 29471 69248 sw
rect 29378 69166 29471 69232
rect 29378 69064 29471 69130
rect 29378 69048 29455 69064
tri 29455 69048 29471 69064 nw
rect 29507 69031 29621 69265
tri 29657 69232 29673 69248 se
rect 29673 69232 29750 69248
rect 29657 69166 29750 69232
rect 29657 69064 29750 69130
tri 29657 69048 29673 69064 ne
rect 29673 69048 29750 69064
rect 29490 68949 29638 69031
rect 29378 68916 29455 68932
tri 29455 68916 29471 68932 sw
rect 29378 68850 29471 68916
rect 29507 68791 29621 68949
tri 29657 68916 29673 68932 se
rect 29673 68916 29750 68932
rect 29657 68850 29750 68916
rect 29378 68715 29750 68791
rect 29378 68590 29471 68656
rect 29378 68574 29455 68590
tri 29455 68574 29471 68590 nw
rect 29507 68557 29621 68715
rect 29657 68590 29750 68656
tri 29657 68574 29673 68590 ne
rect 29673 68574 29750 68590
rect 29490 68475 29638 68557
rect 29378 68442 29455 68458
tri 29455 68442 29471 68458 sw
rect 29378 68376 29471 68442
rect 29378 68274 29471 68340
rect 29378 68258 29455 68274
tri 29455 68258 29471 68274 nw
rect 29507 68241 29621 68475
tri 29657 68442 29673 68458 se
rect 29673 68442 29750 68458
rect 29657 68376 29750 68442
rect 29657 68274 29750 68340
tri 29657 68258 29673 68274 ne
rect 29673 68258 29750 68274
rect 29490 68159 29638 68241
rect 29378 68126 29455 68142
tri 29455 68126 29471 68142 sw
rect 29378 68060 29471 68126
rect 29507 68001 29621 68159
tri 29657 68126 29673 68142 se
rect 29673 68126 29750 68142
rect 29657 68060 29750 68126
rect 29378 67925 29750 68001
rect 29378 67800 29471 67866
rect 29378 67784 29455 67800
tri 29455 67784 29471 67800 nw
rect 29507 67767 29621 67925
rect 29657 67800 29750 67866
tri 29657 67784 29673 67800 ne
rect 29673 67784 29750 67800
rect 29490 67685 29638 67767
rect 29378 67652 29455 67668
tri 29455 67652 29471 67668 sw
rect 29378 67586 29471 67652
rect 29378 67484 29471 67550
rect 29378 67468 29455 67484
tri 29455 67468 29471 67484 nw
rect 29507 67451 29621 67685
tri 29657 67652 29673 67668 se
rect 29673 67652 29750 67668
rect 29657 67586 29750 67652
rect 29657 67484 29750 67550
tri 29657 67468 29673 67484 ne
rect 29673 67468 29750 67484
rect 29490 67369 29638 67451
rect 29378 67336 29455 67352
tri 29455 67336 29471 67352 sw
rect 29378 67270 29471 67336
rect 29507 67211 29621 67369
tri 29657 67336 29673 67352 se
rect 29673 67336 29750 67352
rect 29657 67270 29750 67336
rect 29378 67135 29750 67211
rect 29378 67010 29471 67076
rect 29378 66994 29455 67010
tri 29455 66994 29471 67010 nw
rect 29507 66977 29621 67135
rect 29657 67010 29750 67076
tri 29657 66994 29673 67010 ne
rect 29673 66994 29750 67010
rect 29490 66895 29638 66977
rect 29378 66862 29455 66878
tri 29455 66862 29471 66878 sw
rect 29378 66796 29471 66862
rect 29378 66694 29471 66760
rect 29378 66678 29455 66694
tri 29455 66678 29471 66694 nw
rect 29507 66661 29621 66895
tri 29657 66862 29673 66878 se
rect 29673 66862 29750 66878
rect 29657 66796 29750 66862
rect 29657 66694 29750 66760
tri 29657 66678 29673 66694 ne
rect 29673 66678 29750 66694
rect 29490 66579 29638 66661
rect 29378 66546 29455 66562
tri 29455 66546 29471 66562 sw
rect 29378 66480 29471 66546
rect 29507 66421 29621 66579
tri 29657 66546 29673 66562 se
rect 29673 66546 29750 66562
rect 29657 66480 29750 66546
rect 29378 66345 29750 66421
rect 29378 66220 29471 66286
rect 29378 66204 29455 66220
tri 29455 66204 29471 66220 nw
rect 29507 66187 29621 66345
rect 29657 66220 29750 66286
tri 29657 66204 29673 66220 ne
rect 29673 66204 29750 66220
rect 29490 66105 29638 66187
rect 29378 66072 29455 66088
tri 29455 66072 29471 66088 sw
rect 29378 66006 29471 66072
rect 29378 65904 29471 65970
rect 29378 65888 29455 65904
tri 29455 65888 29471 65904 nw
rect 29507 65871 29621 66105
tri 29657 66072 29673 66088 se
rect 29673 66072 29750 66088
rect 29657 66006 29750 66072
rect 29657 65904 29750 65970
tri 29657 65888 29673 65904 ne
rect 29673 65888 29750 65904
rect 29490 65789 29638 65871
rect 29378 65756 29455 65772
tri 29455 65756 29471 65772 sw
rect 29378 65690 29471 65756
rect 29507 65631 29621 65789
tri 29657 65756 29673 65772 se
rect 29673 65756 29750 65772
rect 29657 65690 29750 65756
rect 29378 65555 29750 65631
rect 29378 65430 29471 65496
rect 29378 65414 29455 65430
tri 29455 65414 29471 65430 nw
rect 29507 65397 29621 65555
rect 29657 65430 29750 65496
tri 29657 65414 29673 65430 ne
rect 29673 65414 29750 65430
rect 29490 65315 29638 65397
rect 29378 65282 29455 65298
tri 29455 65282 29471 65298 sw
rect 29378 65216 29471 65282
rect 29378 65114 29471 65180
rect 29378 65098 29455 65114
tri 29455 65098 29471 65114 nw
rect 29507 65081 29621 65315
tri 29657 65282 29673 65298 se
rect 29673 65282 29750 65298
rect 29657 65216 29750 65282
rect 29657 65114 29750 65180
tri 29657 65098 29673 65114 ne
rect 29673 65098 29750 65114
rect 29490 64999 29638 65081
rect 29378 64966 29455 64982
tri 29455 64966 29471 64982 sw
rect 29378 64900 29471 64966
rect 29507 64841 29621 64999
tri 29657 64966 29673 64982 se
rect 29673 64966 29750 64982
rect 29657 64900 29750 64966
rect 29378 64765 29750 64841
rect 29378 64640 29471 64706
rect 29378 64624 29455 64640
tri 29455 64624 29471 64640 nw
rect 29507 64607 29621 64765
rect 29657 64640 29750 64706
tri 29657 64624 29673 64640 ne
rect 29673 64624 29750 64640
rect 29490 64525 29638 64607
rect 29378 64492 29455 64508
tri 29455 64492 29471 64508 sw
rect 29378 64426 29471 64492
rect 29378 64324 29471 64390
rect 29378 64308 29455 64324
tri 29455 64308 29471 64324 nw
rect 29507 64291 29621 64525
tri 29657 64492 29673 64508 se
rect 29673 64492 29750 64508
rect 29657 64426 29750 64492
rect 29657 64324 29750 64390
tri 29657 64308 29673 64324 ne
rect 29673 64308 29750 64324
rect 29490 64209 29638 64291
rect 29378 64176 29455 64192
tri 29455 64176 29471 64192 sw
rect 29378 64110 29471 64176
rect 29507 64051 29621 64209
tri 29657 64176 29673 64192 se
rect 29673 64176 29750 64192
rect 29657 64110 29750 64176
rect 29378 63975 29750 64051
rect 29378 63850 29471 63916
rect 29378 63834 29455 63850
tri 29455 63834 29471 63850 nw
rect 29507 63817 29621 63975
rect 29657 63850 29750 63916
tri 29657 63834 29673 63850 ne
rect 29673 63834 29750 63850
rect 29490 63735 29638 63817
rect 29378 63702 29455 63718
tri 29455 63702 29471 63718 sw
rect 29378 63636 29471 63702
rect 29378 63534 29471 63600
rect 29378 63518 29455 63534
tri 29455 63518 29471 63534 nw
rect 29507 63501 29621 63735
tri 29657 63702 29673 63718 se
rect 29673 63702 29750 63718
rect 29657 63636 29750 63702
rect 29657 63534 29750 63600
tri 29657 63518 29673 63534 ne
rect 29673 63518 29750 63534
rect 29490 63419 29638 63501
rect 29378 63386 29455 63402
tri 29455 63386 29471 63402 sw
rect 29378 63320 29471 63386
rect 29507 63261 29621 63419
tri 29657 63386 29673 63402 se
rect 29673 63386 29750 63402
rect 29657 63320 29750 63386
rect 29378 63185 29750 63261
rect 29378 63060 29471 63126
rect 29378 63044 29455 63060
tri 29455 63044 29471 63060 nw
rect 29507 63027 29621 63185
rect 29657 63060 29750 63126
tri 29657 63044 29673 63060 ne
rect 29673 63044 29750 63060
rect 29490 62945 29638 63027
rect 29378 62912 29455 62928
tri 29455 62912 29471 62928 sw
rect 29378 62846 29471 62912
rect 29378 62744 29471 62810
rect 29378 62728 29455 62744
tri 29455 62728 29471 62744 nw
rect 29507 62711 29621 62945
tri 29657 62912 29673 62928 se
rect 29673 62912 29750 62928
rect 29657 62846 29750 62912
rect 29657 62744 29750 62810
tri 29657 62728 29673 62744 ne
rect 29673 62728 29750 62744
rect 29490 62629 29638 62711
rect 29378 62596 29455 62612
tri 29455 62596 29471 62612 sw
rect 29378 62530 29471 62596
rect 29507 62471 29621 62629
tri 29657 62596 29673 62612 se
rect 29673 62596 29750 62612
rect 29657 62530 29750 62596
rect 29378 62395 29750 62471
rect 29378 62270 29471 62336
rect 29378 62254 29455 62270
tri 29455 62254 29471 62270 nw
rect 29507 62237 29621 62395
rect 29657 62270 29750 62336
tri 29657 62254 29673 62270 ne
rect 29673 62254 29750 62270
rect 29490 62155 29638 62237
rect 29378 62122 29455 62138
tri 29455 62122 29471 62138 sw
rect 29378 62056 29471 62122
rect 29378 61954 29471 62020
rect 29378 61938 29455 61954
tri 29455 61938 29471 61954 nw
rect 29507 61921 29621 62155
tri 29657 62122 29673 62138 se
rect 29673 62122 29750 62138
rect 29657 62056 29750 62122
rect 29657 61954 29750 62020
tri 29657 61938 29673 61954 ne
rect 29673 61938 29750 61954
rect 29490 61839 29638 61921
rect 29378 61806 29455 61822
tri 29455 61806 29471 61822 sw
rect 29378 61740 29471 61806
rect 29507 61681 29621 61839
tri 29657 61806 29673 61822 se
rect 29673 61806 29750 61822
rect 29657 61740 29750 61806
rect 29378 61605 29750 61681
rect 29378 61480 29471 61546
rect 29378 61464 29455 61480
tri 29455 61464 29471 61480 nw
rect 29507 61447 29621 61605
rect 29657 61480 29750 61546
tri 29657 61464 29673 61480 ne
rect 29673 61464 29750 61480
rect 29490 61365 29638 61447
rect 29378 61332 29455 61348
tri 29455 61332 29471 61348 sw
rect 29378 61266 29471 61332
rect 29378 61164 29471 61230
rect 29378 61148 29455 61164
tri 29455 61148 29471 61164 nw
rect 29507 61131 29621 61365
tri 29657 61332 29673 61348 se
rect 29673 61332 29750 61348
rect 29657 61266 29750 61332
rect 29657 61164 29750 61230
tri 29657 61148 29673 61164 ne
rect 29673 61148 29750 61164
rect 29490 61049 29638 61131
rect 29378 61016 29455 61032
tri 29455 61016 29471 61032 sw
rect 29378 60950 29471 61016
rect 29507 60891 29621 61049
tri 29657 61016 29673 61032 se
rect 29673 61016 29750 61032
rect 29657 60950 29750 61016
rect 29378 60815 29750 60891
rect 29378 60690 29471 60756
rect 29378 60674 29455 60690
tri 29455 60674 29471 60690 nw
rect 29507 60657 29621 60815
rect 29657 60690 29750 60756
tri 29657 60674 29673 60690 ne
rect 29673 60674 29750 60690
rect 29490 60575 29638 60657
rect 29378 60542 29455 60558
tri 29455 60542 29471 60558 sw
rect 29378 60476 29471 60542
rect 29378 60374 29471 60440
rect 29378 60358 29455 60374
tri 29455 60358 29471 60374 nw
rect 29507 60341 29621 60575
tri 29657 60542 29673 60558 se
rect 29673 60542 29750 60558
rect 29657 60476 29750 60542
rect 29657 60374 29750 60440
tri 29657 60358 29673 60374 ne
rect 29673 60358 29750 60374
rect 29490 60259 29638 60341
rect 29378 60226 29455 60242
tri 29455 60226 29471 60242 sw
rect 29378 60160 29471 60226
rect 29507 60101 29621 60259
tri 29657 60226 29673 60242 se
rect 29673 60226 29750 60242
rect 29657 60160 29750 60226
rect 29378 60025 29750 60101
rect 29378 59900 29471 59966
rect 29378 59884 29455 59900
tri 29455 59884 29471 59900 nw
rect 29507 59867 29621 60025
rect 29657 59900 29750 59966
tri 29657 59884 29673 59900 ne
rect 29673 59884 29750 59900
rect 29490 59785 29638 59867
rect 29378 59752 29455 59768
tri 29455 59752 29471 59768 sw
rect 29378 59686 29471 59752
rect 29378 59584 29471 59650
rect 29378 59568 29455 59584
tri 29455 59568 29471 59584 nw
rect 29507 59551 29621 59785
tri 29657 59752 29673 59768 se
rect 29673 59752 29750 59768
rect 29657 59686 29750 59752
rect 29657 59584 29750 59650
tri 29657 59568 29673 59584 ne
rect 29673 59568 29750 59584
rect 29490 59469 29638 59551
rect 29378 59436 29455 59452
tri 29455 59436 29471 59452 sw
rect 29378 59370 29471 59436
rect 29507 59311 29621 59469
tri 29657 59436 29673 59452 se
rect 29673 59436 29750 59452
rect 29657 59370 29750 59436
rect 29378 59235 29750 59311
rect 29378 59110 29471 59176
rect 29378 59094 29455 59110
tri 29455 59094 29471 59110 nw
rect 29507 59077 29621 59235
rect 29657 59110 29750 59176
tri 29657 59094 29673 59110 ne
rect 29673 59094 29750 59110
rect 29490 58995 29638 59077
rect 29378 58962 29455 58978
tri 29455 58962 29471 58978 sw
rect 29378 58896 29471 58962
rect 29378 58794 29471 58860
rect 29378 58778 29455 58794
tri 29455 58778 29471 58794 nw
rect 29507 58761 29621 58995
tri 29657 58962 29673 58978 se
rect 29673 58962 29750 58978
rect 29657 58896 29750 58962
rect 29657 58794 29750 58860
tri 29657 58778 29673 58794 ne
rect 29673 58778 29750 58794
rect 29490 58679 29638 58761
rect 29378 58646 29455 58662
tri 29455 58646 29471 58662 sw
rect 29378 58580 29471 58646
rect 29507 58521 29621 58679
tri 29657 58646 29673 58662 se
rect 29673 58646 29750 58662
rect 29657 58580 29750 58646
rect 29378 58445 29750 58521
rect 29378 58320 29471 58386
rect 29378 58304 29455 58320
tri 29455 58304 29471 58320 nw
rect 29507 58287 29621 58445
rect 29657 58320 29750 58386
tri 29657 58304 29673 58320 ne
rect 29673 58304 29750 58320
rect 29490 58205 29638 58287
rect 29378 58172 29455 58188
tri 29455 58172 29471 58188 sw
rect 29378 58106 29471 58172
rect 29378 58004 29471 58070
rect 29378 57988 29455 58004
tri 29455 57988 29471 58004 nw
rect 29507 57971 29621 58205
tri 29657 58172 29673 58188 se
rect 29673 58172 29750 58188
rect 29657 58106 29750 58172
rect 29657 58004 29750 58070
tri 29657 57988 29673 58004 ne
rect 29673 57988 29750 58004
rect 29490 57889 29638 57971
rect 29378 57856 29455 57872
tri 29455 57856 29471 57872 sw
rect 29378 57790 29471 57856
rect 29507 57731 29621 57889
tri 29657 57856 29673 57872 se
rect 29673 57856 29750 57872
rect 29657 57790 29750 57856
rect 29378 57655 29750 57731
rect 29378 57530 29471 57596
rect 29378 57514 29455 57530
tri 29455 57514 29471 57530 nw
rect 29507 57497 29621 57655
rect 29657 57530 29750 57596
tri 29657 57514 29673 57530 ne
rect 29673 57514 29750 57530
rect 29490 57415 29638 57497
rect 29378 57382 29455 57398
tri 29455 57382 29471 57398 sw
rect 29378 57316 29471 57382
rect 29378 57214 29471 57280
rect 29378 57198 29455 57214
tri 29455 57198 29471 57214 nw
rect 29507 57181 29621 57415
tri 29657 57382 29673 57398 se
rect 29673 57382 29750 57398
rect 29657 57316 29750 57382
rect 29657 57214 29750 57280
tri 29657 57198 29673 57214 ne
rect 29673 57198 29750 57214
rect 29490 57099 29638 57181
rect 29378 57066 29455 57082
tri 29455 57066 29471 57082 sw
rect 29378 57000 29471 57066
rect 29507 56941 29621 57099
tri 29657 57066 29673 57082 se
rect 29673 57066 29750 57082
rect 29657 57000 29750 57066
rect 29378 56865 29750 56941
rect 29378 56740 29471 56806
rect 29378 56724 29455 56740
tri 29455 56724 29471 56740 nw
rect 29507 56707 29621 56865
rect 29657 56740 29750 56806
tri 29657 56724 29673 56740 ne
rect 29673 56724 29750 56740
rect 29490 56625 29638 56707
rect 29378 56592 29455 56608
tri 29455 56592 29471 56608 sw
rect 29378 56526 29471 56592
rect 29378 56424 29471 56490
rect 29378 56408 29455 56424
tri 29455 56408 29471 56424 nw
rect 29507 56391 29621 56625
tri 29657 56592 29673 56608 se
rect 29673 56592 29750 56608
rect 29657 56526 29750 56592
rect 29657 56424 29750 56490
tri 29657 56408 29673 56424 ne
rect 29673 56408 29750 56424
rect 29490 56309 29638 56391
rect 29378 56276 29455 56292
tri 29455 56276 29471 56292 sw
rect 29378 56210 29471 56276
rect 29507 56151 29621 56309
tri 29657 56276 29673 56292 se
rect 29673 56276 29750 56292
rect 29657 56210 29750 56276
rect 29378 56075 29750 56151
rect 29378 55950 29471 56016
rect 29378 55934 29455 55950
tri 29455 55934 29471 55950 nw
rect 29507 55917 29621 56075
rect 29657 55950 29750 56016
tri 29657 55934 29673 55950 ne
rect 29673 55934 29750 55950
rect 29490 55835 29638 55917
rect 29378 55802 29455 55818
tri 29455 55802 29471 55818 sw
rect 29378 55736 29471 55802
rect 29378 55634 29471 55700
rect 29378 55618 29455 55634
tri 29455 55618 29471 55634 nw
rect 29507 55601 29621 55835
tri 29657 55802 29673 55818 se
rect 29673 55802 29750 55818
rect 29657 55736 29750 55802
rect 29657 55634 29750 55700
tri 29657 55618 29673 55634 ne
rect 29673 55618 29750 55634
rect 29490 55519 29638 55601
rect 29378 55486 29455 55502
tri 29455 55486 29471 55502 sw
rect 29378 55420 29471 55486
rect 29507 55361 29621 55519
tri 29657 55486 29673 55502 se
rect 29673 55486 29750 55502
rect 29657 55420 29750 55486
rect 29378 55285 29750 55361
rect 29378 55160 29471 55226
rect 29378 55144 29455 55160
tri 29455 55144 29471 55160 nw
rect 29507 55127 29621 55285
rect 29657 55160 29750 55226
tri 29657 55144 29673 55160 ne
rect 29673 55144 29750 55160
rect 29490 55045 29638 55127
rect 29378 55012 29455 55028
tri 29455 55012 29471 55028 sw
rect 29378 54946 29471 55012
rect 29378 54844 29471 54910
rect 29378 54828 29455 54844
tri 29455 54828 29471 54844 nw
rect 29507 54811 29621 55045
tri 29657 55012 29673 55028 se
rect 29673 55012 29750 55028
rect 29657 54946 29750 55012
rect 29657 54844 29750 54910
tri 29657 54828 29673 54844 ne
rect 29673 54828 29750 54844
rect 29490 54729 29638 54811
rect 29378 54696 29455 54712
tri 29455 54696 29471 54712 sw
rect 29378 54630 29471 54696
rect 29507 54571 29621 54729
tri 29657 54696 29673 54712 se
rect 29673 54696 29750 54712
rect 29657 54630 29750 54696
rect 29378 54495 29750 54571
rect 29378 54370 29471 54436
rect 29378 54354 29455 54370
tri 29455 54354 29471 54370 nw
rect 29507 54337 29621 54495
rect 29657 54370 29750 54436
tri 29657 54354 29673 54370 ne
rect 29673 54354 29750 54370
rect 29490 54255 29638 54337
rect 29378 54222 29455 54238
tri 29455 54222 29471 54238 sw
rect 29378 54156 29471 54222
rect 29378 54054 29471 54120
rect 29378 54038 29455 54054
tri 29455 54038 29471 54054 nw
rect 29507 54021 29621 54255
tri 29657 54222 29673 54238 se
rect 29673 54222 29750 54238
rect 29657 54156 29750 54222
rect 29657 54054 29750 54120
tri 29657 54038 29673 54054 ne
rect 29673 54038 29750 54054
rect 29490 53939 29638 54021
rect 29378 53906 29455 53922
tri 29455 53906 29471 53922 sw
rect 29378 53840 29471 53906
rect 29507 53781 29621 53939
tri 29657 53906 29673 53922 se
rect 29673 53906 29750 53922
rect 29657 53840 29750 53906
rect 29378 53705 29750 53781
rect 29378 53580 29471 53646
rect 29378 53564 29455 53580
tri 29455 53564 29471 53580 nw
rect 29507 53547 29621 53705
rect 29657 53580 29750 53646
tri 29657 53564 29673 53580 ne
rect 29673 53564 29750 53580
rect 29490 53465 29638 53547
rect 29378 53432 29455 53448
tri 29455 53432 29471 53448 sw
rect 29378 53366 29471 53432
rect 29378 53264 29471 53330
rect 29378 53248 29455 53264
tri 29455 53248 29471 53264 nw
rect 29507 53231 29621 53465
tri 29657 53432 29673 53448 se
rect 29673 53432 29750 53448
rect 29657 53366 29750 53432
rect 29657 53264 29750 53330
tri 29657 53248 29673 53264 ne
rect 29673 53248 29750 53264
rect 29490 53149 29638 53231
rect 29378 53116 29455 53132
tri 29455 53116 29471 53132 sw
rect 29378 53050 29471 53116
rect 29507 52991 29621 53149
tri 29657 53116 29673 53132 se
rect 29673 53116 29750 53132
rect 29657 53050 29750 53116
rect 29378 52915 29750 52991
rect 29378 52790 29471 52856
rect 29378 52774 29455 52790
tri 29455 52774 29471 52790 nw
rect 29507 52757 29621 52915
rect 29657 52790 29750 52856
tri 29657 52774 29673 52790 ne
rect 29673 52774 29750 52790
rect 29490 52675 29638 52757
rect 29378 52642 29455 52658
tri 29455 52642 29471 52658 sw
rect 29378 52576 29471 52642
rect 29378 52474 29471 52540
rect 29378 52458 29455 52474
tri 29455 52458 29471 52474 nw
rect 29507 52441 29621 52675
tri 29657 52642 29673 52658 se
rect 29673 52642 29750 52658
rect 29657 52576 29750 52642
rect 29657 52474 29750 52540
tri 29657 52458 29673 52474 ne
rect 29673 52458 29750 52474
rect 29490 52359 29638 52441
rect 29378 52326 29455 52342
tri 29455 52326 29471 52342 sw
rect 29378 52260 29471 52326
rect 29507 52201 29621 52359
tri 29657 52326 29673 52342 se
rect 29673 52326 29750 52342
rect 29657 52260 29750 52326
rect 29378 52125 29750 52201
rect 29378 52000 29471 52066
rect 29378 51984 29455 52000
tri 29455 51984 29471 52000 nw
rect 29507 51967 29621 52125
rect 29657 52000 29750 52066
tri 29657 51984 29673 52000 ne
rect 29673 51984 29750 52000
rect 29490 51885 29638 51967
rect 29378 51852 29455 51868
tri 29455 51852 29471 51868 sw
rect 29378 51786 29471 51852
rect 29378 51684 29471 51750
rect 29378 51668 29455 51684
tri 29455 51668 29471 51684 nw
rect 29507 51651 29621 51885
tri 29657 51852 29673 51868 se
rect 29673 51852 29750 51868
rect 29657 51786 29750 51852
rect 29657 51684 29750 51750
tri 29657 51668 29673 51684 ne
rect 29673 51668 29750 51684
rect 29490 51569 29638 51651
rect 29378 51536 29455 51552
tri 29455 51536 29471 51552 sw
rect 29378 51470 29471 51536
rect 29507 51411 29621 51569
tri 29657 51536 29673 51552 se
rect 29673 51536 29750 51552
rect 29657 51470 29750 51536
rect 29378 51335 29750 51411
rect 29378 51210 29471 51276
rect 29378 51194 29455 51210
tri 29455 51194 29471 51210 nw
rect 29507 51177 29621 51335
rect 29657 51210 29750 51276
tri 29657 51194 29673 51210 ne
rect 29673 51194 29750 51210
rect 29490 51095 29638 51177
rect 29378 51062 29455 51078
tri 29455 51062 29471 51078 sw
rect 29378 50996 29471 51062
rect 29378 50894 29471 50960
rect 29378 50878 29455 50894
tri 29455 50878 29471 50894 nw
rect 29507 50861 29621 51095
tri 29657 51062 29673 51078 se
rect 29673 51062 29750 51078
rect 29657 50996 29750 51062
rect 29657 50894 29750 50960
tri 29657 50878 29673 50894 ne
rect 29673 50878 29750 50894
rect 29490 50779 29638 50861
rect 29378 50746 29455 50762
tri 29455 50746 29471 50762 sw
rect 29378 50680 29471 50746
rect 29507 50621 29621 50779
tri 29657 50746 29673 50762 se
rect 29673 50746 29750 50762
rect 29657 50680 29750 50746
rect 29378 50545 29750 50621
rect 29378 50420 29471 50486
rect 29378 50404 29455 50420
tri 29455 50404 29471 50420 nw
rect 29507 50387 29621 50545
rect 29657 50420 29750 50486
tri 29657 50404 29673 50420 ne
rect 29673 50404 29750 50420
rect 29490 50305 29638 50387
rect 29378 50272 29455 50288
tri 29455 50272 29471 50288 sw
rect 29378 50206 29471 50272
rect 29378 50104 29471 50170
rect 29378 50088 29455 50104
tri 29455 50088 29471 50104 nw
rect 29507 50071 29621 50305
tri 29657 50272 29673 50288 se
rect 29673 50272 29750 50288
rect 29657 50206 29750 50272
rect 29657 50104 29750 50170
tri 29657 50088 29673 50104 ne
rect 29673 50088 29750 50104
rect 29490 49989 29638 50071
rect 29378 49956 29455 49972
tri 29455 49956 29471 49972 sw
rect 29378 49890 29471 49956
rect 29507 49831 29621 49989
tri 29657 49956 29673 49972 se
rect 29673 49956 29750 49972
rect 29657 49890 29750 49956
rect 29378 49755 29750 49831
rect 29378 49630 29471 49696
rect 29378 49614 29455 49630
tri 29455 49614 29471 49630 nw
rect 29507 49597 29621 49755
rect 29657 49630 29750 49696
tri 29657 49614 29673 49630 ne
rect 29673 49614 29750 49630
rect 29490 49515 29638 49597
rect 29378 49482 29455 49498
tri 29455 49482 29471 49498 sw
rect 29378 49416 29471 49482
rect 29378 49314 29471 49380
rect 29378 49298 29455 49314
tri 29455 49298 29471 49314 nw
rect 29507 49281 29621 49515
tri 29657 49482 29673 49498 se
rect 29673 49482 29750 49498
rect 29657 49416 29750 49482
rect 29657 49314 29750 49380
tri 29657 49298 29673 49314 ne
rect 29673 49298 29750 49314
rect 29490 49199 29638 49281
rect 29378 49166 29455 49182
tri 29455 49166 29471 49182 sw
rect 29378 49100 29471 49166
rect 29507 49041 29621 49199
tri 29657 49166 29673 49182 se
rect 29673 49166 29750 49182
rect 29657 49100 29750 49166
rect 29378 48965 29750 49041
rect 29378 48840 29471 48906
rect 29378 48824 29455 48840
tri 29455 48824 29471 48840 nw
rect 29507 48807 29621 48965
rect 29657 48840 29750 48906
tri 29657 48824 29673 48840 ne
rect 29673 48824 29750 48840
rect 29490 48725 29638 48807
rect 29378 48692 29455 48708
tri 29455 48692 29471 48708 sw
rect 29378 48626 29471 48692
rect 29378 48524 29471 48590
rect 29378 48508 29455 48524
tri 29455 48508 29471 48524 nw
rect 29507 48491 29621 48725
tri 29657 48692 29673 48708 se
rect 29673 48692 29750 48708
rect 29657 48626 29750 48692
rect 29657 48524 29750 48590
tri 29657 48508 29673 48524 ne
rect 29673 48508 29750 48524
rect 29490 48409 29638 48491
rect 29378 48376 29455 48392
tri 29455 48376 29471 48392 sw
rect 29378 48310 29471 48376
rect 29507 48251 29621 48409
tri 29657 48376 29673 48392 se
rect 29673 48376 29750 48392
rect 29657 48310 29750 48376
rect 29378 48175 29750 48251
rect 29378 48050 29471 48116
rect 29378 48034 29455 48050
tri 29455 48034 29471 48050 nw
rect 29507 48017 29621 48175
rect 29657 48050 29750 48116
tri 29657 48034 29673 48050 ne
rect 29673 48034 29750 48050
rect 29490 47935 29638 48017
rect 29378 47902 29455 47918
tri 29455 47902 29471 47918 sw
rect 29378 47836 29471 47902
rect 29378 47734 29471 47800
rect 29378 47718 29455 47734
tri 29455 47718 29471 47734 nw
rect 29507 47701 29621 47935
tri 29657 47902 29673 47918 se
rect 29673 47902 29750 47918
rect 29657 47836 29750 47902
rect 29657 47734 29750 47800
tri 29657 47718 29673 47734 ne
rect 29673 47718 29750 47734
rect 29490 47619 29638 47701
rect 29378 47586 29455 47602
tri 29455 47586 29471 47602 sw
rect 29378 47520 29471 47586
rect 29507 47461 29621 47619
tri 29657 47586 29673 47602 se
rect 29673 47586 29750 47602
rect 29657 47520 29750 47586
rect 29378 47385 29750 47461
rect 29378 47260 29471 47326
rect 29378 47244 29455 47260
tri 29455 47244 29471 47260 nw
rect 29507 47227 29621 47385
rect 29657 47260 29750 47326
tri 29657 47244 29673 47260 ne
rect 29673 47244 29750 47260
rect 29490 47145 29638 47227
rect 29378 47112 29455 47128
tri 29455 47112 29471 47128 sw
rect 29378 47046 29471 47112
rect 29378 46944 29471 47010
rect 29378 46928 29455 46944
tri 29455 46928 29471 46944 nw
rect 29507 46911 29621 47145
tri 29657 47112 29673 47128 se
rect 29673 47112 29750 47128
rect 29657 47046 29750 47112
rect 29657 46944 29750 47010
tri 29657 46928 29673 46944 ne
rect 29673 46928 29750 46944
rect 29490 46829 29638 46911
rect 29378 46796 29455 46812
tri 29455 46796 29471 46812 sw
rect 29378 46730 29471 46796
rect 29507 46671 29621 46829
tri 29657 46796 29673 46812 se
rect 29673 46796 29750 46812
rect 29657 46730 29750 46796
rect 29378 46595 29750 46671
rect 29378 46470 29471 46536
rect 29378 46454 29455 46470
tri 29455 46454 29471 46470 nw
rect 29507 46437 29621 46595
rect 29657 46470 29750 46536
tri 29657 46454 29673 46470 ne
rect 29673 46454 29750 46470
rect 29490 46355 29638 46437
rect 29378 46322 29455 46338
tri 29455 46322 29471 46338 sw
rect 29378 46256 29471 46322
rect 29378 46154 29471 46220
rect 29378 46138 29455 46154
tri 29455 46138 29471 46154 nw
rect 29507 46121 29621 46355
tri 29657 46322 29673 46338 se
rect 29673 46322 29750 46338
rect 29657 46256 29750 46322
rect 29657 46154 29750 46220
tri 29657 46138 29673 46154 ne
rect 29673 46138 29750 46154
rect 29490 46039 29638 46121
rect 29378 46006 29455 46022
tri 29455 46006 29471 46022 sw
rect 29378 45940 29471 46006
rect 29507 45881 29621 46039
tri 29657 46006 29673 46022 se
rect 29673 46006 29750 46022
rect 29657 45940 29750 46006
rect 29378 45805 29750 45881
rect 29378 45680 29471 45746
rect 29378 45664 29455 45680
tri 29455 45664 29471 45680 nw
rect 29507 45647 29621 45805
rect 29657 45680 29750 45746
tri 29657 45664 29673 45680 ne
rect 29673 45664 29750 45680
rect 29490 45565 29638 45647
rect 29378 45532 29455 45548
tri 29455 45532 29471 45548 sw
rect 29378 45466 29471 45532
rect 29378 45364 29471 45430
rect 29378 45348 29455 45364
tri 29455 45348 29471 45364 nw
rect 29507 45331 29621 45565
tri 29657 45532 29673 45548 se
rect 29673 45532 29750 45548
rect 29657 45466 29750 45532
rect 29657 45364 29750 45430
tri 29657 45348 29673 45364 ne
rect 29673 45348 29750 45364
rect 29490 45249 29638 45331
rect 29378 45216 29455 45232
tri 29455 45216 29471 45232 sw
rect 29378 45150 29471 45216
rect 29507 45091 29621 45249
tri 29657 45216 29673 45232 se
rect 29673 45216 29750 45232
rect 29657 45150 29750 45216
rect 29378 45015 29750 45091
rect 29378 44890 29471 44956
rect 29378 44874 29455 44890
tri 29455 44874 29471 44890 nw
rect 29507 44857 29621 45015
rect 29657 44890 29750 44956
tri 29657 44874 29673 44890 ne
rect 29673 44874 29750 44890
rect 29490 44775 29638 44857
rect 29378 44742 29455 44758
tri 29455 44742 29471 44758 sw
rect 29378 44676 29471 44742
rect 29378 44574 29471 44640
rect 29378 44558 29455 44574
tri 29455 44558 29471 44574 nw
rect 29507 44541 29621 44775
tri 29657 44742 29673 44758 se
rect 29673 44742 29750 44758
rect 29657 44676 29750 44742
rect 29657 44574 29750 44640
tri 29657 44558 29673 44574 ne
rect 29673 44558 29750 44574
rect 29490 44459 29638 44541
rect 29378 44426 29455 44442
tri 29455 44426 29471 44442 sw
rect 29378 44360 29471 44426
rect 29507 44301 29621 44459
tri 29657 44426 29673 44442 se
rect 29673 44426 29750 44442
rect 29657 44360 29750 44426
rect 29378 44225 29750 44301
rect 29378 44100 29471 44166
rect 29378 44084 29455 44100
tri 29455 44084 29471 44100 nw
rect 29507 44067 29621 44225
rect 29657 44100 29750 44166
tri 29657 44084 29673 44100 ne
rect 29673 44084 29750 44100
rect 29490 43985 29638 44067
rect 29378 43952 29455 43968
tri 29455 43952 29471 43968 sw
rect 29378 43886 29471 43952
rect 29378 43784 29471 43850
rect 29378 43768 29455 43784
tri 29455 43768 29471 43784 nw
rect 29507 43751 29621 43985
tri 29657 43952 29673 43968 se
rect 29673 43952 29750 43968
rect 29657 43886 29750 43952
rect 29657 43784 29750 43850
tri 29657 43768 29673 43784 ne
rect 29673 43768 29750 43784
rect 29490 43669 29638 43751
rect 29378 43636 29455 43652
tri 29455 43636 29471 43652 sw
rect 29378 43570 29471 43636
rect 29507 43511 29621 43669
tri 29657 43636 29673 43652 se
rect 29673 43636 29750 43652
rect 29657 43570 29750 43636
rect 29378 43435 29750 43511
rect 29378 43310 29471 43376
rect 29378 43294 29455 43310
tri 29455 43294 29471 43310 nw
rect 29507 43277 29621 43435
rect 29657 43310 29750 43376
tri 29657 43294 29673 43310 ne
rect 29673 43294 29750 43310
rect 29490 43195 29638 43277
rect 29378 43162 29455 43178
tri 29455 43162 29471 43178 sw
rect 29378 43096 29471 43162
rect 29378 42994 29471 43060
rect 29378 42978 29455 42994
tri 29455 42978 29471 42994 nw
rect 29507 42961 29621 43195
tri 29657 43162 29673 43178 se
rect 29673 43162 29750 43178
rect 29657 43096 29750 43162
rect 29657 42994 29750 43060
tri 29657 42978 29673 42994 ne
rect 29673 42978 29750 42994
rect 29490 42879 29638 42961
rect 29378 42846 29455 42862
tri 29455 42846 29471 42862 sw
rect 29378 42780 29471 42846
rect 29507 42721 29621 42879
tri 29657 42846 29673 42862 se
rect 29673 42846 29750 42862
rect 29657 42780 29750 42846
rect 29378 42645 29750 42721
rect 29378 42520 29471 42586
rect 29378 42504 29455 42520
tri 29455 42504 29471 42520 nw
rect 29507 42487 29621 42645
rect 29657 42520 29750 42586
tri 29657 42504 29673 42520 ne
rect 29673 42504 29750 42520
rect 29490 42405 29638 42487
rect 29378 42372 29455 42388
tri 29455 42372 29471 42388 sw
rect 29378 42306 29471 42372
rect 29378 42204 29471 42270
rect 29378 42188 29455 42204
tri 29455 42188 29471 42204 nw
rect 29507 42171 29621 42405
tri 29657 42372 29673 42388 se
rect 29673 42372 29750 42388
rect 29657 42306 29750 42372
rect 29657 42204 29750 42270
tri 29657 42188 29673 42204 ne
rect 29673 42188 29750 42204
rect 29490 42089 29638 42171
rect 29378 42056 29455 42072
tri 29455 42056 29471 42072 sw
rect 29378 41990 29471 42056
rect 29507 41931 29621 42089
tri 29657 42056 29673 42072 se
rect 29673 42056 29750 42072
rect 29657 41990 29750 42056
rect 29378 41855 29750 41931
rect 29378 41730 29471 41796
rect 29378 41714 29455 41730
tri 29455 41714 29471 41730 nw
rect 29507 41697 29621 41855
rect 29657 41730 29750 41796
tri 29657 41714 29673 41730 ne
rect 29673 41714 29750 41730
rect 29490 41615 29638 41697
rect 29378 41582 29455 41598
tri 29455 41582 29471 41598 sw
rect 29378 41516 29471 41582
rect 29378 41414 29471 41480
rect 29378 41398 29455 41414
tri 29455 41398 29471 41414 nw
rect 29507 41381 29621 41615
tri 29657 41582 29673 41598 se
rect 29673 41582 29750 41598
rect 29657 41516 29750 41582
rect 29657 41414 29750 41480
tri 29657 41398 29673 41414 ne
rect 29673 41398 29750 41414
rect 29490 41299 29638 41381
rect 29378 41266 29455 41282
tri 29455 41266 29471 41282 sw
rect 29378 41200 29471 41266
rect 29507 41141 29621 41299
tri 29657 41266 29673 41282 se
rect 29673 41266 29750 41282
rect 29657 41200 29750 41266
rect 29378 41065 29750 41141
rect 29378 40940 29471 41006
rect 29378 40924 29455 40940
tri 29455 40924 29471 40940 nw
rect 29507 40907 29621 41065
rect 29657 40940 29750 41006
tri 29657 40924 29673 40940 ne
rect 29673 40924 29750 40940
rect 29490 40825 29638 40907
rect 29378 40792 29455 40808
tri 29455 40792 29471 40808 sw
rect 29378 40726 29471 40792
rect 29378 40624 29471 40690
rect 29378 40608 29455 40624
tri 29455 40608 29471 40624 nw
rect 29507 40591 29621 40825
tri 29657 40792 29673 40808 se
rect 29673 40792 29750 40808
rect 29657 40726 29750 40792
rect 29657 40624 29750 40690
tri 29657 40608 29673 40624 ne
rect 29673 40608 29750 40624
rect 29490 40509 29638 40591
rect 29378 40476 29455 40492
tri 29455 40476 29471 40492 sw
rect 29378 40410 29471 40476
rect 29507 40351 29621 40509
tri 29657 40476 29673 40492 se
rect 29673 40476 29750 40492
rect 29657 40410 29750 40476
rect 29378 40275 29750 40351
rect 29378 40150 29471 40216
rect 29378 40134 29455 40150
tri 29455 40134 29471 40150 nw
rect 29507 40117 29621 40275
rect 29657 40150 29750 40216
tri 29657 40134 29673 40150 ne
rect 29673 40134 29750 40150
rect 29490 40035 29638 40117
rect 29378 40002 29455 40018
tri 29455 40002 29471 40018 sw
rect 29378 39936 29471 40002
rect 29378 39834 29471 39900
rect 29378 39818 29455 39834
tri 29455 39818 29471 39834 nw
rect 29507 39801 29621 40035
tri 29657 40002 29673 40018 se
rect 29673 40002 29750 40018
rect 29657 39936 29750 40002
rect 29657 39834 29750 39900
tri 29657 39818 29673 39834 ne
rect 29673 39818 29750 39834
rect 29490 39719 29638 39801
rect 29378 39686 29455 39702
tri 29455 39686 29471 39702 sw
rect 29378 39620 29471 39686
rect 29507 39561 29621 39719
tri 29657 39686 29673 39702 se
rect 29673 39686 29750 39702
rect 29657 39620 29750 39686
rect 29378 39485 29750 39561
rect 29378 39360 29471 39426
rect 29378 39344 29455 39360
tri 29455 39344 29471 39360 nw
rect 29507 39327 29621 39485
rect 29657 39360 29750 39426
tri 29657 39344 29673 39360 ne
rect 29673 39344 29750 39360
rect 29490 39245 29638 39327
rect 29378 39212 29455 39228
tri 29455 39212 29471 39228 sw
rect 29378 39146 29471 39212
rect 29378 39044 29471 39110
rect 29378 39028 29455 39044
tri 29455 39028 29471 39044 nw
rect 29507 39011 29621 39245
tri 29657 39212 29673 39228 se
rect 29673 39212 29750 39228
rect 29657 39146 29750 39212
rect 29657 39044 29750 39110
tri 29657 39028 29673 39044 ne
rect 29673 39028 29750 39044
rect 29490 38929 29638 39011
rect 29378 38896 29455 38912
tri 29455 38896 29471 38912 sw
rect 29378 38830 29471 38896
rect 29507 38771 29621 38929
tri 29657 38896 29673 38912 se
rect 29673 38896 29750 38912
rect 29657 38830 29750 38896
rect 29378 38695 29750 38771
rect 29378 38570 29471 38636
rect 29378 38554 29455 38570
tri 29455 38554 29471 38570 nw
rect 29507 38537 29621 38695
rect 29657 38570 29750 38636
tri 29657 38554 29673 38570 ne
rect 29673 38554 29750 38570
rect 29490 38455 29638 38537
rect 29378 38422 29455 38438
tri 29455 38422 29471 38438 sw
rect 29378 38356 29471 38422
rect 29378 38254 29471 38320
rect 29378 38238 29455 38254
tri 29455 38238 29471 38254 nw
rect 29507 38221 29621 38455
tri 29657 38422 29673 38438 se
rect 29673 38422 29750 38438
rect 29657 38356 29750 38422
rect 29657 38254 29750 38320
tri 29657 38238 29673 38254 ne
rect 29673 38238 29750 38254
rect 29490 38139 29638 38221
rect 29378 38106 29455 38122
tri 29455 38106 29471 38122 sw
rect 29378 38040 29471 38106
rect 29507 37981 29621 38139
tri 29657 38106 29673 38122 se
rect 29673 38106 29750 38122
rect 29657 38040 29750 38106
rect 29378 37905 29750 37981
rect 29378 37780 29471 37846
rect 29378 37764 29455 37780
tri 29455 37764 29471 37780 nw
rect 29507 37747 29621 37905
rect 29657 37780 29750 37846
tri 29657 37764 29673 37780 ne
rect 29673 37764 29750 37780
rect 29490 37665 29638 37747
rect 29378 37632 29455 37648
tri 29455 37632 29471 37648 sw
rect 29378 37566 29471 37632
rect 29378 37464 29471 37530
rect 29378 37448 29455 37464
tri 29455 37448 29471 37464 nw
rect 29507 37431 29621 37665
tri 29657 37632 29673 37648 se
rect 29673 37632 29750 37648
rect 29657 37566 29750 37632
rect 29657 37464 29750 37530
tri 29657 37448 29673 37464 ne
rect 29673 37448 29750 37464
rect 29490 37349 29638 37431
rect 29378 37316 29455 37332
tri 29455 37316 29471 37332 sw
rect 29378 37250 29471 37316
rect 29507 37191 29621 37349
tri 29657 37316 29673 37332 se
rect 29673 37316 29750 37332
rect 29657 37250 29750 37316
rect 29378 37115 29750 37191
rect 29378 36990 29471 37056
rect 29378 36974 29455 36990
tri 29455 36974 29471 36990 nw
rect 29507 36957 29621 37115
rect 29657 36990 29750 37056
tri 29657 36974 29673 36990 ne
rect 29673 36974 29750 36990
rect 29490 36875 29638 36957
rect 29378 36842 29455 36858
tri 29455 36842 29471 36858 sw
rect 29378 36776 29471 36842
rect 29378 36674 29471 36740
rect 29378 36658 29455 36674
tri 29455 36658 29471 36674 nw
rect 29507 36641 29621 36875
tri 29657 36842 29673 36858 se
rect 29673 36842 29750 36858
rect 29657 36776 29750 36842
rect 29657 36674 29750 36740
tri 29657 36658 29673 36674 ne
rect 29673 36658 29750 36674
rect 29490 36559 29638 36641
rect 29378 36526 29455 36542
tri 29455 36526 29471 36542 sw
rect 29378 36460 29471 36526
rect 29507 36401 29621 36559
tri 29657 36526 29673 36542 se
rect 29673 36526 29750 36542
rect 29657 36460 29750 36526
rect 29378 36325 29750 36401
rect 29378 36200 29471 36266
rect 29378 36184 29455 36200
tri 29455 36184 29471 36200 nw
rect 29507 36167 29621 36325
rect 29657 36200 29750 36266
tri 29657 36184 29673 36200 ne
rect 29673 36184 29750 36200
rect 29490 36085 29638 36167
rect 29378 36052 29455 36068
tri 29455 36052 29471 36068 sw
rect 29378 35986 29471 36052
rect 29378 35884 29471 35950
rect 29378 35868 29455 35884
tri 29455 35868 29471 35884 nw
rect 29507 35851 29621 36085
tri 29657 36052 29673 36068 se
rect 29673 36052 29750 36068
rect 29657 35986 29750 36052
rect 29657 35884 29750 35950
tri 29657 35868 29673 35884 ne
rect 29673 35868 29750 35884
rect 29490 35769 29638 35851
rect 29378 35736 29455 35752
tri 29455 35736 29471 35752 sw
rect 29378 35670 29471 35736
rect 29507 35611 29621 35769
tri 29657 35736 29673 35752 se
rect 29673 35736 29750 35752
rect 29657 35670 29750 35736
rect 29378 35535 29750 35611
rect 29378 35410 29471 35476
rect 29378 35394 29455 35410
tri 29455 35394 29471 35410 nw
rect 29507 35377 29621 35535
rect 29657 35410 29750 35476
tri 29657 35394 29673 35410 ne
rect 29673 35394 29750 35410
rect 29490 35295 29638 35377
rect 29378 35262 29455 35278
tri 29455 35262 29471 35278 sw
rect 29378 35196 29471 35262
rect 29378 35094 29471 35160
rect 29378 35078 29455 35094
tri 29455 35078 29471 35094 nw
rect 29507 35061 29621 35295
tri 29657 35262 29673 35278 se
rect 29673 35262 29750 35278
rect 29657 35196 29750 35262
rect 29657 35094 29750 35160
tri 29657 35078 29673 35094 ne
rect 29673 35078 29750 35094
rect 29490 34979 29638 35061
rect 29378 34946 29455 34962
tri 29455 34946 29471 34962 sw
rect 29378 34880 29471 34946
rect 29507 34821 29621 34979
tri 29657 34946 29673 34962 se
rect 29673 34946 29750 34962
rect 29657 34880 29750 34946
rect 29378 34745 29750 34821
rect 29378 34620 29471 34686
rect 29378 34604 29455 34620
tri 29455 34604 29471 34620 nw
rect 29507 34587 29621 34745
rect 29657 34620 29750 34686
tri 29657 34604 29673 34620 ne
rect 29673 34604 29750 34620
rect 29490 34505 29638 34587
rect 29378 34472 29455 34488
tri 29455 34472 29471 34488 sw
rect 29378 34406 29471 34472
rect 29378 34304 29471 34370
rect 29378 34288 29455 34304
tri 29455 34288 29471 34304 nw
rect 29507 34271 29621 34505
tri 29657 34472 29673 34488 se
rect 29673 34472 29750 34488
rect 29657 34406 29750 34472
rect 29657 34304 29750 34370
tri 29657 34288 29673 34304 ne
rect 29673 34288 29750 34304
rect 29490 34189 29638 34271
rect 29378 34156 29455 34172
tri 29455 34156 29471 34172 sw
rect 29378 34090 29471 34156
rect 29507 34031 29621 34189
tri 29657 34156 29673 34172 se
rect 29673 34156 29750 34172
rect 29657 34090 29750 34156
rect 29378 33955 29750 34031
rect 29378 33830 29471 33896
rect 29378 33814 29455 33830
tri 29455 33814 29471 33830 nw
rect 29507 33797 29621 33955
rect 29657 33830 29750 33896
tri 29657 33814 29673 33830 ne
rect 29673 33814 29750 33830
rect 29490 33715 29638 33797
rect 29378 33682 29455 33698
tri 29455 33682 29471 33698 sw
rect 29378 33616 29471 33682
rect 29378 33514 29471 33580
rect 29378 33498 29455 33514
tri 29455 33498 29471 33514 nw
rect 29507 33481 29621 33715
tri 29657 33682 29673 33698 se
rect 29673 33682 29750 33698
rect 29657 33616 29750 33682
rect 29657 33514 29750 33580
tri 29657 33498 29673 33514 ne
rect 29673 33498 29750 33514
rect 29490 33399 29638 33481
rect 29378 33366 29455 33382
tri 29455 33366 29471 33382 sw
rect 29378 33300 29471 33366
rect 29507 33241 29621 33399
tri 29657 33366 29673 33382 se
rect 29673 33366 29750 33382
rect 29657 33300 29750 33366
rect 29378 33165 29750 33241
rect 29378 33040 29471 33106
rect 29378 33024 29455 33040
tri 29455 33024 29471 33040 nw
rect 29507 33007 29621 33165
rect 29657 33040 29750 33106
tri 29657 33024 29673 33040 ne
rect 29673 33024 29750 33040
rect 29490 32925 29638 33007
rect 29378 32892 29455 32908
tri 29455 32892 29471 32908 sw
rect 29378 32826 29471 32892
rect 29378 32724 29471 32790
rect 29378 32708 29455 32724
tri 29455 32708 29471 32724 nw
rect 29507 32691 29621 32925
tri 29657 32892 29673 32908 se
rect 29673 32892 29750 32908
rect 29657 32826 29750 32892
rect 29657 32724 29750 32790
tri 29657 32708 29673 32724 ne
rect 29673 32708 29750 32724
rect 29490 32609 29638 32691
rect 29378 32576 29455 32592
tri 29455 32576 29471 32592 sw
rect 29378 32510 29471 32576
rect 29507 32451 29621 32609
tri 29657 32576 29673 32592 se
rect 29673 32576 29750 32592
rect 29657 32510 29750 32576
rect 29378 32375 29750 32451
rect 29378 32250 29471 32316
rect 29378 32234 29455 32250
tri 29455 32234 29471 32250 nw
rect 29507 32217 29621 32375
rect 29657 32250 29750 32316
tri 29657 32234 29673 32250 ne
rect 29673 32234 29750 32250
rect 29490 32135 29638 32217
rect 29378 32102 29455 32118
tri 29455 32102 29471 32118 sw
rect 29378 32036 29471 32102
rect 29378 31934 29471 32000
rect 29378 31918 29455 31934
tri 29455 31918 29471 31934 nw
rect 29507 31901 29621 32135
tri 29657 32102 29673 32118 se
rect 29673 32102 29750 32118
rect 29657 32036 29750 32102
rect 29657 31934 29750 32000
tri 29657 31918 29673 31934 ne
rect 29673 31918 29750 31934
rect 29490 31819 29638 31901
rect 29378 31786 29455 31802
tri 29455 31786 29471 31802 sw
rect 29378 31720 29471 31786
rect 29507 31661 29621 31819
tri 29657 31786 29673 31802 se
rect 29673 31786 29750 31802
rect 29657 31720 29750 31786
rect 29378 31585 29750 31661
rect 29378 31460 29471 31526
rect 29378 31444 29455 31460
tri 29455 31444 29471 31460 nw
rect 29507 31427 29621 31585
rect 29657 31460 29750 31526
tri 29657 31444 29673 31460 ne
rect 29673 31444 29750 31460
rect 29490 31345 29638 31427
rect 29378 31312 29455 31328
tri 29455 31312 29471 31328 sw
rect 29378 31246 29471 31312
rect 29378 31144 29471 31210
rect 29378 31128 29455 31144
tri 29455 31128 29471 31144 nw
rect 29507 31111 29621 31345
tri 29657 31312 29673 31328 se
rect 29673 31312 29750 31328
rect 29657 31246 29750 31312
rect 29657 31144 29750 31210
tri 29657 31128 29673 31144 ne
rect 29673 31128 29750 31144
rect 29490 31029 29638 31111
rect 29378 30996 29455 31012
tri 29455 30996 29471 31012 sw
rect 29378 30930 29471 30996
rect 29507 30871 29621 31029
tri 29657 30996 29673 31012 se
rect 29673 30996 29750 31012
rect 29657 30930 29750 30996
rect 29378 30795 29750 30871
rect 29378 30670 29471 30736
rect 29378 30654 29455 30670
tri 29455 30654 29471 30670 nw
rect 29507 30637 29621 30795
rect 29657 30670 29750 30736
tri 29657 30654 29673 30670 ne
rect 29673 30654 29750 30670
rect 29490 30555 29638 30637
rect 29378 30522 29455 30538
tri 29455 30522 29471 30538 sw
rect 29378 30456 29471 30522
rect 29378 30354 29471 30420
rect 29378 30338 29455 30354
tri 29455 30338 29471 30354 nw
rect 29507 30321 29621 30555
tri 29657 30522 29673 30538 se
rect 29673 30522 29750 30538
rect 29657 30456 29750 30522
rect 29657 30354 29750 30420
tri 29657 30338 29673 30354 ne
rect 29673 30338 29750 30354
rect 29490 30239 29638 30321
rect 29378 30206 29455 30222
tri 29455 30206 29471 30222 sw
rect 29378 30140 29471 30206
rect 29507 30081 29621 30239
tri 29657 30206 29673 30222 se
rect 29673 30206 29750 30222
rect 29657 30140 29750 30206
rect 29378 30005 29750 30081
rect 29378 29880 29471 29946
rect 29378 29864 29455 29880
tri 29455 29864 29471 29880 nw
rect 29507 29847 29621 30005
rect 29657 29880 29750 29946
tri 29657 29864 29673 29880 ne
rect 29673 29864 29750 29880
rect 29490 29765 29638 29847
rect 29378 29732 29455 29748
tri 29455 29732 29471 29748 sw
rect 29378 29666 29471 29732
rect 29378 29564 29471 29630
rect 29378 29548 29455 29564
tri 29455 29548 29471 29564 nw
rect 29507 29531 29621 29765
tri 29657 29732 29673 29748 se
rect 29673 29732 29750 29748
rect 29657 29666 29750 29732
rect 29657 29564 29750 29630
tri 29657 29548 29673 29564 ne
rect 29673 29548 29750 29564
rect 29490 29449 29638 29531
rect 29378 29416 29455 29432
tri 29455 29416 29471 29432 sw
rect 29378 29350 29471 29416
rect 29507 29291 29621 29449
tri 29657 29416 29673 29432 se
rect 29673 29416 29750 29432
rect 29657 29350 29750 29416
rect 29378 29215 29750 29291
rect 29378 29090 29471 29156
rect 29378 29074 29455 29090
tri 29455 29074 29471 29090 nw
rect 29507 29057 29621 29215
rect 29657 29090 29750 29156
tri 29657 29074 29673 29090 ne
rect 29673 29074 29750 29090
rect 29490 28975 29638 29057
rect 29378 28942 29455 28958
tri 29455 28942 29471 28958 sw
rect 29378 28876 29471 28942
rect 29507 28833 29621 28975
tri 29657 28942 29673 28958 se
rect 29673 28942 29750 28958
rect 29657 28876 29750 28942
rect 29786 28463 29822 80603
rect 29858 28463 29894 80603
rect 29930 80445 29966 80603
rect 29922 80303 29974 80445
rect 29930 28763 29966 80303
rect 29922 28621 29974 28763
rect 29930 28463 29966 28621
rect 30002 28463 30038 80603
rect 30074 28463 30110 80603
rect 30146 28833 30230 80233
rect 30266 28463 30302 80603
rect 30338 28463 30374 80603
rect 30410 80445 30446 80603
rect 30402 80303 30454 80445
rect 30410 28763 30446 80303
rect 30402 28621 30454 28763
rect 30410 28463 30446 28621
rect 30482 28463 30518 80603
rect 30554 28463 30590 80603
rect 30626 80124 30719 80190
rect 30626 80108 30703 80124
tri 30703 80108 30719 80124 nw
rect 30755 80091 30869 80233
rect 30905 80124 30998 80190
tri 30905 80108 30921 80124 ne
rect 30921 80108 30998 80124
rect 30738 80009 30886 80091
rect 30626 79976 30703 79992
tri 30703 79976 30719 79992 sw
rect 30626 79910 30719 79976
rect 30755 79851 30869 80009
tri 30905 79976 30921 79992 se
rect 30921 79976 30998 79992
rect 30905 79910 30998 79976
rect 30626 79775 30998 79851
rect 30626 79650 30719 79716
rect 30626 79634 30703 79650
tri 30703 79634 30719 79650 nw
rect 30755 79617 30869 79775
rect 30905 79650 30998 79716
tri 30905 79634 30921 79650 ne
rect 30921 79634 30998 79650
rect 30738 79535 30886 79617
rect 30626 79502 30703 79518
tri 30703 79502 30719 79518 sw
rect 30626 79436 30719 79502
rect 30626 79334 30719 79400
rect 30626 79318 30703 79334
tri 30703 79318 30719 79334 nw
rect 30755 79301 30869 79535
tri 30905 79502 30921 79518 se
rect 30921 79502 30998 79518
rect 30905 79436 30998 79502
rect 30905 79334 30998 79400
tri 30905 79318 30921 79334 ne
rect 30921 79318 30998 79334
rect 30738 79219 30886 79301
rect 30626 79186 30703 79202
tri 30703 79186 30719 79202 sw
rect 30626 79120 30719 79186
rect 30755 79061 30869 79219
tri 30905 79186 30921 79202 se
rect 30921 79186 30998 79202
rect 30905 79120 30998 79186
rect 30626 78985 30998 79061
rect 30626 78860 30719 78926
rect 30626 78844 30703 78860
tri 30703 78844 30719 78860 nw
rect 30755 78827 30869 78985
rect 30905 78860 30998 78926
tri 30905 78844 30921 78860 ne
rect 30921 78844 30998 78860
rect 30738 78745 30886 78827
rect 30626 78712 30703 78728
tri 30703 78712 30719 78728 sw
rect 30626 78646 30719 78712
rect 30626 78544 30719 78610
rect 30626 78528 30703 78544
tri 30703 78528 30719 78544 nw
rect 30755 78511 30869 78745
tri 30905 78712 30921 78728 se
rect 30921 78712 30998 78728
rect 30905 78646 30998 78712
rect 30905 78544 30998 78610
tri 30905 78528 30921 78544 ne
rect 30921 78528 30998 78544
rect 30738 78429 30886 78511
rect 30626 78396 30703 78412
tri 30703 78396 30719 78412 sw
rect 30626 78330 30719 78396
rect 30755 78271 30869 78429
tri 30905 78396 30921 78412 se
rect 30921 78396 30998 78412
rect 30905 78330 30998 78396
rect 30626 78195 30998 78271
rect 30626 78070 30719 78136
rect 30626 78054 30703 78070
tri 30703 78054 30719 78070 nw
rect 30755 78037 30869 78195
rect 30905 78070 30998 78136
tri 30905 78054 30921 78070 ne
rect 30921 78054 30998 78070
rect 30738 77955 30886 78037
rect 30626 77922 30703 77938
tri 30703 77922 30719 77938 sw
rect 30626 77856 30719 77922
rect 30626 77754 30719 77820
rect 30626 77738 30703 77754
tri 30703 77738 30719 77754 nw
rect 30755 77721 30869 77955
tri 30905 77922 30921 77938 se
rect 30921 77922 30998 77938
rect 30905 77856 30998 77922
rect 30905 77754 30998 77820
tri 30905 77738 30921 77754 ne
rect 30921 77738 30998 77754
rect 30738 77639 30886 77721
rect 30626 77606 30703 77622
tri 30703 77606 30719 77622 sw
rect 30626 77540 30719 77606
rect 30755 77481 30869 77639
tri 30905 77606 30921 77622 se
rect 30921 77606 30998 77622
rect 30905 77540 30998 77606
rect 30626 77405 30998 77481
rect 30626 77280 30719 77346
rect 30626 77264 30703 77280
tri 30703 77264 30719 77280 nw
rect 30755 77247 30869 77405
rect 30905 77280 30998 77346
tri 30905 77264 30921 77280 ne
rect 30921 77264 30998 77280
rect 30738 77165 30886 77247
rect 30626 77132 30703 77148
tri 30703 77132 30719 77148 sw
rect 30626 77066 30719 77132
rect 30626 76964 30719 77030
rect 30626 76948 30703 76964
tri 30703 76948 30719 76964 nw
rect 30755 76931 30869 77165
tri 30905 77132 30921 77148 se
rect 30921 77132 30998 77148
rect 30905 77066 30998 77132
rect 30905 76964 30998 77030
tri 30905 76948 30921 76964 ne
rect 30921 76948 30998 76964
rect 30738 76849 30886 76931
rect 30626 76816 30703 76832
tri 30703 76816 30719 76832 sw
rect 30626 76750 30719 76816
rect 30755 76691 30869 76849
tri 30905 76816 30921 76832 se
rect 30921 76816 30998 76832
rect 30905 76750 30998 76816
rect 30626 76615 30998 76691
rect 30626 76490 30719 76556
rect 30626 76474 30703 76490
tri 30703 76474 30719 76490 nw
rect 30755 76457 30869 76615
rect 30905 76490 30998 76556
tri 30905 76474 30921 76490 ne
rect 30921 76474 30998 76490
rect 30738 76375 30886 76457
rect 30626 76342 30703 76358
tri 30703 76342 30719 76358 sw
rect 30626 76276 30719 76342
rect 30626 76174 30719 76240
rect 30626 76158 30703 76174
tri 30703 76158 30719 76174 nw
rect 30755 76141 30869 76375
tri 30905 76342 30921 76358 se
rect 30921 76342 30998 76358
rect 30905 76276 30998 76342
rect 30905 76174 30998 76240
tri 30905 76158 30921 76174 ne
rect 30921 76158 30998 76174
rect 30738 76059 30886 76141
rect 30626 76026 30703 76042
tri 30703 76026 30719 76042 sw
rect 30626 75960 30719 76026
rect 30755 75901 30869 76059
tri 30905 76026 30921 76042 se
rect 30921 76026 30998 76042
rect 30905 75960 30998 76026
rect 30626 75825 30998 75901
rect 30626 75700 30719 75766
rect 30626 75684 30703 75700
tri 30703 75684 30719 75700 nw
rect 30755 75667 30869 75825
rect 30905 75700 30998 75766
tri 30905 75684 30921 75700 ne
rect 30921 75684 30998 75700
rect 30738 75585 30886 75667
rect 30626 75552 30703 75568
tri 30703 75552 30719 75568 sw
rect 30626 75486 30719 75552
rect 30626 75384 30719 75450
rect 30626 75368 30703 75384
tri 30703 75368 30719 75384 nw
rect 30755 75351 30869 75585
tri 30905 75552 30921 75568 se
rect 30921 75552 30998 75568
rect 30905 75486 30998 75552
rect 30905 75384 30998 75450
tri 30905 75368 30921 75384 ne
rect 30921 75368 30998 75384
rect 30738 75269 30886 75351
rect 30626 75236 30703 75252
tri 30703 75236 30719 75252 sw
rect 30626 75170 30719 75236
rect 30755 75111 30869 75269
tri 30905 75236 30921 75252 se
rect 30921 75236 30998 75252
rect 30905 75170 30998 75236
rect 30626 75035 30998 75111
rect 30626 74910 30719 74976
rect 30626 74894 30703 74910
tri 30703 74894 30719 74910 nw
rect 30755 74877 30869 75035
rect 30905 74910 30998 74976
tri 30905 74894 30921 74910 ne
rect 30921 74894 30998 74910
rect 30738 74795 30886 74877
rect 30626 74762 30703 74778
tri 30703 74762 30719 74778 sw
rect 30626 74696 30719 74762
rect 30626 74594 30719 74660
rect 30626 74578 30703 74594
tri 30703 74578 30719 74594 nw
rect 30755 74561 30869 74795
tri 30905 74762 30921 74778 se
rect 30921 74762 30998 74778
rect 30905 74696 30998 74762
rect 30905 74594 30998 74660
tri 30905 74578 30921 74594 ne
rect 30921 74578 30998 74594
rect 30738 74479 30886 74561
rect 30626 74446 30703 74462
tri 30703 74446 30719 74462 sw
rect 30626 74380 30719 74446
rect 30755 74321 30869 74479
tri 30905 74446 30921 74462 se
rect 30921 74446 30998 74462
rect 30905 74380 30998 74446
rect 30626 74245 30998 74321
rect 30626 74120 30719 74186
rect 30626 74104 30703 74120
tri 30703 74104 30719 74120 nw
rect 30755 74087 30869 74245
rect 30905 74120 30998 74186
tri 30905 74104 30921 74120 ne
rect 30921 74104 30998 74120
rect 30738 74005 30886 74087
rect 30626 73972 30703 73988
tri 30703 73972 30719 73988 sw
rect 30626 73906 30719 73972
rect 30626 73804 30719 73870
rect 30626 73788 30703 73804
tri 30703 73788 30719 73804 nw
rect 30755 73771 30869 74005
tri 30905 73972 30921 73988 se
rect 30921 73972 30998 73988
rect 30905 73906 30998 73972
rect 30905 73804 30998 73870
tri 30905 73788 30921 73804 ne
rect 30921 73788 30998 73804
rect 30738 73689 30886 73771
rect 30626 73656 30703 73672
tri 30703 73656 30719 73672 sw
rect 30626 73590 30719 73656
rect 30755 73531 30869 73689
tri 30905 73656 30921 73672 se
rect 30921 73656 30998 73672
rect 30905 73590 30998 73656
rect 30626 73455 30998 73531
rect 30626 73330 30719 73396
rect 30626 73314 30703 73330
tri 30703 73314 30719 73330 nw
rect 30755 73297 30869 73455
rect 30905 73330 30998 73396
tri 30905 73314 30921 73330 ne
rect 30921 73314 30998 73330
rect 30738 73215 30886 73297
rect 30626 73182 30703 73198
tri 30703 73182 30719 73198 sw
rect 30626 73116 30719 73182
rect 30626 73014 30719 73080
rect 30626 72998 30703 73014
tri 30703 72998 30719 73014 nw
rect 30755 72981 30869 73215
tri 30905 73182 30921 73198 se
rect 30921 73182 30998 73198
rect 30905 73116 30998 73182
rect 30905 73014 30998 73080
tri 30905 72998 30921 73014 ne
rect 30921 72998 30998 73014
rect 30738 72899 30886 72981
rect 30626 72866 30703 72882
tri 30703 72866 30719 72882 sw
rect 30626 72800 30719 72866
rect 30755 72741 30869 72899
tri 30905 72866 30921 72882 se
rect 30921 72866 30998 72882
rect 30905 72800 30998 72866
rect 30626 72665 30998 72741
rect 30626 72540 30719 72606
rect 30626 72524 30703 72540
tri 30703 72524 30719 72540 nw
rect 30755 72507 30869 72665
rect 30905 72540 30998 72606
tri 30905 72524 30921 72540 ne
rect 30921 72524 30998 72540
rect 30738 72425 30886 72507
rect 30626 72392 30703 72408
tri 30703 72392 30719 72408 sw
rect 30626 72326 30719 72392
rect 30626 72224 30719 72290
rect 30626 72208 30703 72224
tri 30703 72208 30719 72224 nw
rect 30755 72191 30869 72425
tri 30905 72392 30921 72408 se
rect 30921 72392 30998 72408
rect 30905 72326 30998 72392
rect 30905 72224 30998 72290
tri 30905 72208 30921 72224 ne
rect 30921 72208 30998 72224
rect 30738 72109 30886 72191
rect 30626 72076 30703 72092
tri 30703 72076 30719 72092 sw
rect 30626 72010 30719 72076
rect 30755 71951 30869 72109
tri 30905 72076 30921 72092 se
rect 30921 72076 30998 72092
rect 30905 72010 30998 72076
rect 30626 71875 30998 71951
rect 30626 71750 30719 71816
rect 30626 71734 30703 71750
tri 30703 71734 30719 71750 nw
rect 30755 71717 30869 71875
rect 30905 71750 30998 71816
tri 30905 71734 30921 71750 ne
rect 30921 71734 30998 71750
rect 30738 71635 30886 71717
rect 30626 71602 30703 71618
tri 30703 71602 30719 71618 sw
rect 30626 71536 30719 71602
rect 30626 71434 30719 71500
rect 30626 71418 30703 71434
tri 30703 71418 30719 71434 nw
rect 30755 71401 30869 71635
tri 30905 71602 30921 71618 se
rect 30921 71602 30998 71618
rect 30905 71536 30998 71602
rect 30905 71434 30998 71500
tri 30905 71418 30921 71434 ne
rect 30921 71418 30998 71434
rect 30738 71319 30886 71401
rect 30626 71286 30703 71302
tri 30703 71286 30719 71302 sw
rect 30626 71220 30719 71286
rect 30755 71161 30869 71319
tri 30905 71286 30921 71302 se
rect 30921 71286 30998 71302
rect 30905 71220 30998 71286
rect 30626 71085 30998 71161
rect 30626 70960 30719 71026
rect 30626 70944 30703 70960
tri 30703 70944 30719 70960 nw
rect 30755 70927 30869 71085
rect 30905 70960 30998 71026
tri 30905 70944 30921 70960 ne
rect 30921 70944 30998 70960
rect 30738 70845 30886 70927
rect 30626 70812 30703 70828
tri 30703 70812 30719 70828 sw
rect 30626 70746 30719 70812
rect 30626 70644 30719 70710
rect 30626 70628 30703 70644
tri 30703 70628 30719 70644 nw
rect 30755 70611 30869 70845
tri 30905 70812 30921 70828 se
rect 30921 70812 30998 70828
rect 30905 70746 30998 70812
rect 30905 70644 30998 70710
tri 30905 70628 30921 70644 ne
rect 30921 70628 30998 70644
rect 30738 70529 30886 70611
rect 30626 70496 30703 70512
tri 30703 70496 30719 70512 sw
rect 30626 70430 30719 70496
rect 30755 70371 30869 70529
tri 30905 70496 30921 70512 se
rect 30921 70496 30998 70512
rect 30905 70430 30998 70496
rect 30626 70295 30998 70371
rect 30626 70170 30719 70236
rect 30626 70154 30703 70170
tri 30703 70154 30719 70170 nw
rect 30755 70137 30869 70295
rect 30905 70170 30998 70236
tri 30905 70154 30921 70170 ne
rect 30921 70154 30998 70170
rect 30738 70055 30886 70137
rect 30626 70022 30703 70038
tri 30703 70022 30719 70038 sw
rect 30626 69956 30719 70022
rect 30626 69854 30719 69920
rect 30626 69838 30703 69854
tri 30703 69838 30719 69854 nw
rect 30755 69821 30869 70055
tri 30905 70022 30921 70038 se
rect 30921 70022 30998 70038
rect 30905 69956 30998 70022
rect 30905 69854 30998 69920
tri 30905 69838 30921 69854 ne
rect 30921 69838 30998 69854
rect 30738 69739 30886 69821
rect 30626 69706 30703 69722
tri 30703 69706 30719 69722 sw
rect 30626 69640 30719 69706
rect 30755 69581 30869 69739
tri 30905 69706 30921 69722 se
rect 30921 69706 30998 69722
rect 30905 69640 30998 69706
rect 30626 69505 30998 69581
rect 30626 69380 30719 69446
rect 30626 69364 30703 69380
tri 30703 69364 30719 69380 nw
rect 30755 69347 30869 69505
rect 30905 69380 30998 69446
tri 30905 69364 30921 69380 ne
rect 30921 69364 30998 69380
rect 30738 69265 30886 69347
rect 30626 69232 30703 69248
tri 30703 69232 30719 69248 sw
rect 30626 69166 30719 69232
rect 30626 69064 30719 69130
rect 30626 69048 30703 69064
tri 30703 69048 30719 69064 nw
rect 30755 69031 30869 69265
tri 30905 69232 30921 69248 se
rect 30921 69232 30998 69248
rect 30905 69166 30998 69232
rect 30905 69064 30998 69130
tri 30905 69048 30921 69064 ne
rect 30921 69048 30998 69064
rect 30738 68949 30886 69031
rect 30626 68916 30703 68932
tri 30703 68916 30719 68932 sw
rect 30626 68850 30719 68916
rect 30755 68791 30869 68949
tri 30905 68916 30921 68932 se
rect 30921 68916 30998 68932
rect 30905 68850 30998 68916
rect 30626 68715 30998 68791
rect 30626 68590 30719 68656
rect 30626 68574 30703 68590
tri 30703 68574 30719 68590 nw
rect 30755 68557 30869 68715
rect 30905 68590 30998 68656
tri 30905 68574 30921 68590 ne
rect 30921 68574 30998 68590
rect 30738 68475 30886 68557
rect 30626 68442 30703 68458
tri 30703 68442 30719 68458 sw
rect 30626 68376 30719 68442
rect 30626 68274 30719 68340
rect 30626 68258 30703 68274
tri 30703 68258 30719 68274 nw
rect 30755 68241 30869 68475
tri 30905 68442 30921 68458 se
rect 30921 68442 30998 68458
rect 30905 68376 30998 68442
rect 30905 68274 30998 68340
tri 30905 68258 30921 68274 ne
rect 30921 68258 30998 68274
rect 30738 68159 30886 68241
rect 30626 68126 30703 68142
tri 30703 68126 30719 68142 sw
rect 30626 68060 30719 68126
rect 30755 68001 30869 68159
tri 30905 68126 30921 68142 se
rect 30921 68126 30998 68142
rect 30905 68060 30998 68126
rect 30626 67925 30998 68001
rect 30626 67800 30719 67866
rect 30626 67784 30703 67800
tri 30703 67784 30719 67800 nw
rect 30755 67767 30869 67925
rect 30905 67800 30998 67866
tri 30905 67784 30921 67800 ne
rect 30921 67784 30998 67800
rect 30738 67685 30886 67767
rect 30626 67652 30703 67668
tri 30703 67652 30719 67668 sw
rect 30626 67586 30719 67652
rect 30626 67484 30719 67550
rect 30626 67468 30703 67484
tri 30703 67468 30719 67484 nw
rect 30755 67451 30869 67685
tri 30905 67652 30921 67668 se
rect 30921 67652 30998 67668
rect 30905 67586 30998 67652
rect 30905 67484 30998 67550
tri 30905 67468 30921 67484 ne
rect 30921 67468 30998 67484
rect 30738 67369 30886 67451
rect 30626 67336 30703 67352
tri 30703 67336 30719 67352 sw
rect 30626 67270 30719 67336
rect 30755 67211 30869 67369
tri 30905 67336 30921 67352 se
rect 30921 67336 30998 67352
rect 30905 67270 30998 67336
rect 30626 67135 30998 67211
rect 30626 67010 30719 67076
rect 30626 66994 30703 67010
tri 30703 66994 30719 67010 nw
rect 30755 66977 30869 67135
rect 30905 67010 30998 67076
tri 30905 66994 30921 67010 ne
rect 30921 66994 30998 67010
rect 30738 66895 30886 66977
rect 30626 66862 30703 66878
tri 30703 66862 30719 66878 sw
rect 30626 66796 30719 66862
rect 30626 66694 30719 66760
rect 30626 66678 30703 66694
tri 30703 66678 30719 66694 nw
rect 30755 66661 30869 66895
tri 30905 66862 30921 66878 se
rect 30921 66862 30998 66878
rect 30905 66796 30998 66862
rect 30905 66694 30998 66760
tri 30905 66678 30921 66694 ne
rect 30921 66678 30998 66694
rect 30738 66579 30886 66661
rect 30626 66546 30703 66562
tri 30703 66546 30719 66562 sw
rect 30626 66480 30719 66546
rect 30755 66421 30869 66579
tri 30905 66546 30921 66562 se
rect 30921 66546 30998 66562
rect 30905 66480 30998 66546
rect 30626 66345 30998 66421
rect 30626 66220 30719 66286
rect 30626 66204 30703 66220
tri 30703 66204 30719 66220 nw
rect 30755 66187 30869 66345
rect 30905 66220 30998 66286
tri 30905 66204 30921 66220 ne
rect 30921 66204 30998 66220
rect 30738 66105 30886 66187
rect 30626 66072 30703 66088
tri 30703 66072 30719 66088 sw
rect 30626 66006 30719 66072
rect 30626 65904 30719 65970
rect 30626 65888 30703 65904
tri 30703 65888 30719 65904 nw
rect 30755 65871 30869 66105
tri 30905 66072 30921 66088 se
rect 30921 66072 30998 66088
rect 30905 66006 30998 66072
rect 30905 65904 30998 65970
tri 30905 65888 30921 65904 ne
rect 30921 65888 30998 65904
rect 30738 65789 30886 65871
rect 30626 65756 30703 65772
tri 30703 65756 30719 65772 sw
rect 30626 65690 30719 65756
rect 30755 65631 30869 65789
tri 30905 65756 30921 65772 se
rect 30921 65756 30998 65772
rect 30905 65690 30998 65756
rect 30626 65555 30998 65631
rect 30626 65430 30719 65496
rect 30626 65414 30703 65430
tri 30703 65414 30719 65430 nw
rect 30755 65397 30869 65555
rect 30905 65430 30998 65496
tri 30905 65414 30921 65430 ne
rect 30921 65414 30998 65430
rect 30738 65315 30886 65397
rect 30626 65282 30703 65298
tri 30703 65282 30719 65298 sw
rect 30626 65216 30719 65282
rect 30626 65114 30719 65180
rect 30626 65098 30703 65114
tri 30703 65098 30719 65114 nw
rect 30755 65081 30869 65315
tri 30905 65282 30921 65298 se
rect 30921 65282 30998 65298
rect 30905 65216 30998 65282
rect 30905 65114 30998 65180
tri 30905 65098 30921 65114 ne
rect 30921 65098 30998 65114
rect 30738 64999 30886 65081
rect 30626 64966 30703 64982
tri 30703 64966 30719 64982 sw
rect 30626 64900 30719 64966
rect 30755 64841 30869 64999
tri 30905 64966 30921 64982 se
rect 30921 64966 30998 64982
rect 30905 64900 30998 64966
rect 30626 64765 30998 64841
rect 30626 64640 30719 64706
rect 30626 64624 30703 64640
tri 30703 64624 30719 64640 nw
rect 30755 64607 30869 64765
rect 30905 64640 30998 64706
tri 30905 64624 30921 64640 ne
rect 30921 64624 30998 64640
rect 30738 64525 30886 64607
rect 30626 64492 30703 64508
tri 30703 64492 30719 64508 sw
rect 30626 64426 30719 64492
rect 30626 64324 30719 64390
rect 30626 64308 30703 64324
tri 30703 64308 30719 64324 nw
rect 30755 64291 30869 64525
tri 30905 64492 30921 64508 se
rect 30921 64492 30998 64508
rect 30905 64426 30998 64492
rect 30905 64324 30998 64390
tri 30905 64308 30921 64324 ne
rect 30921 64308 30998 64324
rect 30738 64209 30886 64291
rect 30626 64176 30703 64192
tri 30703 64176 30719 64192 sw
rect 30626 64110 30719 64176
rect 30755 64051 30869 64209
tri 30905 64176 30921 64192 se
rect 30921 64176 30998 64192
rect 30905 64110 30998 64176
rect 30626 63975 30998 64051
rect 30626 63850 30719 63916
rect 30626 63834 30703 63850
tri 30703 63834 30719 63850 nw
rect 30755 63817 30869 63975
rect 30905 63850 30998 63916
tri 30905 63834 30921 63850 ne
rect 30921 63834 30998 63850
rect 30738 63735 30886 63817
rect 30626 63702 30703 63718
tri 30703 63702 30719 63718 sw
rect 30626 63636 30719 63702
rect 30626 63534 30719 63600
rect 30626 63518 30703 63534
tri 30703 63518 30719 63534 nw
rect 30755 63501 30869 63735
tri 30905 63702 30921 63718 se
rect 30921 63702 30998 63718
rect 30905 63636 30998 63702
rect 30905 63534 30998 63600
tri 30905 63518 30921 63534 ne
rect 30921 63518 30998 63534
rect 30738 63419 30886 63501
rect 30626 63386 30703 63402
tri 30703 63386 30719 63402 sw
rect 30626 63320 30719 63386
rect 30755 63261 30869 63419
tri 30905 63386 30921 63402 se
rect 30921 63386 30998 63402
rect 30905 63320 30998 63386
rect 30626 63185 30998 63261
rect 30626 63060 30719 63126
rect 30626 63044 30703 63060
tri 30703 63044 30719 63060 nw
rect 30755 63027 30869 63185
rect 30905 63060 30998 63126
tri 30905 63044 30921 63060 ne
rect 30921 63044 30998 63060
rect 30738 62945 30886 63027
rect 30626 62912 30703 62928
tri 30703 62912 30719 62928 sw
rect 30626 62846 30719 62912
rect 30626 62744 30719 62810
rect 30626 62728 30703 62744
tri 30703 62728 30719 62744 nw
rect 30755 62711 30869 62945
tri 30905 62912 30921 62928 se
rect 30921 62912 30998 62928
rect 30905 62846 30998 62912
rect 30905 62744 30998 62810
tri 30905 62728 30921 62744 ne
rect 30921 62728 30998 62744
rect 30738 62629 30886 62711
rect 30626 62596 30703 62612
tri 30703 62596 30719 62612 sw
rect 30626 62530 30719 62596
rect 30755 62471 30869 62629
tri 30905 62596 30921 62612 se
rect 30921 62596 30998 62612
rect 30905 62530 30998 62596
rect 30626 62395 30998 62471
rect 30626 62270 30719 62336
rect 30626 62254 30703 62270
tri 30703 62254 30719 62270 nw
rect 30755 62237 30869 62395
rect 30905 62270 30998 62336
tri 30905 62254 30921 62270 ne
rect 30921 62254 30998 62270
rect 30738 62155 30886 62237
rect 30626 62122 30703 62138
tri 30703 62122 30719 62138 sw
rect 30626 62056 30719 62122
rect 30626 61954 30719 62020
rect 30626 61938 30703 61954
tri 30703 61938 30719 61954 nw
rect 30755 61921 30869 62155
tri 30905 62122 30921 62138 se
rect 30921 62122 30998 62138
rect 30905 62056 30998 62122
rect 30905 61954 30998 62020
tri 30905 61938 30921 61954 ne
rect 30921 61938 30998 61954
rect 30738 61839 30886 61921
rect 30626 61806 30703 61822
tri 30703 61806 30719 61822 sw
rect 30626 61740 30719 61806
rect 30755 61681 30869 61839
tri 30905 61806 30921 61822 se
rect 30921 61806 30998 61822
rect 30905 61740 30998 61806
rect 30626 61605 30998 61681
rect 30626 61480 30719 61546
rect 30626 61464 30703 61480
tri 30703 61464 30719 61480 nw
rect 30755 61447 30869 61605
rect 30905 61480 30998 61546
tri 30905 61464 30921 61480 ne
rect 30921 61464 30998 61480
rect 30738 61365 30886 61447
rect 30626 61332 30703 61348
tri 30703 61332 30719 61348 sw
rect 30626 61266 30719 61332
rect 30626 61164 30719 61230
rect 30626 61148 30703 61164
tri 30703 61148 30719 61164 nw
rect 30755 61131 30869 61365
tri 30905 61332 30921 61348 se
rect 30921 61332 30998 61348
rect 30905 61266 30998 61332
rect 30905 61164 30998 61230
tri 30905 61148 30921 61164 ne
rect 30921 61148 30998 61164
rect 30738 61049 30886 61131
rect 30626 61016 30703 61032
tri 30703 61016 30719 61032 sw
rect 30626 60950 30719 61016
rect 30755 60891 30869 61049
tri 30905 61016 30921 61032 se
rect 30921 61016 30998 61032
rect 30905 60950 30998 61016
rect 30626 60815 30998 60891
rect 30626 60690 30719 60756
rect 30626 60674 30703 60690
tri 30703 60674 30719 60690 nw
rect 30755 60657 30869 60815
rect 30905 60690 30998 60756
tri 30905 60674 30921 60690 ne
rect 30921 60674 30998 60690
rect 30738 60575 30886 60657
rect 30626 60542 30703 60558
tri 30703 60542 30719 60558 sw
rect 30626 60476 30719 60542
rect 30626 60374 30719 60440
rect 30626 60358 30703 60374
tri 30703 60358 30719 60374 nw
rect 30755 60341 30869 60575
tri 30905 60542 30921 60558 se
rect 30921 60542 30998 60558
rect 30905 60476 30998 60542
rect 30905 60374 30998 60440
tri 30905 60358 30921 60374 ne
rect 30921 60358 30998 60374
rect 30738 60259 30886 60341
rect 30626 60226 30703 60242
tri 30703 60226 30719 60242 sw
rect 30626 60160 30719 60226
rect 30755 60101 30869 60259
tri 30905 60226 30921 60242 se
rect 30921 60226 30998 60242
rect 30905 60160 30998 60226
rect 30626 60025 30998 60101
rect 30626 59900 30719 59966
rect 30626 59884 30703 59900
tri 30703 59884 30719 59900 nw
rect 30755 59867 30869 60025
rect 30905 59900 30998 59966
tri 30905 59884 30921 59900 ne
rect 30921 59884 30998 59900
rect 30738 59785 30886 59867
rect 30626 59752 30703 59768
tri 30703 59752 30719 59768 sw
rect 30626 59686 30719 59752
rect 30626 59584 30719 59650
rect 30626 59568 30703 59584
tri 30703 59568 30719 59584 nw
rect 30755 59551 30869 59785
tri 30905 59752 30921 59768 se
rect 30921 59752 30998 59768
rect 30905 59686 30998 59752
rect 30905 59584 30998 59650
tri 30905 59568 30921 59584 ne
rect 30921 59568 30998 59584
rect 30738 59469 30886 59551
rect 30626 59436 30703 59452
tri 30703 59436 30719 59452 sw
rect 30626 59370 30719 59436
rect 30755 59311 30869 59469
tri 30905 59436 30921 59452 se
rect 30921 59436 30998 59452
rect 30905 59370 30998 59436
rect 30626 59235 30998 59311
rect 30626 59110 30719 59176
rect 30626 59094 30703 59110
tri 30703 59094 30719 59110 nw
rect 30755 59077 30869 59235
rect 30905 59110 30998 59176
tri 30905 59094 30921 59110 ne
rect 30921 59094 30998 59110
rect 30738 58995 30886 59077
rect 30626 58962 30703 58978
tri 30703 58962 30719 58978 sw
rect 30626 58896 30719 58962
rect 30626 58794 30719 58860
rect 30626 58778 30703 58794
tri 30703 58778 30719 58794 nw
rect 30755 58761 30869 58995
tri 30905 58962 30921 58978 se
rect 30921 58962 30998 58978
rect 30905 58896 30998 58962
rect 30905 58794 30998 58860
tri 30905 58778 30921 58794 ne
rect 30921 58778 30998 58794
rect 30738 58679 30886 58761
rect 30626 58646 30703 58662
tri 30703 58646 30719 58662 sw
rect 30626 58580 30719 58646
rect 30755 58521 30869 58679
tri 30905 58646 30921 58662 se
rect 30921 58646 30998 58662
rect 30905 58580 30998 58646
rect 30626 58445 30998 58521
rect 30626 58320 30719 58386
rect 30626 58304 30703 58320
tri 30703 58304 30719 58320 nw
rect 30755 58287 30869 58445
rect 30905 58320 30998 58386
tri 30905 58304 30921 58320 ne
rect 30921 58304 30998 58320
rect 30738 58205 30886 58287
rect 30626 58172 30703 58188
tri 30703 58172 30719 58188 sw
rect 30626 58106 30719 58172
rect 30626 58004 30719 58070
rect 30626 57988 30703 58004
tri 30703 57988 30719 58004 nw
rect 30755 57971 30869 58205
tri 30905 58172 30921 58188 se
rect 30921 58172 30998 58188
rect 30905 58106 30998 58172
rect 30905 58004 30998 58070
tri 30905 57988 30921 58004 ne
rect 30921 57988 30998 58004
rect 30738 57889 30886 57971
rect 30626 57856 30703 57872
tri 30703 57856 30719 57872 sw
rect 30626 57790 30719 57856
rect 30755 57731 30869 57889
tri 30905 57856 30921 57872 se
rect 30921 57856 30998 57872
rect 30905 57790 30998 57856
rect 30626 57655 30998 57731
rect 30626 57530 30719 57596
rect 30626 57514 30703 57530
tri 30703 57514 30719 57530 nw
rect 30755 57497 30869 57655
rect 30905 57530 30998 57596
tri 30905 57514 30921 57530 ne
rect 30921 57514 30998 57530
rect 30738 57415 30886 57497
rect 30626 57382 30703 57398
tri 30703 57382 30719 57398 sw
rect 30626 57316 30719 57382
rect 30626 57214 30719 57280
rect 30626 57198 30703 57214
tri 30703 57198 30719 57214 nw
rect 30755 57181 30869 57415
tri 30905 57382 30921 57398 se
rect 30921 57382 30998 57398
rect 30905 57316 30998 57382
rect 30905 57214 30998 57280
tri 30905 57198 30921 57214 ne
rect 30921 57198 30998 57214
rect 30738 57099 30886 57181
rect 30626 57066 30703 57082
tri 30703 57066 30719 57082 sw
rect 30626 57000 30719 57066
rect 30755 56941 30869 57099
tri 30905 57066 30921 57082 se
rect 30921 57066 30998 57082
rect 30905 57000 30998 57066
rect 30626 56865 30998 56941
rect 30626 56740 30719 56806
rect 30626 56724 30703 56740
tri 30703 56724 30719 56740 nw
rect 30755 56707 30869 56865
rect 30905 56740 30998 56806
tri 30905 56724 30921 56740 ne
rect 30921 56724 30998 56740
rect 30738 56625 30886 56707
rect 30626 56592 30703 56608
tri 30703 56592 30719 56608 sw
rect 30626 56526 30719 56592
rect 30626 56424 30719 56490
rect 30626 56408 30703 56424
tri 30703 56408 30719 56424 nw
rect 30755 56391 30869 56625
tri 30905 56592 30921 56608 se
rect 30921 56592 30998 56608
rect 30905 56526 30998 56592
rect 30905 56424 30998 56490
tri 30905 56408 30921 56424 ne
rect 30921 56408 30998 56424
rect 30738 56309 30886 56391
rect 30626 56276 30703 56292
tri 30703 56276 30719 56292 sw
rect 30626 56210 30719 56276
rect 30755 56151 30869 56309
tri 30905 56276 30921 56292 se
rect 30921 56276 30998 56292
rect 30905 56210 30998 56276
rect 30626 56075 30998 56151
rect 30626 55950 30719 56016
rect 30626 55934 30703 55950
tri 30703 55934 30719 55950 nw
rect 30755 55917 30869 56075
rect 30905 55950 30998 56016
tri 30905 55934 30921 55950 ne
rect 30921 55934 30998 55950
rect 30738 55835 30886 55917
rect 30626 55802 30703 55818
tri 30703 55802 30719 55818 sw
rect 30626 55736 30719 55802
rect 30626 55634 30719 55700
rect 30626 55618 30703 55634
tri 30703 55618 30719 55634 nw
rect 30755 55601 30869 55835
tri 30905 55802 30921 55818 se
rect 30921 55802 30998 55818
rect 30905 55736 30998 55802
rect 30905 55634 30998 55700
tri 30905 55618 30921 55634 ne
rect 30921 55618 30998 55634
rect 30738 55519 30886 55601
rect 30626 55486 30703 55502
tri 30703 55486 30719 55502 sw
rect 30626 55420 30719 55486
rect 30755 55361 30869 55519
tri 30905 55486 30921 55502 se
rect 30921 55486 30998 55502
rect 30905 55420 30998 55486
rect 30626 55285 30998 55361
rect 30626 55160 30719 55226
rect 30626 55144 30703 55160
tri 30703 55144 30719 55160 nw
rect 30755 55127 30869 55285
rect 30905 55160 30998 55226
tri 30905 55144 30921 55160 ne
rect 30921 55144 30998 55160
rect 30738 55045 30886 55127
rect 30626 55012 30703 55028
tri 30703 55012 30719 55028 sw
rect 30626 54946 30719 55012
rect 30626 54844 30719 54910
rect 30626 54828 30703 54844
tri 30703 54828 30719 54844 nw
rect 30755 54811 30869 55045
tri 30905 55012 30921 55028 se
rect 30921 55012 30998 55028
rect 30905 54946 30998 55012
rect 30905 54844 30998 54910
tri 30905 54828 30921 54844 ne
rect 30921 54828 30998 54844
rect 30738 54729 30886 54811
rect 30626 54696 30703 54712
tri 30703 54696 30719 54712 sw
rect 30626 54630 30719 54696
rect 30755 54571 30869 54729
tri 30905 54696 30921 54712 se
rect 30921 54696 30998 54712
rect 30905 54630 30998 54696
rect 30626 54495 30998 54571
rect 30626 54370 30719 54436
rect 30626 54354 30703 54370
tri 30703 54354 30719 54370 nw
rect 30755 54337 30869 54495
rect 30905 54370 30998 54436
tri 30905 54354 30921 54370 ne
rect 30921 54354 30998 54370
rect 30738 54255 30886 54337
rect 30626 54222 30703 54238
tri 30703 54222 30719 54238 sw
rect 30626 54156 30719 54222
rect 30626 54054 30719 54120
rect 30626 54038 30703 54054
tri 30703 54038 30719 54054 nw
rect 30755 54021 30869 54255
tri 30905 54222 30921 54238 se
rect 30921 54222 30998 54238
rect 30905 54156 30998 54222
rect 30905 54054 30998 54120
tri 30905 54038 30921 54054 ne
rect 30921 54038 30998 54054
rect 30738 53939 30886 54021
rect 30626 53906 30703 53922
tri 30703 53906 30719 53922 sw
rect 30626 53840 30719 53906
rect 30755 53781 30869 53939
tri 30905 53906 30921 53922 se
rect 30921 53906 30998 53922
rect 30905 53840 30998 53906
rect 30626 53705 30998 53781
rect 30626 53580 30719 53646
rect 30626 53564 30703 53580
tri 30703 53564 30719 53580 nw
rect 30755 53547 30869 53705
rect 30905 53580 30998 53646
tri 30905 53564 30921 53580 ne
rect 30921 53564 30998 53580
rect 30738 53465 30886 53547
rect 30626 53432 30703 53448
tri 30703 53432 30719 53448 sw
rect 30626 53366 30719 53432
rect 30626 53264 30719 53330
rect 30626 53248 30703 53264
tri 30703 53248 30719 53264 nw
rect 30755 53231 30869 53465
tri 30905 53432 30921 53448 se
rect 30921 53432 30998 53448
rect 30905 53366 30998 53432
rect 30905 53264 30998 53330
tri 30905 53248 30921 53264 ne
rect 30921 53248 30998 53264
rect 30738 53149 30886 53231
rect 30626 53116 30703 53132
tri 30703 53116 30719 53132 sw
rect 30626 53050 30719 53116
rect 30755 52991 30869 53149
tri 30905 53116 30921 53132 se
rect 30921 53116 30998 53132
rect 30905 53050 30998 53116
rect 30626 52915 30998 52991
rect 30626 52790 30719 52856
rect 30626 52774 30703 52790
tri 30703 52774 30719 52790 nw
rect 30755 52757 30869 52915
rect 30905 52790 30998 52856
tri 30905 52774 30921 52790 ne
rect 30921 52774 30998 52790
rect 30738 52675 30886 52757
rect 30626 52642 30703 52658
tri 30703 52642 30719 52658 sw
rect 30626 52576 30719 52642
rect 30626 52474 30719 52540
rect 30626 52458 30703 52474
tri 30703 52458 30719 52474 nw
rect 30755 52441 30869 52675
tri 30905 52642 30921 52658 se
rect 30921 52642 30998 52658
rect 30905 52576 30998 52642
rect 30905 52474 30998 52540
tri 30905 52458 30921 52474 ne
rect 30921 52458 30998 52474
rect 30738 52359 30886 52441
rect 30626 52326 30703 52342
tri 30703 52326 30719 52342 sw
rect 30626 52260 30719 52326
rect 30755 52201 30869 52359
tri 30905 52326 30921 52342 se
rect 30921 52326 30998 52342
rect 30905 52260 30998 52326
rect 30626 52125 30998 52201
rect 30626 52000 30719 52066
rect 30626 51984 30703 52000
tri 30703 51984 30719 52000 nw
rect 30755 51967 30869 52125
rect 30905 52000 30998 52066
tri 30905 51984 30921 52000 ne
rect 30921 51984 30998 52000
rect 30738 51885 30886 51967
rect 30626 51852 30703 51868
tri 30703 51852 30719 51868 sw
rect 30626 51786 30719 51852
rect 30626 51684 30719 51750
rect 30626 51668 30703 51684
tri 30703 51668 30719 51684 nw
rect 30755 51651 30869 51885
tri 30905 51852 30921 51868 se
rect 30921 51852 30998 51868
rect 30905 51786 30998 51852
rect 30905 51684 30998 51750
tri 30905 51668 30921 51684 ne
rect 30921 51668 30998 51684
rect 30738 51569 30886 51651
rect 30626 51536 30703 51552
tri 30703 51536 30719 51552 sw
rect 30626 51470 30719 51536
rect 30755 51411 30869 51569
tri 30905 51536 30921 51552 se
rect 30921 51536 30998 51552
rect 30905 51470 30998 51536
rect 30626 51335 30998 51411
rect 30626 51210 30719 51276
rect 30626 51194 30703 51210
tri 30703 51194 30719 51210 nw
rect 30755 51177 30869 51335
rect 30905 51210 30998 51276
tri 30905 51194 30921 51210 ne
rect 30921 51194 30998 51210
rect 30738 51095 30886 51177
rect 30626 51062 30703 51078
tri 30703 51062 30719 51078 sw
rect 30626 50996 30719 51062
rect 30626 50894 30719 50960
rect 30626 50878 30703 50894
tri 30703 50878 30719 50894 nw
rect 30755 50861 30869 51095
tri 30905 51062 30921 51078 se
rect 30921 51062 30998 51078
rect 30905 50996 30998 51062
rect 30905 50894 30998 50960
tri 30905 50878 30921 50894 ne
rect 30921 50878 30998 50894
rect 30738 50779 30886 50861
rect 30626 50746 30703 50762
tri 30703 50746 30719 50762 sw
rect 30626 50680 30719 50746
rect 30755 50621 30869 50779
tri 30905 50746 30921 50762 se
rect 30921 50746 30998 50762
rect 30905 50680 30998 50746
rect 30626 50545 30998 50621
rect 30626 50420 30719 50486
rect 30626 50404 30703 50420
tri 30703 50404 30719 50420 nw
rect 30755 50387 30869 50545
rect 30905 50420 30998 50486
tri 30905 50404 30921 50420 ne
rect 30921 50404 30998 50420
rect 30738 50305 30886 50387
rect 30626 50272 30703 50288
tri 30703 50272 30719 50288 sw
rect 30626 50206 30719 50272
rect 30626 50104 30719 50170
rect 30626 50088 30703 50104
tri 30703 50088 30719 50104 nw
rect 30755 50071 30869 50305
tri 30905 50272 30921 50288 se
rect 30921 50272 30998 50288
rect 30905 50206 30998 50272
rect 30905 50104 30998 50170
tri 30905 50088 30921 50104 ne
rect 30921 50088 30998 50104
rect 30738 49989 30886 50071
rect 30626 49956 30703 49972
tri 30703 49956 30719 49972 sw
rect 30626 49890 30719 49956
rect 30755 49831 30869 49989
tri 30905 49956 30921 49972 se
rect 30921 49956 30998 49972
rect 30905 49890 30998 49956
rect 30626 49755 30998 49831
rect 30626 49630 30719 49696
rect 30626 49614 30703 49630
tri 30703 49614 30719 49630 nw
rect 30755 49597 30869 49755
rect 30905 49630 30998 49696
tri 30905 49614 30921 49630 ne
rect 30921 49614 30998 49630
rect 30738 49515 30886 49597
rect 30626 49482 30703 49498
tri 30703 49482 30719 49498 sw
rect 30626 49416 30719 49482
rect 30626 49314 30719 49380
rect 30626 49298 30703 49314
tri 30703 49298 30719 49314 nw
rect 30755 49281 30869 49515
tri 30905 49482 30921 49498 se
rect 30921 49482 30998 49498
rect 30905 49416 30998 49482
rect 30905 49314 30998 49380
tri 30905 49298 30921 49314 ne
rect 30921 49298 30998 49314
rect 30738 49199 30886 49281
rect 30626 49166 30703 49182
tri 30703 49166 30719 49182 sw
rect 30626 49100 30719 49166
rect 30755 49041 30869 49199
tri 30905 49166 30921 49182 se
rect 30921 49166 30998 49182
rect 30905 49100 30998 49166
rect 30626 48965 30998 49041
rect 30626 48840 30719 48906
rect 30626 48824 30703 48840
tri 30703 48824 30719 48840 nw
rect 30755 48807 30869 48965
rect 30905 48840 30998 48906
tri 30905 48824 30921 48840 ne
rect 30921 48824 30998 48840
rect 30738 48725 30886 48807
rect 30626 48692 30703 48708
tri 30703 48692 30719 48708 sw
rect 30626 48626 30719 48692
rect 30626 48524 30719 48590
rect 30626 48508 30703 48524
tri 30703 48508 30719 48524 nw
rect 30755 48491 30869 48725
tri 30905 48692 30921 48708 se
rect 30921 48692 30998 48708
rect 30905 48626 30998 48692
rect 30905 48524 30998 48590
tri 30905 48508 30921 48524 ne
rect 30921 48508 30998 48524
rect 30738 48409 30886 48491
rect 30626 48376 30703 48392
tri 30703 48376 30719 48392 sw
rect 30626 48310 30719 48376
rect 30755 48251 30869 48409
tri 30905 48376 30921 48392 se
rect 30921 48376 30998 48392
rect 30905 48310 30998 48376
rect 30626 48175 30998 48251
rect 30626 48050 30719 48116
rect 30626 48034 30703 48050
tri 30703 48034 30719 48050 nw
rect 30755 48017 30869 48175
rect 30905 48050 30998 48116
tri 30905 48034 30921 48050 ne
rect 30921 48034 30998 48050
rect 30738 47935 30886 48017
rect 30626 47902 30703 47918
tri 30703 47902 30719 47918 sw
rect 30626 47836 30719 47902
rect 30626 47734 30719 47800
rect 30626 47718 30703 47734
tri 30703 47718 30719 47734 nw
rect 30755 47701 30869 47935
tri 30905 47902 30921 47918 se
rect 30921 47902 30998 47918
rect 30905 47836 30998 47902
rect 30905 47734 30998 47800
tri 30905 47718 30921 47734 ne
rect 30921 47718 30998 47734
rect 30738 47619 30886 47701
rect 30626 47586 30703 47602
tri 30703 47586 30719 47602 sw
rect 30626 47520 30719 47586
rect 30755 47461 30869 47619
tri 30905 47586 30921 47602 se
rect 30921 47586 30998 47602
rect 30905 47520 30998 47586
rect 30626 47385 30998 47461
rect 30626 47260 30719 47326
rect 30626 47244 30703 47260
tri 30703 47244 30719 47260 nw
rect 30755 47227 30869 47385
rect 30905 47260 30998 47326
tri 30905 47244 30921 47260 ne
rect 30921 47244 30998 47260
rect 30738 47145 30886 47227
rect 30626 47112 30703 47128
tri 30703 47112 30719 47128 sw
rect 30626 47046 30719 47112
rect 30626 46944 30719 47010
rect 30626 46928 30703 46944
tri 30703 46928 30719 46944 nw
rect 30755 46911 30869 47145
tri 30905 47112 30921 47128 se
rect 30921 47112 30998 47128
rect 30905 47046 30998 47112
rect 30905 46944 30998 47010
tri 30905 46928 30921 46944 ne
rect 30921 46928 30998 46944
rect 30738 46829 30886 46911
rect 30626 46796 30703 46812
tri 30703 46796 30719 46812 sw
rect 30626 46730 30719 46796
rect 30755 46671 30869 46829
tri 30905 46796 30921 46812 se
rect 30921 46796 30998 46812
rect 30905 46730 30998 46796
rect 30626 46595 30998 46671
rect 30626 46470 30719 46536
rect 30626 46454 30703 46470
tri 30703 46454 30719 46470 nw
rect 30755 46437 30869 46595
rect 30905 46470 30998 46536
tri 30905 46454 30921 46470 ne
rect 30921 46454 30998 46470
rect 30738 46355 30886 46437
rect 30626 46322 30703 46338
tri 30703 46322 30719 46338 sw
rect 30626 46256 30719 46322
rect 30626 46154 30719 46220
rect 30626 46138 30703 46154
tri 30703 46138 30719 46154 nw
rect 30755 46121 30869 46355
tri 30905 46322 30921 46338 se
rect 30921 46322 30998 46338
rect 30905 46256 30998 46322
rect 30905 46154 30998 46220
tri 30905 46138 30921 46154 ne
rect 30921 46138 30998 46154
rect 30738 46039 30886 46121
rect 30626 46006 30703 46022
tri 30703 46006 30719 46022 sw
rect 30626 45940 30719 46006
rect 30755 45881 30869 46039
tri 30905 46006 30921 46022 se
rect 30921 46006 30998 46022
rect 30905 45940 30998 46006
rect 30626 45805 30998 45881
rect 30626 45680 30719 45746
rect 30626 45664 30703 45680
tri 30703 45664 30719 45680 nw
rect 30755 45647 30869 45805
rect 30905 45680 30998 45746
tri 30905 45664 30921 45680 ne
rect 30921 45664 30998 45680
rect 30738 45565 30886 45647
rect 30626 45532 30703 45548
tri 30703 45532 30719 45548 sw
rect 30626 45466 30719 45532
rect 30626 45364 30719 45430
rect 30626 45348 30703 45364
tri 30703 45348 30719 45364 nw
rect 30755 45331 30869 45565
tri 30905 45532 30921 45548 se
rect 30921 45532 30998 45548
rect 30905 45466 30998 45532
rect 30905 45364 30998 45430
tri 30905 45348 30921 45364 ne
rect 30921 45348 30998 45364
rect 30738 45249 30886 45331
rect 30626 45216 30703 45232
tri 30703 45216 30719 45232 sw
rect 30626 45150 30719 45216
rect 30755 45091 30869 45249
tri 30905 45216 30921 45232 se
rect 30921 45216 30998 45232
rect 30905 45150 30998 45216
rect 30626 45015 30998 45091
rect 30626 44890 30719 44956
rect 30626 44874 30703 44890
tri 30703 44874 30719 44890 nw
rect 30755 44857 30869 45015
rect 30905 44890 30998 44956
tri 30905 44874 30921 44890 ne
rect 30921 44874 30998 44890
rect 30738 44775 30886 44857
rect 30626 44742 30703 44758
tri 30703 44742 30719 44758 sw
rect 30626 44676 30719 44742
rect 30626 44574 30719 44640
rect 30626 44558 30703 44574
tri 30703 44558 30719 44574 nw
rect 30755 44541 30869 44775
tri 30905 44742 30921 44758 se
rect 30921 44742 30998 44758
rect 30905 44676 30998 44742
rect 30905 44574 30998 44640
tri 30905 44558 30921 44574 ne
rect 30921 44558 30998 44574
rect 30738 44459 30886 44541
rect 30626 44426 30703 44442
tri 30703 44426 30719 44442 sw
rect 30626 44360 30719 44426
rect 30755 44301 30869 44459
tri 30905 44426 30921 44442 se
rect 30921 44426 30998 44442
rect 30905 44360 30998 44426
rect 30626 44225 30998 44301
rect 30626 44100 30719 44166
rect 30626 44084 30703 44100
tri 30703 44084 30719 44100 nw
rect 30755 44067 30869 44225
rect 30905 44100 30998 44166
tri 30905 44084 30921 44100 ne
rect 30921 44084 30998 44100
rect 30738 43985 30886 44067
rect 30626 43952 30703 43968
tri 30703 43952 30719 43968 sw
rect 30626 43886 30719 43952
rect 30626 43784 30719 43850
rect 30626 43768 30703 43784
tri 30703 43768 30719 43784 nw
rect 30755 43751 30869 43985
tri 30905 43952 30921 43968 se
rect 30921 43952 30998 43968
rect 30905 43886 30998 43952
rect 30905 43784 30998 43850
tri 30905 43768 30921 43784 ne
rect 30921 43768 30998 43784
rect 30738 43669 30886 43751
rect 30626 43636 30703 43652
tri 30703 43636 30719 43652 sw
rect 30626 43570 30719 43636
rect 30755 43511 30869 43669
tri 30905 43636 30921 43652 se
rect 30921 43636 30998 43652
rect 30905 43570 30998 43636
rect 30626 43435 30998 43511
rect 30626 43310 30719 43376
rect 30626 43294 30703 43310
tri 30703 43294 30719 43310 nw
rect 30755 43277 30869 43435
rect 30905 43310 30998 43376
tri 30905 43294 30921 43310 ne
rect 30921 43294 30998 43310
rect 30738 43195 30886 43277
rect 30626 43162 30703 43178
tri 30703 43162 30719 43178 sw
rect 30626 43096 30719 43162
rect 30626 42994 30719 43060
rect 30626 42978 30703 42994
tri 30703 42978 30719 42994 nw
rect 30755 42961 30869 43195
tri 30905 43162 30921 43178 se
rect 30921 43162 30998 43178
rect 30905 43096 30998 43162
rect 30905 42994 30998 43060
tri 30905 42978 30921 42994 ne
rect 30921 42978 30998 42994
rect 30738 42879 30886 42961
rect 30626 42846 30703 42862
tri 30703 42846 30719 42862 sw
rect 30626 42780 30719 42846
rect 30755 42721 30869 42879
tri 30905 42846 30921 42862 se
rect 30921 42846 30998 42862
rect 30905 42780 30998 42846
rect 30626 42645 30998 42721
rect 30626 42520 30719 42586
rect 30626 42504 30703 42520
tri 30703 42504 30719 42520 nw
rect 30755 42487 30869 42645
rect 30905 42520 30998 42586
tri 30905 42504 30921 42520 ne
rect 30921 42504 30998 42520
rect 30738 42405 30886 42487
rect 30626 42372 30703 42388
tri 30703 42372 30719 42388 sw
rect 30626 42306 30719 42372
rect 30626 42204 30719 42270
rect 30626 42188 30703 42204
tri 30703 42188 30719 42204 nw
rect 30755 42171 30869 42405
tri 30905 42372 30921 42388 se
rect 30921 42372 30998 42388
rect 30905 42306 30998 42372
rect 30905 42204 30998 42270
tri 30905 42188 30921 42204 ne
rect 30921 42188 30998 42204
rect 30738 42089 30886 42171
rect 30626 42056 30703 42072
tri 30703 42056 30719 42072 sw
rect 30626 41990 30719 42056
rect 30755 41931 30869 42089
tri 30905 42056 30921 42072 se
rect 30921 42056 30998 42072
rect 30905 41990 30998 42056
rect 30626 41855 30998 41931
rect 30626 41730 30719 41796
rect 30626 41714 30703 41730
tri 30703 41714 30719 41730 nw
rect 30755 41697 30869 41855
rect 30905 41730 30998 41796
tri 30905 41714 30921 41730 ne
rect 30921 41714 30998 41730
rect 30738 41615 30886 41697
rect 30626 41582 30703 41598
tri 30703 41582 30719 41598 sw
rect 30626 41516 30719 41582
rect 30626 41414 30719 41480
rect 30626 41398 30703 41414
tri 30703 41398 30719 41414 nw
rect 30755 41381 30869 41615
tri 30905 41582 30921 41598 se
rect 30921 41582 30998 41598
rect 30905 41516 30998 41582
rect 30905 41414 30998 41480
tri 30905 41398 30921 41414 ne
rect 30921 41398 30998 41414
rect 30738 41299 30886 41381
rect 30626 41266 30703 41282
tri 30703 41266 30719 41282 sw
rect 30626 41200 30719 41266
rect 30755 41141 30869 41299
tri 30905 41266 30921 41282 se
rect 30921 41266 30998 41282
rect 30905 41200 30998 41266
rect 30626 41065 30998 41141
rect 30626 40940 30719 41006
rect 30626 40924 30703 40940
tri 30703 40924 30719 40940 nw
rect 30755 40907 30869 41065
rect 30905 40940 30998 41006
tri 30905 40924 30921 40940 ne
rect 30921 40924 30998 40940
rect 30738 40825 30886 40907
rect 30626 40792 30703 40808
tri 30703 40792 30719 40808 sw
rect 30626 40726 30719 40792
rect 30626 40624 30719 40690
rect 30626 40608 30703 40624
tri 30703 40608 30719 40624 nw
rect 30755 40591 30869 40825
tri 30905 40792 30921 40808 se
rect 30921 40792 30998 40808
rect 30905 40726 30998 40792
rect 30905 40624 30998 40690
tri 30905 40608 30921 40624 ne
rect 30921 40608 30998 40624
rect 30738 40509 30886 40591
rect 30626 40476 30703 40492
tri 30703 40476 30719 40492 sw
rect 30626 40410 30719 40476
rect 30755 40351 30869 40509
tri 30905 40476 30921 40492 se
rect 30921 40476 30998 40492
rect 30905 40410 30998 40476
rect 30626 40275 30998 40351
rect 30626 40150 30719 40216
rect 30626 40134 30703 40150
tri 30703 40134 30719 40150 nw
rect 30755 40117 30869 40275
rect 30905 40150 30998 40216
tri 30905 40134 30921 40150 ne
rect 30921 40134 30998 40150
rect 30738 40035 30886 40117
rect 30626 40002 30703 40018
tri 30703 40002 30719 40018 sw
rect 30626 39936 30719 40002
rect 30626 39834 30719 39900
rect 30626 39818 30703 39834
tri 30703 39818 30719 39834 nw
rect 30755 39801 30869 40035
tri 30905 40002 30921 40018 se
rect 30921 40002 30998 40018
rect 30905 39936 30998 40002
rect 30905 39834 30998 39900
tri 30905 39818 30921 39834 ne
rect 30921 39818 30998 39834
rect 30738 39719 30886 39801
rect 30626 39686 30703 39702
tri 30703 39686 30719 39702 sw
rect 30626 39620 30719 39686
rect 30755 39561 30869 39719
tri 30905 39686 30921 39702 se
rect 30921 39686 30998 39702
rect 30905 39620 30998 39686
rect 30626 39485 30998 39561
rect 30626 39360 30719 39426
rect 30626 39344 30703 39360
tri 30703 39344 30719 39360 nw
rect 30755 39327 30869 39485
rect 30905 39360 30998 39426
tri 30905 39344 30921 39360 ne
rect 30921 39344 30998 39360
rect 30738 39245 30886 39327
rect 30626 39212 30703 39228
tri 30703 39212 30719 39228 sw
rect 30626 39146 30719 39212
rect 30626 39044 30719 39110
rect 30626 39028 30703 39044
tri 30703 39028 30719 39044 nw
rect 30755 39011 30869 39245
tri 30905 39212 30921 39228 se
rect 30921 39212 30998 39228
rect 30905 39146 30998 39212
rect 30905 39044 30998 39110
tri 30905 39028 30921 39044 ne
rect 30921 39028 30998 39044
rect 30738 38929 30886 39011
rect 30626 38896 30703 38912
tri 30703 38896 30719 38912 sw
rect 30626 38830 30719 38896
rect 30755 38771 30869 38929
tri 30905 38896 30921 38912 se
rect 30921 38896 30998 38912
rect 30905 38830 30998 38896
rect 30626 38695 30998 38771
rect 30626 38570 30719 38636
rect 30626 38554 30703 38570
tri 30703 38554 30719 38570 nw
rect 30755 38537 30869 38695
rect 30905 38570 30998 38636
tri 30905 38554 30921 38570 ne
rect 30921 38554 30998 38570
rect 30738 38455 30886 38537
rect 30626 38422 30703 38438
tri 30703 38422 30719 38438 sw
rect 30626 38356 30719 38422
rect 30626 38254 30719 38320
rect 30626 38238 30703 38254
tri 30703 38238 30719 38254 nw
rect 30755 38221 30869 38455
tri 30905 38422 30921 38438 se
rect 30921 38422 30998 38438
rect 30905 38356 30998 38422
rect 30905 38254 30998 38320
tri 30905 38238 30921 38254 ne
rect 30921 38238 30998 38254
rect 30738 38139 30886 38221
rect 30626 38106 30703 38122
tri 30703 38106 30719 38122 sw
rect 30626 38040 30719 38106
rect 30755 37981 30869 38139
tri 30905 38106 30921 38122 se
rect 30921 38106 30998 38122
rect 30905 38040 30998 38106
rect 30626 37905 30998 37981
rect 30626 37780 30719 37846
rect 30626 37764 30703 37780
tri 30703 37764 30719 37780 nw
rect 30755 37747 30869 37905
rect 30905 37780 30998 37846
tri 30905 37764 30921 37780 ne
rect 30921 37764 30998 37780
rect 30738 37665 30886 37747
rect 30626 37632 30703 37648
tri 30703 37632 30719 37648 sw
rect 30626 37566 30719 37632
rect 30626 37464 30719 37530
rect 30626 37448 30703 37464
tri 30703 37448 30719 37464 nw
rect 30755 37431 30869 37665
tri 30905 37632 30921 37648 se
rect 30921 37632 30998 37648
rect 30905 37566 30998 37632
rect 30905 37464 30998 37530
tri 30905 37448 30921 37464 ne
rect 30921 37448 30998 37464
rect 30738 37349 30886 37431
rect 30626 37316 30703 37332
tri 30703 37316 30719 37332 sw
rect 30626 37250 30719 37316
rect 30755 37191 30869 37349
tri 30905 37316 30921 37332 se
rect 30921 37316 30998 37332
rect 30905 37250 30998 37316
rect 30626 37115 30998 37191
rect 30626 36990 30719 37056
rect 30626 36974 30703 36990
tri 30703 36974 30719 36990 nw
rect 30755 36957 30869 37115
rect 30905 36990 30998 37056
tri 30905 36974 30921 36990 ne
rect 30921 36974 30998 36990
rect 30738 36875 30886 36957
rect 30626 36842 30703 36858
tri 30703 36842 30719 36858 sw
rect 30626 36776 30719 36842
rect 30626 36674 30719 36740
rect 30626 36658 30703 36674
tri 30703 36658 30719 36674 nw
rect 30755 36641 30869 36875
tri 30905 36842 30921 36858 se
rect 30921 36842 30998 36858
rect 30905 36776 30998 36842
rect 30905 36674 30998 36740
tri 30905 36658 30921 36674 ne
rect 30921 36658 30998 36674
rect 30738 36559 30886 36641
rect 30626 36526 30703 36542
tri 30703 36526 30719 36542 sw
rect 30626 36460 30719 36526
rect 30755 36401 30869 36559
tri 30905 36526 30921 36542 se
rect 30921 36526 30998 36542
rect 30905 36460 30998 36526
rect 30626 36325 30998 36401
rect 30626 36200 30719 36266
rect 30626 36184 30703 36200
tri 30703 36184 30719 36200 nw
rect 30755 36167 30869 36325
rect 30905 36200 30998 36266
tri 30905 36184 30921 36200 ne
rect 30921 36184 30998 36200
rect 30738 36085 30886 36167
rect 30626 36052 30703 36068
tri 30703 36052 30719 36068 sw
rect 30626 35986 30719 36052
rect 30626 35884 30719 35950
rect 30626 35868 30703 35884
tri 30703 35868 30719 35884 nw
rect 30755 35851 30869 36085
tri 30905 36052 30921 36068 se
rect 30921 36052 30998 36068
rect 30905 35986 30998 36052
rect 30905 35884 30998 35950
tri 30905 35868 30921 35884 ne
rect 30921 35868 30998 35884
rect 30738 35769 30886 35851
rect 30626 35736 30703 35752
tri 30703 35736 30719 35752 sw
rect 30626 35670 30719 35736
rect 30755 35611 30869 35769
tri 30905 35736 30921 35752 se
rect 30921 35736 30998 35752
rect 30905 35670 30998 35736
rect 30626 35535 30998 35611
rect 30626 35410 30719 35476
rect 30626 35394 30703 35410
tri 30703 35394 30719 35410 nw
rect 30755 35377 30869 35535
rect 30905 35410 30998 35476
tri 30905 35394 30921 35410 ne
rect 30921 35394 30998 35410
rect 30738 35295 30886 35377
rect 30626 35262 30703 35278
tri 30703 35262 30719 35278 sw
rect 30626 35196 30719 35262
rect 30626 35094 30719 35160
rect 30626 35078 30703 35094
tri 30703 35078 30719 35094 nw
rect 30755 35061 30869 35295
tri 30905 35262 30921 35278 se
rect 30921 35262 30998 35278
rect 30905 35196 30998 35262
rect 30905 35094 30998 35160
tri 30905 35078 30921 35094 ne
rect 30921 35078 30998 35094
rect 30738 34979 30886 35061
rect 30626 34946 30703 34962
tri 30703 34946 30719 34962 sw
rect 30626 34880 30719 34946
rect 30755 34821 30869 34979
tri 30905 34946 30921 34962 se
rect 30921 34946 30998 34962
rect 30905 34880 30998 34946
rect 30626 34745 30998 34821
rect 30626 34620 30719 34686
rect 30626 34604 30703 34620
tri 30703 34604 30719 34620 nw
rect 30755 34587 30869 34745
rect 30905 34620 30998 34686
tri 30905 34604 30921 34620 ne
rect 30921 34604 30998 34620
rect 30738 34505 30886 34587
rect 30626 34472 30703 34488
tri 30703 34472 30719 34488 sw
rect 30626 34406 30719 34472
rect 30626 34304 30719 34370
rect 30626 34288 30703 34304
tri 30703 34288 30719 34304 nw
rect 30755 34271 30869 34505
tri 30905 34472 30921 34488 se
rect 30921 34472 30998 34488
rect 30905 34406 30998 34472
rect 30905 34304 30998 34370
tri 30905 34288 30921 34304 ne
rect 30921 34288 30998 34304
rect 30738 34189 30886 34271
rect 30626 34156 30703 34172
tri 30703 34156 30719 34172 sw
rect 30626 34090 30719 34156
rect 30755 34031 30869 34189
tri 30905 34156 30921 34172 se
rect 30921 34156 30998 34172
rect 30905 34090 30998 34156
rect 30626 33955 30998 34031
rect 30626 33830 30719 33896
rect 30626 33814 30703 33830
tri 30703 33814 30719 33830 nw
rect 30755 33797 30869 33955
rect 30905 33830 30998 33896
tri 30905 33814 30921 33830 ne
rect 30921 33814 30998 33830
rect 30738 33715 30886 33797
rect 30626 33682 30703 33698
tri 30703 33682 30719 33698 sw
rect 30626 33616 30719 33682
rect 30626 33514 30719 33580
rect 30626 33498 30703 33514
tri 30703 33498 30719 33514 nw
rect 30755 33481 30869 33715
tri 30905 33682 30921 33698 se
rect 30921 33682 30998 33698
rect 30905 33616 30998 33682
rect 30905 33514 30998 33580
tri 30905 33498 30921 33514 ne
rect 30921 33498 30998 33514
rect 30738 33399 30886 33481
rect 30626 33366 30703 33382
tri 30703 33366 30719 33382 sw
rect 30626 33300 30719 33366
rect 30755 33241 30869 33399
tri 30905 33366 30921 33382 se
rect 30921 33366 30998 33382
rect 30905 33300 30998 33366
rect 30626 33165 30998 33241
rect 30626 33040 30719 33106
rect 30626 33024 30703 33040
tri 30703 33024 30719 33040 nw
rect 30755 33007 30869 33165
rect 30905 33040 30998 33106
tri 30905 33024 30921 33040 ne
rect 30921 33024 30998 33040
rect 30738 32925 30886 33007
rect 30626 32892 30703 32908
tri 30703 32892 30719 32908 sw
rect 30626 32826 30719 32892
rect 30626 32724 30719 32790
rect 30626 32708 30703 32724
tri 30703 32708 30719 32724 nw
rect 30755 32691 30869 32925
tri 30905 32892 30921 32908 se
rect 30921 32892 30998 32908
rect 30905 32826 30998 32892
rect 30905 32724 30998 32790
tri 30905 32708 30921 32724 ne
rect 30921 32708 30998 32724
rect 30738 32609 30886 32691
rect 30626 32576 30703 32592
tri 30703 32576 30719 32592 sw
rect 30626 32510 30719 32576
rect 30755 32451 30869 32609
tri 30905 32576 30921 32592 se
rect 30921 32576 30998 32592
rect 30905 32510 30998 32576
rect 30626 32375 30998 32451
rect 30626 32250 30719 32316
rect 30626 32234 30703 32250
tri 30703 32234 30719 32250 nw
rect 30755 32217 30869 32375
rect 30905 32250 30998 32316
tri 30905 32234 30921 32250 ne
rect 30921 32234 30998 32250
rect 30738 32135 30886 32217
rect 30626 32102 30703 32118
tri 30703 32102 30719 32118 sw
rect 30626 32036 30719 32102
rect 30626 31934 30719 32000
rect 30626 31918 30703 31934
tri 30703 31918 30719 31934 nw
rect 30755 31901 30869 32135
tri 30905 32102 30921 32118 se
rect 30921 32102 30998 32118
rect 30905 32036 30998 32102
rect 30905 31934 30998 32000
tri 30905 31918 30921 31934 ne
rect 30921 31918 30998 31934
rect 30738 31819 30886 31901
rect 30626 31786 30703 31802
tri 30703 31786 30719 31802 sw
rect 30626 31720 30719 31786
rect 30755 31661 30869 31819
tri 30905 31786 30921 31802 se
rect 30921 31786 30998 31802
rect 30905 31720 30998 31786
rect 30626 31585 30998 31661
rect 30626 31460 30719 31526
rect 30626 31444 30703 31460
tri 30703 31444 30719 31460 nw
rect 30755 31427 30869 31585
rect 30905 31460 30998 31526
tri 30905 31444 30921 31460 ne
rect 30921 31444 30998 31460
rect 30738 31345 30886 31427
rect 30626 31312 30703 31328
tri 30703 31312 30719 31328 sw
rect 30626 31246 30719 31312
rect 30626 31144 30719 31210
rect 30626 31128 30703 31144
tri 30703 31128 30719 31144 nw
rect 30755 31111 30869 31345
tri 30905 31312 30921 31328 se
rect 30921 31312 30998 31328
rect 30905 31246 30998 31312
rect 30905 31144 30998 31210
tri 30905 31128 30921 31144 ne
rect 30921 31128 30998 31144
rect 30738 31029 30886 31111
rect 30626 30996 30703 31012
tri 30703 30996 30719 31012 sw
rect 30626 30930 30719 30996
rect 30755 30871 30869 31029
tri 30905 30996 30921 31012 se
rect 30921 30996 30998 31012
rect 30905 30930 30998 30996
rect 30626 30795 30998 30871
rect 30626 30670 30719 30736
rect 30626 30654 30703 30670
tri 30703 30654 30719 30670 nw
rect 30755 30637 30869 30795
rect 30905 30670 30998 30736
tri 30905 30654 30921 30670 ne
rect 30921 30654 30998 30670
rect 30738 30555 30886 30637
rect 30626 30522 30703 30538
tri 30703 30522 30719 30538 sw
rect 30626 30456 30719 30522
rect 30626 30354 30719 30420
rect 30626 30338 30703 30354
tri 30703 30338 30719 30354 nw
rect 30755 30321 30869 30555
tri 30905 30522 30921 30538 se
rect 30921 30522 30998 30538
rect 30905 30456 30998 30522
rect 30905 30354 30998 30420
tri 30905 30338 30921 30354 ne
rect 30921 30338 30998 30354
rect 30738 30239 30886 30321
rect 30626 30206 30703 30222
tri 30703 30206 30719 30222 sw
rect 30626 30140 30719 30206
rect 30755 30081 30869 30239
tri 30905 30206 30921 30222 se
rect 30921 30206 30998 30222
rect 30905 30140 30998 30206
rect 30626 30005 30998 30081
rect 30626 29880 30719 29946
rect 30626 29864 30703 29880
tri 30703 29864 30719 29880 nw
rect 30755 29847 30869 30005
rect 30905 29880 30998 29946
tri 30905 29864 30921 29880 ne
rect 30921 29864 30998 29880
rect 30738 29765 30886 29847
rect 30626 29732 30703 29748
tri 30703 29732 30719 29748 sw
rect 30626 29666 30719 29732
rect 30626 29564 30719 29630
rect 30626 29548 30703 29564
tri 30703 29548 30719 29564 nw
rect 30755 29531 30869 29765
tri 30905 29732 30921 29748 se
rect 30921 29732 30998 29748
rect 30905 29666 30998 29732
rect 30905 29564 30998 29630
tri 30905 29548 30921 29564 ne
rect 30921 29548 30998 29564
rect 30738 29449 30886 29531
rect 30626 29416 30703 29432
tri 30703 29416 30719 29432 sw
rect 30626 29350 30719 29416
rect 30755 29291 30869 29449
tri 30905 29416 30921 29432 se
rect 30921 29416 30998 29432
rect 30905 29350 30998 29416
rect 30626 29215 30998 29291
rect 30626 29090 30719 29156
rect 30626 29074 30703 29090
tri 30703 29074 30719 29090 nw
rect 30755 29057 30869 29215
rect 30905 29090 30998 29156
tri 30905 29074 30921 29090 ne
rect 30921 29074 30998 29090
rect 30738 28975 30886 29057
rect 30626 28942 30703 28958
tri 30703 28942 30719 28958 sw
rect 30626 28876 30719 28942
rect 30755 28833 30869 28975
tri 30905 28942 30921 28958 se
rect 30921 28942 30998 28958
rect 30905 28876 30998 28942
rect 31034 28463 31070 80603
rect 31106 28463 31142 80603
rect 31178 80445 31214 80603
rect 31170 80303 31222 80445
rect 31178 28763 31214 80303
rect 31170 28621 31222 28763
rect 31178 28463 31214 28621
rect 31250 28463 31286 80603
rect 31322 28463 31358 80603
rect 31394 28833 31478 80233
rect 31514 28463 31550 80603
rect 31586 28463 31622 80603
rect 31658 80445 31694 80603
rect 31650 80303 31702 80445
rect 31658 28763 31694 80303
rect 31650 28621 31702 28763
rect 31658 28463 31694 28621
rect 31730 28463 31766 80603
rect 31802 28463 31838 80603
rect 31874 80124 31967 80190
rect 31874 80108 31951 80124
tri 31951 80108 31967 80124 nw
rect 32003 80091 32117 80233
rect 32153 80124 32246 80190
tri 32153 80108 32169 80124 ne
rect 32169 80108 32246 80124
rect 31986 80009 32134 80091
rect 31874 79976 31951 79992
tri 31951 79976 31967 79992 sw
rect 31874 79910 31967 79976
rect 32003 79851 32117 80009
tri 32153 79976 32169 79992 se
rect 32169 79976 32246 79992
rect 32153 79910 32246 79976
rect 31874 79775 32246 79851
rect 31874 79650 31967 79716
rect 31874 79634 31951 79650
tri 31951 79634 31967 79650 nw
rect 32003 79617 32117 79775
rect 32153 79650 32246 79716
tri 32153 79634 32169 79650 ne
rect 32169 79634 32246 79650
rect 31986 79535 32134 79617
rect 31874 79502 31951 79518
tri 31951 79502 31967 79518 sw
rect 31874 79436 31967 79502
rect 31874 79334 31967 79400
rect 31874 79318 31951 79334
tri 31951 79318 31967 79334 nw
rect 32003 79301 32117 79535
tri 32153 79502 32169 79518 se
rect 32169 79502 32246 79518
rect 32153 79436 32246 79502
rect 32153 79334 32246 79400
tri 32153 79318 32169 79334 ne
rect 32169 79318 32246 79334
rect 31986 79219 32134 79301
rect 31874 79186 31951 79202
tri 31951 79186 31967 79202 sw
rect 31874 79120 31967 79186
rect 32003 79061 32117 79219
tri 32153 79186 32169 79202 se
rect 32169 79186 32246 79202
rect 32153 79120 32246 79186
rect 31874 78985 32246 79061
rect 31874 78860 31967 78926
rect 31874 78844 31951 78860
tri 31951 78844 31967 78860 nw
rect 32003 78827 32117 78985
rect 32153 78860 32246 78926
tri 32153 78844 32169 78860 ne
rect 32169 78844 32246 78860
rect 31986 78745 32134 78827
rect 31874 78712 31951 78728
tri 31951 78712 31967 78728 sw
rect 31874 78646 31967 78712
rect 31874 78544 31967 78610
rect 31874 78528 31951 78544
tri 31951 78528 31967 78544 nw
rect 32003 78511 32117 78745
tri 32153 78712 32169 78728 se
rect 32169 78712 32246 78728
rect 32153 78646 32246 78712
rect 32153 78544 32246 78610
tri 32153 78528 32169 78544 ne
rect 32169 78528 32246 78544
rect 31986 78429 32134 78511
rect 31874 78396 31951 78412
tri 31951 78396 31967 78412 sw
rect 31874 78330 31967 78396
rect 32003 78271 32117 78429
tri 32153 78396 32169 78412 se
rect 32169 78396 32246 78412
rect 32153 78330 32246 78396
rect 31874 78195 32246 78271
rect 31874 78070 31967 78136
rect 31874 78054 31951 78070
tri 31951 78054 31967 78070 nw
rect 32003 78037 32117 78195
rect 32153 78070 32246 78136
tri 32153 78054 32169 78070 ne
rect 32169 78054 32246 78070
rect 31986 77955 32134 78037
rect 31874 77922 31951 77938
tri 31951 77922 31967 77938 sw
rect 31874 77856 31967 77922
rect 31874 77754 31967 77820
rect 31874 77738 31951 77754
tri 31951 77738 31967 77754 nw
rect 32003 77721 32117 77955
tri 32153 77922 32169 77938 se
rect 32169 77922 32246 77938
rect 32153 77856 32246 77922
rect 32153 77754 32246 77820
tri 32153 77738 32169 77754 ne
rect 32169 77738 32246 77754
rect 31986 77639 32134 77721
rect 31874 77606 31951 77622
tri 31951 77606 31967 77622 sw
rect 31874 77540 31967 77606
rect 32003 77481 32117 77639
tri 32153 77606 32169 77622 se
rect 32169 77606 32246 77622
rect 32153 77540 32246 77606
rect 31874 77405 32246 77481
rect 31874 77280 31967 77346
rect 31874 77264 31951 77280
tri 31951 77264 31967 77280 nw
rect 32003 77247 32117 77405
rect 32153 77280 32246 77346
tri 32153 77264 32169 77280 ne
rect 32169 77264 32246 77280
rect 31986 77165 32134 77247
rect 31874 77132 31951 77148
tri 31951 77132 31967 77148 sw
rect 31874 77066 31967 77132
rect 31874 76964 31967 77030
rect 31874 76948 31951 76964
tri 31951 76948 31967 76964 nw
rect 32003 76931 32117 77165
tri 32153 77132 32169 77148 se
rect 32169 77132 32246 77148
rect 32153 77066 32246 77132
rect 32153 76964 32246 77030
tri 32153 76948 32169 76964 ne
rect 32169 76948 32246 76964
rect 31986 76849 32134 76931
rect 31874 76816 31951 76832
tri 31951 76816 31967 76832 sw
rect 31874 76750 31967 76816
rect 32003 76691 32117 76849
tri 32153 76816 32169 76832 se
rect 32169 76816 32246 76832
rect 32153 76750 32246 76816
rect 31874 76615 32246 76691
rect 31874 76490 31967 76556
rect 31874 76474 31951 76490
tri 31951 76474 31967 76490 nw
rect 32003 76457 32117 76615
rect 32153 76490 32246 76556
tri 32153 76474 32169 76490 ne
rect 32169 76474 32246 76490
rect 31986 76375 32134 76457
rect 31874 76342 31951 76358
tri 31951 76342 31967 76358 sw
rect 31874 76276 31967 76342
rect 31874 76174 31967 76240
rect 31874 76158 31951 76174
tri 31951 76158 31967 76174 nw
rect 32003 76141 32117 76375
tri 32153 76342 32169 76358 se
rect 32169 76342 32246 76358
rect 32153 76276 32246 76342
rect 32153 76174 32246 76240
tri 32153 76158 32169 76174 ne
rect 32169 76158 32246 76174
rect 31986 76059 32134 76141
rect 31874 76026 31951 76042
tri 31951 76026 31967 76042 sw
rect 31874 75960 31967 76026
rect 32003 75901 32117 76059
tri 32153 76026 32169 76042 se
rect 32169 76026 32246 76042
rect 32153 75960 32246 76026
rect 31874 75825 32246 75901
rect 31874 75700 31967 75766
rect 31874 75684 31951 75700
tri 31951 75684 31967 75700 nw
rect 32003 75667 32117 75825
rect 32153 75700 32246 75766
tri 32153 75684 32169 75700 ne
rect 32169 75684 32246 75700
rect 31986 75585 32134 75667
rect 31874 75552 31951 75568
tri 31951 75552 31967 75568 sw
rect 31874 75486 31967 75552
rect 31874 75384 31967 75450
rect 31874 75368 31951 75384
tri 31951 75368 31967 75384 nw
rect 32003 75351 32117 75585
tri 32153 75552 32169 75568 se
rect 32169 75552 32246 75568
rect 32153 75486 32246 75552
rect 32153 75384 32246 75450
tri 32153 75368 32169 75384 ne
rect 32169 75368 32246 75384
rect 31986 75269 32134 75351
rect 31874 75236 31951 75252
tri 31951 75236 31967 75252 sw
rect 31874 75170 31967 75236
rect 32003 75111 32117 75269
tri 32153 75236 32169 75252 se
rect 32169 75236 32246 75252
rect 32153 75170 32246 75236
rect 31874 75035 32246 75111
rect 31874 74910 31967 74976
rect 31874 74894 31951 74910
tri 31951 74894 31967 74910 nw
rect 32003 74877 32117 75035
rect 32153 74910 32246 74976
tri 32153 74894 32169 74910 ne
rect 32169 74894 32246 74910
rect 31986 74795 32134 74877
rect 31874 74762 31951 74778
tri 31951 74762 31967 74778 sw
rect 31874 74696 31967 74762
rect 31874 74594 31967 74660
rect 31874 74578 31951 74594
tri 31951 74578 31967 74594 nw
rect 32003 74561 32117 74795
tri 32153 74762 32169 74778 se
rect 32169 74762 32246 74778
rect 32153 74696 32246 74762
rect 32153 74594 32246 74660
tri 32153 74578 32169 74594 ne
rect 32169 74578 32246 74594
rect 31986 74479 32134 74561
rect 31874 74446 31951 74462
tri 31951 74446 31967 74462 sw
rect 31874 74380 31967 74446
rect 32003 74321 32117 74479
tri 32153 74446 32169 74462 se
rect 32169 74446 32246 74462
rect 32153 74380 32246 74446
rect 31874 74245 32246 74321
rect 31874 74120 31967 74186
rect 31874 74104 31951 74120
tri 31951 74104 31967 74120 nw
rect 32003 74087 32117 74245
rect 32153 74120 32246 74186
tri 32153 74104 32169 74120 ne
rect 32169 74104 32246 74120
rect 31986 74005 32134 74087
rect 31874 73972 31951 73988
tri 31951 73972 31967 73988 sw
rect 31874 73906 31967 73972
rect 31874 73804 31967 73870
rect 31874 73788 31951 73804
tri 31951 73788 31967 73804 nw
rect 32003 73771 32117 74005
tri 32153 73972 32169 73988 se
rect 32169 73972 32246 73988
rect 32153 73906 32246 73972
rect 32153 73804 32246 73870
tri 32153 73788 32169 73804 ne
rect 32169 73788 32246 73804
rect 31986 73689 32134 73771
rect 31874 73656 31951 73672
tri 31951 73656 31967 73672 sw
rect 31874 73590 31967 73656
rect 32003 73531 32117 73689
tri 32153 73656 32169 73672 se
rect 32169 73656 32246 73672
rect 32153 73590 32246 73656
rect 31874 73455 32246 73531
rect 31874 73330 31967 73396
rect 31874 73314 31951 73330
tri 31951 73314 31967 73330 nw
rect 32003 73297 32117 73455
rect 32153 73330 32246 73396
tri 32153 73314 32169 73330 ne
rect 32169 73314 32246 73330
rect 31986 73215 32134 73297
rect 31874 73182 31951 73198
tri 31951 73182 31967 73198 sw
rect 31874 73116 31967 73182
rect 31874 73014 31967 73080
rect 31874 72998 31951 73014
tri 31951 72998 31967 73014 nw
rect 32003 72981 32117 73215
tri 32153 73182 32169 73198 se
rect 32169 73182 32246 73198
rect 32153 73116 32246 73182
rect 32153 73014 32246 73080
tri 32153 72998 32169 73014 ne
rect 32169 72998 32246 73014
rect 31986 72899 32134 72981
rect 31874 72866 31951 72882
tri 31951 72866 31967 72882 sw
rect 31874 72800 31967 72866
rect 32003 72741 32117 72899
tri 32153 72866 32169 72882 se
rect 32169 72866 32246 72882
rect 32153 72800 32246 72866
rect 31874 72665 32246 72741
rect 31874 72540 31967 72606
rect 31874 72524 31951 72540
tri 31951 72524 31967 72540 nw
rect 32003 72507 32117 72665
rect 32153 72540 32246 72606
tri 32153 72524 32169 72540 ne
rect 32169 72524 32246 72540
rect 31986 72425 32134 72507
rect 31874 72392 31951 72408
tri 31951 72392 31967 72408 sw
rect 31874 72326 31967 72392
rect 31874 72224 31967 72290
rect 31874 72208 31951 72224
tri 31951 72208 31967 72224 nw
rect 32003 72191 32117 72425
tri 32153 72392 32169 72408 se
rect 32169 72392 32246 72408
rect 32153 72326 32246 72392
rect 32153 72224 32246 72290
tri 32153 72208 32169 72224 ne
rect 32169 72208 32246 72224
rect 31986 72109 32134 72191
rect 31874 72076 31951 72092
tri 31951 72076 31967 72092 sw
rect 31874 72010 31967 72076
rect 32003 71951 32117 72109
tri 32153 72076 32169 72092 se
rect 32169 72076 32246 72092
rect 32153 72010 32246 72076
rect 31874 71875 32246 71951
rect 31874 71750 31967 71816
rect 31874 71734 31951 71750
tri 31951 71734 31967 71750 nw
rect 32003 71717 32117 71875
rect 32153 71750 32246 71816
tri 32153 71734 32169 71750 ne
rect 32169 71734 32246 71750
rect 31986 71635 32134 71717
rect 31874 71602 31951 71618
tri 31951 71602 31967 71618 sw
rect 31874 71536 31967 71602
rect 31874 71434 31967 71500
rect 31874 71418 31951 71434
tri 31951 71418 31967 71434 nw
rect 32003 71401 32117 71635
tri 32153 71602 32169 71618 se
rect 32169 71602 32246 71618
rect 32153 71536 32246 71602
rect 32153 71434 32246 71500
tri 32153 71418 32169 71434 ne
rect 32169 71418 32246 71434
rect 31986 71319 32134 71401
rect 31874 71286 31951 71302
tri 31951 71286 31967 71302 sw
rect 31874 71220 31967 71286
rect 32003 71161 32117 71319
tri 32153 71286 32169 71302 se
rect 32169 71286 32246 71302
rect 32153 71220 32246 71286
rect 31874 71085 32246 71161
rect 31874 70960 31967 71026
rect 31874 70944 31951 70960
tri 31951 70944 31967 70960 nw
rect 32003 70927 32117 71085
rect 32153 70960 32246 71026
tri 32153 70944 32169 70960 ne
rect 32169 70944 32246 70960
rect 31986 70845 32134 70927
rect 31874 70812 31951 70828
tri 31951 70812 31967 70828 sw
rect 31874 70746 31967 70812
rect 31874 70644 31967 70710
rect 31874 70628 31951 70644
tri 31951 70628 31967 70644 nw
rect 32003 70611 32117 70845
tri 32153 70812 32169 70828 se
rect 32169 70812 32246 70828
rect 32153 70746 32246 70812
rect 32153 70644 32246 70710
tri 32153 70628 32169 70644 ne
rect 32169 70628 32246 70644
rect 31986 70529 32134 70611
rect 31874 70496 31951 70512
tri 31951 70496 31967 70512 sw
rect 31874 70430 31967 70496
rect 32003 70371 32117 70529
tri 32153 70496 32169 70512 se
rect 32169 70496 32246 70512
rect 32153 70430 32246 70496
rect 31874 70295 32246 70371
rect 31874 70170 31967 70236
rect 31874 70154 31951 70170
tri 31951 70154 31967 70170 nw
rect 32003 70137 32117 70295
rect 32153 70170 32246 70236
tri 32153 70154 32169 70170 ne
rect 32169 70154 32246 70170
rect 31986 70055 32134 70137
rect 31874 70022 31951 70038
tri 31951 70022 31967 70038 sw
rect 31874 69956 31967 70022
rect 31874 69854 31967 69920
rect 31874 69838 31951 69854
tri 31951 69838 31967 69854 nw
rect 32003 69821 32117 70055
tri 32153 70022 32169 70038 se
rect 32169 70022 32246 70038
rect 32153 69956 32246 70022
rect 32153 69854 32246 69920
tri 32153 69838 32169 69854 ne
rect 32169 69838 32246 69854
rect 31986 69739 32134 69821
rect 31874 69706 31951 69722
tri 31951 69706 31967 69722 sw
rect 31874 69640 31967 69706
rect 32003 69581 32117 69739
tri 32153 69706 32169 69722 se
rect 32169 69706 32246 69722
rect 32153 69640 32246 69706
rect 31874 69505 32246 69581
rect 31874 69380 31967 69446
rect 31874 69364 31951 69380
tri 31951 69364 31967 69380 nw
rect 32003 69347 32117 69505
rect 32153 69380 32246 69446
tri 32153 69364 32169 69380 ne
rect 32169 69364 32246 69380
rect 31986 69265 32134 69347
rect 31874 69232 31951 69248
tri 31951 69232 31967 69248 sw
rect 31874 69166 31967 69232
rect 31874 69064 31967 69130
rect 31874 69048 31951 69064
tri 31951 69048 31967 69064 nw
rect 32003 69031 32117 69265
tri 32153 69232 32169 69248 se
rect 32169 69232 32246 69248
rect 32153 69166 32246 69232
rect 32153 69064 32246 69130
tri 32153 69048 32169 69064 ne
rect 32169 69048 32246 69064
rect 31986 68949 32134 69031
rect 31874 68916 31951 68932
tri 31951 68916 31967 68932 sw
rect 31874 68850 31967 68916
rect 32003 68791 32117 68949
tri 32153 68916 32169 68932 se
rect 32169 68916 32246 68932
rect 32153 68850 32246 68916
rect 31874 68715 32246 68791
rect 31874 68590 31967 68656
rect 31874 68574 31951 68590
tri 31951 68574 31967 68590 nw
rect 32003 68557 32117 68715
rect 32153 68590 32246 68656
tri 32153 68574 32169 68590 ne
rect 32169 68574 32246 68590
rect 31986 68475 32134 68557
rect 31874 68442 31951 68458
tri 31951 68442 31967 68458 sw
rect 31874 68376 31967 68442
rect 31874 68274 31967 68340
rect 31874 68258 31951 68274
tri 31951 68258 31967 68274 nw
rect 32003 68241 32117 68475
tri 32153 68442 32169 68458 se
rect 32169 68442 32246 68458
rect 32153 68376 32246 68442
rect 32153 68274 32246 68340
tri 32153 68258 32169 68274 ne
rect 32169 68258 32246 68274
rect 31986 68159 32134 68241
rect 31874 68126 31951 68142
tri 31951 68126 31967 68142 sw
rect 31874 68060 31967 68126
rect 32003 68001 32117 68159
tri 32153 68126 32169 68142 se
rect 32169 68126 32246 68142
rect 32153 68060 32246 68126
rect 31874 67925 32246 68001
rect 31874 67800 31967 67866
rect 31874 67784 31951 67800
tri 31951 67784 31967 67800 nw
rect 32003 67767 32117 67925
rect 32153 67800 32246 67866
tri 32153 67784 32169 67800 ne
rect 32169 67784 32246 67800
rect 31986 67685 32134 67767
rect 31874 67652 31951 67668
tri 31951 67652 31967 67668 sw
rect 31874 67586 31967 67652
rect 31874 67484 31967 67550
rect 31874 67468 31951 67484
tri 31951 67468 31967 67484 nw
rect 32003 67451 32117 67685
tri 32153 67652 32169 67668 se
rect 32169 67652 32246 67668
rect 32153 67586 32246 67652
rect 32153 67484 32246 67550
tri 32153 67468 32169 67484 ne
rect 32169 67468 32246 67484
rect 31986 67369 32134 67451
rect 31874 67336 31951 67352
tri 31951 67336 31967 67352 sw
rect 31874 67270 31967 67336
rect 32003 67211 32117 67369
tri 32153 67336 32169 67352 se
rect 32169 67336 32246 67352
rect 32153 67270 32246 67336
rect 31874 67135 32246 67211
rect 31874 67010 31967 67076
rect 31874 66994 31951 67010
tri 31951 66994 31967 67010 nw
rect 32003 66977 32117 67135
rect 32153 67010 32246 67076
tri 32153 66994 32169 67010 ne
rect 32169 66994 32246 67010
rect 31986 66895 32134 66977
rect 31874 66862 31951 66878
tri 31951 66862 31967 66878 sw
rect 31874 66796 31967 66862
rect 31874 66694 31967 66760
rect 31874 66678 31951 66694
tri 31951 66678 31967 66694 nw
rect 32003 66661 32117 66895
tri 32153 66862 32169 66878 se
rect 32169 66862 32246 66878
rect 32153 66796 32246 66862
rect 32153 66694 32246 66760
tri 32153 66678 32169 66694 ne
rect 32169 66678 32246 66694
rect 31986 66579 32134 66661
rect 31874 66546 31951 66562
tri 31951 66546 31967 66562 sw
rect 31874 66480 31967 66546
rect 32003 66421 32117 66579
tri 32153 66546 32169 66562 se
rect 32169 66546 32246 66562
rect 32153 66480 32246 66546
rect 31874 66345 32246 66421
rect 31874 66220 31967 66286
rect 31874 66204 31951 66220
tri 31951 66204 31967 66220 nw
rect 32003 66187 32117 66345
rect 32153 66220 32246 66286
tri 32153 66204 32169 66220 ne
rect 32169 66204 32246 66220
rect 31986 66105 32134 66187
rect 31874 66072 31951 66088
tri 31951 66072 31967 66088 sw
rect 31874 66006 31967 66072
rect 31874 65904 31967 65970
rect 31874 65888 31951 65904
tri 31951 65888 31967 65904 nw
rect 32003 65871 32117 66105
tri 32153 66072 32169 66088 se
rect 32169 66072 32246 66088
rect 32153 66006 32246 66072
rect 32153 65904 32246 65970
tri 32153 65888 32169 65904 ne
rect 32169 65888 32246 65904
rect 31986 65789 32134 65871
rect 31874 65756 31951 65772
tri 31951 65756 31967 65772 sw
rect 31874 65690 31967 65756
rect 32003 65631 32117 65789
tri 32153 65756 32169 65772 se
rect 32169 65756 32246 65772
rect 32153 65690 32246 65756
rect 31874 65555 32246 65631
rect 31874 65430 31967 65496
rect 31874 65414 31951 65430
tri 31951 65414 31967 65430 nw
rect 32003 65397 32117 65555
rect 32153 65430 32246 65496
tri 32153 65414 32169 65430 ne
rect 32169 65414 32246 65430
rect 31986 65315 32134 65397
rect 31874 65282 31951 65298
tri 31951 65282 31967 65298 sw
rect 31874 65216 31967 65282
rect 31874 65114 31967 65180
rect 31874 65098 31951 65114
tri 31951 65098 31967 65114 nw
rect 32003 65081 32117 65315
tri 32153 65282 32169 65298 se
rect 32169 65282 32246 65298
rect 32153 65216 32246 65282
rect 32153 65114 32246 65180
tri 32153 65098 32169 65114 ne
rect 32169 65098 32246 65114
rect 31986 64999 32134 65081
rect 31874 64966 31951 64982
tri 31951 64966 31967 64982 sw
rect 31874 64900 31967 64966
rect 32003 64841 32117 64999
tri 32153 64966 32169 64982 se
rect 32169 64966 32246 64982
rect 32153 64900 32246 64966
rect 31874 64765 32246 64841
rect 31874 64640 31967 64706
rect 31874 64624 31951 64640
tri 31951 64624 31967 64640 nw
rect 32003 64607 32117 64765
rect 32153 64640 32246 64706
tri 32153 64624 32169 64640 ne
rect 32169 64624 32246 64640
rect 31986 64525 32134 64607
rect 31874 64492 31951 64508
tri 31951 64492 31967 64508 sw
rect 31874 64426 31967 64492
rect 31874 64324 31967 64390
rect 31874 64308 31951 64324
tri 31951 64308 31967 64324 nw
rect 32003 64291 32117 64525
tri 32153 64492 32169 64508 se
rect 32169 64492 32246 64508
rect 32153 64426 32246 64492
rect 32153 64324 32246 64390
tri 32153 64308 32169 64324 ne
rect 32169 64308 32246 64324
rect 31986 64209 32134 64291
rect 31874 64176 31951 64192
tri 31951 64176 31967 64192 sw
rect 31874 64110 31967 64176
rect 32003 64051 32117 64209
tri 32153 64176 32169 64192 se
rect 32169 64176 32246 64192
rect 32153 64110 32246 64176
rect 31874 63975 32246 64051
rect 31874 63850 31967 63916
rect 31874 63834 31951 63850
tri 31951 63834 31967 63850 nw
rect 32003 63817 32117 63975
rect 32153 63850 32246 63916
tri 32153 63834 32169 63850 ne
rect 32169 63834 32246 63850
rect 31986 63735 32134 63817
rect 31874 63702 31951 63718
tri 31951 63702 31967 63718 sw
rect 31874 63636 31967 63702
rect 31874 63534 31967 63600
rect 31874 63518 31951 63534
tri 31951 63518 31967 63534 nw
rect 32003 63501 32117 63735
tri 32153 63702 32169 63718 se
rect 32169 63702 32246 63718
rect 32153 63636 32246 63702
rect 32153 63534 32246 63600
tri 32153 63518 32169 63534 ne
rect 32169 63518 32246 63534
rect 31986 63419 32134 63501
rect 31874 63386 31951 63402
tri 31951 63386 31967 63402 sw
rect 31874 63320 31967 63386
rect 32003 63261 32117 63419
tri 32153 63386 32169 63402 se
rect 32169 63386 32246 63402
rect 32153 63320 32246 63386
rect 31874 63185 32246 63261
rect 31874 63060 31967 63126
rect 31874 63044 31951 63060
tri 31951 63044 31967 63060 nw
rect 32003 63027 32117 63185
rect 32153 63060 32246 63126
tri 32153 63044 32169 63060 ne
rect 32169 63044 32246 63060
rect 31986 62945 32134 63027
rect 31874 62912 31951 62928
tri 31951 62912 31967 62928 sw
rect 31874 62846 31967 62912
rect 31874 62744 31967 62810
rect 31874 62728 31951 62744
tri 31951 62728 31967 62744 nw
rect 32003 62711 32117 62945
tri 32153 62912 32169 62928 se
rect 32169 62912 32246 62928
rect 32153 62846 32246 62912
rect 32153 62744 32246 62810
tri 32153 62728 32169 62744 ne
rect 32169 62728 32246 62744
rect 31986 62629 32134 62711
rect 31874 62596 31951 62612
tri 31951 62596 31967 62612 sw
rect 31874 62530 31967 62596
rect 32003 62471 32117 62629
tri 32153 62596 32169 62612 se
rect 32169 62596 32246 62612
rect 32153 62530 32246 62596
rect 31874 62395 32246 62471
rect 31874 62270 31967 62336
rect 31874 62254 31951 62270
tri 31951 62254 31967 62270 nw
rect 32003 62237 32117 62395
rect 32153 62270 32246 62336
tri 32153 62254 32169 62270 ne
rect 32169 62254 32246 62270
rect 31986 62155 32134 62237
rect 31874 62122 31951 62138
tri 31951 62122 31967 62138 sw
rect 31874 62056 31967 62122
rect 31874 61954 31967 62020
rect 31874 61938 31951 61954
tri 31951 61938 31967 61954 nw
rect 32003 61921 32117 62155
tri 32153 62122 32169 62138 se
rect 32169 62122 32246 62138
rect 32153 62056 32246 62122
rect 32153 61954 32246 62020
tri 32153 61938 32169 61954 ne
rect 32169 61938 32246 61954
rect 31986 61839 32134 61921
rect 31874 61806 31951 61822
tri 31951 61806 31967 61822 sw
rect 31874 61740 31967 61806
rect 32003 61681 32117 61839
tri 32153 61806 32169 61822 se
rect 32169 61806 32246 61822
rect 32153 61740 32246 61806
rect 31874 61605 32246 61681
rect 31874 61480 31967 61546
rect 31874 61464 31951 61480
tri 31951 61464 31967 61480 nw
rect 32003 61447 32117 61605
rect 32153 61480 32246 61546
tri 32153 61464 32169 61480 ne
rect 32169 61464 32246 61480
rect 31986 61365 32134 61447
rect 31874 61332 31951 61348
tri 31951 61332 31967 61348 sw
rect 31874 61266 31967 61332
rect 31874 61164 31967 61230
rect 31874 61148 31951 61164
tri 31951 61148 31967 61164 nw
rect 32003 61131 32117 61365
tri 32153 61332 32169 61348 se
rect 32169 61332 32246 61348
rect 32153 61266 32246 61332
rect 32153 61164 32246 61230
tri 32153 61148 32169 61164 ne
rect 32169 61148 32246 61164
rect 31986 61049 32134 61131
rect 31874 61016 31951 61032
tri 31951 61016 31967 61032 sw
rect 31874 60950 31967 61016
rect 32003 60891 32117 61049
tri 32153 61016 32169 61032 se
rect 32169 61016 32246 61032
rect 32153 60950 32246 61016
rect 31874 60815 32246 60891
rect 31874 60690 31967 60756
rect 31874 60674 31951 60690
tri 31951 60674 31967 60690 nw
rect 32003 60657 32117 60815
rect 32153 60690 32246 60756
tri 32153 60674 32169 60690 ne
rect 32169 60674 32246 60690
rect 31986 60575 32134 60657
rect 31874 60542 31951 60558
tri 31951 60542 31967 60558 sw
rect 31874 60476 31967 60542
rect 31874 60374 31967 60440
rect 31874 60358 31951 60374
tri 31951 60358 31967 60374 nw
rect 32003 60341 32117 60575
tri 32153 60542 32169 60558 se
rect 32169 60542 32246 60558
rect 32153 60476 32246 60542
rect 32153 60374 32246 60440
tri 32153 60358 32169 60374 ne
rect 32169 60358 32246 60374
rect 31986 60259 32134 60341
rect 31874 60226 31951 60242
tri 31951 60226 31967 60242 sw
rect 31874 60160 31967 60226
rect 32003 60101 32117 60259
tri 32153 60226 32169 60242 se
rect 32169 60226 32246 60242
rect 32153 60160 32246 60226
rect 31874 60025 32246 60101
rect 31874 59900 31967 59966
rect 31874 59884 31951 59900
tri 31951 59884 31967 59900 nw
rect 32003 59867 32117 60025
rect 32153 59900 32246 59966
tri 32153 59884 32169 59900 ne
rect 32169 59884 32246 59900
rect 31986 59785 32134 59867
rect 31874 59752 31951 59768
tri 31951 59752 31967 59768 sw
rect 31874 59686 31967 59752
rect 31874 59584 31967 59650
rect 31874 59568 31951 59584
tri 31951 59568 31967 59584 nw
rect 32003 59551 32117 59785
tri 32153 59752 32169 59768 se
rect 32169 59752 32246 59768
rect 32153 59686 32246 59752
rect 32153 59584 32246 59650
tri 32153 59568 32169 59584 ne
rect 32169 59568 32246 59584
rect 31986 59469 32134 59551
rect 31874 59436 31951 59452
tri 31951 59436 31967 59452 sw
rect 31874 59370 31967 59436
rect 32003 59311 32117 59469
tri 32153 59436 32169 59452 se
rect 32169 59436 32246 59452
rect 32153 59370 32246 59436
rect 31874 59235 32246 59311
rect 31874 59110 31967 59176
rect 31874 59094 31951 59110
tri 31951 59094 31967 59110 nw
rect 32003 59077 32117 59235
rect 32153 59110 32246 59176
tri 32153 59094 32169 59110 ne
rect 32169 59094 32246 59110
rect 31986 58995 32134 59077
rect 31874 58962 31951 58978
tri 31951 58962 31967 58978 sw
rect 31874 58896 31967 58962
rect 31874 58794 31967 58860
rect 31874 58778 31951 58794
tri 31951 58778 31967 58794 nw
rect 32003 58761 32117 58995
tri 32153 58962 32169 58978 se
rect 32169 58962 32246 58978
rect 32153 58896 32246 58962
rect 32153 58794 32246 58860
tri 32153 58778 32169 58794 ne
rect 32169 58778 32246 58794
rect 31986 58679 32134 58761
rect 31874 58646 31951 58662
tri 31951 58646 31967 58662 sw
rect 31874 58580 31967 58646
rect 32003 58521 32117 58679
tri 32153 58646 32169 58662 se
rect 32169 58646 32246 58662
rect 32153 58580 32246 58646
rect 31874 58445 32246 58521
rect 31874 58320 31967 58386
rect 31874 58304 31951 58320
tri 31951 58304 31967 58320 nw
rect 32003 58287 32117 58445
rect 32153 58320 32246 58386
tri 32153 58304 32169 58320 ne
rect 32169 58304 32246 58320
rect 31986 58205 32134 58287
rect 31874 58172 31951 58188
tri 31951 58172 31967 58188 sw
rect 31874 58106 31967 58172
rect 31874 58004 31967 58070
rect 31874 57988 31951 58004
tri 31951 57988 31967 58004 nw
rect 32003 57971 32117 58205
tri 32153 58172 32169 58188 se
rect 32169 58172 32246 58188
rect 32153 58106 32246 58172
rect 32153 58004 32246 58070
tri 32153 57988 32169 58004 ne
rect 32169 57988 32246 58004
rect 31986 57889 32134 57971
rect 31874 57856 31951 57872
tri 31951 57856 31967 57872 sw
rect 31874 57790 31967 57856
rect 32003 57731 32117 57889
tri 32153 57856 32169 57872 se
rect 32169 57856 32246 57872
rect 32153 57790 32246 57856
rect 31874 57655 32246 57731
rect 31874 57530 31967 57596
rect 31874 57514 31951 57530
tri 31951 57514 31967 57530 nw
rect 32003 57497 32117 57655
rect 32153 57530 32246 57596
tri 32153 57514 32169 57530 ne
rect 32169 57514 32246 57530
rect 31986 57415 32134 57497
rect 31874 57382 31951 57398
tri 31951 57382 31967 57398 sw
rect 31874 57316 31967 57382
rect 31874 57214 31967 57280
rect 31874 57198 31951 57214
tri 31951 57198 31967 57214 nw
rect 32003 57181 32117 57415
tri 32153 57382 32169 57398 se
rect 32169 57382 32246 57398
rect 32153 57316 32246 57382
rect 32153 57214 32246 57280
tri 32153 57198 32169 57214 ne
rect 32169 57198 32246 57214
rect 31986 57099 32134 57181
rect 31874 57066 31951 57082
tri 31951 57066 31967 57082 sw
rect 31874 57000 31967 57066
rect 32003 56941 32117 57099
tri 32153 57066 32169 57082 se
rect 32169 57066 32246 57082
rect 32153 57000 32246 57066
rect 31874 56865 32246 56941
rect 31874 56740 31967 56806
rect 31874 56724 31951 56740
tri 31951 56724 31967 56740 nw
rect 32003 56707 32117 56865
rect 32153 56740 32246 56806
tri 32153 56724 32169 56740 ne
rect 32169 56724 32246 56740
rect 31986 56625 32134 56707
rect 31874 56592 31951 56608
tri 31951 56592 31967 56608 sw
rect 31874 56526 31967 56592
rect 31874 56424 31967 56490
rect 31874 56408 31951 56424
tri 31951 56408 31967 56424 nw
rect 32003 56391 32117 56625
tri 32153 56592 32169 56608 se
rect 32169 56592 32246 56608
rect 32153 56526 32246 56592
rect 32153 56424 32246 56490
tri 32153 56408 32169 56424 ne
rect 32169 56408 32246 56424
rect 31986 56309 32134 56391
rect 31874 56276 31951 56292
tri 31951 56276 31967 56292 sw
rect 31874 56210 31967 56276
rect 32003 56151 32117 56309
tri 32153 56276 32169 56292 se
rect 32169 56276 32246 56292
rect 32153 56210 32246 56276
rect 31874 56075 32246 56151
rect 31874 55950 31967 56016
rect 31874 55934 31951 55950
tri 31951 55934 31967 55950 nw
rect 32003 55917 32117 56075
rect 32153 55950 32246 56016
tri 32153 55934 32169 55950 ne
rect 32169 55934 32246 55950
rect 31986 55835 32134 55917
rect 31874 55802 31951 55818
tri 31951 55802 31967 55818 sw
rect 31874 55736 31967 55802
rect 31874 55634 31967 55700
rect 31874 55618 31951 55634
tri 31951 55618 31967 55634 nw
rect 32003 55601 32117 55835
tri 32153 55802 32169 55818 se
rect 32169 55802 32246 55818
rect 32153 55736 32246 55802
rect 32153 55634 32246 55700
tri 32153 55618 32169 55634 ne
rect 32169 55618 32246 55634
rect 31986 55519 32134 55601
rect 31874 55486 31951 55502
tri 31951 55486 31967 55502 sw
rect 31874 55420 31967 55486
rect 32003 55361 32117 55519
tri 32153 55486 32169 55502 se
rect 32169 55486 32246 55502
rect 32153 55420 32246 55486
rect 31874 55285 32246 55361
rect 31874 55160 31967 55226
rect 31874 55144 31951 55160
tri 31951 55144 31967 55160 nw
rect 32003 55127 32117 55285
rect 32153 55160 32246 55226
tri 32153 55144 32169 55160 ne
rect 32169 55144 32246 55160
rect 31986 55045 32134 55127
rect 31874 55012 31951 55028
tri 31951 55012 31967 55028 sw
rect 31874 54946 31967 55012
rect 31874 54844 31967 54910
rect 31874 54828 31951 54844
tri 31951 54828 31967 54844 nw
rect 32003 54811 32117 55045
tri 32153 55012 32169 55028 se
rect 32169 55012 32246 55028
rect 32153 54946 32246 55012
rect 32153 54844 32246 54910
tri 32153 54828 32169 54844 ne
rect 32169 54828 32246 54844
rect 31986 54729 32134 54811
rect 31874 54696 31951 54712
tri 31951 54696 31967 54712 sw
rect 31874 54630 31967 54696
rect 32003 54571 32117 54729
tri 32153 54696 32169 54712 se
rect 32169 54696 32246 54712
rect 32153 54630 32246 54696
rect 31874 54495 32246 54571
rect 31874 54370 31967 54436
rect 31874 54354 31951 54370
tri 31951 54354 31967 54370 nw
rect 32003 54337 32117 54495
rect 32153 54370 32246 54436
tri 32153 54354 32169 54370 ne
rect 32169 54354 32246 54370
rect 31986 54255 32134 54337
rect 31874 54222 31951 54238
tri 31951 54222 31967 54238 sw
rect 31874 54156 31967 54222
rect 31874 54054 31967 54120
rect 31874 54038 31951 54054
tri 31951 54038 31967 54054 nw
rect 32003 54021 32117 54255
tri 32153 54222 32169 54238 se
rect 32169 54222 32246 54238
rect 32153 54156 32246 54222
rect 32153 54054 32246 54120
tri 32153 54038 32169 54054 ne
rect 32169 54038 32246 54054
rect 31986 53939 32134 54021
rect 31874 53906 31951 53922
tri 31951 53906 31967 53922 sw
rect 31874 53840 31967 53906
rect 32003 53781 32117 53939
tri 32153 53906 32169 53922 se
rect 32169 53906 32246 53922
rect 32153 53840 32246 53906
rect 31874 53705 32246 53781
rect 31874 53580 31967 53646
rect 31874 53564 31951 53580
tri 31951 53564 31967 53580 nw
rect 32003 53547 32117 53705
rect 32153 53580 32246 53646
tri 32153 53564 32169 53580 ne
rect 32169 53564 32246 53580
rect 31986 53465 32134 53547
rect 31874 53432 31951 53448
tri 31951 53432 31967 53448 sw
rect 31874 53366 31967 53432
rect 31874 53264 31967 53330
rect 31874 53248 31951 53264
tri 31951 53248 31967 53264 nw
rect 32003 53231 32117 53465
tri 32153 53432 32169 53448 se
rect 32169 53432 32246 53448
rect 32153 53366 32246 53432
rect 32153 53264 32246 53330
tri 32153 53248 32169 53264 ne
rect 32169 53248 32246 53264
rect 31986 53149 32134 53231
rect 31874 53116 31951 53132
tri 31951 53116 31967 53132 sw
rect 31874 53050 31967 53116
rect 32003 52991 32117 53149
tri 32153 53116 32169 53132 se
rect 32169 53116 32246 53132
rect 32153 53050 32246 53116
rect 31874 52915 32246 52991
rect 31874 52790 31967 52856
rect 31874 52774 31951 52790
tri 31951 52774 31967 52790 nw
rect 32003 52757 32117 52915
rect 32153 52790 32246 52856
tri 32153 52774 32169 52790 ne
rect 32169 52774 32246 52790
rect 31986 52675 32134 52757
rect 31874 52642 31951 52658
tri 31951 52642 31967 52658 sw
rect 31874 52576 31967 52642
rect 31874 52474 31967 52540
rect 31874 52458 31951 52474
tri 31951 52458 31967 52474 nw
rect 32003 52441 32117 52675
tri 32153 52642 32169 52658 se
rect 32169 52642 32246 52658
rect 32153 52576 32246 52642
rect 32153 52474 32246 52540
tri 32153 52458 32169 52474 ne
rect 32169 52458 32246 52474
rect 31986 52359 32134 52441
rect 31874 52326 31951 52342
tri 31951 52326 31967 52342 sw
rect 31874 52260 31967 52326
rect 32003 52201 32117 52359
tri 32153 52326 32169 52342 se
rect 32169 52326 32246 52342
rect 32153 52260 32246 52326
rect 31874 52125 32246 52201
rect 31874 52000 31967 52066
rect 31874 51984 31951 52000
tri 31951 51984 31967 52000 nw
rect 32003 51967 32117 52125
rect 32153 52000 32246 52066
tri 32153 51984 32169 52000 ne
rect 32169 51984 32246 52000
rect 31986 51885 32134 51967
rect 31874 51852 31951 51868
tri 31951 51852 31967 51868 sw
rect 31874 51786 31967 51852
rect 31874 51684 31967 51750
rect 31874 51668 31951 51684
tri 31951 51668 31967 51684 nw
rect 32003 51651 32117 51885
tri 32153 51852 32169 51868 se
rect 32169 51852 32246 51868
rect 32153 51786 32246 51852
rect 32153 51684 32246 51750
tri 32153 51668 32169 51684 ne
rect 32169 51668 32246 51684
rect 31986 51569 32134 51651
rect 31874 51536 31951 51552
tri 31951 51536 31967 51552 sw
rect 31874 51470 31967 51536
rect 32003 51411 32117 51569
tri 32153 51536 32169 51552 se
rect 32169 51536 32246 51552
rect 32153 51470 32246 51536
rect 31874 51335 32246 51411
rect 31874 51210 31967 51276
rect 31874 51194 31951 51210
tri 31951 51194 31967 51210 nw
rect 32003 51177 32117 51335
rect 32153 51210 32246 51276
tri 32153 51194 32169 51210 ne
rect 32169 51194 32246 51210
rect 31986 51095 32134 51177
rect 31874 51062 31951 51078
tri 31951 51062 31967 51078 sw
rect 31874 50996 31967 51062
rect 31874 50894 31967 50960
rect 31874 50878 31951 50894
tri 31951 50878 31967 50894 nw
rect 32003 50861 32117 51095
tri 32153 51062 32169 51078 se
rect 32169 51062 32246 51078
rect 32153 50996 32246 51062
rect 32153 50894 32246 50960
tri 32153 50878 32169 50894 ne
rect 32169 50878 32246 50894
rect 31986 50779 32134 50861
rect 31874 50746 31951 50762
tri 31951 50746 31967 50762 sw
rect 31874 50680 31967 50746
rect 32003 50621 32117 50779
tri 32153 50746 32169 50762 se
rect 32169 50746 32246 50762
rect 32153 50680 32246 50746
rect 31874 50545 32246 50621
rect 31874 50420 31967 50486
rect 31874 50404 31951 50420
tri 31951 50404 31967 50420 nw
rect 32003 50387 32117 50545
rect 32153 50420 32246 50486
tri 32153 50404 32169 50420 ne
rect 32169 50404 32246 50420
rect 31986 50305 32134 50387
rect 31874 50272 31951 50288
tri 31951 50272 31967 50288 sw
rect 31874 50206 31967 50272
rect 31874 50104 31967 50170
rect 31874 50088 31951 50104
tri 31951 50088 31967 50104 nw
rect 32003 50071 32117 50305
tri 32153 50272 32169 50288 se
rect 32169 50272 32246 50288
rect 32153 50206 32246 50272
rect 32153 50104 32246 50170
tri 32153 50088 32169 50104 ne
rect 32169 50088 32246 50104
rect 31986 49989 32134 50071
rect 31874 49956 31951 49972
tri 31951 49956 31967 49972 sw
rect 31874 49890 31967 49956
rect 32003 49831 32117 49989
tri 32153 49956 32169 49972 se
rect 32169 49956 32246 49972
rect 32153 49890 32246 49956
rect 31874 49755 32246 49831
rect 31874 49630 31967 49696
rect 31874 49614 31951 49630
tri 31951 49614 31967 49630 nw
rect 32003 49597 32117 49755
rect 32153 49630 32246 49696
tri 32153 49614 32169 49630 ne
rect 32169 49614 32246 49630
rect 31986 49515 32134 49597
rect 31874 49482 31951 49498
tri 31951 49482 31967 49498 sw
rect 31874 49416 31967 49482
rect 31874 49314 31967 49380
rect 31874 49298 31951 49314
tri 31951 49298 31967 49314 nw
rect 32003 49281 32117 49515
tri 32153 49482 32169 49498 se
rect 32169 49482 32246 49498
rect 32153 49416 32246 49482
rect 32153 49314 32246 49380
tri 32153 49298 32169 49314 ne
rect 32169 49298 32246 49314
rect 31986 49199 32134 49281
rect 31874 49166 31951 49182
tri 31951 49166 31967 49182 sw
rect 31874 49100 31967 49166
rect 32003 49041 32117 49199
tri 32153 49166 32169 49182 se
rect 32169 49166 32246 49182
rect 32153 49100 32246 49166
rect 31874 48965 32246 49041
rect 31874 48840 31967 48906
rect 31874 48824 31951 48840
tri 31951 48824 31967 48840 nw
rect 32003 48807 32117 48965
rect 32153 48840 32246 48906
tri 32153 48824 32169 48840 ne
rect 32169 48824 32246 48840
rect 31986 48725 32134 48807
rect 31874 48692 31951 48708
tri 31951 48692 31967 48708 sw
rect 31874 48626 31967 48692
rect 31874 48524 31967 48590
rect 31874 48508 31951 48524
tri 31951 48508 31967 48524 nw
rect 32003 48491 32117 48725
tri 32153 48692 32169 48708 se
rect 32169 48692 32246 48708
rect 32153 48626 32246 48692
rect 32153 48524 32246 48590
tri 32153 48508 32169 48524 ne
rect 32169 48508 32246 48524
rect 31986 48409 32134 48491
rect 31874 48376 31951 48392
tri 31951 48376 31967 48392 sw
rect 31874 48310 31967 48376
rect 32003 48251 32117 48409
tri 32153 48376 32169 48392 se
rect 32169 48376 32246 48392
rect 32153 48310 32246 48376
rect 31874 48175 32246 48251
rect 31874 48050 31967 48116
rect 31874 48034 31951 48050
tri 31951 48034 31967 48050 nw
rect 32003 48017 32117 48175
rect 32153 48050 32246 48116
tri 32153 48034 32169 48050 ne
rect 32169 48034 32246 48050
rect 31986 47935 32134 48017
rect 31874 47902 31951 47918
tri 31951 47902 31967 47918 sw
rect 31874 47836 31967 47902
rect 31874 47734 31967 47800
rect 31874 47718 31951 47734
tri 31951 47718 31967 47734 nw
rect 32003 47701 32117 47935
tri 32153 47902 32169 47918 se
rect 32169 47902 32246 47918
rect 32153 47836 32246 47902
rect 32153 47734 32246 47800
tri 32153 47718 32169 47734 ne
rect 32169 47718 32246 47734
rect 31986 47619 32134 47701
rect 31874 47586 31951 47602
tri 31951 47586 31967 47602 sw
rect 31874 47520 31967 47586
rect 32003 47461 32117 47619
tri 32153 47586 32169 47602 se
rect 32169 47586 32246 47602
rect 32153 47520 32246 47586
rect 31874 47385 32246 47461
rect 31874 47260 31967 47326
rect 31874 47244 31951 47260
tri 31951 47244 31967 47260 nw
rect 32003 47227 32117 47385
rect 32153 47260 32246 47326
tri 32153 47244 32169 47260 ne
rect 32169 47244 32246 47260
rect 31986 47145 32134 47227
rect 31874 47112 31951 47128
tri 31951 47112 31967 47128 sw
rect 31874 47046 31967 47112
rect 31874 46944 31967 47010
rect 31874 46928 31951 46944
tri 31951 46928 31967 46944 nw
rect 32003 46911 32117 47145
tri 32153 47112 32169 47128 se
rect 32169 47112 32246 47128
rect 32153 47046 32246 47112
rect 32153 46944 32246 47010
tri 32153 46928 32169 46944 ne
rect 32169 46928 32246 46944
rect 31986 46829 32134 46911
rect 31874 46796 31951 46812
tri 31951 46796 31967 46812 sw
rect 31874 46730 31967 46796
rect 32003 46671 32117 46829
tri 32153 46796 32169 46812 se
rect 32169 46796 32246 46812
rect 32153 46730 32246 46796
rect 31874 46595 32246 46671
rect 31874 46470 31967 46536
rect 31874 46454 31951 46470
tri 31951 46454 31967 46470 nw
rect 32003 46437 32117 46595
rect 32153 46470 32246 46536
tri 32153 46454 32169 46470 ne
rect 32169 46454 32246 46470
rect 31986 46355 32134 46437
rect 31874 46322 31951 46338
tri 31951 46322 31967 46338 sw
rect 31874 46256 31967 46322
rect 31874 46154 31967 46220
rect 31874 46138 31951 46154
tri 31951 46138 31967 46154 nw
rect 32003 46121 32117 46355
tri 32153 46322 32169 46338 se
rect 32169 46322 32246 46338
rect 32153 46256 32246 46322
rect 32153 46154 32246 46220
tri 32153 46138 32169 46154 ne
rect 32169 46138 32246 46154
rect 31986 46039 32134 46121
rect 31874 46006 31951 46022
tri 31951 46006 31967 46022 sw
rect 31874 45940 31967 46006
rect 32003 45881 32117 46039
tri 32153 46006 32169 46022 se
rect 32169 46006 32246 46022
rect 32153 45940 32246 46006
rect 31874 45805 32246 45881
rect 31874 45680 31967 45746
rect 31874 45664 31951 45680
tri 31951 45664 31967 45680 nw
rect 32003 45647 32117 45805
rect 32153 45680 32246 45746
tri 32153 45664 32169 45680 ne
rect 32169 45664 32246 45680
rect 31986 45565 32134 45647
rect 31874 45532 31951 45548
tri 31951 45532 31967 45548 sw
rect 31874 45466 31967 45532
rect 31874 45364 31967 45430
rect 31874 45348 31951 45364
tri 31951 45348 31967 45364 nw
rect 32003 45331 32117 45565
tri 32153 45532 32169 45548 se
rect 32169 45532 32246 45548
rect 32153 45466 32246 45532
rect 32153 45364 32246 45430
tri 32153 45348 32169 45364 ne
rect 32169 45348 32246 45364
rect 31986 45249 32134 45331
rect 31874 45216 31951 45232
tri 31951 45216 31967 45232 sw
rect 31874 45150 31967 45216
rect 32003 45091 32117 45249
tri 32153 45216 32169 45232 se
rect 32169 45216 32246 45232
rect 32153 45150 32246 45216
rect 31874 45015 32246 45091
rect 31874 44890 31967 44956
rect 31874 44874 31951 44890
tri 31951 44874 31967 44890 nw
rect 32003 44857 32117 45015
rect 32153 44890 32246 44956
tri 32153 44874 32169 44890 ne
rect 32169 44874 32246 44890
rect 31986 44775 32134 44857
rect 31874 44742 31951 44758
tri 31951 44742 31967 44758 sw
rect 31874 44676 31967 44742
rect 31874 44574 31967 44640
rect 31874 44558 31951 44574
tri 31951 44558 31967 44574 nw
rect 32003 44541 32117 44775
tri 32153 44742 32169 44758 se
rect 32169 44742 32246 44758
rect 32153 44676 32246 44742
rect 32153 44574 32246 44640
tri 32153 44558 32169 44574 ne
rect 32169 44558 32246 44574
rect 31986 44459 32134 44541
rect 31874 44426 31951 44442
tri 31951 44426 31967 44442 sw
rect 31874 44360 31967 44426
rect 32003 44301 32117 44459
tri 32153 44426 32169 44442 se
rect 32169 44426 32246 44442
rect 32153 44360 32246 44426
rect 31874 44225 32246 44301
rect 31874 44100 31967 44166
rect 31874 44084 31951 44100
tri 31951 44084 31967 44100 nw
rect 32003 44067 32117 44225
rect 32153 44100 32246 44166
tri 32153 44084 32169 44100 ne
rect 32169 44084 32246 44100
rect 31986 43985 32134 44067
rect 31874 43952 31951 43968
tri 31951 43952 31967 43968 sw
rect 31874 43886 31967 43952
rect 31874 43784 31967 43850
rect 31874 43768 31951 43784
tri 31951 43768 31967 43784 nw
rect 32003 43751 32117 43985
tri 32153 43952 32169 43968 se
rect 32169 43952 32246 43968
rect 32153 43886 32246 43952
rect 32153 43784 32246 43850
tri 32153 43768 32169 43784 ne
rect 32169 43768 32246 43784
rect 31986 43669 32134 43751
rect 31874 43636 31951 43652
tri 31951 43636 31967 43652 sw
rect 31874 43570 31967 43636
rect 32003 43511 32117 43669
tri 32153 43636 32169 43652 se
rect 32169 43636 32246 43652
rect 32153 43570 32246 43636
rect 31874 43435 32246 43511
rect 31874 43310 31967 43376
rect 31874 43294 31951 43310
tri 31951 43294 31967 43310 nw
rect 32003 43277 32117 43435
rect 32153 43310 32246 43376
tri 32153 43294 32169 43310 ne
rect 32169 43294 32246 43310
rect 31986 43195 32134 43277
rect 31874 43162 31951 43178
tri 31951 43162 31967 43178 sw
rect 31874 43096 31967 43162
rect 31874 42994 31967 43060
rect 31874 42978 31951 42994
tri 31951 42978 31967 42994 nw
rect 32003 42961 32117 43195
tri 32153 43162 32169 43178 se
rect 32169 43162 32246 43178
rect 32153 43096 32246 43162
rect 32153 42994 32246 43060
tri 32153 42978 32169 42994 ne
rect 32169 42978 32246 42994
rect 31986 42879 32134 42961
rect 31874 42846 31951 42862
tri 31951 42846 31967 42862 sw
rect 31874 42780 31967 42846
rect 32003 42721 32117 42879
tri 32153 42846 32169 42862 se
rect 32169 42846 32246 42862
rect 32153 42780 32246 42846
rect 31874 42645 32246 42721
rect 31874 42520 31967 42586
rect 31874 42504 31951 42520
tri 31951 42504 31967 42520 nw
rect 32003 42487 32117 42645
rect 32153 42520 32246 42586
tri 32153 42504 32169 42520 ne
rect 32169 42504 32246 42520
rect 31986 42405 32134 42487
rect 31874 42372 31951 42388
tri 31951 42372 31967 42388 sw
rect 31874 42306 31967 42372
rect 31874 42204 31967 42270
rect 31874 42188 31951 42204
tri 31951 42188 31967 42204 nw
rect 32003 42171 32117 42405
tri 32153 42372 32169 42388 se
rect 32169 42372 32246 42388
rect 32153 42306 32246 42372
rect 32153 42204 32246 42270
tri 32153 42188 32169 42204 ne
rect 32169 42188 32246 42204
rect 31986 42089 32134 42171
rect 31874 42056 31951 42072
tri 31951 42056 31967 42072 sw
rect 31874 41990 31967 42056
rect 32003 41931 32117 42089
tri 32153 42056 32169 42072 se
rect 32169 42056 32246 42072
rect 32153 41990 32246 42056
rect 31874 41855 32246 41931
rect 31874 41730 31967 41796
rect 31874 41714 31951 41730
tri 31951 41714 31967 41730 nw
rect 32003 41697 32117 41855
rect 32153 41730 32246 41796
tri 32153 41714 32169 41730 ne
rect 32169 41714 32246 41730
rect 31986 41615 32134 41697
rect 31874 41582 31951 41598
tri 31951 41582 31967 41598 sw
rect 31874 41516 31967 41582
rect 31874 41414 31967 41480
rect 31874 41398 31951 41414
tri 31951 41398 31967 41414 nw
rect 32003 41381 32117 41615
tri 32153 41582 32169 41598 se
rect 32169 41582 32246 41598
rect 32153 41516 32246 41582
rect 32153 41414 32246 41480
tri 32153 41398 32169 41414 ne
rect 32169 41398 32246 41414
rect 31986 41299 32134 41381
rect 31874 41266 31951 41282
tri 31951 41266 31967 41282 sw
rect 31874 41200 31967 41266
rect 32003 41141 32117 41299
tri 32153 41266 32169 41282 se
rect 32169 41266 32246 41282
rect 32153 41200 32246 41266
rect 31874 41065 32246 41141
rect 31874 40940 31967 41006
rect 31874 40924 31951 40940
tri 31951 40924 31967 40940 nw
rect 32003 40907 32117 41065
rect 32153 40940 32246 41006
tri 32153 40924 32169 40940 ne
rect 32169 40924 32246 40940
rect 31986 40825 32134 40907
rect 31874 40792 31951 40808
tri 31951 40792 31967 40808 sw
rect 31874 40726 31967 40792
rect 31874 40624 31967 40690
rect 31874 40608 31951 40624
tri 31951 40608 31967 40624 nw
rect 32003 40591 32117 40825
tri 32153 40792 32169 40808 se
rect 32169 40792 32246 40808
rect 32153 40726 32246 40792
rect 32153 40624 32246 40690
tri 32153 40608 32169 40624 ne
rect 32169 40608 32246 40624
rect 31986 40509 32134 40591
rect 31874 40476 31951 40492
tri 31951 40476 31967 40492 sw
rect 31874 40410 31967 40476
rect 32003 40351 32117 40509
tri 32153 40476 32169 40492 se
rect 32169 40476 32246 40492
rect 32153 40410 32246 40476
rect 31874 40275 32246 40351
rect 31874 40150 31967 40216
rect 31874 40134 31951 40150
tri 31951 40134 31967 40150 nw
rect 32003 40117 32117 40275
rect 32153 40150 32246 40216
tri 32153 40134 32169 40150 ne
rect 32169 40134 32246 40150
rect 31986 40035 32134 40117
rect 31874 40002 31951 40018
tri 31951 40002 31967 40018 sw
rect 31874 39936 31967 40002
rect 31874 39834 31967 39900
rect 31874 39818 31951 39834
tri 31951 39818 31967 39834 nw
rect 32003 39801 32117 40035
tri 32153 40002 32169 40018 se
rect 32169 40002 32246 40018
rect 32153 39936 32246 40002
rect 32153 39834 32246 39900
tri 32153 39818 32169 39834 ne
rect 32169 39818 32246 39834
rect 31986 39719 32134 39801
rect 31874 39686 31951 39702
tri 31951 39686 31967 39702 sw
rect 31874 39620 31967 39686
rect 32003 39561 32117 39719
tri 32153 39686 32169 39702 se
rect 32169 39686 32246 39702
rect 32153 39620 32246 39686
rect 31874 39485 32246 39561
rect 31874 39360 31967 39426
rect 31874 39344 31951 39360
tri 31951 39344 31967 39360 nw
rect 32003 39327 32117 39485
rect 32153 39360 32246 39426
tri 32153 39344 32169 39360 ne
rect 32169 39344 32246 39360
rect 31986 39245 32134 39327
rect 31874 39212 31951 39228
tri 31951 39212 31967 39228 sw
rect 31874 39146 31967 39212
rect 31874 39044 31967 39110
rect 31874 39028 31951 39044
tri 31951 39028 31967 39044 nw
rect 32003 39011 32117 39245
tri 32153 39212 32169 39228 se
rect 32169 39212 32246 39228
rect 32153 39146 32246 39212
rect 32153 39044 32246 39110
tri 32153 39028 32169 39044 ne
rect 32169 39028 32246 39044
rect 31986 38929 32134 39011
rect 31874 38896 31951 38912
tri 31951 38896 31967 38912 sw
rect 31874 38830 31967 38896
rect 32003 38771 32117 38929
tri 32153 38896 32169 38912 se
rect 32169 38896 32246 38912
rect 32153 38830 32246 38896
rect 31874 38695 32246 38771
rect 31874 38570 31967 38636
rect 31874 38554 31951 38570
tri 31951 38554 31967 38570 nw
rect 32003 38537 32117 38695
rect 32153 38570 32246 38636
tri 32153 38554 32169 38570 ne
rect 32169 38554 32246 38570
rect 31986 38455 32134 38537
rect 31874 38422 31951 38438
tri 31951 38422 31967 38438 sw
rect 31874 38356 31967 38422
rect 31874 38254 31967 38320
rect 31874 38238 31951 38254
tri 31951 38238 31967 38254 nw
rect 32003 38221 32117 38455
tri 32153 38422 32169 38438 se
rect 32169 38422 32246 38438
rect 32153 38356 32246 38422
rect 32153 38254 32246 38320
tri 32153 38238 32169 38254 ne
rect 32169 38238 32246 38254
rect 31986 38139 32134 38221
rect 31874 38106 31951 38122
tri 31951 38106 31967 38122 sw
rect 31874 38040 31967 38106
rect 32003 37981 32117 38139
tri 32153 38106 32169 38122 se
rect 32169 38106 32246 38122
rect 32153 38040 32246 38106
rect 31874 37905 32246 37981
rect 31874 37780 31967 37846
rect 31874 37764 31951 37780
tri 31951 37764 31967 37780 nw
rect 32003 37747 32117 37905
rect 32153 37780 32246 37846
tri 32153 37764 32169 37780 ne
rect 32169 37764 32246 37780
rect 31986 37665 32134 37747
rect 31874 37632 31951 37648
tri 31951 37632 31967 37648 sw
rect 31874 37566 31967 37632
rect 31874 37464 31967 37530
rect 31874 37448 31951 37464
tri 31951 37448 31967 37464 nw
rect 32003 37431 32117 37665
tri 32153 37632 32169 37648 se
rect 32169 37632 32246 37648
rect 32153 37566 32246 37632
rect 32153 37464 32246 37530
tri 32153 37448 32169 37464 ne
rect 32169 37448 32246 37464
rect 31986 37349 32134 37431
rect 31874 37316 31951 37332
tri 31951 37316 31967 37332 sw
rect 31874 37250 31967 37316
rect 32003 37191 32117 37349
tri 32153 37316 32169 37332 se
rect 32169 37316 32246 37332
rect 32153 37250 32246 37316
rect 31874 37115 32246 37191
rect 31874 36990 31967 37056
rect 31874 36974 31951 36990
tri 31951 36974 31967 36990 nw
rect 32003 36957 32117 37115
rect 32153 36990 32246 37056
tri 32153 36974 32169 36990 ne
rect 32169 36974 32246 36990
rect 31986 36875 32134 36957
rect 31874 36842 31951 36858
tri 31951 36842 31967 36858 sw
rect 31874 36776 31967 36842
rect 31874 36674 31967 36740
rect 31874 36658 31951 36674
tri 31951 36658 31967 36674 nw
rect 32003 36641 32117 36875
tri 32153 36842 32169 36858 se
rect 32169 36842 32246 36858
rect 32153 36776 32246 36842
rect 32153 36674 32246 36740
tri 32153 36658 32169 36674 ne
rect 32169 36658 32246 36674
rect 31986 36559 32134 36641
rect 31874 36526 31951 36542
tri 31951 36526 31967 36542 sw
rect 31874 36460 31967 36526
rect 32003 36401 32117 36559
tri 32153 36526 32169 36542 se
rect 32169 36526 32246 36542
rect 32153 36460 32246 36526
rect 31874 36325 32246 36401
rect 31874 36200 31967 36266
rect 31874 36184 31951 36200
tri 31951 36184 31967 36200 nw
rect 32003 36167 32117 36325
rect 32153 36200 32246 36266
tri 32153 36184 32169 36200 ne
rect 32169 36184 32246 36200
rect 31986 36085 32134 36167
rect 31874 36052 31951 36068
tri 31951 36052 31967 36068 sw
rect 31874 35986 31967 36052
rect 31874 35884 31967 35950
rect 31874 35868 31951 35884
tri 31951 35868 31967 35884 nw
rect 32003 35851 32117 36085
tri 32153 36052 32169 36068 se
rect 32169 36052 32246 36068
rect 32153 35986 32246 36052
rect 32153 35884 32246 35950
tri 32153 35868 32169 35884 ne
rect 32169 35868 32246 35884
rect 31986 35769 32134 35851
rect 31874 35736 31951 35752
tri 31951 35736 31967 35752 sw
rect 31874 35670 31967 35736
rect 32003 35611 32117 35769
tri 32153 35736 32169 35752 se
rect 32169 35736 32246 35752
rect 32153 35670 32246 35736
rect 31874 35535 32246 35611
rect 31874 35410 31967 35476
rect 31874 35394 31951 35410
tri 31951 35394 31967 35410 nw
rect 32003 35377 32117 35535
rect 32153 35410 32246 35476
tri 32153 35394 32169 35410 ne
rect 32169 35394 32246 35410
rect 31986 35295 32134 35377
rect 31874 35262 31951 35278
tri 31951 35262 31967 35278 sw
rect 31874 35196 31967 35262
rect 31874 35094 31967 35160
rect 31874 35078 31951 35094
tri 31951 35078 31967 35094 nw
rect 32003 35061 32117 35295
tri 32153 35262 32169 35278 se
rect 32169 35262 32246 35278
rect 32153 35196 32246 35262
rect 32153 35094 32246 35160
tri 32153 35078 32169 35094 ne
rect 32169 35078 32246 35094
rect 31986 34979 32134 35061
rect 31874 34946 31951 34962
tri 31951 34946 31967 34962 sw
rect 31874 34880 31967 34946
rect 32003 34821 32117 34979
tri 32153 34946 32169 34962 se
rect 32169 34946 32246 34962
rect 32153 34880 32246 34946
rect 31874 34745 32246 34821
rect 31874 34620 31967 34686
rect 31874 34604 31951 34620
tri 31951 34604 31967 34620 nw
rect 32003 34587 32117 34745
rect 32153 34620 32246 34686
tri 32153 34604 32169 34620 ne
rect 32169 34604 32246 34620
rect 31986 34505 32134 34587
rect 31874 34472 31951 34488
tri 31951 34472 31967 34488 sw
rect 31874 34406 31967 34472
rect 31874 34304 31967 34370
rect 31874 34288 31951 34304
tri 31951 34288 31967 34304 nw
rect 32003 34271 32117 34505
tri 32153 34472 32169 34488 se
rect 32169 34472 32246 34488
rect 32153 34406 32246 34472
rect 32153 34304 32246 34370
tri 32153 34288 32169 34304 ne
rect 32169 34288 32246 34304
rect 31986 34189 32134 34271
rect 31874 34156 31951 34172
tri 31951 34156 31967 34172 sw
rect 31874 34090 31967 34156
rect 32003 34031 32117 34189
tri 32153 34156 32169 34172 se
rect 32169 34156 32246 34172
rect 32153 34090 32246 34156
rect 31874 33955 32246 34031
rect 31874 33830 31967 33896
rect 31874 33814 31951 33830
tri 31951 33814 31967 33830 nw
rect 32003 33797 32117 33955
rect 32153 33830 32246 33896
tri 32153 33814 32169 33830 ne
rect 32169 33814 32246 33830
rect 31986 33715 32134 33797
rect 31874 33682 31951 33698
tri 31951 33682 31967 33698 sw
rect 31874 33616 31967 33682
rect 31874 33514 31967 33580
rect 31874 33498 31951 33514
tri 31951 33498 31967 33514 nw
rect 32003 33481 32117 33715
tri 32153 33682 32169 33698 se
rect 32169 33682 32246 33698
rect 32153 33616 32246 33682
rect 32153 33514 32246 33580
tri 32153 33498 32169 33514 ne
rect 32169 33498 32246 33514
rect 31986 33399 32134 33481
rect 31874 33366 31951 33382
tri 31951 33366 31967 33382 sw
rect 31874 33300 31967 33366
rect 32003 33241 32117 33399
tri 32153 33366 32169 33382 se
rect 32169 33366 32246 33382
rect 32153 33300 32246 33366
rect 31874 33165 32246 33241
rect 31874 33040 31967 33106
rect 31874 33024 31951 33040
tri 31951 33024 31967 33040 nw
rect 32003 33007 32117 33165
rect 32153 33040 32246 33106
tri 32153 33024 32169 33040 ne
rect 32169 33024 32246 33040
rect 31986 32925 32134 33007
rect 31874 32892 31951 32908
tri 31951 32892 31967 32908 sw
rect 31874 32826 31967 32892
rect 31874 32724 31967 32790
rect 31874 32708 31951 32724
tri 31951 32708 31967 32724 nw
rect 32003 32691 32117 32925
tri 32153 32892 32169 32908 se
rect 32169 32892 32246 32908
rect 32153 32826 32246 32892
rect 32153 32724 32246 32790
tri 32153 32708 32169 32724 ne
rect 32169 32708 32246 32724
rect 31986 32609 32134 32691
rect 31874 32576 31951 32592
tri 31951 32576 31967 32592 sw
rect 31874 32510 31967 32576
rect 32003 32451 32117 32609
tri 32153 32576 32169 32592 se
rect 32169 32576 32246 32592
rect 32153 32510 32246 32576
rect 31874 32375 32246 32451
rect 31874 32250 31967 32316
rect 31874 32234 31951 32250
tri 31951 32234 31967 32250 nw
rect 32003 32217 32117 32375
rect 32153 32250 32246 32316
tri 32153 32234 32169 32250 ne
rect 32169 32234 32246 32250
rect 31986 32135 32134 32217
rect 31874 32102 31951 32118
tri 31951 32102 31967 32118 sw
rect 31874 32036 31967 32102
rect 31874 31934 31967 32000
rect 31874 31918 31951 31934
tri 31951 31918 31967 31934 nw
rect 32003 31901 32117 32135
tri 32153 32102 32169 32118 se
rect 32169 32102 32246 32118
rect 32153 32036 32246 32102
rect 32153 31934 32246 32000
tri 32153 31918 32169 31934 ne
rect 32169 31918 32246 31934
rect 31986 31819 32134 31901
rect 31874 31786 31951 31802
tri 31951 31786 31967 31802 sw
rect 31874 31720 31967 31786
rect 32003 31661 32117 31819
tri 32153 31786 32169 31802 se
rect 32169 31786 32246 31802
rect 32153 31720 32246 31786
rect 31874 31585 32246 31661
rect 31874 31460 31967 31526
rect 31874 31444 31951 31460
tri 31951 31444 31967 31460 nw
rect 32003 31427 32117 31585
rect 32153 31460 32246 31526
tri 32153 31444 32169 31460 ne
rect 32169 31444 32246 31460
rect 31986 31345 32134 31427
rect 31874 31312 31951 31328
tri 31951 31312 31967 31328 sw
rect 31874 31246 31967 31312
rect 31874 31144 31967 31210
rect 31874 31128 31951 31144
tri 31951 31128 31967 31144 nw
rect 32003 31111 32117 31345
tri 32153 31312 32169 31328 se
rect 32169 31312 32246 31328
rect 32153 31246 32246 31312
rect 32153 31144 32246 31210
tri 32153 31128 32169 31144 ne
rect 32169 31128 32246 31144
rect 31986 31029 32134 31111
rect 31874 30996 31951 31012
tri 31951 30996 31967 31012 sw
rect 31874 30930 31967 30996
rect 32003 30871 32117 31029
tri 32153 30996 32169 31012 se
rect 32169 30996 32246 31012
rect 32153 30930 32246 30996
rect 31874 30795 32246 30871
rect 31874 30670 31967 30736
rect 31874 30654 31951 30670
tri 31951 30654 31967 30670 nw
rect 32003 30637 32117 30795
rect 32153 30670 32246 30736
tri 32153 30654 32169 30670 ne
rect 32169 30654 32246 30670
rect 31986 30555 32134 30637
rect 31874 30522 31951 30538
tri 31951 30522 31967 30538 sw
rect 31874 30456 31967 30522
rect 31874 30354 31967 30420
rect 31874 30338 31951 30354
tri 31951 30338 31967 30354 nw
rect 32003 30321 32117 30555
tri 32153 30522 32169 30538 se
rect 32169 30522 32246 30538
rect 32153 30456 32246 30522
rect 32153 30354 32246 30420
tri 32153 30338 32169 30354 ne
rect 32169 30338 32246 30354
rect 31986 30239 32134 30321
rect 31874 30206 31951 30222
tri 31951 30206 31967 30222 sw
rect 31874 30140 31967 30206
rect 32003 30081 32117 30239
tri 32153 30206 32169 30222 se
rect 32169 30206 32246 30222
rect 32153 30140 32246 30206
rect 31874 30005 32246 30081
rect 31874 29880 31967 29946
rect 31874 29864 31951 29880
tri 31951 29864 31967 29880 nw
rect 32003 29847 32117 30005
rect 32153 29880 32246 29946
tri 32153 29864 32169 29880 ne
rect 32169 29864 32246 29880
rect 31986 29765 32134 29847
rect 31874 29732 31951 29748
tri 31951 29732 31967 29748 sw
rect 31874 29666 31967 29732
rect 31874 29564 31967 29630
rect 31874 29548 31951 29564
tri 31951 29548 31967 29564 nw
rect 32003 29531 32117 29765
tri 32153 29732 32169 29748 se
rect 32169 29732 32246 29748
rect 32153 29666 32246 29732
rect 32153 29564 32246 29630
tri 32153 29548 32169 29564 ne
rect 32169 29548 32246 29564
rect 31986 29449 32134 29531
rect 31874 29416 31951 29432
tri 31951 29416 31967 29432 sw
rect 31874 29350 31967 29416
rect 32003 29291 32117 29449
tri 32153 29416 32169 29432 se
rect 32169 29416 32246 29432
rect 32153 29350 32246 29416
rect 31874 29215 32246 29291
rect 31874 29090 31967 29156
rect 31874 29074 31951 29090
tri 31951 29074 31967 29090 nw
rect 32003 29057 32117 29215
rect 32153 29090 32246 29156
tri 32153 29074 32169 29090 ne
rect 32169 29074 32246 29090
rect 31986 28975 32134 29057
rect 31874 28942 31951 28958
tri 31951 28942 31967 28958 sw
rect 31874 28876 31967 28942
rect 32003 28833 32117 28975
tri 32153 28942 32169 28958 se
rect 32169 28942 32246 28958
rect 32153 28876 32246 28942
rect 32282 28463 32318 80603
rect 32354 28463 32390 80603
rect 32426 80445 32462 80603
rect 32418 80303 32470 80445
rect 32426 28763 32462 80303
rect 32418 28621 32470 28763
rect 32426 28463 32462 28621
rect 32498 28463 32534 80603
rect 32570 28463 32606 80603
rect 32642 28833 32726 80233
rect 32762 28463 32798 80603
rect 32834 28463 32870 80603
rect 32906 80445 32942 80603
rect 32898 80303 32950 80445
rect 32906 28763 32942 80303
rect 32898 28621 32950 28763
rect 32906 28463 32942 28621
rect 32978 28463 33014 80603
rect 33050 28463 33086 80603
rect 33122 80124 33215 80190
rect 33122 80108 33199 80124
tri 33199 80108 33215 80124 nw
rect 33251 80091 33365 80233
rect 33401 80124 33494 80190
tri 33401 80108 33417 80124 ne
rect 33417 80108 33494 80124
rect 33234 80009 33382 80091
rect 33122 79976 33199 79992
tri 33199 79976 33215 79992 sw
rect 33122 79910 33215 79976
rect 33251 79851 33365 80009
tri 33401 79976 33417 79992 se
rect 33417 79976 33494 79992
rect 33401 79910 33494 79976
rect 33122 79775 33494 79851
rect 33122 79650 33215 79716
rect 33122 79634 33199 79650
tri 33199 79634 33215 79650 nw
rect 33251 79617 33365 79775
rect 33401 79650 33494 79716
tri 33401 79634 33417 79650 ne
rect 33417 79634 33494 79650
rect 33234 79535 33382 79617
rect 33122 79502 33199 79518
tri 33199 79502 33215 79518 sw
rect 33122 79436 33215 79502
rect 33122 79334 33215 79400
rect 33122 79318 33199 79334
tri 33199 79318 33215 79334 nw
rect 33251 79301 33365 79535
tri 33401 79502 33417 79518 se
rect 33417 79502 33494 79518
rect 33401 79436 33494 79502
rect 33401 79334 33494 79400
tri 33401 79318 33417 79334 ne
rect 33417 79318 33494 79334
rect 33234 79219 33382 79301
rect 33122 79186 33199 79202
tri 33199 79186 33215 79202 sw
rect 33122 79120 33215 79186
rect 33251 79061 33365 79219
tri 33401 79186 33417 79202 se
rect 33417 79186 33494 79202
rect 33401 79120 33494 79186
rect 33122 78985 33494 79061
rect 33122 78860 33215 78926
rect 33122 78844 33199 78860
tri 33199 78844 33215 78860 nw
rect 33251 78827 33365 78985
rect 33401 78860 33494 78926
tri 33401 78844 33417 78860 ne
rect 33417 78844 33494 78860
rect 33234 78745 33382 78827
rect 33122 78712 33199 78728
tri 33199 78712 33215 78728 sw
rect 33122 78646 33215 78712
rect 33122 78544 33215 78610
rect 33122 78528 33199 78544
tri 33199 78528 33215 78544 nw
rect 33251 78511 33365 78745
tri 33401 78712 33417 78728 se
rect 33417 78712 33494 78728
rect 33401 78646 33494 78712
rect 33401 78544 33494 78610
tri 33401 78528 33417 78544 ne
rect 33417 78528 33494 78544
rect 33234 78429 33382 78511
rect 33122 78396 33199 78412
tri 33199 78396 33215 78412 sw
rect 33122 78330 33215 78396
rect 33251 78271 33365 78429
tri 33401 78396 33417 78412 se
rect 33417 78396 33494 78412
rect 33401 78330 33494 78396
rect 33122 78195 33494 78271
rect 33122 78070 33215 78136
rect 33122 78054 33199 78070
tri 33199 78054 33215 78070 nw
rect 33251 78037 33365 78195
rect 33401 78070 33494 78136
tri 33401 78054 33417 78070 ne
rect 33417 78054 33494 78070
rect 33234 77955 33382 78037
rect 33122 77922 33199 77938
tri 33199 77922 33215 77938 sw
rect 33122 77856 33215 77922
rect 33122 77754 33215 77820
rect 33122 77738 33199 77754
tri 33199 77738 33215 77754 nw
rect 33251 77721 33365 77955
tri 33401 77922 33417 77938 se
rect 33417 77922 33494 77938
rect 33401 77856 33494 77922
rect 33401 77754 33494 77820
tri 33401 77738 33417 77754 ne
rect 33417 77738 33494 77754
rect 33234 77639 33382 77721
rect 33122 77606 33199 77622
tri 33199 77606 33215 77622 sw
rect 33122 77540 33215 77606
rect 33251 77481 33365 77639
tri 33401 77606 33417 77622 se
rect 33417 77606 33494 77622
rect 33401 77540 33494 77606
rect 33122 77405 33494 77481
rect 33122 77280 33215 77346
rect 33122 77264 33199 77280
tri 33199 77264 33215 77280 nw
rect 33251 77247 33365 77405
rect 33401 77280 33494 77346
tri 33401 77264 33417 77280 ne
rect 33417 77264 33494 77280
rect 33234 77165 33382 77247
rect 33122 77132 33199 77148
tri 33199 77132 33215 77148 sw
rect 33122 77066 33215 77132
rect 33122 76964 33215 77030
rect 33122 76948 33199 76964
tri 33199 76948 33215 76964 nw
rect 33251 76931 33365 77165
tri 33401 77132 33417 77148 se
rect 33417 77132 33494 77148
rect 33401 77066 33494 77132
rect 33401 76964 33494 77030
tri 33401 76948 33417 76964 ne
rect 33417 76948 33494 76964
rect 33234 76849 33382 76931
rect 33122 76816 33199 76832
tri 33199 76816 33215 76832 sw
rect 33122 76750 33215 76816
rect 33251 76691 33365 76849
tri 33401 76816 33417 76832 se
rect 33417 76816 33494 76832
rect 33401 76750 33494 76816
rect 33122 76615 33494 76691
rect 33122 76490 33215 76556
rect 33122 76474 33199 76490
tri 33199 76474 33215 76490 nw
rect 33251 76457 33365 76615
rect 33401 76490 33494 76556
tri 33401 76474 33417 76490 ne
rect 33417 76474 33494 76490
rect 33234 76375 33382 76457
rect 33122 76342 33199 76358
tri 33199 76342 33215 76358 sw
rect 33122 76276 33215 76342
rect 33122 76174 33215 76240
rect 33122 76158 33199 76174
tri 33199 76158 33215 76174 nw
rect 33251 76141 33365 76375
tri 33401 76342 33417 76358 se
rect 33417 76342 33494 76358
rect 33401 76276 33494 76342
rect 33401 76174 33494 76240
tri 33401 76158 33417 76174 ne
rect 33417 76158 33494 76174
rect 33234 76059 33382 76141
rect 33122 76026 33199 76042
tri 33199 76026 33215 76042 sw
rect 33122 75960 33215 76026
rect 33251 75901 33365 76059
tri 33401 76026 33417 76042 se
rect 33417 76026 33494 76042
rect 33401 75960 33494 76026
rect 33122 75825 33494 75901
rect 33122 75700 33215 75766
rect 33122 75684 33199 75700
tri 33199 75684 33215 75700 nw
rect 33251 75667 33365 75825
rect 33401 75700 33494 75766
tri 33401 75684 33417 75700 ne
rect 33417 75684 33494 75700
rect 33234 75585 33382 75667
rect 33122 75552 33199 75568
tri 33199 75552 33215 75568 sw
rect 33122 75486 33215 75552
rect 33122 75384 33215 75450
rect 33122 75368 33199 75384
tri 33199 75368 33215 75384 nw
rect 33251 75351 33365 75585
tri 33401 75552 33417 75568 se
rect 33417 75552 33494 75568
rect 33401 75486 33494 75552
rect 33401 75384 33494 75450
tri 33401 75368 33417 75384 ne
rect 33417 75368 33494 75384
rect 33234 75269 33382 75351
rect 33122 75236 33199 75252
tri 33199 75236 33215 75252 sw
rect 33122 75170 33215 75236
rect 33251 75111 33365 75269
tri 33401 75236 33417 75252 se
rect 33417 75236 33494 75252
rect 33401 75170 33494 75236
rect 33122 75035 33494 75111
rect 33122 74910 33215 74976
rect 33122 74894 33199 74910
tri 33199 74894 33215 74910 nw
rect 33251 74877 33365 75035
rect 33401 74910 33494 74976
tri 33401 74894 33417 74910 ne
rect 33417 74894 33494 74910
rect 33234 74795 33382 74877
rect 33122 74762 33199 74778
tri 33199 74762 33215 74778 sw
rect 33122 74696 33215 74762
rect 33122 74594 33215 74660
rect 33122 74578 33199 74594
tri 33199 74578 33215 74594 nw
rect 33251 74561 33365 74795
tri 33401 74762 33417 74778 se
rect 33417 74762 33494 74778
rect 33401 74696 33494 74762
rect 33401 74594 33494 74660
tri 33401 74578 33417 74594 ne
rect 33417 74578 33494 74594
rect 33234 74479 33382 74561
rect 33122 74446 33199 74462
tri 33199 74446 33215 74462 sw
rect 33122 74380 33215 74446
rect 33251 74321 33365 74479
tri 33401 74446 33417 74462 se
rect 33417 74446 33494 74462
rect 33401 74380 33494 74446
rect 33122 74245 33494 74321
rect 33122 74120 33215 74186
rect 33122 74104 33199 74120
tri 33199 74104 33215 74120 nw
rect 33251 74087 33365 74245
rect 33401 74120 33494 74186
tri 33401 74104 33417 74120 ne
rect 33417 74104 33494 74120
rect 33234 74005 33382 74087
rect 33122 73972 33199 73988
tri 33199 73972 33215 73988 sw
rect 33122 73906 33215 73972
rect 33122 73804 33215 73870
rect 33122 73788 33199 73804
tri 33199 73788 33215 73804 nw
rect 33251 73771 33365 74005
tri 33401 73972 33417 73988 se
rect 33417 73972 33494 73988
rect 33401 73906 33494 73972
rect 33401 73804 33494 73870
tri 33401 73788 33417 73804 ne
rect 33417 73788 33494 73804
rect 33234 73689 33382 73771
rect 33122 73656 33199 73672
tri 33199 73656 33215 73672 sw
rect 33122 73590 33215 73656
rect 33251 73531 33365 73689
tri 33401 73656 33417 73672 se
rect 33417 73656 33494 73672
rect 33401 73590 33494 73656
rect 33122 73455 33494 73531
rect 33122 73330 33215 73396
rect 33122 73314 33199 73330
tri 33199 73314 33215 73330 nw
rect 33251 73297 33365 73455
rect 33401 73330 33494 73396
tri 33401 73314 33417 73330 ne
rect 33417 73314 33494 73330
rect 33234 73215 33382 73297
rect 33122 73182 33199 73198
tri 33199 73182 33215 73198 sw
rect 33122 73116 33215 73182
rect 33122 73014 33215 73080
rect 33122 72998 33199 73014
tri 33199 72998 33215 73014 nw
rect 33251 72981 33365 73215
tri 33401 73182 33417 73198 se
rect 33417 73182 33494 73198
rect 33401 73116 33494 73182
rect 33401 73014 33494 73080
tri 33401 72998 33417 73014 ne
rect 33417 72998 33494 73014
rect 33234 72899 33382 72981
rect 33122 72866 33199 72882
tri 33199 72866 33215 72882 sw
rect 33122 72800 33215 72866
rect 33251 72741 33365 72899
tri 33401 72866 33417 72882 se
rect 33417 72866 33494 72882
rect 33401 72800 33494 72866
rect 33122 72665 33494 72741
rect 33122 72540 33215 72606
rect 33122 72524 33199 72540
tri 33199 72524 33215 72540 nw
rect 33251 72507 33365 72665
rect 33401 72540 33494 72606
tri 33401 72524 33417 72540 ne
rect 33417 72524 33494 72540
rect 33234 72425 33382 72507
rect 33122 72392 33199 72408
tri 33199 72392 33215 72408 sw
rect 33122 72326 33215 72392
rect 33122 72224 33215 72290
rect 33122 72208 33199 72224
tri 33199 72208 33215 72224 nw
rect 33251 72191 33365 72425
tri 33401 72392 33417 72408 se
rect 33417 72392 33494 72408
rect 33401 72326 33494 72392
rect 33401 72224 33494 72290
tri 33401 72208 33417 72224 ne
rect 33417 72208 33494 72224
rect 33234 72109 33382 72191
rect 33122 72076 33199 72092
tri 33199 72076 33215 72092 sw
rect 33122 72010 33215 72076
rect 33251 71951 33365 72109
tri 33401 72076 33417 72092 se
rect 33417 72076 33494 72092
rect 33401 72010 33494 72076
rect 33122 71875 33494 71951
rect 33122 71750 33215 71816
rect 33122 71734 33199 71750
tri 33199 71734 33215 71750 nw
rect 33251 71717 33365 71875
rect 33401 71750 33494 71816
tri 33401 71734 33417 71750 ne
rect 33417 71734 33494 71750
rect 33234 71635 33382 71717
rect 33122 71602 33199 71618
tri 33199 71602 33215 71618 sw
rect 33122 71536 33215 71602
rect 33122 71434 33215 71500
rect 33122 71418 33199 71434
tri 33199 71418 33215 71434 nw
rect 33251 71401 33365 71635
tri 33401 71602 33417 71618 se
rect 33417 71602 33494 71618
rect 33401 71536 33494 71602
rect 33401 71434 33494 71500
tri 33401 71418 33417 71434 ne
rect 33417 71418 33494 71434
rect 33234 71319 33382 71401
rect 33122 71286 33199 71302
tri 33199 71286 33215 71302 sw
rect 33122 71220 33215 71286
rect 33251 71161 33365 71319
tri 33401 71286 33417 71302 se
rect 33417 71286 33494 71302
rect 33401 71220 33494 71286
rect 33122 71085 33494 71161
rect 33122 70960 33215 71026
rect 33122 70944 33199 70960
tri 33199 70944 33215 70960 nw
rect 33251 70927 33365 71085
rect 33401 70960 33494 71026
tri 33401 70944 33417 70960 ne
rect 33417 70944 33494 70960
rect 33234 70845 33382 70927
rect 33122 70812 33199 70828
tri 33199 70812 33215 70828 sw
rect 33122 70746 33215 70812
rect 33122 70644 33215 70710
rect 33122 70628 33199 70644
tri 33199 70628 33215 70644 nw
rect 33251 70611 33365 70845
tri 33401 70812 33417 70828 se
rect 33417 70812 33494 70828
rect 33401 70746 33494 70812
rect 33401 70644 33494 70710
tri 33401 70628 33417 70644 ne
rect 33417 70628 33494 70644
rect 33234 70529 33382 70611
rect 33122 70496 33199 70512
tri 33199 70496 33215 70512 sw
rect 33122 70430 33215 70496
rect 33251 70371 33365 70529
tri 33401 70496 33417 70512 se
rect 33417 70496 33494 70512
rect 33401 70430 33494 70496
rect 33122 70295 33494 70371
rect 33122 70170 33215 70236
rect 33122 70154 33199 70170
tri 33199 70154 33215 70170 nw
rect 33251 70137 33365 70295
rect 33401 70170 33494 70236
tri 33401 70154 33417 70170 ne
rect 33417 70154 33494 70170
rect 33234 70055 33382 70137
rect 33122 70022 33199 70038
tri 33199 70022 33215 70038 sw
rect 33122 69956 33215 70022
rect 33122 69854 33215 69920
rect 33122 69838 33199 69854
tri 33199 69838 33215 69854 nw
rect 33251 69821 33365 70055
tri 33401 70022 33417 70038 se
rect 33417 70022 33494 70038
rect 33401 69956 33494 70022
rect 33401 69854 33494 69920
tri 33401 69838 33417 69854 ne
rect 33417 69838 33494 69854
rect 33234 69739 33382 69821
rect 33122 69706 33199 69722
tri 33199 69706 33215 69722 sw
rect 33122 69640 33215 69706
rect 33251 69581 33365 69739
tri 33401 69706 33417 69722 se
rect 33417 69706 33494 69722
rect 33401 69640 33494 69706
rect 33122 69505 33494 69581
rect 33122 69380 33215 69446
rect 33122 69364 33199 69380
tri 33199 69364 33215 69380 nw
rect 33251 69347 33365 69505
rect 33401 69380 33494 69446
tri 33401 69364 33417 69380 ne
rect 33417 69364 33494 69380
rect 33234 69265 33382 69347
rect 33122 69232 33199 69248
tri 33199 69232 33215 69248 sw
rect 33122 69166 33215 69232
rect 33122 69064 33215 69130
rect 33122 69048 33199 69064
tri 33199 69048 33215 69064 nw
rect 33251 69031 33365 69265
tri 33401 69232 33417 69248 se
rect 33417 69232 33494 69248
rect 33401 69166 33494 69232
rect 33401 69064 33494 69130
tri 33401 69048 33417 69064 ne
rect 33417 69048 33494 69064
rect 33234 68949 33382 69031
rect 33122 68916 33199 68932
tri 33199 68916 33215 68932 sw
rect 33122 68850 33215 68916
rect 33251 68791 33365 68949
tri 33401 68916 33417 68932 se
rect 33417 68916 33494 68932
rect 33401 68850 33494 68916
rect 33122 68715 33494 68791
rect 33122 68590 33215 68656
rect 33122 68574 33199 68590
tri 33199 68574 33215 68590 nw
rect 33251 68557 33365 68715
rect 33401 68590 33494 68656
tri 33401 68574 33417 68590 ne
rect 33417 68574 33494 68590
rect 33234 68475 33382 68557
rect 33122 68442 33199 68458
tri 33199 68442 33215 68458 sw
rect 33122 68376 33215 68442
rect 33122 68274 33215 68340
rect 33122 68258 33199 68274
tri 33199 68258 33215 68274 nw
rect 33251 68241 33365 68475
tri 33401 68442 33417 68458 se
rect 33417 68442 33494 68458
rect 33401 68376 33494 68442
rect 33401 68274 33494 68340
tri 33401 68258 33417 68274 ne
rect 33417 68258 33494 68274
rect 33234 68159 33382 68241
rect 33122 68126 33199 68142
tri 33199 68126 33215 68142 sw
rect 33122 68060 33215 68126
rect 33251 68001 33365 68159
tri 33401 68126 33417 68142 se
rect 33417 68126 33494 68142
rect 33401 68060 33494 68126
rect 33122 67925 33494 68001
rect 33122 67800 33215 67866
rect 33122 67784 33199 67800
tri 33199 67784 33215 67800 nw
rect 33251 67767 33365 67925
rect 33401 67800 33494 67866
tri 33401 67784 33417 67800 ne
rect 33417 67784 33494 67800
rect 33234 67685 33382 67767
rect 33122 67652 33199 67668
tri 33199 67652 33215 67668 sw
rect 33122 67586 33215 67652
rect 33122 67484 33215 67550
rect 33122 67468 33199 67484
tri 33199 67468 33215 67484 nw
rect 33251 67451 33365 67685
tri 33401 67652 33417 67668 se
rect 33417 67652 33494 67668
rect 33401 67586 33494 67652
rect 33401 67484 33494 67550
tri 33401 67468 33417 67484 ne
rect 33417 67468 33494 67484
rect 33234 67369 33382 67451
rect 33122 67336 33199 67352
tri 33199 67336 33215 67352 sw
rect 33122 67270 33215 67336
rect 33251 67211 33365 67369
tri 33401 67336 33417 67352 se
rect 33417 67336 33494 67352
rect 33401 67270 33494 67336
rect 33122 67135 33494 67211
rect 33122 67010 33215 67076
rect 33122 66994 33199 67010
tri 33199 66994 33215 67010 nw
rect 33251 66977 33365 67135
rect 33401 67010 33494 67076
tri 33401 66994 33417 67010 ne
rect 33417 66994 33494 67010
rect 33234 66895 33382 66977
rect 33122 66862 33199 66878
tri 33199 66862 33215 66878 sw
rect 33122 66796 33215 66862
rect 33122 66694 33215 66760
rect 33122 66678 33199 66694
tri 33199 66678 33215 66694 nw
rect 33251 66661 33365 66895
tri 33401 66862 33417 66878 se
rect 33417 66862 33494 66878
rect 33401 66796 33494 66862
rect 33401 66694 33494 66760
tri 33401 66678 33417 66694 ne
rect 33417 66678 33494 66694
rect 33234 66579 33382 66661
rect 33122 66546 33199 66562
tri 33199 66546 33215 66562 sw
rect 33122 66480 33215 66546
rect 33251 66421 33365 66579
tri 33401 66546 33417 66562 se
rect 33417 66546 33494 66562
rect 33401 66480 33494 66546
rect 33122 66345 33494 66421
rect 33122 66220 33215 66286
rect 33122 66204 33199 66220
tri 33199 66204 33215 66220 nw
rect 33251 66187 33365 66345
rect 33401 66220 33494 66286
tri 33401 66204 33417 66220 ne
rect 33417 66204 33494 66220
rect 33234 66105 33382 66187
rect 33122 66072 33199 66088
tri 33199 66072 33215 66088 sw
rect 33122 66006 33215 66072
rect 33122 65904 33215 65970
rect 33122 65888 33199 65904
tri 33199 65888 33215 65904 nw
rect 33251 65871 33365 66105
tri 33401 66072 33417 66088 se
rect 33417 66072 33494 66088
rect 33401 66006 33494 66072
rect 33401 65904 33494 65970
tri 33401 65888 33417 65904 ne
rect 33417 65888 33494 65904
rect 33234 65789 33382 65871
rect 33122 65756 33199 65772
tri 33199 65756 33215 65772 sw
rect 33122 65690 33215 65756
rect 33251 65631 33365 65789
tri 33401 65756 33417 65772 se
rect 33417 65756 33494 65772
rect 33401 65690 33494 65756
rect 33122 65555 33494 65631
rect 33122 65430 33215 65496
rect 33122 65414 33199 65430
tri 33199 65414 33215 65430 nw
rect 33251 65397 33365 65555
rect 33401 65430 33494 65496
tri 33401 65414 33417 65430 ne
rect 33417 65414 33494 65430
rect 33234 65315 33382 65397
rect 33122 65282 33199 65298
tri 33199 65282 33215 65298 sw
rect 33122 65216 33215 65282
rect 33122 65114 33215 65180
rect 33122 65098 33199 65114
tri 33199 65098 33215 65114 nw
rect 33251 65081 33365 65315
tri 33401 65282 33417 65298 se
rect 33417 65282 33494 65298
rect 33401 65216 33494 65282
rect 33401 65114 33494 65180
tri 33401 65098 33417 65114 ne
rect 33417 65098 33494 65114
rect 33234 64999 33382 65081
rect 33122 64966 33199 64982
tri 33199 64966 33215 64982 sw
rect 33122 64900 33215 64966
rect 33251 64841 33365 64999
tri 33401 64966 33417 64982 se
rect 33417 64966 33494 64982
rect 33401 64900 33494 64966
rect 33122 64765 33494 64841
rect 33122 64640 33215 64706
rect 33122 64624 33199 64640
tri 33199 64624 33215 64640 nw
rect 33251 64607 33365 64765
rect 33401 64640 33494 64706
tri 33401 64624 33417 64640 ne
rect 33417 64624 33494 64640
rect 33234 64525 33382 64607
rect 33122 64492 33199 64508
tri 33199 64492 33215 64508 sw
rect 33122 64426 33215 64492
rect 33122 64324 33215 64390
rect 33122 64308 33199 64324
tri 33199 64308 33215 64324 nw
rect 33251 64291 33365 64525
tri 33401 64492 33417 64508 se
rect 33417 64492 33494 64508
rect 33401 64426 33494 64492
rect 33401 64324 33494 64390
tri 33401 64308 33417 64324 ne
rect 33417 64308 33494 64324
rect 33234 64209 33382 64291
rect 33122 64176 33199 64192
tri 33199 64176 33215 64192 sw
rect 33122 64110 33215 64176
rect 33251 64051 33365 64209
tri 33401 64176 33417 64192 se
rect 33417 64176 33494 64192
rect 33401 64110 33494 64176
rect 33122 63975 33494 64051
rect 33122 63850 33215 63916
rect 33122 63834 33199 63850
tri 33199 63834 33215 63850 nw
rect 33251 63817 33365 63975
rect 33401 63850 33494 63916
tri 33401 63834 33417 63850 ne
rect 33417 63834 33494 63850
rect 33234 63735 33382 63817
rect 33122 63702 33199 63718
tri 33199 63702 33215 63718 sw
rect 33122 63636 33215 63702
rect 33122 63534 33215 63600
rect 33122 63518 33199 63534
tri 33199 63518 33215 63534 nw
rect 33251 63501 33365 63735
tri 33401 63702 33417 63718 se
rect 33417 63702 33494 63718
rect 33401 63636 33494 63702
rect 33401 63534 33494 63600
tri 33401 63518 33417 63534 ne
rect 33417 63518 33494 63534
rect 33234 63419 33382 63501
rect 33122 63386 33199 63402
tri 33199 63386 33215 63402 sw
rect 33122 63320 33215 63386
rect 33251 63261 33365 63419
tri 33401 63386 33417 63402 se
rect 33417 63386 33494 63402
rect 33401 63320 33494 63386
rect 33122 63185 33494 63261
rect 33122 63060 33215 63126
rect 33122 63044 33199 63060
tri 33199 63044 33215 63060 nw
rect 33251 63027 33365 63185
rect 33401 63060 33494 63126
tri 33401 63044 33417 63060 ne
rect 33417 63044 33494 63060
rect 33234 62945 33382 63027
rect 33122 62912 33199 62928
tri 33199 62912 33215 62928 sw
rect 33122 62846 33215 62912
rect 33122 62744 33215 62810
rect 33122 62728 33199 62744
tri 33199 62728 33215 62744 nw
rect 33251 62711 33365 62945
tri 33401 62912 33417 62928 se
rect 33417 62912 33494 62928
rect 33401 62846 33494 62912
rect 33401 62744 33494 62810
tri 33401 62728 33417 62744 ne
rect 33417 62728 33494 62744
rect 33234 62629 33382 62711
rect 33122 62596 33199 62612
tri 33199 62596 33215 62612 sw
rect 33122 62530 33215 62596
rect 33251 62471 33365 62629
tri 33401 62596 33417 62612 se
rect 33417 62596 33494 62612
rect 33401 62530 33494 62596
rect 33122 62395 33494 62471
rect 33122 62270 33215 62336
rect 33122 62254 33199 62270
tri 33199 62254 33215 62270 nw
rect 33251 62237 33365 62395
rect 33401 62270 33494 62336
tri 33401 62254 33417 62270 ne
rect 33417 62254 33494 62270
rect 33234 62155 33382 62237
rect 33122 62122 33199 62138
tri 33199 62122 33215 62138 sw
rect 33122 62056 33215 62122
rect 33122 61954 33215 62020
rect 33122 61938 33199 61954
tri 33199 61938 33215 61954 nw
rect 33251 61921 33365 62155
tri 33401 62122 33417 62138 se
rect 33417 62122 33494 62138
rect 33401 62056 33494 62122
rect 33401 61954 33494 62020
tri 33401 61938 33417 61954 ne
rect 33417 61938 33494 61954
rect 33234 61839 33382 61921
rect 33122 61806 33199 61822
tri 33199 61806 33215 61822 sw
rect 33122 61740 33215 61806
rect 33251 61681 33365 61839
tri 33401 61806 33417 61822 se
rect 33417 61806 33494 61822
rect 33401 61740 33494 61806
rect 33122 61605 33494 61681
rect 33122 61480 33215 61546
rect 33122 61464 33199 61480
tri 33199 61464 33215 61480 nw
rect 33251 61447 33365 61605
rect 33401 61480 33494 61546
tri 33401 61464 33417 61480 ne
rect 33417 61464 33494 61480
rect 33234 61365 33382 61447
rect 33122 61332 33199 61348
tri 33199 61332 33215 61348 sw
rect 33122 61266 33215 61332
rect 33122 61164 33215 61230
rect 33122 61148 33199 61164
tri 33199 61148 33215 61164 nw
rect 33251 61131 33365 61365
tri 33401 61332 33417 61348 se
rect 33417 61332 33494 61348
rect 33401 61266 33494 61332
rect 33401 61164 33494 61230
tri 33401 61148 33417 61164 ne
rect 33417 61148 33494 61164
rect 33234 61049 33382 61131
rect 33122 61016 33199 61032
tri 33199 61016 33215 61032 sw
rect 33122 60950 33215 61016
rect 33251 60891 33365 61049
tri 33401 61016 33417 61032 se
rect 33417 61016 33494 61032
rect 33401 60950 33494 61016
rect 33122 60815 33494 60891
rect 33122 60690 33215 60756
rect 33122 60674 33199 60690
tri 33199 60674 33215 60690 nw
rect 33251 60657 33365 60815
rect 33401 60690 33494 60756
tri 33401 60674 33417 60690 ne
rect 33417 60674 33494 60690
rect 33234 60575 33382 60657
rect 33122 60542 33199 60558
tri 33199 60542 33215 60558 sw
rect 33122 60476 33215 60542
rect 33122 60374 33215 60440
rect 33122 60358 33199 60374
tri 33199 60358 33215 60374 nw
rect 33251 60341 33365 60575
tri 33401 60542 33417 60558 se
rect 33417 60542 33494 60558
rect 33401 60476 33494 60542
rect 33401 60374 33494 60440
tri 33401 60358 33417 60374 ne
rect 33417 60358 33494 60374
rect 33234 60259 33382 60341
rect 33122 60226 33199 60242
tri 33199 60226 33215 60242 sw
rect 33122 60160 33215 60226
rect 33251 60101 33365 60259
tri 33401 60226 33417 60242 se
rect 33417 60226 33494 60242
rect 33401 60160 33494 60226
rect 33122 60025 33494 60101
rect 33122 59900 33215 59966
rect 33122 59884 33199 59900
tri 33199 59884 33215 59900 nw
rect 33251 59867 33365 60025
rect 33401 59900 33494 59966
tri 33401 59884 33417 59900 ne
rect 33417 59884 33494 59900
rect 33234 59785 33382 59867
rect 33122 59752 33199 59768
tri 33199 59752 33215 59768 sw
rect 33122 59686 33215 59752
rect 33122 59584 33215 59650
rect 33122 59568 33199 59584
tri 33199 59568 33215 59584 nw
rect 33251 59551 33365 59785
tri 33401 59752 33417 59768 se
rect 33417 59752 33494 59768
rect 33401 59686 33494 59752
rect 33401 59584 33494 59650
tri 33401 59568 33417 59584 ne
rect 33417 59568 33494 59584
rect 33234 59469 33382 59551
rect 33122 59436 33199 59452
tri 33199 59436 33215 59452 sw
rect 33122 59370 33215 59436
rect 33251 59311 33365 59469
tri 33401 59436 33417 59452 se
rect 33417 59436 33494 59452
rect 33401 59370 33494 59436
rect 33122 59235 33494 59311
rect 33122 59110 33215 59176
rect 33122 59094 33199 59110
tri 33199 59094 33215 59110 nw
rect 33251 59077 33365 59235
rect 33401 59110 33494 59176
tri 33401 59094 33417 59110 ne
rect 33417 59094 33494 59110
rect 33234 58995 33382 59077
rect 33122 58962 33199 58978
tri 33199 58962 33215 58978 sw
rect 33122 58896 33215 58962
rect 33122 58794 33215 58860
rect 33122 58778 33199 58794
tri 33199 58778 33215 58794 nw
rect 33251 58761 33365 58995
tri 33401 58962 33417 58978 se
rect 33417 58962 33494 58978
rect 33401 58896 33494 58962
rect 33401 58794 33494 58860
tri 33401 58778 33417 58794 ne
rect 33417 58778 33494 58794
rect 33234 58679 33382 58761
rect 33122 58646 33199 58662
tri 33199 58646 33215 58662 sw
rect 33122 58580 33215 58646
rect 33251 58521 33365 58679
tri 33401 58646 33417 58662 se
rect 33417 58646 33494 58662
rect 33401 58580 33494 58646
rect 33122 58445 33494 58521
rect 33122 58320 33215 58386
rect 33122 58304 33199 58320
tri 33199 58304 33215 58320 nw
rect 33251 58287 33365 58445
rect 33401 58320 33494 58386
tri 33401 58304 33417 58320 ne
rect 33417 58304 33494 58320
rect 33234 58205 33382 58287
rect 33122 58172 33199 58188
tri 33199 58172 33215 58188 sw
rect 33122 58106 33215 58172
rect 33122 58004 33215 58070
rect 33122 57988 33199 58004
tri 33199 57988 33215 58004 nw
rect 33251 57971 33365 58205
tri 33401 58172 33417 58188 se
rect 33417 58172 33494 58188
rect 33401 58106 33494 58172
rect 33401 58004 33494 58070
tri 33401 57988 33417 58004 ne
rect 33417 57988 33494 58004
rect 33234 57889 33382 57971
rect 33122 57856 33199 57872
tri 33199 57856 33215 57872 sw
rect 33122 57790 33215 57856
rect 33251 57731 33365 57889
tri 33401 57856 33417 57872 se
rect 33417 57856 33494 57872
rect 33401 57790 33494 57856
rect 33122 57655 33494 57731
rect 33122 57530 33215 57596
rect 33122 57514 33199 57530
tri 33199 57514 33215 57530 nw
rect 33251 57497 33365 57655
rect 33401 57530 33494 57596
tri 33401 57514 33417 57530 ne
rect 33417 57514 33494 57530
rect 33234 57415 33382 57497
rect 33122 57382 33199 57398
tri 33199 57382 33215 57398 sw
rect 33122 57316 33215 57382
rect 33122 57214 33215 57280
rect 33122 57198 33199 57214
tri 33199 57198 33215 57214 nw
rect 33251 57181 33365 57415
tri 33401 57382 33417 57398 se
rect 33417 57382 33494 57398
rect 33401 57316 33494 57382
rect 33401 57214 33494 57280
tri 33401 57198 33417 57214 ne
rect 33417 57198 33494 57214
rect 33234 57099 33382 57181
rect 33122 57066 33199 57082
tri 33199 57066 33215 57082 sw
rect 33122 57000 33215 57066
rect 33251 56941 33365 57099
tri 33401 57066 33417 57082 se
rect 33417 57066 33494 57082
rect 33401 57000 33494 57066
rect 33122 56865 33494 56941
rect 33122 56740 33215 56806
rect 33122 56724 33199 56740
tri 33199 56724 33215 56740 nw
rect 33251 56707 33365 56865
rect 33401 56740 33494 56806
tri 33401 56724 33417 56740 ne
rect 33417 56724 33494 56740
rect 33234 56625 33382 56707
rect 33122 56592 33199 56608
tri 33199 56592 33215 56608 sw
rect 33122 56526 33215 56592
rect 33122 56424 33215 56490
rect 33122 56408 33199 56424
tri 33199 56408 33215 56424 nw
rect 33251 56391 33365 56625
tri 33401 56592 33417 56608 se
rect 33417 56592 33494 56608
rect 33401 56526 33494 56592
rect 33401 56424 33494 56490
tri 33401 56408 33417 56424 ne
rect 33417 56408 33494 56424
rect 33234 56309 33382 56391
rect 33122 56276 33199 56292
tri 33199 56276 33215 56292 sw
rect 33122 56210 33215 56276
rect 33251 56151 33365 56309
tri 33401 56276 33417 56292 se
rect 33417 56276 33494 56292
rect 33401 56210 33494 56276
rect 33122 56075 33494 56151
rect 33122 55950 33215 56016
rect 33122 55934 33199 55950
tri 33199 55934 33215 55950 nw
rect 33251 55917 33365 56075
rect 33401 55950 33494 56016
tri 33401 55934 33417 55950 ne
rect 33417 55934 33494 55950
rect 33234 55835 33382 55917
rect 33122 55802 33199 55818
tri 33199 55802 33215 55818 sw
rect 33122 55736 33215 55802
rect 33122 55634 33215 55700
rect 33122 55618 33199 55634
tri 33199 55618 33215 55634 nw
rect 33251 55601 33365 55835
tri 33401 55802 33417 55818 se
rect 33417 55802 33494 55818
rect 33401 55736 33494 55802
rect 33401 55634 33494 55700
tri 33401 55618 33417 55634 ne
rect 33417 55618 33494 55634
rect 33234 55519 33382 55601
rect 33122 55486 33199 55502
tri 33199 55486 33215 55502 sw
rect 33122 55420 33215 55486
rect 33251 55361 33365 55519
tri 33401 55486 33417 55502 se
rect 33417 55486 33494 55502
rect 33401 55420 33494 55486
rect 33122 55285 33494 55361
rect 33122 55160 33215 55226
rect 33122 55144 33199 55160
tri 33199 55144 33215 55160 nw
rect 33251 55127 33365 55285
rect 33401 55160 33494 55226
tri 33401 55144 33417 55160 ne
rect 33417 55144 33494 55160
rect 33234 55045 33382 55127
rect 33122 55012 33199 55028
tri 33199 55012 33215 55028 sw
rect 33122 54946 33215 55012
rect 33122 54844 33215 54910
rect 33122 54828 33199 54844
tri 33199 54828 33215 54844 nw
rect 33251 54811 33365 55045
tri 33401 55012 33417 55028 se
rect 33417 55012 33494 55028
rect 33401 54946 33494 55012
rect 33401 54844 33494 54910
tri 33401 54828 33417 54844 ne
rect 33417 54828 33494 54844
rect 33234 54729 33382 54811
rect 33122 54696 33199 54712
tri 33199 54696 33215 54712 sw
rect 33122 54630 33215 54696
rect 33251 54571 33365 54729
tri 33401 54696 33417 54712 se
rect 33417 54696 33494 54712
rect 33401 54630 33494 54696
rect 33122 54495 33494 54571
rect 33122 54370 33215 54436
rect 33122 54354 33199 54370
tri 33199 54354 33215 54370 nw
rect 33251 54337 33365 54495
rect 33401 54370 33494 54436
tri 33401 54354 33417 54370 ne
rect 33417 54354 33494 54370
rect 33234 54255 33382 54337
rect 33122 54222 33199 54238
tri 33199 54222 33215 54238 sw
rect 33122 54156 33215 54222
rect 33122 54054 33215 54120
rect 33122 54038 33199 54054
tri 33199 54038 33215 54054 nw
rect 33251 54021 33365 54255
tri 33401 54222 33417 54238 se
rect 33417 54222 33494 54238
rect 33401 54156 33494 54222
rect 33401 54054 33494 54120
tri 33401 54038 33417 54054 ne
rect 33417 54038 33494 54054
rect 33234 53939 33382 54021
rect 33122 53906 33199 53922
tri 33199 53906 33215 53922 sw
rect 33122 53840 33215 53906
rect 33251 53781 33365 53939
tri 33401 53906 33417 53922 se
rect 33417 53906 33494 53922
rect 33401 53840 33494 53906
rect 33122 53705 33494 53781
rect 33122 53580 33215 53646
rect 33122 53564 33199 53580
tri 33199 53564 33215 53580 nw
rect 33251 53547 33365 53705
rect 33401 53580 33494 53646
tri 33401 53564 33417 53580 ne
rect 33417 53564 33494 53580
rect 33234 53465 33382 53547
rect 33122 53432 33199 53448
tri 33199 53432 33215 53448 sw
rect 33122 53366 33215 53432
rect 33122 53264 33215 53330
rect 33122 53248 33199 53264
tri 33199 53248 33215 53264 nw
rect 33251 53231 33365 53465
tri 33401 53432 33417 53448 se
rect 33417 53432 33494 53448
rect 33401 53366 33494 53432
rect 33401 53264 33494 53330
tri 33401 53248 33417 53264 ne
rect 33417 53248 33494 53264
rect 33234 53149 33382 53231
rect 33122 53116 33199 53132
tri 33199 53116 33215 53132 sw
rect 33122 53050 33215 53116
rect 33251 52991 33365 53149
tri 33401 53116 33417 53132 se
rect 33417 53116 33494 53132
rect 33401 53050 33494 53116
rect 33122 52915 33494 52991
rect 33122 52790 33215 52856
rect 33122 52774 33199 52790
tri 33199 52774 33215 52790 nw
rect 33251 52757 33365 52915
rect 33401 52790 33494 52856
tri 33401 52774 33417 52790 ne
rect 33417 52774 33494 52790
rect 33234 52675 33382 52757
rect 33122 52642 33199 52658
tri 33199 52642 33215 52658 sw
rect 33122 52576 33215 52642
rect 33122 52474 33215 52540
rect 33122 52458 33199 52474
tri 33199 52458 33215 52474 nw
rect 33251 52441 33365 52675
tri 33401 52642 33417 52658 se
rect 33417 52642 33494 52658
rect 33401 52576 33494 52642
rect 33401 52474 33494 52540
tri 33401 52458 33417 52474 ne
rect 33417 52458 33494 52474
rect 33234 52359 33382 52441
rect 33122 52326 33199 52342
tri 33199 52326 33215 52342 sw
rect 33122 52260 33215 52326
rect 33251 52201 33365 52359
tri 33401 52326 33417 52342 se
rect 33417 52326 33494 52342
rect 33401 52260 33494 52326
rect 33122 52125 33494 52201
rect 33122 52000 33215 52066
rect 33122 51984 33199 52000
tri 33199 51984 33215 52000 nw
rect 33251 51967 33365 52125
rect 33401 52000 33494 52066
tri 33401 51984 33417 52000 ne
rect 33417 51984 33494 52000
rect 33234 51885 33382 51967
rect 33122 51852 33199 51868
tri 33199 51852 33215 51868 sw
rect 33122 51786 33215 51852
rect 33122 51684 33215 51750
rect 33122 51668 33199 51684
tri 33199 51668 33215 51684 nw
rect 33251 51651 33365 51885
tri 33401 51852 33417 51868 se
rect 33417 51852 33494 51868
rect 33401 51786 33494 51852
rect 33401 51684 33494 51750
tri 33401 51668 33417 51684 ne
rect 33417 51668 33494 51684
rect 33234 51569 33382 51651
rect 33122 51536 33199 51552
tri 33199 51536 33215 51552 sw
rect 33122 51470 33215 51536
rect 33251 51411 33365 51569
tri 33401 51536 33417 51552 se
rect 33417 51536 33494 51552
rect 33401 51470 33494 51536
rect 33122 51335 33494 51411
rect 33122 51210 33215 51276
rect 33122 51194 33199 51210
tri 33199 51194 33215 51210 nw
rect 33251 51177 33365 51335
rect 33401 51210 33494 51276
tri 33401 51194 33417 51210 ne
rect 33417 51194 33494 51210
rect 33234 51095 33382 51177
rect 33122 51062 33199 51078
tri 33199 51062 33215 51078 sw
rect 33122 50996 33215 51062
rect 33122 50894 33215 50960
rect 33122 50878 33199 50894
tri 33199 50878 33215 50894 nw
rect 33251 50861 33365 51095
tri 33401 51062 33417 51078 se
rect 33417 51062 33494 51078
rect 33401 50996 33494 51062
rect 33401 50894 33494 50960
tri 33401 50878 33417 50894 ne
rect 33417 50878 33494 50894
rect 33234 50779 33382 50861
rect 33122 50746 33199 50762
tri 33199 50746 33215 50762 sw
rect 33122 50680 33215 50746
rect 33251 50621 33365 50779
tri 33401 50746 33417 50762 se
rect 33417 50746 33494 50762
rect 33401 50680 33494 50746
rect 33122 50545 33494 50621
rect 33122 50420 33215 50486
rect 33122 50404 33199 50420
tri 33199 50404 33215 50420 nw
rect 33251 50387 33365 50545
rect 33401 50420 33494 50486
tri 33401 50404 33417 50420 ne
rect 33417 50404 33494 50420
rect 33234 50305 33382 50387
rect 33122 50272 33199 50288
tri 33199 50272 33215 50288 sw
rect 33122 50206 33215 50272
rect 33122 50104 33215 50170
rect 33122 50088 33199 50104
tri 33199 50088 33215 50104 nw
rect 33251 50071 33365 50305
tri 33401 50272 33417 50288 se
rect 33417 50272 33494 50288
rect 33401 50206 33494 50272
rect 33401 50104 33494 50170
tri 33401 50088 33417 50104 ne
rect 33417 50088 33494 50104
rect 33234 49989 33382 50071
rect 33122 49956 33199 49972
tri 33199 49956 33215 49972 sw
rect 33122 49890 33215 49956
rect 33251 49831 33365 49989
tri 33401 49956 33417 49972 se
rect 33417 49956 33494 49972
rect 33401 49890 33494 49956
rect 33122 49755 33494 49831
rect 33122 49630 33215 49696
rect 33122 49614 33199 49630
tri 33199 49614 33215 49630 nw
rect 33251 49597 33365 49755
rect 33401 49630 33494 49696
tri 33401 49614 33417 49630 ne
rect 33417 49614 33494 49630
rect 33234 49515 33382 49597
rect 33122 49482 33199 49498
tri 33199 49482 33215 49498 sw
rect 33122 49416 33215 49482
rect 33122 49314 33215 49380
rect 33122 49298 33199 49314
tri 33199 49298 33215 49314 nw
rect 33251 49281 33365 49515
tri 33401 49482 33417 49498 se
rect 33417 49482 33494 49498
rect 33401 49416 33494 49482
rect 33401 49314 33494 49380
tri 33401 49298 33417 49314 ne
rect 33417 49298 33494 49314
rect 33234 49199 33382 49281
rect 33122 49166 33199 49182
tri 33199 49166 33215 49182 sw
rect 33122 49100 33215 49166
rect 33251 49041 33365 49199
tri 33401 49166 33417 49182 se
rect 33417 49166 33494 49182
rect 33401 49100 33494 49166
rect 33122 48965 33494 49041
rect 33122 48840 33215 48906
rect 33122 48824 33199 48840
tri 33199 48824 33215 48840 nw
rect 33251 48807 33365 48965
rect 33401 48840 33494 48906
tri 33401 48824 33417 48840 ne
rect 33417 48824 33494 48840
rect 33234 48725 33382 48807
rect 33122 48692 33199 48708
tri 33199 48692 33215 48708 sw
rect 33122 48626 33215 48692
rect 33122 48524 33215 48590
rect 33122 48508 33199 48524
tri 33199 48508 33215 48524 nw
rect 33251 48491 33365 48725
tri 33401 48692 33417 48708 se
rect 33417 48692 33494 48708
rect 33401 48626 33494 48692
rect 33401 48524 33494 48590
tri 33401 48508 33417 48524 ne
rect 33417 48508 33494 48524
rect 33234 48409 33382 48491
rect 33122 48376 33199 48392
tri 33199 48376 33215 48392 sw
rect 33122 48310 33215 48376
rect 33251 48251 33365 48409
tri 33401 48376 33417 48392 se
rect 33417 48376 33494 48392
rect 33401 48310 33494 48376
rect 33122 48175 33494 48251
rect 33122 48050 33215 48116
rect 33122 48034 33199 48050
tri 33199 48034 33215 48050 nw
rect 33251 48017 33365 48175
rect 33401 48050 33494 48116
tri 33401 48034 33417 48050 ne
rect 33417 48034 33494 48050
rect 33234 47935 33382 48017
rect 33122 47902 33199 47918
tri 33199 47902 33215 47918 sw
rect 33122 47836 33215 47902
rect 33122 47734 33215 47800
rect 33122 47718 33199 47734
tri 33199 47718 33215 47734 nw
rect 33251 47701 33365 47935
tri 33401 47902 33417 47918 se
rect 33417 47902 33494 47918
rect 33401 47836 33494 47902
rect 33401 47734 33494 47800
tri 33401 47718 33417 47734 ne
rect 33417 47718 33494 47734
rect 33234 47619 33382 47701
rect 33122 47586 33199 47602
tri 33199 47586 33215 47602 sw
rect 33122 47520 33215 47586
rect 33251 47461 33365 47619
tri 33401 47586 33417 47602 se
rect 33417 47586 33494 47602
rect 33401 47520 33494 47586
rect 33122 47385 33494 47461
rect 33122 47260 33215 47326
rect 33122 47244 33199 47260
tri 33199 47244 33215 47260 nw
rect 33251 47227 33365 47385
rect 33401 47260 33494 47326
tri 33401 47244 33417 47260 ne
rect 33417 47244 33494 47260
rect 33234 47145 33382 47227
rect 33122 47112 33199 47128
tri 33199 47112 33215 47128 sw
rect 33122 47046 33215 47112
rect 33122 46944 33215 47010
rect 33122 46928 33199 46944
tri 33199 46928 33215 46944 nw
rect 33251 46911 33365 47145
tri 33401 47112 33417 47128 se
rect 33417 47112 33494 47128
rect 33401 47046 33494 47112
rect 33401 46944 33494 47010
tri 33401 46928 33417 46944 ne
rect 33417 46928 33494 46944
rect 33234 46829 33382 46911
rect 33122 46796 33199 46812
tri 33199 46796 33215 46812 sw
rect 33122 46730 33215 46796
rect 33251 46671 33365 46829
tri 33401 46796 33417 46812 se
rect 33417 46796 33494 46812
rect 33401 46730 33494 46796
rect 33122 46595 33494 46671
rect 33122 46470 33215 46536
rect 33122 46454 33199 46470
tri 33199 46454 33215 46470 nw
rect 33251 46437 33365 46595
rect 33401 46470 33494 46536
tri 33401 46454 33417 46470 ne
rect 33417 46454 33494 46470
rect 33234 46355 33382 46437
rect 33122 46322 33199 46338
tri 33199 46322 33215 46338 sw
rect 33122 46256 33215 46322
rect 33122 46154 33215 46220
rect 33122 46138 33199 46154
tri 33199 46138 33215 46154 nw
rect 33251 46121 33365 46355
tri 33401 46322 33417 46338 se
rect 33417 46322 33494 46338
rect 33401 46256 33494 46322
rect 33401 46154 33494 46220
tri 33401 46138 33417 46154 ne
rect 33417 46138 33494 46154
rect 33234 46039 33382 46121
rect 33122 46006 33199 46022
tri 33199 46006 33215 46022 sw
rect 33122 45940 33215 46006
rect 33251 45881 33365 46039
tri 33401 46006 33417 46022 se
rect 33417 46006 33494 46022
rect 33401 45940 33494 46006
rect 33122 45805 33494 45881
rect 33122 45680 33215 45746
rect 33122 45664 33199 45680
tri 33199 45664 33215 45680 nw
rect 33251 45647 33365 45805
rect 33401 45680 33494 45746
tri 33401 45664 33417 45680 ne
rect 33417 45664 33494 45680
rect 33234 45565 33382 45647
rect 33122 45532 33199 45548
tri 33199 45532 33215 45548 sw
rect 33122 45466 33215 45532
rect 33122 45364 33215 45430
rect 33122 45348 33199 45364
tri 33199 45348 33215 45364 nw
rect 33251 45331 33365 45565
tri 33401 45532 33417 45548 se
rect 33417 45532 33494 45548
rect 33401 45466 33494 45532
rect 33401 45364 33494 45430
tri 33401 45348 33417 45364 ne
rect 33417 45348 33494 45364
rect 33234 45249 33382 45331
rect 33122 45216 33199 45232
tri 33199 45216 33215 45232 sw
rect 33122 45150 33215 45216
rect 33251 45091 33365 45249
tri 33401 45216 33417 45232 se
rect 33417 45216 33494 45232
rect 33401 45150 33494 45216
rect 33122 45015 33494 45091
rect 33122 44890 33215 44956
rect 33122 44874 33199 44890
tri 33199 44874 33215 44890 nw
rect 33251 44857 33365 45015
rect 33401 44890 33494 44956
tri 33401 44874 33417 44890 ne
rect 33417 44874 33494 44890
rect 33234 44775 33382 44857
rect 33122 44742 33199 44758
tri 33199 44742 33215 44758 sw
rect 33122 44676 33215 44742
rect 33122 44574 33215 44640
rect 33122 44558 33199 44574
tri 33199 44558 33215 44574 nw
rect 33251 44541 33365 44775
tri 33401 44742 33417 44758 se
rect 33417 44742 33494 44758
rect 33401 44676 33494 44742
rect 33401 44574 33494 44640
tri 33401 44558 33417 44574 ne
rect 33417 44558 33494 44574
rect 33234 44459 33382 44541
rect 33122 44426 33199 44442
tri 33199 44426 33215 44442 sw
rect 33122 44360 33215 44426
rect 33251 44301 33365 44459
tri 33401 44426 33417 44442 se
rect 33417 44426 33494 44442
rect 33401 44360 33494 44426
rect 33122 44225 33494 44301
rect 33122 44100 33215 44166
rect 33122 44084 33199 44100
tri 33199 44084 33215 44100 nw
rect 33251 44067 33365 44225
rect 33401 44100 33494 44166
tri 33401 44084 33417 44100 ne
rect 33417 44084 33494 44100
rect 33234 43985 33382 44067
rect 33122 43952 33199 43968
tri 33199 43952 33215 43968 sw
rect 33122 43886 33215 43952
rect 33122 43784 33215 43850
rect 33122 43768 33199 43784
tri 33199 43768 33215 43784 nw
rect 33251 43751 33365 43985
tri 33401 43952 33417 43968 se
rect 33417 43952 33494 43968
rect 33401 43886 33494 43952
rect 33401 43784 33494 43850
tri 33401 43768 33417 43784 ne
rect 33417 43768 33494 43784
rect 33234 43669 33382 43751
rect 33122 43636 33199 43652
tri 33199 43636 33215 43652 sw
rect 33122 43570 33215 43636
rect 33251 43511 33365 43669
tri 33401 43636 33417 43652 se
rect 33417 43636 33494 43652
rect 33401 43570 33494 43636
rect 33122 43435 33494 43511
rect 33122 43310 33215 43376
rect 33122 43294 33199 43310
tri 33199 43294 33215 43310 nw
rect 33251 43277 33365 43435
rect 33401 43310 33494 43376
tri 33401 43294 33417 43310 ne
rect 33417 43294 33494 43310
rect 33234 43195 33382 43277
rect 33122 43162 33199 43178
tri 33199 43162 33215 43178 sw
rect 33122 43096 33215 43162
rect 33122 42994 33215 43060
rect 33122 42978 33199 42994
tri 33199 42978 33215 42994 nw
rect 33251 42961 33365 43195
tri 33401 43162 33417 43178 se
rect 33417 43162 33494 43178
rect 33401 43096 33494 43162
rect 33401 42994 33494 43060
tri 33401 42978 33417 42994 ne
rect 33417 42978 33494 42994
rect 33234 42879 33382 42961
rect 33122 42846 33199 42862
tri 33199 42846 33215 42862 sw
rect 33122 42780 33215 42846
rect 33251 42721 33365 42879
tri 33401 42846 33417 42862 se
rect 33417 42846 33494 42862
rect 33401 42780 33494 42846
rect 33122 42645 33494 42721
rect 33122 42520 33215 42586
rect 33122 42504 33199 42520
tri 33199 42504 33215 42520 nw
rect 33251 42487 33365 42645
rect 33401 42520 33494 42586
tri 33401 42504 33417 42520 ne
rect 33417 42504 33494 42520
rect 33234 42405 33382 42487
rect 33122 42372 33199 42388
tri 33199 42372 33215 42388 sw
rect 33122 42306 33215 42372
rect 33122 42204 33215 42270
rect 33122 42188 33199 42204
tri 33199 42188 33215 42204 nw
rect 33251 42171 33365 42405
tri 33401 42372 33417 42388 se
rect 33417 42372 33494 42388
rect 33401 42306 33494 42372
rect 33401 42204 33494 42270
tri 33401 42188 33417 42204 ne
rect 33417 42188 33494 42204
rect 33234 42089 33382 42171
rect 33122 42056 33199 42072
tri 33199 42056 33215 42072 sw
rect 33122 41990 33215 42056
rect 33251 41931 33365 42089
tri 33401 42056 33417 42072 se
rect 33417 42056 33494 42072
rect 33401 41990 33494 42056
rect 33122 41855 33494 41931
rect 33122 41730 33215 41796
rect 33122 41714 33199 41730
tri 33199 41714 33215 41730 nw
rect 33251 41697 33365 41855
rect 33401 41730 33494 41796
tri 33401 41714 33417 41730 ne
rect 33417 41714 33494 41730
rect 33234 41615 33382 41697
rect 33122 41582 33199 41598
tri 33199 41582 33215 41598 sw
rect 33122 41516 33215 41582
rect 33122 41414 33215 41480
rect 33122 41398 33199 41414
tri 33199 41398 33215 41414 nw
rect 33251 41381 33365 41615
tri 33401 41582 33417 41598 se
rect 33417 41582 33494 41598
rect 33401 41516 33494 41582
rect 33401 41414 33494 41480
tri 33401 41398 33417 41414 ne
rect 33417 41398 33494 41414
rect 33234 41299 33382 41381
rect 33122 41266 33199 41282
tri 33199 41266 33215 41282 sw
rect 33122 41200 33215 41266
rect 33251 41141 33365 41299
tri 33401 41266 33417 41282 se
rect 33417 41266 33494 41282
rect 33401 41200 33494 41266
rect 33122 41065 33494 41141
rect 33122 40940 33215 41006
rect 33122 40924 33199 40940
tri 33199 40924 33215 40940 nw
rect 33251 40907 33365 41065
rect 33401 40940 33494 41006
tri 33401 40924 33417 40940 ne
rect 33417 40924 33494 40940
rect 33234 40825 33382 40907
rect 33122 40792 33199 40808
tri 33199 40792 33215 40808 sw
rect 33122 40726 33215 40792
rect 33122 40624 33215 40690
rect 33122 40608 33199 40624
tri 33199 40608 33215 40624 nw
rect 33251 40591 33365 40825
tri 33401 40792 33417 40808 se
rect 33417 40792 33494 40808
rect 33401 40726 33494 40792
rect 33401 40624 33494 40690
tri 33401 40608 33417 40624 ne
rect 33417 40608 33494 40624
rect 33234 40509 33382 40591
rect 33122 40476 33199 40492
tri 33199 40476 33215 40492 sw
rect 33122 40410 33215 40476
rect 33251 40351 33365 40509
tri 33401 40476 33417 40492 se
rect 33417 40476 33494 40492
rect 33401 40410 33494 40476
rect 33122 40275 33494 40351
rect 33122 40150 33215 40216
rect 33122 40134 33199 40150
tri 33199 40134 33215 40150 nw
rect 33251 40117 33365 40275
rect 33401 40150 33494 40216
tri 33401 40134 33417 40150 ne
rect 33417 40134 33494 40150
rect 33234 40035 33382 40117
rect 33122 40002 33199 40018
tri 33199 40002 33215 40018 sw
rect 33122 39936 33215 40002
rect 33122 39834 33215 39900
rect 33122 39818 33199 39834
tri 33199 39818 33215 39834 nw
rect 33251 39801 33365 40035
tri 33401 40002 33417 40018 se
rect 33417 40002 33494 40018
rect 33401 39936 33494 40002
rect 33401 39834 33494 39900
tri 33401 39818 33417 39834 ne
rect 33417 39818 33494 39834
rect 33234 39719 33382 39801
rect 33122 39686 33199 39702
tri 33199 39686 33215 39702 sw
rect 33122 39620 33215 39686
rect 33251 39561 33365 39719
tri 33401 39686 33417 39702 se
rect 33417 39686 33494 39702
rect 33401 39620 33494 39686
rect 33122 39485 33494 39561
rect 33122 39360 33215 39426
rect 33122 39344 33199 39360
tri 33199 39344 33215 39360 nw
rect 33251 39327 33365 39485
rect 33401 39360 33494 39426
tri 33401 39344 33417 39360 ne
rect 33417 39344 33494 39360
rect 33234 39245 33382 39327
rect 33122 39212 33199 39228
tri 33199 39212 33215 39228 sw
rect 33122 39146 33215 39212
rect 33122 39044 33215 39110
rect 33122 39028 33199 39044
tri 33199 39028 33215 39044 nw
rect 33251 39011 33365 39245
tri 33401 39212 33417 39228 se
rect 33417 39212 33494 39228
rect 33401 39146 33494 39212
rect 33401 39044 33494 39110
tri 33401 39028 33417 39044 ne
rect 33417 39028 33494 39044
rect 33234 38929 33382 39011
rect 33122 38896 33199 38912
tri 33199 38896 33215 38912 sw
rect 33122 38830 33215 38896
rect 33251 38771 33365 38929
tri 33401 38896 33417 38912 se
rect 33417 38896 33494 38912
rect 33401 38830 33494 38896
rect 33122 38695 33494 38771
rect 33122 38570 33215 38636
rect 33122 38554 33199 38570
tri 33199 38554 33215 38570 nw
rect 33251 38537 33365 38695
rect 33401 38570 33494 38636
tri 33401 38554 33417 38570 ne
rect 33417 38554 33494 38570
rect 33234 38455 33382 38537
rect 33122 38422 33199 38438
tri 33199 38422 33215 38438 sw
rect 33122 38356 33215 38422
rect 33122 38254 33215 38320
rect 33122 38238 33199 38254
tri 33199 38238 33215 38254 nw
rect 33251 38221 33365 38455
tri 33401 38422 33417 38438 se
rect 33417 38422 33494 38438
rect 33401 38356 33494 38422
rect 33401 38254 33494 38320
tri 33401 38238 33417 38254 ne
rect 33417 38238 33494 38254
rect 33234 38139 33382 38221
rect 33122 38106 33199 38122
tri 33199 38106 33215 38122 sw
rect 33122 38040 33215 38106
rect 33251 37981 33365 38139
tri 33401 38106 33417 38122 se
rect 33417 38106 33494 38122
rect 33401 38040 33494 38106
rect 33122 37905 33494 37981
rect 33122 37780 33215 37846
rect 33122 37764 33199 37780
tri 33199 37764 33215 37780 nw
rect 33251 37747 33365 37905
rect 33401 37780 33494 37846
tri 33401 37764 33417 37780 ne
rect 33417 37764 33494 37780
rect 33234 37665 33382 37747
rect 33122 37632 33199 37648
tri 33199 37632 33215 37648 sw
rect 33122 37566 33215 37632
rect 33122 37464 33215 37530
rect 33122 37448 33199 37464
tri 33199 37448 33215 37464 nw
rect 33251 37431 33365 37665
tri 33401 37632 33417 37648 se
rect 33417 37632 33494 37648
rect 33401 37566 33494 37632
rect 33401 37464 33494 37530
tri 33401 37448 33417 37464 ne
rect 33417 37448 33494 37464
rect 33234 37349 33382 37431
rect 33122 37316 33199 37332
tri 33199 37316 33215 37332 sw
rect 33122 37250 33215 37316
rect 33251 37191 33365 37349
tri 33401 37316 33417 37332 se
rect 33417 37316 33494 37332
rect 33401 37250 33494 37316
rect 33122 37115 33494 37191
rect 33122 36990 33215 37056
rect 33122 36974 33199 36990
tri 33199 36974 33215 36990 nw
rect 33251 36957 33365 37115
rect 33401 36990 33494 37056
tri 33401 36974 33417 36990 ne
rect 33417 36974 33494 36990
rect 33234 36875 33382 36957
rect 33122 36842 33199 36858
tri 33199 36842 33215 36858 sw
rect 33122 36776 33215 36842
rect 33122 36674 33215 36740
rect 33122 36658 33199 36674
tri 33199 36658 33215 36674 nw
rect 33251 36641 33365 36875
tri 33401 36842 33417 36858 se
rect 33417 36842 33494 36858
rect 33401 36776 33494 36842
rect 33401 36674 33494 36740
tri 33401 36658 33417 36674 ne
rect 33417 36658 33494 36674
rect 33234 36559 33382 36641
rect 33122 36526 33199 36542
tri 33199 36526 33215 36542 sw
rect 33122 36460 33215 36526
rect 33251 36401 33365 36559
tri 33401 36526 33417 36542 se
rect 33417 36526 33494 36542
rect 33401 36460 33494 36526
rect 33122 36325 33494 36401
rect 33122 36200 33215 36266
rect 33122 36184 33199 36200
tri 33199 36184 33215 36200 nw
rect 33251 36167 33365 36325
rect 33401 36200 33494 36266
tri 33401 36184 33417 36200 ne
rect 33417 36184 33494 36200
rect 33234 36085 33382 36167
rect 33122 36052 33199 36068
tri 33199 36052 33215 36068 sw
rect 33122 35986 33215 36052
rect 33122 35884 33215 35950
rect 33122 35868 33199 35884
tri 33199 35868 33215 35884 nw
rect 33251 35851 33365 36085
tri 33401 36052 33417 36068 se
rect 33417 36052 33494 36068
rect 33401 35986 33494 36052
rect 33401 35884 33494 35950
tri 33401 35868 33417 35884 ne
rect 33417 35868 33494 35884
rect 33234 35769 33382 35851
rect 33122 35736 33199 35752
tri 33199 35736 33215 35752 sw
rect 33122 35670 33215 35736
rect 33251 35611 33365 35769
tri 33401 35736 33417 35752 se
rect 33417 35736 33494 35752
rect 33401 35670 33494 35736
rect 33122 35535 33494 35611
rect 33122 35410 33215 35476
rect 33122 35394 33199 35410
tri 33199 35394 33215 35410 nw
rect 33251 35377 33365 35535
rect 33401 35410 33494 35476
tri 33401 35394 33417 35410 ne
rect 33417 35394 33494 35410
rect 33234 35295 33382 35377
rect 33122 35262 33199 35278
tri 33199 35262 33215 35278 sw
rect 33122 35196 33215 35262
rect 33122 35094 33215 35160
rect 33122 35078 33199 35094
tri 33199 35078 33215 35094 nw
rect 33251 35061 33365 35295
tri 33401 35262 33417 35278 se
rect 33417 35262 33494 35278
rect 33401 35196 33494 35262
rect 33401 35094 33494 35160
tri 33401 35078 33417 35094 ne
rect 33417 35078 33494 35094
rect 33234 34979 33382 35061
rect 33122 34946 33199 34962
tri 33199 34946 33215 34962 sw
rect 33122 34880 33215 34946
rect 33251 34821 33365 34979
tri 33401 34946 33417 34962 se
rect 33417 34946 33494 34962
rect 33401 34880 33494 34946
rect 33122 34745 33494 34821
rect 33122 34620 33215 34686
rect 33122 34604 33199 34620
tri 33199 34604 33215 34620 nw
rect 33251 34587 33365 34745
rect 33401 34620 33494 34686
tri 33401 34604 33417 34620 ne
rect 33417 34604 33494 34620
rect 33234 34505 33382 34587
rect 33122 34472 33199 34488
tri 33199 34472 33215 34488 sw
rect 33122 34406 33215 34472
rect 33122 34304 33215 34370
rect 33122 34288 33199 34304
tri 33199 34288 33215 34304 nw
rect 33251 34271 33365 34505
tri 33401 34472 33417 34488 se
rect 33417 34472 33494 34488
rect 33401 34406 33494 34472
rect 33401 34304 33494 34370
tri 33401 34288 33417 34304 ne
rect 33417 34288 33494 34304
rect 33234 34189 33382 34271
rect 33122 34156 33199 34172
tri 33199 34156 33215 34172 sw
rect 33122 34090 33215 34156
rect 33251 34031 33365 34189
tri 33401 34156 33417 34172 se
rect 33417 34156 33494 34172
rect 33401 34090 33494 34156
rect 33122 33955 33494 34031
rect 33122 33830 33215 33896
rect 33122 33814 33199 33830
tri 33199 33814 33215 33830 nw
rect 33251 33797 33365 33955
rect 33401 33830 33494 33896
tri 33401 33814 33417 33830 ne
rect 33417 33814 33494 33830
rect 33234 33715 33382 33797
rect 33122 33682 33199 33698
tri 33199 33682 33215 33698 sw
rect 33122 33616 33215 33682
rect 33122 33514 33215 33580
rect 33122 33498 33199 33514
tri 33199 33498 33215 33514 nw
rect 33251 33481 33365 33715
tri 33401 33682 33417 33698 se
rect 33417 33682 33494 33698
rect 33401 33616 33494 33682
rect 33401 33514 33494 33580
tri 33401 33498 33417 33514 ne
rect 33417 33498 33494 33514
rect 33234 33399 33382 33481
rect 33122 33366 33199 33382
tri 33199 33366 33215 33382 sw
rect 33122 33300 33215 33366
rect 33251 33241 33365 33399
tri 33401 33366 33417 33382 se
rect 33417 33366 33494 33382
rect 33401 33300 33494 33366
rect 33122 33165 33494 33241
rect 33122 33040 33215 33106
rect 33122 33024 33199 33040
tri 33199 33024 33215 33040 nw
rect 33251 33007 33365 33165
rect 33401 33040 33494 33106
tri 33401 33024 33417 33040 ne
rect 33417 33024 33494 33040
rect 33234 32925 33382 33007
rect 33122 32892 33199 32908
tri 33199 32892 33215 32908 sw
rect 33122 32826 33215 32892
rect 33122 32724 33215 32790
rect 33122 32708 33199 32724
tri 33199 32708 33215 32724 nw
rect 33251 32691 33365 32925
tri 33401 32892 33417 32908 se
rect 33417 32892 33494 32908
rect 33401 32826 33494 32892
rect 33401 32724 33494 32790
tri 33401 32708 33417 32724 ne
rect 33417 32708 33494 32724
rect 33234 32609 33382 32691
rect 33122 32576 33199 32592
tri 33199 32576 33215 32592 sw
rect 33122 32510 33215 32576
rect 33251 32451 33365 32609
tri 33401 32576 33417 32592 se
rect 33417 32576 33494 32592
rect 33401 32510 33494 32576
rect 33122 32375 33494 32451
rect 33122 32250 33215 32316
rect 33122 32234 33199 32250
tri 33199 32234 33215 32250 nw
rect 33251 32217 33365 32375
rect 33401 32250 33494 32316
tri 33401 32234 33417 32250 ne
rect 33417 32234 33494 32250
rect 33234 32135 33382 32217
rect 33122 32102 33199 32118
tri 33199 32102 33215 32118 sw
rect 33122 32036 33215 32102
rect 33122 31934 33215 32000
rect 33122 31918 33199 31934
tri 33199 31918 33215 31934 nw
rect 33251 31901 33365 32135
tri 33401 32102 33417 32118 se
rect 33417 32102 33494 32118
rect 33401 32036 33494 32102
rect 33401 31934 33494 32000
tri 33401 31918 33417 31934 ne
rect 33417 31918 33494 31934
rect 33234 31819 33382 31901
rect 33122 31786 33199 31802
tri 33199 31786 33215 31802 sw
rect 33122 31720 33215 31786
rect 33251 31661 33365 31819
tri 33401 31786 33417 31802 se
rect 33417 31786 33494 31802
rect 33401 31720 33494 31786
rect 33122 31585 33494 31661
rect 33122 31460 33215 31526
rect 33122 31444 33199 31460
tri 33199 31444 33215 31460 nw
rect 33251 31427 33365 31585
rect 33401 31460 33494 31526
tri 33401 31444 33417 31460 ne
rect 33417 31444 33494 31460
rect 33234 31345 33382 31427
rect 33122 31312 33199 31328
tri 33199 31312 33215 31328 sw
rect 33122 31246 33215 31312
rect 33122 31144 33215 31210
rect 33122 31128 33199 31144
tri 33199 31128 33215 31144 nw
rect 33251 31111 33365 31345
tri 33401 31312 33417 31328 se
rect 33417 31312 33494 31328
rect 33401 31246 33494 31312
rect 33401 31144 33494 31210
tri 33401 31128 33417 31144 ne
rect 33417 31128 33494 31144
rect 33234 31029 33382 31111
rect 33122 30996 33199 31012
tri 33199 30996 33215 31012 sw
rect 33122 30930 33215 30996
rect 33251 30871 33365 31029
tri 33401 30996 33417 31012 se
rect 33417 30996 33494 31012
rect 33401 30930 33494 30996
rect 33122 30795 33494 30871
rect 33122 30670 33215 30736
rect 33122 30654 33199 30670
tri 33199 30654 33215 30670 nw
rect 33251 30637 33365 30795
rect 33401 30670 33494 30736
tri 33401 30654 33417 30670 ne
rect 33417 30654 33494 30670
rect 33234 30555 33382 30637
rect 33122 30522 33199 30538
tri 33199 30522 33215 30538 sw
rect 33122 30456 33215 30522
rect 33122 30354 33215 30420
rect 33122 30338 33199 30354
tri 33199 30338 33215 30354 nw
rect 33251 30321 33365 30555
tri 33401 30522 33417 30538 se
rect 33417 30522 33494 30538
rect 33401 30456 33494 30522
rect 33401 30354 33494 30420
tri 33401 30338 33417 30354 ne
rect 33417 30338 33494 30354
rect 33234 30239 33382 30321
rect 33122 30206 33199 30222
tri 33199 30206 33215 30222 sw
rect 33122 30140 33215 30206
rect 33251 30081 33365 30239
tri 33401 30206 33417 30222 se
rect 33417 30206 33494 30222
rect 33401 30140 33494 30206
rect 33122 30005 33494 30081
rect 33122 29880 33215 29946
rect 33122 29864 33199 29880
tri 33199 29864 33215 29880 nw
rect 33251 29847 33365 30005
rect 33401 29880 33494 29946
tri 33401 29864 33417 29880 ne
rect 33417 29864 33494 29880
rect 33234 29765 33382 29847
rect 33122 29732 33199 29748
tri 33199 29732 33215 29748 sw
rect 33122 29666 33215 29732
rect 33122 29564 33215 29630
rect 33122 29548 33199 29564
tri 33199 29548 33215 29564 nw
rect 33251 29531 33365 29765
tri 33401 29732 33417 29748 se
rect 33417 29732 33494 29748
rect 33401 29666 33494 29732
rect 33401 29564 33494 29630
tri 33401 29548 33417 29564 ne
rect 33417 29548 33494 29564
rect 33234 29449 33382 29531
rect 33122 29416 33199 29432
tri 33199 29416 33215 29432 sw
rect 33122 29350 33215 29416
rect 33251 29291 33365 29449
tri 33401 29416 33417 29432 se
rect 33417 29416 33494 29432
rect 33401 29350 33494 29416
rect 33122 29215 33494 29291
rect 33122 29090 33215 29156
rect 33122 29074 33199 29090
tri 33199 29074 33215 29090 nw
rect 33251 29057 33365 29215
rect 33401 29090 33494 29156
tri 33401 29074 33417 29090 ne
rect 33417 29074 33494 29090
rect 33234 28975 33382 29057
rect 33122 28942 33199 28958
tri 33199 28942 33215 28958 sw
rect 33122 28876 33215 28942
rect 33251 28833 33365 28975
tri 33401 28942 33417 28958 se
rect 33417 28942 33494 28958
rect 33401 28876 33494 28942
rect 33530 28463 33566 80603
rect 33602 28463 33638 80603
rect 33674 80445 33710 80603
rect 33666 80303 33718 80445
rect 33674 28763 33710 80303
rect 33666 28621 33718 28763
rect 33674 28463 33710 28621
rect 33746 28463 33782 80603
rect 33818 28463 33854 80603
rect 33890 28833 33974 80233
rect 34010 28463 34046 80603
rect 34082 28463 34118 80603
rect 34154 80445 34190 80603
rect 34146 80303 34198 80445
rect 34154 28763 34190 80303
rect 34146 28621 34198 28763
rect 34154 28463 34190 28621
rect 34226 28463 34262 80603
rect 34298 28463 34334 80603
rect 34370 80124 34463 80190
rect 34370 80108 34447 80124
tri 34447 80108 34463 80124 nw
rect 34499 80091 34613 80233
rect 34649 80124 34742 80190
tri 34649 80108 34665 80124 ne
rect 34665 80108 34742 80124
rect 34482 80009 34630 80091
rect 34370 79976 34447 79992
tri 34447 79976 34463 79992 sw
rect 34370 79910 34463 79976
rect 34499 79851 34613 80009
tri 34649 79976 34665 79992 se
rect 34665 79976 34742 79992
rect 34649 79910 34742 79976
rect 34370 79775 34742 79851
rect 34370 79650 34463 79716
rect 34370 79634 34447 79650
tri 34447 79634 34463 79650 nw
rect 34499 79617 34613 79775
rect 34649 79650 34742 79716
tri 34649 79634 34665 79650 ne
rect 34665 79634 34742 79650
rect 34482 79535 34630 79617
rect 34370 79502 34447 79518
tri 34447 79502 34463 79518 sw
rect 34370 79436 34463 79502
rect 34370 79334 34463 79400
rect 34370 79318 34447 79334
tri 34447 79318 34463 79334 nw
rect 34499 79301 34613 79535
tri 34649 79502 34665 79518 se
rect 34665 79502 34742 79518
rect 34649 79436 34742 79502
rect 34649 79334 34742 79400
tri 34649 79318 34665 79334 ne
rect 34665 79318 34742 79334
rect 34482 79219 34630 79301
rect 34370 79186 34447 79202
tri 34447 79186 34463 79202 sw
rect 34370 79120 34463 79186
rect 34499 79061 34613 79219
tri 34649 79186 34665 79202 se
rect 34665 79186 34742 79202
rect 34649 79120 34742 79186
rect 34370 78985 34742 79061
rect 34370 78860 34463 78926
rect 34370 78844 34447 78860
tri 34447 78844 34463 78860 nw
rect 34499 78827 34613 78985
rect 34649 78860 34742 78926
tri 34649 78844 34665 78860 ne
rect 34665 78844 34742 78860
rect 34482 78745 34630 78827
rect 34370 78712 34447 78728
tri 34447 78712 34463 78728 sw
rect 34370 78646 34463 78712
rect 34370 78544 34463 78610
rect 34370 78528 34447 78544
tri 34447 78528 34463 78544 nw
rect 34499 78511 34613 78745
tri 34649 78712 34665 78728 se
rect 34665 78712 34742 78728
rect 34649 78646 34742 78712
rect 34649 78544 34742 78610
tri 34649 78528 34665 78544 ne
rect 34665 78528 34742 78544
rect 34482 78429 34630 78511
rect 34370 78396 34447 78412
tri 34447 78396 34463 78412 sw
rect 34370 78330 34463 78396
rect 34499 78271 34613 78429
tri 34649 78396 34665 78412 se
rect 34665 78396 34742 78412
rect 34649 78330 34742 78396
rect 34370 78195 34742 78271
rect 34370 78070 34463 78136
rect 34370 78054 34447 78070
tri 34447 78054 34463 78070 nw
rect 34499 78037 34613 78195
rect 34649 78070 34742 78136
tri 34649 78054 34665 78070 ne
rect 34665 78054 34742 78070
rect 34482 77955 34630 78037
rect 34370 77922 34447 77938
tri 34447 77922 34463 77938 sw
rect 34370 77856 34463 77922
rect 34370 77754 34463 77820
rect 34370 77738 34447 77754
tri 34447 77738 34463 77754 nw
rect 34499 77721 34613 77955
tri 34649 77922 34665 77938 se
rect 34665 77922 34742 77938
rect 34649 77856 34742 77922
rect 34649 77754 34742 77820
tri 34649 77738 34665 77754 ne
rect 34665 77738 34742 77754
rect 34482 77639 34630 77721
rect 34370 77606 34447 77622
tri 34447 77606 34463 77622 sw
rect 34370 77540 34463 77606
rect 34499 77481 34613 77639
tri 34649 77606 34665 77622 se
rect 34665 77606 34742 77622
rect 34649 77540 34742 77606
rect 34370 77405 34742 77481
rect 34370 77280 34463 77346
rect 34370 77264 34447 77280
tri 34447 77264 34463 77280 nw
rect 34499 77247 34613 77405
rect 34649 77280 34742 77346
tri 34649 77264 34665 77280 ne
rect 34665 77264 34742 77280
rect 34482 77165 34630 77247
rect 34370 77132 34447 77148
tri 34447 77132 34463 77148 sw
rect 34370 77066 34463 77132
rect 34370 76964 34463 77030
rect 34370 76948 34447 76964
tri 34447 76948 34463 76964 nw
rect 34499 76931 34613 77165
tri 34649 77132 34665 77148 se
rect 34665 77132 34742 77148
rect 34649 77066 34742 77132
rect 34649 76964 34742 77030
tri 34649 76948 34665 76964 ne
rect 34665 76948 34742 76964
rect 34482 76849 34630 76931
rect 34370 76816 34447 76832
tri 34447 76816 34463 76832 sw
rect 34370 76750 34463 76816
rect 34499 76691 34613 76849
tri 34649 76816 34665 76832 se
rect 34665 76816 34742 76832
rect 34649 76750 34742 76816
rect 34370 76615 34742 76691
rect 34370 76490 34463 76556
rect 34370 76474 34447 76490
tri 34447 76474 34463 76490 nw
rect 34499 76457 34613 76615
rect 34649 76490 34742 76556
tri 34649 76474 34665 76490 ne
rect 34665 76474 34742 76490
rect 34482 76375 34630 76457
rect 34370 76342 34447 76358
tri 34447 76342 34463 76358 sw
rect 34370 76276 34463 76342
rect 34370 76174 34463 76240
rect 34370 76158 34447 76174
tri 34447 76158 34463 76174 nw
rect 34499 76141 34613 76375
tri 34649 76342 34665 76358 se
rect 34665 76342 34742 76358
rect 34649 76276 34742 76342
rect 34649 76174 34742 76240
tri 34649 76158 34665 76174 ne
rect 34665 76158 34742 76174
rect 34482 76059 34630 76141
rect 34370 76026 34447 76042
tri 34447 76026 34463 76042 sw
rect 34370 75960 34463 76026
rect 34499 75901 34613 76059
tri 34649 76026 34665 76042 se
rect 34665 76026 34742 76042
rect 34649 75960 34742 76026
rect 34370 75825 34742 75901
rect 34370 75700 34463 75766
rect 34370 75684 34447 75700
tri 34447 75684 34463 75700 nw
rect 34499 75667 34613 75825
rect 34649 75700 34742 75766
tri 34649 75684 34665 75700 ne
rect 34665 75684 34742 75700
rect 34482 75585 34630 75667
rect 34370 75552 34447 75568
tri 34447 75552 34463 75568 sw
rect 34370 75486 34463 75552
rect 34370 75384 34463 75450
rect 34370 75368 34447 75384
tri 34447 75368 34463 75384 nw
rect 34499 75351 34613 75585
tri 34649 75552 34665 75568 se
rect 34665 75552 34742 75568
rect 34649 75486 34742 75552
rect 34649 75384 34742 75450
tri 34649 75368 34665 75384 ne
rect 34665 75368 34742 75384
rect 34482 75269 34630 75351
rect 34370 75236 34447 75252
tri 34447 75236 34463 75252 sw
rect 34370 75170 34463 75236
rect 34499 75111 34613 75269
tri 34649 75236 34665 75252 se
rect 34665 75236 34742 75252
rect 34649 75170 34742 75236
rect 34370 75035 34742 75111
rect 34370 74910 34463 74976
rect 34370 74894 34447 74910
tri 34447 74894 34463 74910 nw
rect 34499 74877 34613 75035
rect 34649 74910 34742 74976
tri 34649 74894 34665 74910 ne
rect 34665 74894 34742 74910
rect 34482 74795 34630 74877
rect 34370 74762 34447 74778
tri 34447 74762 34463 74778 sw
rect 34370 74696 34463 74762
rect 34370 74594 34463 74660
rect 34370 74578 34447 74594
tri 34447 74578 34463 74594 nw
rect 34499 74561 34613 74795
tri 34649 74762 34665 74778 se
rect 34665 74762 34742 74778
rect 34649 74696 34742 74762
rect 34649 74594 34742 74660
tri 34649 74578 34665 74594 ne
rect 34665 74578 34742 74594
rect 34482 74479 34630 74561
rect 34370 74446 34447 74462
tri 34447 74446 34463 74462 sw
rect 34370 74380 34463 74446
rect 34499 74321 34613 74479
tri 34649 74446 34665 74462 se
rect 34665 74446 34742 74462
rect 34649 74380 34742 74446
rect 34370 74245 34742 74321
rect 34370 74120 34463 74186
rect 34370 74104 34447 74120
tri 34447 74104 34463 74120 nw
rect 34499 74087 34613 74245
rect 34649 74120 34742 74186
tri 34649 74104 34665 74120 ne
rect 34665 74104 34742 74120
rect 34482 74005 34630 74087
rect 34370 73972 34447 73988
tri 34447 73972 34463 73988 sw
rect 34370 73906 34463 73972
rect 34370 73804 34463 73870
rect 34370 73788 34447 73804
tri 34447 73788 34463 73804 nw
rect 34499 73771 34613 74005
tri 34649 73972 34665 73988 se
rect 34665 73972 34742 73988
rect 34649 73906 34742 73972
rect 34649 73804 34742 73870
tri 34649 73788 34665 73804 ne
rect 34665 73788 34742 73804
rect 34482 73689 34630 73771
rect 34370 73656 34447 73672
tri 34447 73656 34463 73672 sw
rect 34370 73590 34463 73656
rect 34499 73531 34613 73689
tri 34649 73656 34665 73672 se
rect 34665 73656 34742 73672
rect 34649 73590 34742 73656
rect 34370 73455 34742 73531
rect 34370 73330 34463 73396
rect 34370 73314 34447 73330
tri 34447 73314 34463 73330 nw
rect 34499 73297 34613 73455
rect 34649 73330 34742 73396
tri 34649 73314 34665 73330 ne
rect 34665 73314 34742 73330
rect 34482 73215 34630 73297
rect 34370 73182 34447 73198
tri 34447 73182 34463 73198 sw
rect 34370 73116 34463 73182
rect 34370 73014 34463 73080
rect 34370 72998 34447 73014
tri 34447 72998 34463 73014 nw
rect 34499 72981 34613 73215
tri 34649 73182 34665 73198 se
rect 34665 73182 34742 73198
rect 34649 73116 34742 73182
rect 34649 73014 34742 73080
tri 34649 72998 34665 73014 ne
rect 34665 72998 34742 73014
rect 34482 72899 34630 72981
rect 34370 72866 34447 72882
tri 34447 72866 34463 72882 sw
rect 34370 72800 34463 72866
rect 34499 72741 34613 72899
tri 34649 72866 34665 72882 se
rect 34665 72866 34742 72882
rect 34649 72800 34742 72866
rect 34370 72665 34742 72741
rect 34370 72540 34463 72606
rect 34370 72524 34447 72540
tri 34447 72524 34463 72540 nw
rect 34499 72507 34613 72665
rect 34649 72540 34742 72606
tri 34649 72524 34665 72540 ne
rect 34665 72524 34742 72540
rect 34482 72425 34630 72507
rect 34370 72392 34447 72408
tri 34447 72392 34463 72408 sw
rect 34370 72326 34463 72392
rect 34370 72224 34463 72290
rect 34370 72208 34447 72224
tri 34447 72208 34463 72224 nw
rect 34499 72191 34613 72425
tri 34649 72392 34665 72408 se
rect 34665 72392 34742 72408
rect 34649 72326 34742 72392
rect 34649 72224 34742 72290
tri 34649 72208 34665 72224 ne
rect 34665 72208 34742 72224
rect 34482 72109 34630 72191
rect 34370 72076 34447 72092
tri 34447 72076 34463 72092 sw
rect 34370 72010 34463 72076
rect 34499 71951 34613 72109
tri 34649 72076 34665 72092 se
rect 34665 72076 34742 72092
rect 34649 72010 34742 72076
rect 34370 71875 34742 71951
rect 34370 71750 34463 71816
rect 34370 71734 34447 71750
tri 34447 71734 34463 71750 nw
rect 34499 71717 34613 71875
rect 34649 71750 34742 71816
tri 34649 71734 34665 71750 ne
rect 34665 71734 34742 71750
rect 34482 71635 34630 71717
rect 34370 71602 34447 71618
tri 34447 71602 34463 71618 sw
rect 34370 71536 34463 71602
rect 34370 71434 34463 71500
rect 34370 71418 34447 71434
tri 34447 71418 34463 71434 nw
rect 34499 71401 34613 71635
tri 34649 71602 34665 71618 se
rect 34665 71602 34742 71618
rect 34649 71536 34742 71602
rect 34649 71434 34742 71500
tri 34649 71418 34665 71434 ne
rect 34665 71418 34742 71434
rect 34482 71319 34630 71401
rect 34370 71286 34447 71302
tri 34447 71286 34463 71302 sw
rect 34370 71220 34463 71286
rect 34499 71161 34613 71319
tri 34649 71286 34665 71302 se
rect 34665 71286 34742 71302
rect 34649 71220 34742 71286
rect 34370 71085 34742 71161
rect 34370 70960 34463 71026
rect 34370 70944 34447 70960
tri 34447 70944 34463 70960 nw
rect 34499 70927 34613 71085
rect 34649 70960 34742 71026
tri 34649 70944 34665 70960 ne
rect 34665 70944 34742 70960
rect 34482 70845 34630 70927
rect 34370 70812 34447 70828
tri 34447 70812 34463 70828 sw
rect 34370 70746 34463 70812
rect 34370 70644 34463 70710
rect 34370 70628 34447 70644
tri 34447 70628 34463 70644 nw
rect 34499 70611 34613 70845
tri 34649 70812 34665 70828 se
rect 34665 70812 34742 70828
rect 34649 70746 34742 70812
rect 34649 70644 34742 70710
tri 34649 70628 34665 70644 ne
rect 34665 70628 34742 70644
rect 34482 70529 34630 70611
rect 34370 70496 34447 70512
tri 34447 70496 34463 70512 sw
rect 34370 70430 34463 70496
rect 34499 70371 34613 70529
tri 34649 70496 34665 70512 se
rect 34665 70496 34742 70512
rect 34649 70430 34742 70496
rect 34370 70295 34742 70371
rect 34370 70170 34463 70236
rect 34370 70154 34447 70170
tri 34447 70154 34463 70170 nw
rect 34499 70137 34613 70295
rect 34649 70170 34742 70236
tri 34649 70154 34665 70170 ne
rect 34665 70154 34742 70170
rect 34482 70055 34630 70137
rect 34370 70022 34447 70038
tri 34447 70022 34463 70038 sw
rect 34370 69956 34463 70022
rect 34370 69854 34463 69920
rect 34370 69838 34447 69854
tri 34447 69838 34463 69854 nw
rect 34499 69821 34613 70055
tri 34649 70022 34665 70038 se
rect 34665 70022 34742 70038
rect 34649 69956 34742 70022
rect 34649 69854 34742 69920
tri 34649 69838 34665 69854 ne
rect 34665 69838 34742 69854
rect 34482 69739 34630 69821
rect 34370 69706 34447 69722
tri 34447 69706 34463 69722 sw
rect 34370 69640 34463 69706
rect 34499 69581 34613 69739
tri 34649 69706 34665 69722 se
rect 34665 69706 34742 69722
rect 34649 69640 34742 69706
rect 34370 69505 34742 69581
rect 34370 69380 34463 69446
rect 34370 69364 34447 69380
tri 34447 69364 34463 69380 nw
rect 34499 69347 34613 69505
rect 34649 69380 34742 69446
tri 34649 69364 34665 69380 ne
rect 34665 69364 34742 69380
rect 34482 69265 34630 69347
rect 34370 69232 34447 69248
tri 34447 69232 34463 69248 sw
rect 34370 69166 34463 69232
rect 34370 69064 34463 69130
rect 34370 69048 34447 69064
tri 34447 69048 34463 69064 nw
rect 34499 69031 34613 69265
tri 34649 69232 34665 69248 se
rect 34665 69232 34742 69248
rect 34649 69166 34742 69232
rect 34649 69064 34742 69130
tri 34649 69048 34665 69064 ne
rect 34665 69048 34742 69064
rect 34482 68949 34630 69031
rect 34370 68916 34447 68932
tri 34447 68916 34463 68932 sw
rect 34370 68850 34463 68916
rect 34499 68791 34613 68949
tri 34649 68916 34665 68932 se
rect 34665 68916 34742 68932
rect 34649 68850 34742 68916
rect 34370 68715 34742 68791
rect 34370 68590 34463 68656
rect 34370 68574 34447 68590
tri 34447 68574 34463 68590 nw
rect 34499 68557 34613 68715
rect 34649 68590 34742 68656
tri 34649 68574 34665 68590 ne
rect 34665 68574 34742 68590
rect 34482 68475 34630 68557
rect 34370 68442 34447 68458
tri 34447 68442 34463 68458 sw
rect 34370 68376 34463 68442
rect 34370 68274 34463 68340
rect 34370 68258 34447 68274
tri 34447 68258 34463 68274 nw
rect 34499 68241 34613 68475
tri 34649 68442 34665 68458 se
rect 34665 68442 34742 68458
rect 34649 68376 34742 68442
rect 34649 68274 34742 68340
tri 34649 68258 34665 68274 ne
rect 34665 68258 34742 68274
rect 34482 68159 34630 68241
rect 34370 68126 34447 68142
tri 34447 68126 34463 68142 sw
rect 34370 68060 34463 68126
rect 34499 68001 34613 68159
tri 34649 68126 34665 68142 se
rect 34665 68126 34742 68142
rect 34649 68060 34742 68126
rect 34370 67925 34742 68001
rect 34370 67800 34463 67866
rect 34370 67784 34447 67800
tri 34447 67784 34463 67800 nw
rect 34499 67767 34613 67925
rect 34649 67800 34742 67866
tri 34649 67784 34665 67800 ne
rect 34665 67784 34742 67800
rect 34482 67685 34630 67767
rect 34370 67652 34447 67668
tri 34447 67652 34463 67668 sw
rect 34370 67586 34463 67652
rect 34370 67484 34463 67550
rect 34370 67468 34447 67484
tri 34447 67468 34463 67484 nw
rect 34499 67451 34613 67685
tri 34649 67652 34665 67668 se
rect 34665 67652 34742 67668
rect 34649 67586 34742 67652
rect 34649 67484 34742 67550
tri 34649 67468 34665 67484 ne
rect 34665 67468 34742 67484
rect 34482 67369 34630 67451
rect 34370 67336 34447 67352
tri 34447 67336 34463 67352 sw
rect 34370 67270 34463 67336
rect 34499 67211 34613 67369
tri 34649 67336 34665 67352 se
rect 34665 67336 34742 67352
rect 34649 67270 34742 67336
rect 34370 67135 34742 67211
rect 34370 67010 34463 67076
rect 34370 66994 34447 67010
tri 34447 66994 34463 67010 nw
rect 34499 66977 34613 67135
rect 34649 67010 34742 67076
tri 34649 66994 34665 67010 ne
rect 34665 66994 34742 67010
rect 34482 66895 34630 66977
rect 34370 66862 34447 66878
tri 34447 66862 34463 66878 sw
rect 34370 66796 34463 66862
rect 34370 66694 34463 66760
rect 34370 66678 34447 66694
tri 34447 66678 34463 66694 nw
rect 34499 66661 34613 66895
tri 34649 66862 34665 66878 se
rect 34665 66862 34742 66878
rect 34649 66796 34742 66862
rect 34649 66694 34742 66760
tri 34649 66678 34665 66694 ne
rect 34665 66678 34742 66694
rect 34482 66579 34630 66661
rect 34370 66546 34447 66562
tri 34447 66546 34463 66562 sw
rect 34370 66480 34463 66546
rect 34499 66421 34613 66579
tri 34649 66546 34665 66562 se
rect 34665 66546 34742 66562
rect 34649 66480 34742 66546
rect 34370 66345 34742 66421
rect 34370 66220 34463 66286
rect 34370 66204 34447 66220
tri 34447 66204 34463 66220 nw
rect 34499 66187 34613 66345
rect 34649 66220 34742 66286
tri 34649 66204 34665 66220 ne
rect 34665 66204 34742 66220
rect 34482 66105 34630 66187
rect 34370 66072 34447 66088
tri 34447 66072 34463 66088 sw
rect 34370 66006 34463 66072
rect 34370 65904 34463 65970
rect 34370 65888 34447 65904
tri 34447 65888 34463 65904 nw
rect 34499 65871 34613 66105
tri 34649 66072 34665 66088 se
rect 34665 66072 34742 66088
rect 34649 66006 34742 66072
rect 34649 65904 34742 65970
tri 34649 65888 34665 65904 ne
rect 34665 65888 34742 65904
rect 34482 65789 34630 65871
rect 34370 65756 34447 65772
tri 34447 65756 34463 65772 sw
rect 34370 65690 34463 65756
rect 34499 65631 34613 65789
tri 34649 65756 34665 65772 se
rect 34665 65756 34742 65772
rect 34649 65690 34742 65756
rect 34370 65555 34742 65631
rect 34370 65430 34463 65496
rect 34370 65414 34447 65430
tri 34447 65414 34463 65430 nw
rect 34499 65397 34613 65555
rect 34649 65430 34742 65496
tri 34649 65414 34665 65430 ne
rect 34665 65414 34742 65430
rect 34482 65315 34630 65397
rect 34370 65282 34447 65298
tri 34447 65282 34463 65298 sw
rect 34370 65216 34463 65282
rect 34370 65114 34463 65180
rect 34370 65098 34447 65114
tri 34447 65098 34463 65114 nw
rect 34499 65081 34613 65315
tri 34649 65282 34665 65298 se
rect 34665 65282 34742 65298
rect 34649 65216 34742 65282
rect 34649 65114 34742 65180
tri 34649 65098 34665 65114 ne
rect 34665 65098 34742 65114
rect 34482 64999 34630 65081
rect 34370 64966 34447 64982
tri 34447 64966 34463 64982 sw
rect 34370 64900 34463 64966
rect 34499 64841 34613 64999
tri 34649 64966 34665 64982 se
rect 34665 64966 34742 64982
rect 34649 64900 34742 64966
rect 34370 64765 34742 64841
rect 34370 64640 34463 64706
rect 34370 64624 34447 64640
tri 34447 64624 34463 64640 nw
rect 34499 64607 34613 64765
rect 34649 64640 34742 64706
tri 34649 64624 34665 64640 ne
rect 34665 64624 34742 64640
rect 34482 64525 34630 64607
rect 34370 64492 34447 64508
tri 34447 64492 34463 64508 sw
rect 34370 64426 34463 64492
rect 34370 64324 34463 64390
rect 34370 64308 34447 64324
tri 34447 64308 34463 64324 nw
rect 34499 64291 34613 64525
tri 34649 64492 34665 64508 se
rect 34665 64492 34742 64508
rect 34649 64426 34742 64492
rect 34649 64324 34742 64390
tri 34649 64308 34665 64324 ne
rect 34665 64308 34742 64324
rect 34482 64209 34630 64291
rect 34370 64176 34447 64192
tri 34447 64176 34463 64192 sw
rect 34370 64110 34463 64176
rect 34499 64051 34613 64209
tri 34649 64176 34665 64192 se
rect 34665 64176 34742 64192
rect 34649 64110 34742 64176
rect 34370 63975 34742 64051
rect 34370 63850 34463 63916
rect 34370 63834 34447 63850
tri 34447 63834 34463 63850 nw
rect 34499 63817 34613 63975
rect 34649 63850 34742 63916
tri 34649 63834 34665 63850 ne
rect 34665 63834 34742 63850
rect 34482 63735 34630 63817
rect 34370 63702 34447 63718
tri 34447 63702 34463 63718 sw
rect 34370 63636 34463 63702
rect 34370 63534 34463 63600
rect 34370 63518 34447 63534
tri 34447 63518 34463 63534 nw
rect 34499 63501 34613 63735
tri 34649 63702 34665 63718 se
rect 34665 63702 34742 63718
rect 34649 63636 34742 63702
rect 34649 63534 34742 63600
tri 34649 63518 34665 63534 ne
rect 34665 63518 34742 63534
rect 34482 63419 34630 63501
rect 34370 63386 34447 63402
tri 34447 63386 34463 63402 sw
rect 34370 63320 34463 63386
rect 34499 63261 34613 63419
tri 34649 63386 34665 63402 se
rect 34665 63386 34742 63402
rect 34649 63320 34742 63386
rect 34370 63185 34742 63261
rect 34370 63060 34463 63126
rect 34370 63044 34447 63060
tri 34447 63044 34463 63060 nw
rect 34499 63027 34613 63185
rect 34649 63060 34742 63126
tri 34649 63044 34665 63060 ne
rect 34665 63044 34742 63060
rect 34482 62945 34630 63027
rect 34370 62912 34447 62928
tri 34447 62912 34463 62928 sw
rect 34370 62846 34463 62912
rect 34370 62744 34463 62810
rect 34370 62728 34447 62744
tri 34447 62728 34463 62744 nw
rect 34499 62711 34613 62945
tri 34649 62912 34665 62928 se
rect 34665 62912 34742 62928
rect 34649 62846 34742 62912
rect 34649 62744 34742 62810
tri 34649 62728 34665 62744 ne
rect 34665 62728 34742 62744
rect 34482 62629 34630 62711
rect 34370 62596 34447 62612
tri 34447 62596 34463 62612 sw
rect 34370 62530 34463 62596
rect 34499 62471 34613 62629
tri 34649 62596 34665 62612 se
rect 34665 62596 34742 62612
rect 34649 62530 34742 62596
rect 34370 62395 34742 62471
rect 34370 62270 34463 62336
rect 34370 62254 34447 62270
tri 34447 62254 34463 62270 nw
rect 34499 62237 34613 62395
rect 34649 62270 34742 62336
tri 34649 62254 34665 62270 ne
rect 34665 62254 34742 62270
rect 34482 62155 34630 62237
rect 34370 62122 34447 62138
tri 34447 62122 34463 62138 sw
rect 34370 62056 34463 62122
rect 34370 61954 34463 62020
rect 34370 61938 34447 61954
tri 34447 61938 34463 61954 nw
rect 34499 61921 34613 62155
tri 34649 62122 34665 62138 se
rect 34665 62122 34742 62138
rect 34649 62056 34742 62122
rect 34649 61954 34742 62020
tri 34649 61938 34665 61954 ne
rect 34665 61938 34742 61954
rect 34482 61839 34630 61921
rect 34370 61806 34447 61822
tri 34447 61806 34463 61822 sw
rect 34370 61740 34463 61806
rect 34499 61681 34613 61839
tri 34649 61806 34665 61822 se
rect 34665 61806 34742 61822
rect 34649 61740 34742 61806
rect 34370 61605 34742 61681
rect 34370 61480 34463 61546
rect 34370 61464 34447 61480
tri 34447 61464 34463 61480 nw
rect 34499 61447 34613 61605
rect 34649 61480 34742 61546
tri 34649 61464 34665 61480 ne
rect 34665 61464 34742 61480
rect 34482 61365 34630 61447
rect 34370 61332 34447 61348
tri 34447 61332 34463 61348 sw
rect 34370 61266 34463 61332
rect 34370 61164 34463 61230
rect 34370 61148 34447 61164
tri 34447 61148 34463 61164 nw
rect 34499 61131 34613 61365
tri 34649 61332 34665 61348 se
rect 34665 61332 34742 61348
rect 34649 61266 34742 61332
rect 34649 61164 34742 61230
tri 34649 61148 34665 61164 ne
rect 34665 61148 34742 61164
rect 34482 61049 34630 61131
rect 34370 61016 34447 61032
tri 34447 61016 34463 61032 sw
rect 34370 60950 34463 61016
rect 34499 60891 34613 61049
tri 34649 61016 34665 61032 se
rect 34665 61016 34742 61032
rect 34649 60950 34742 61016
rect 34370 60815 34742 60891
rect 34370 60690 34463 60756
rect 34370 60674 34447 60690
tri 34447 60674 34463 60690 nw
rect 34499 60657 34613 60815
rect 34649 60690 34742 60756
tri 34649 60674 34665 60690 ne
rect 34665 60674 34742 60690
rect 34482 60575 34630 60657
rect 34370 60542 34447 60558
tri 34447 60542 34463 60558 sw
rect 34370 60476 34463 60542
rect 34370 60374 34463 60440
rect 34370 60358 34447 60374
tri 34447 60358 34463 60374 nw
rect 34499 60341 34613 60575
tri 34649 60542 34665 60558 se
rect 34665 60542 34742 60558
rect 34649 60476 34742 60542
rect 34649 60374 34742 60440
tri 34649 60358 34665 60374 ne
rect 34665 60358 34742 60374
rect 34482 60259 34630 60341
rect 34370 60226 34447 60242
tri 34447 60226 34463 60242 sw
rect 34370 60160 34463 60226
rect 34499 60101 34613 60259
tri 34649 60226 34665 60242 se
rect 34665 60226 34742 60242
rect 34649 60160 34742 60226
rect 34370 60025 34742 60101
rect 34370 59900 34463 59966
rect 34370 59884 34447 59900
tri 34447 59884 34463 59900 nw
rect 34499 59867 34613 60025
rect 34649 59900 34742 59966
tri 34649 59884 34665 59900 ne
rect 34665 59884 34742 59900
rect 34482 59785 34630 59867
rect 34370 59752 34447 59768
tri 34447 59752 34463 59768 sw
rect 34370 59686 34463 59752
rect 34370 59584 34463 59650
rect 34370 59568 34447 59584
tri 34447 59568 34463 59584 nw
rect 34499 59551 34613 59785
tri 34649 59752 34665 59768 se
rect 34665 59752 34742 59768
rect 34649 59686 34742 59752
rect 34649 59584 34742 59650
tri 34649 59568 34665 59584 ne
rect 34665 59568 34742 59584
rect 34482 59469 34630 59551
rect 34370 59436 34447 59452
tri 34447 59436 34463 59452 sw
rect 34370 59370 34463 59436
rect 34499 59311 34613 59469
tri 34649 59436 34665 59452 se
rect 34665 59436 34742 59452
rect 34649 59370 34742 59436
rect 34370 59235 34742 59311
rect 34370 59110 34463 59176
rect 34370 59094 34447 59110
tri 34447 59094 34463 59110 nw
rect 34499 59077 34613 59235
rect 34649 59110 34742 59176
tri 34649 59094 34665 59110 ne
rect 34665 59094 34742 59110
rect 34482 58995 34630 59077
rect 34370 58962 34447 58978
tri 34447 58962 34463 58978 sw
rect 34370 58896 34463 58962
rect 34370 58794 34463 58860
rect 34370 58778 34447 58794
tri 34447 58778 34463 58794 nw
rect 34499 58761 34613 58995
tri 34649 58962 34665 58978 se
rect 34665 58962 34742 58978
rect 34649 58896 34742 58962
rect 34649 58794 34742 58860
tri 34649 58778 34665 58794 ne
rect 34665 58778 34742 58794
rect 34482 58679 34630 58761
rect 34370 58646 34447 58662
tri 34447 58646 34463 58662 sw
rect 34370 58580 34463 58646
rect 34499 58521 34613 58679
tri 34649 58646 34665 58662 se
rect 34665 58646 34742 58662
rect 34649 58580 34742 58646
rect 34370 58445 34742 58521
rect 34370 58320 34463 58386
rect 34370 58304 34447 58320
tri 34447 58304 34463 58320 nw
rect 34499 58287 34613 58445
rect 34649 58320 34742 58386
tri 34649 58304 34665 58320 ne
rect 34665 58304 34742 58320
rect 34482 58205 34630 58287
rect 34370 58172 34447 58188
tri 34447 58172 34463 58188 sw
rect 34370 58106 34463 58172
rect 34370 58004 34463 58070
rect 34370 57988 34447 58004
tri 34447 57988 34463 58004 nw
rect 34499 57971 34613 58205
tri 34649 58172 34665 58188 se
rect 34665 58172 34742 58188
rect 34649 58106 34742 58172
rect 34649 58004 34742 58070
tri 34649 57988 34665 58004 ne
rect 34665 57988 34742 58004
rect 34482 57889 34630 57971
rect 34370 57856 34447 57872
tri 34447 57856 34463 57872 sw
rect 34370 57790 34463 57856
rect 34499 57731 34613 57889
tri 34649 57856 34665 57872 se
rect 34665 57856 34742 57872
rect 34649 57790 34742 57856
rect 34370 57655 34742 57731
rect 34370 57530 34463 57596
rect 34370 57514 34447 57530
tri 34447 57514 34463 57530 nw
rect 34499 57497 34613 57655
rect 34649 57530 34742 57596
tri 34649 57514 34665 57530 ne
rect 34665 57514 34742 57530
rect 34482 57415 34630 57497
rect 34370 57382 34447 57398
tri 34447 57382 34463 57398 sw
rect 34370 57316 34463 57382
rect 34370 57214 34463 57280
rect 34370 57198 34447 57214
tri 34447 57198 34463 57214 nw
rect 34499 57181 34613 57415
tri 34649 57382 34665 57398 se
rect 34665 57382 34742 57398
rect 34649 57316 34742 57382
rect 34649 57214 34742 57280
tri 34649 57198 34665 57214 ne
rect 34665 57198 34742 57214
rect 34482 57099 34630 57181
rect 34370 57066 34447 57082
tri 34447 57066 34463 57082 sw
rect 34370 57000 34463 57066
rect 34499 56941 34613 57099
tri 34649 57066 34665 57082 se
rect 34665 57066 34742 57082
rect 34649 57000 34742 57066
rect 34370 56865 34742 56941
rect 34370 56740 34463 56806
rect 34370 56724 34447 56740
tri 34447 56724 34463 56740 nw
rect 34499 56707 34613 56865
rect 34649 56740 34742 56806
tri 34649 56724 34665 56740 ne
rect 34665 56724 34742 56740
rect 34482 56625 34630 56707
rect 34370 56592 34447 56608
tri 34447 56592 34463 56608 sw
rect 34370 56526 34463 56592
rect 34370 56424 34463 56490
rect 34370 56408 34447 56424
tri 34447 56408 34463 56424 nw
rect 34499 56391 34613 56625
tri 34649 56592 34665 56608 se
rect 34665 56592 34742 56608
rect 34649 56526 34742 56592
rect 34649 56424 34742 56490
tri 34649 56408 34665 56424 ne
rect 34665 56408 34742 56424
rect 34482 56309 34630 56391
rect 34370 56276 34447 56292
tri 34447 56276 34463 56292 sw
rect 34370 56210 34463 56276
rect 34499 56151 34613 56309
tri 34649 56276 34665 56292 se
rect 34665 56276 34742 56292
rect 34649 56210 34742 56276
rect 34370 56075 34742 56151
rect 34370 55950 34463 56016
rect 34370 55934 34447 55950
tri 34447 55934 34463 55950 nw
rect 34499 55917 34613 56075
rect 34649 55950 34742 56016
tri 34649 55934 34665 55950 ne
rect 34665 55934 34742 55950
rect 34482 55835 34630 55917
rect 34370 55802 34447 55818
tri 34447 55802 34463 55818 sw
rect 34370 55736 34463 55802
rect 34370 55634 34463 55700
rect 34370 55618 34447 55634
tri 34447 55618 34463 55634 nw
rect 34499 55601 34613 55835
tri 34649 55802 34665 55818 se
rect 34665 55802 34742 55818
rect 34649 55736 34742 55802
rect 34649 55634 34742 55700
tri 34649 55618 34665 55634 ne
rect 34665 55618 34742 55634
rect 34482 55519 34630 55601
rect 34370 55486 34447 55502
tri 34447 55486 34463 55502 sw
rect 34370 55420 34463 55486
rect 34499 55361 34613 55519
tri 34649 55486 34665 55502 se
rect 34665 55486 34742 55502
rect 34649 55420 34742 55486
rect 34370 55285 34742 55361
rect 34370 55160 34463 55226
rect 34370 55144 34447 55160
tri 34447 55144 34463 55160 nw
rect 34499 55127 34613 55285
rect 34649 55160 34742 55226
tri 34649 55144 34665 55160 ne
rect 34665 55144 34742 55160
rect 34482 55045 34630 55127
rect 34370 55012 34447 55028
tri 34447 55012 34463 55028 sw
rect 34370 54946 34463 55012
rect 34370 54844 34463 54910
rect 34370 54828 34447 54844
tri 34447 54828 34463 54844 nw
rect 34499 54811 34613 55045
tri 34649 55012 34665 55028 se
rect 34665 55012 34742 55028
rect 34649 54946 34742 55012
rect 34649 54844 34742 54910
tri 34649 54828 34665 54844 ne
rect 34665 54828 34742 54844
rect 34482 54729 34630 54811
rect 34370 54696 34447 54712
tri 34447 54696 34463 54712 sw
rect 34370 54630 34463 54696
rect 34499 54571 34613 54729
tri 34649 54696 34665 54712 se
rect 34665 54696 34742 54712
rect 34649 54630 34742 54696
rect 34370 54495 34742 54571
rect 34370 54370 34463 54436
rect 34370 54354 34447 54370
tri 34447 54354 34463 54370 nw
rect 34499 54337 34613 54495
rect 34649 54370 34742 54436
tri 34649 54354 34665 54370 ne
rect 34665 54354 34742 54370
rect 34482 54255 34630 54337
rect 34370 54222 34447 54238
tri 34447 54222 34463 54238 sw
rect 34370 54156 34463 54222
rect 34370 54054 34463 54120
rect 34370 54038 34447 54054
tri 34447 54038 34463 54054 nw
rect 34499 54021 34613 54255
tri 34649 54222 34665 54238 se
rect 34665 54222 34742 54238
rect 34649 54156 34742 54222
rect 34649 54054 34742 54120
tri 34649 54038 34665 54054 ne
rect 34665 54038 34742 54054
rect 34482 53939 34630 54021
rect 34370 53906 34447 53922
tri 34447 53906 34463 53922 sw
rect 34370 53840 34463 53906
rect 34499 53781 34613 53939
tri 34649 53906 34665 53922 se
rect 34665 53906 34742 53922
rect 34649 53840 34742 53906
rect 34370 53705 34742 53781
rect 34370 53580 34463 53646
rect 34370 53564 34447 53580
tri 34447 53564 34463 53580 nw
rect 34499 53547 34613 53705
rect 34649 53580 34742 53646
tri 34649 53564 34665 53580 ne
rect 34665 53564 34742 53580
rect 34482 53465 34630 53547
rect 34370 53432 34447 53448
tri 34447 53432 34463 53448 sw
rect 34370 53366 34463 53432
rect 34370 53264 34463 53330
rect 34370 53248 34447 53264
tri 34447 53248 34463 53264 nw
rect 34499 53231 34613 53465
tri 34649 53432 34665 53448 se
rect 34665 53432 34742 53448
rect 34649 53366 34742 53432
rect 34649 53264 34742 53330
tri 34649 53248 34665 53264 ne
rect 34665 53248 34742 53264
rect 34482 53149 34630 53231
rect 34370 53116 34447 53132
tri 34447 53116 34463 53132 sw
rect 34370 53050 34463 53116
rect 34499 52991 34613 53149
tri 34649 53116 34665 53132 se
rect 34665 53116 34742 53132
rect 34649 53050 34742 53116
rect 34370 52915 34742 52991
rect 34370 52790 34463 52856
rect 34370 52774 34447 52790
tri 34447 52774 34463 52790 nw
rect 34499 52757 34613 52915
rect 34649 52790 34742 52856
tri 34649 52774 34665 52790 ne
rect 34665 52774 34742 52790
rect 34482 52675 34630 52757
rect 34370 52642 34447 52658
tri 34447 52642 34463 52658 sw
rect 34370 52576 34463 52642
rect 34370 52474 34463 52540
rect 34370 52458 34447 52474
tri 34447 52458 34463 52474 nw
rect 34499 52441 34613 52675
tri 34649 52642 34665 52658 se
rect 34665 52642 34742 52658
rect 34649 52576 34742 52642
rect 34649 52474 34742 52540
tri 34649 52458 34665 52474 ne
rect 34665 52458 34742 52474
rect 34482 52359 34630 52441
rect 34370 52326 34447 52342
tri 34447 52326 34463 52342 sw
rect 34370 52260 34463 52326
rect 34499 52201 34613 52359
tri 34649 52326 34665 52342 se
rect 34665 52326 34742 52342
rect 34649 52260 34742 52326
rect 34370 52125 34742 52201
rect 34370 52000 34463 52066
rect 34370 51984 34447 52000
tri 34447 51984 34463 52000 nw
rect 34499 51967 34613 52125
rect 34649 52000 34742 52066
tri 34649 51984 34665 52000 ne
rect 34665 51984 34742 52000
rect 34482 51885 34630 51967
rect 34370 51852 34447 51868
tri 34447 51852 34463 51868 sw
rect 34370 51786 34463 51852
rect 34370 51684 34463 51750
rect 34370 51668 34447 51684
tri 34447 51668 34463 51684 nw
rect 34499 51651 34613 51885
tri 34649 51852 34665 51868 se
rect 34665 51852 34742 51868
rect 34649 51786 34742 51852
rect 34649 51684 34742 51750
tri 34649 51668 34665 51684 ne
rect 34665 51668 34742 51684
rect 34482 51569 34630 51651
rect 34370 51536 34447 51552
tri 34447 51536 34463 51552 sw
rect 34370 51470 34463 51536
rect 34499 51411 34613 51569
tri 34649 51536 34665 51552 se
rect 34665 51536 34742 51552
rect 34649 51470 34742 51536
rect 34370 51335 34742 51411
rect 34370 51210 34463 51276
rect 34370 51194 34447 51210
tri 34447 51194 34463 51210 nw
rect 34499 51177 34613 51335
rect 34649 51210 34742 51276
tri 34649 51194 34665 51210 ne
rect 34665 51194 34742 51210
rect 34482 51095 34630 51177
rect 34370 51062 34447 51078
tri 34447 51062 34463 51078 sw
rect 34370 50996 34463 51062
rect 34370 50894 34463 50960
rect 34370 50878 34447 50894
tri 34447 50878 34463 50894 nw
rect 34499 50861 34613 51095
tri 34649 51062 34665 51078 se
rect 34665 51062 34742 51078
rect 34649 50996 34742 51062
rect 34649 50894 34742 50960
tri 34649 50878 34665 50894 ne
rect 34665 50878 34742 50894
rect 34482 50779 34630 50861
rect 34370 50746 34447 50762
tri 34447 50746 34463 50762 sw
rect 34370 50680 34463 50746
rect 34499 50621 34613 50779
tri 34649 50746 34665 50762 se
rect 34665 50746 34742 50762
rect 34649 50680 34742 50746
rect 34370 50545 34742 50621
rect 34370 50420 34463 50486
rect 34370 50404 34447 50420
tri 34447 50404 34463 50420 nw
rect 34499 50387 34613 50545
rect 34649 50420 34742 50486
tri 34649 50404 34665 50420 ne
rect 34665 50404 34742 50420
rect 34482 50305 34630 50387
rect 34370 50272 34447 50288
tri 34447 50272 34463 50288 sw
rect 34370 50206 34463 50272
rect 34370 50104 34463 50170
rect 34370 50088 34447 50104
tri 34447 50088 34463 50104 nw
rect 34499 50071 34613 50305
tri 34649 50272 34665 50288 se
rect 34665 50272 34742 50288
rect 34649 50206 34742 50272
rect 34649 50104 34742 50170
tri 34649 50088 34665 50104 ne
rect 34665 50088 34742 50104
rect 34482 49989 34630 50071
rect 34370 49956 34447 49972
tri 34447 49956 34463 49972 sw
rect 34370 49890 34463 49956
rect 34499 49831 34613 49989
tri 34649 49956 34665 49972 se
rect 34665 49956 34742 49972
rect 34649 49890 34742 49956
rect 34370 49755 34742 49831
rect 34370 49630 34463 49696
rect 34370 49614 34447 49630
tri 34447 49614 34463 49630 nw
rect 34499 49597 34613 49755
rect 34649 49630 34742 49696
tri 34649 49614 34665 49630 ne
rect 34665 49614 34742 49630
rect 34482 49515 34630 49597
rect 34370 49482 34447 49498
tri 34447 49482 34463 49498 sw
rect 34370 49416 34463 49482
rect 34370 49314 34463 49380
rect 34370 49298 34447 49314
tri 34447 49298 34463 49314 nw
rect 34499 49281 34613 49515
tri 34649 49482 34665 49498 se
rect 34665 49482 34742 49498
rect 34649 49416 34742 49482
rect 34649 49314 34742 49380
tri 34649 49298 34665 49314 ne
rect 34665 49298 34742 49314
rect 34482 49199 34630 49281
rect 34370 49166 34447 49182
tri 34447 49166 34463 49182 sw
rect 34370 49100 34463 49166
rect 34499 49041 34613 49199
tri 34649 49166 34665 49182 se
rect 34665 49166 34742 49182
rect 34649 49100 34742 49166
rect 34370 48965 34742 49041
rect 34370 48840 34463 48906
rect 34370 48824 34447 48840
tri 34447 48824 34463 48840 nw
rect 34499 48807 34613 48965
rect 34649 48840 34742 48906
tri 34649 48824 34665 48840 ne
rect 34665 48824 34742 48840
rect 34482 48725 34630 48807
rect 34370 48692 34447 48708
tri 34447 48692 34463 48708 sw
rect 34370 48626 34463 48692
rect 34370 48524 34463 48590
rect 34370 48508 34447 48524
tri 34447 48508 34463 48524 nw
rect 34499 48491 34613 48725
tri 34649 48692 34665 48708 se
rect 34665 48692 34742 48708
rect 34649 48626 34742 48692
rect 34649 48524 34742 48590
tri 34649 48508 34665 48524 ne
rect 34665 48508 34742 48524
rect 34482 48409 34630 48491
rect 34370 48376 34447 48392
tri 34447 48376 34463 48392 sw
rect 34370 48310 34463 48376
rect 34499 48251 34613 48409
tri 34649 48376 34665 48392 se
rect 34665 48376 34742 48392
rect 34649 48310 34742 48376
rect 34370 48175 34742 48251
rect 34370 48050 34463 48116
rect 34370 48034 34447 48050
tri 34447 48034 34463 48050 nw
rect 34499 48017 34613 48175
rect 34649 48050 34742 48116
tri 34649 48034 34665 48050 ne
rect 34665 48034 34742 48050
rect 34482 47935 34630 48017
rect 34370 47902 34447 47918
tri 34447 47902 34463 47918 sw
rect 34370 47836 34463 47902
rect 34370 47734 34463 47800
rect 34370 47718 34447 47734
tri 34447 47718 34463 47734 nw
rect 34499 47701 34613 47935
tri 34649 47902 34665 47918 se
rect 34665 47902 34742 47918
rect 34649 47836 34742 47902
rect 34649 47734 34742 47800
tri 34649 47718 34665 47734 ne
rect 34665 47718 34742 47734
rect 34482 47619 34630 47701
rect 34370 47586 34447 47602
tri 34447 47586 34463 47602 sw
rect 34370 47520 34463 47586
rect 34499 47461 34613 47619
tri 34649 47586 34665 47602 se
rect 34665 47586 34742 47602
rect 34649 47520 34742 47586
rect 34370 47385 34742 47461
rect 34370 47260 34463 47326
rect 34370 47244 34447 47260
tri 34447 47244 34463 47260 nw
rect 34499 47227 34613 47385
rect 34649 47260 34742 47326
tri 34649 47244 34665 47260 ne
rect 34665 47244 34742 47260
rect 34482 47145 34630 47227
rect 34370 47112 34447 47128
tri 34447 47112 34463 47128 sw
rect 34370 47046 34463 47112
rect 34370 46944 34463 47010
rect 34370 46928 34447 46944
tri 34447 46928 34463 46944 nw
rect 34499 46911 34613 47145
tri 34649 47112 34665 47128 se
rect 34665 47112 34742 47128
rect 34649 47046 34742 47112
rect 34649 46944 34742 47010
tri 34649 46928 34665 46944 ne
rect 34665 46928 34742 46944
rect 34482 46829 34630 46911
rect 34370 46796 34447 46812
tri 34447 46796 34463 46812 sw
rect 34370 46730 34463 46796
rect 34499 46671 34613 46829
tri 34649 46796 34665 46812 se
rect 34665 46796 34742 46812
rect 34649 46730 34742 46796
rect 34370 46595 34742 46671
rect 34370 46470 34463 46536
rect 34370 46454 34447 46470
tri 34447 46454 34463 46470 nw
rect 34499 46437 34613 46595
rect 34649 46470 34742 46536
tri 34649 46454 34665 46470 ne
rect 34665 46454 34742 46470
rect 34482 46355 34630 46437
rect 34370 46322 34447 46338
tri 34447 46322 34463 46338 sw
rect 34370 46256 34463 46322
rect 34370 46154 34463 46220
rect 34370 46138 34447 46154
tri 34447 46138 34463 46154 nw
rect 34499 46121 34613 46355
tri 34649 46322 34665 46338 se
rect 34665 46322 34742 46338
rect 34649 46256 34742 46322
rect 34649 46154 34742 46220
tri 34649 46138 34665 46154 ne
rect 34665 46138 34742 46154
rect 34482 46039 34630 46121
rect 34370 46006 34447 46022
tri 34447 46006 34463 46022 sw
rect 34370 45940 34463 46006
rect 34499 45881 34613 46039
tri 34649 46006 34665 46022 se
rect 34665 46006 34742 46022
rect 34649 45940 34742 46006
rect 34370 45805 34742 45881
rect 34370 45680 34463 45746
rect 34370 45664 34447 45680
tri 34447 45664 34463 45680 nw
rect 34499 45647 34613 45805
rect 34649 45680 34742 45746
tri 34649 45664 34665 45680 ne
rect 34665 45664 34742 45680
rect 34482 45565 34630 45647
rect 34370 45532 34447 45548
tri 34447 45532 34463 45548 sw
rect 34370 45466 34463 45532
rect 34370 45364 34463 45430
rect 34370 45348 34447 45364
tri 34447 45348 34463 45364 nw
rect 34499 45331 34613 45565
tri 34649 45532 34665 45548 se
rect 34665 45532 34742 45548
rect 34649 45466 34742 45532
rect 34649 45364 34742 45430
tri 34649 45348 34665 45364 ne
rect 34665 45348 34742 45364
rect 34482 45249 34630 45331
rect 34370 45216 34447 45232
tri 34447 45216 34463 45232 sw
rect 34370 45150 34463 45216
rect 34499 45091 34613 45249
tri 34649 45216 34665 45232 se
rect 34665 45216 34742 45232
rect 34649 45150 34742 45216
rect 34370 45015 34742 45091
rect 34370 44890 34463 44956
rect 34370 44874 34447 44890
tri 34447 44874 34463 44890 nw
rect 34499 44857 34613 45015
rect 34649 44890 34742 44956
tri 34649 44874 34665 44890 ne
rect 34665 44874 34742 44890
rect 34482 44775 34630 44857
rect 34370 44742 34447 44758
tri 34447 44742 34463 44758 sw
rect 34370 44676 34463 44742
rect 34370 44574 34463 44640
rect 34370 44558 34447 44574
tri 34447 44558 34463 44574 nw
rect 34499 44541 34613 44775
tri 34649 44742 34665 44758 se
rect 34665 44742 34742 44758
rect 34649 44676 34742 44742
rect 34649 44574 34742 44640
tri 34649 44558 34665 44574 ne
rect 34665 44558 34742 44574
rect 34482 44459 34630 44541
rect 34370 44426 34447 44442
tri 34447 44426 34463 44442 sw
rect 34370 44360 34463 44426
rect 34499 44301 34613 44459
tri 34649 44426 34665 44442 se
rect 34665 44426 34742 44442
rect 34649 44360 34742 44426
rect 34370 44225 34742 44301
rect 34370 44100 34463 44166
rect 34370 44084 34447 44100
tri 34447 44084 34463 44100 nw
rect 34499 44067 34613 44225
rect 34649 44100 34742 44166
tri 34649 44084 34665 44100 ne
rect 34665 44084 34742 44100
rect 34482 43985 34630 44067
rect 34370 43952 34447 43968
tri 34447 43952 34463 43968 sw
rect 34370 43886 34463 43952
rect 34370 43784 34463 43850
rect 34370 43768 34447 43784
tri 34447 43768 34463 43784 nw
rect 34499 43751 34613 43985
tri 34649 43952 34665 43968 se
rect 34665 43952 34742 43968
rect 34649 43886 34742 43952
rect 34649 43784 34742 43850
tri 34649 43768 34665 43784 ne
rect 34665 43768 34742 43784
rect 34482 43669 34630 43751
rect 34370 43636 34447 43652
tri 34447 43636 34463 43652 sw
rect 34370 43570 34463 43636
rect 34499 43511 34613 43669
tri 34649 43636 34665 43652 se
rect 34665 43636 34742 43652
rect 34649 43570 34742 43636
rect 34370 43435 34742 43511
rect 34370 43310 34463 43376
rect 34370 43294 34447 43310
tri 34447 43294 34463 43310 nw
rect 34499 43277 34613 43435
rect 34649 43310 34742 43376
tri 34649 43294 34665 43310 ne
rect 34665 43294 34742 43310
rect 34482 43195 34630 43277
rect 34370 43162 34447 43178
tri 34447 43162 34463 43178 sw
rect 34370 43096 34463 43162
rect 34370 42994 34463 43060
rect 34370 42978 34447 42994
tri 34447 42978 34463 42994 nw
rect 34499 42961 34613 43195
tri 34649 43162 34665 43178 se
rect 34665 43162 34742 43178
rect 34649 43096 34742 43162
rect 34649 42994 34742 43060
tri 34649 42978 34665 42994 ne
rect 34665 42978 34742 42994
rect 34482 42879 34630 42961
rect 34370 42846 34447 42862
tri 34447 42846 34463 42862 sw
rect 34370 42780 34463 42846
rect 34499 42721 34613 42879
tri 34649 42846 34665 42862 se
rect 34665 42846 34742 42862
rect 34649 42780 34742 42846
rect 34370 42645 34742 42721
rect 34370 42520 34463 42586
rect 34370 42504 34447 42520
tri 34447 42504 34463 42520 nw
rect 34499 42487 34613 42645
rect 34649 42520 34742 42586
tri 34649 42504 34665 42520 ne
rect 34665 42504 34742 42520
rect 34482 42405 34630 42487
rect 34370 42372 34447 42388
tri 34447 42372 34463 42388 sw
rect 34370 42306 34463 42372
rect 34370 42204 34463 42270
rect 34370 42188 34447 42204
tri 34447 42188 34463 42204 nw
rect 34499 42171 34613 42405
tri 34649 42372 34665 42388 se
rect 34665 42372 34742 42388
rect 34649 42306 34742 42372
rect 34649 42204 34742 42270
tri 34649 42188 34665 42204 ne
rect 34665 42188 34742 42204
rect 34482 42089 34630 42171
rect 34370 42056 34447 42072
tri 34447 42056 34463 42072 sw
rect 34370 41990 34463 42056
rect 34499 41931 34613 42089
tri 34649 42056 34665 42072 se
rect 34665 42056 34742 42072
rect 34649 41990 34742 42056
rect 34370 41855 34742 41931
rect 34370 41730 34463 41796
rect 34370 41714 34447 41730
tri 34447 41714 34463 41730 nw
rect 34499 41697 34613 41855
rect 34649 41730 34742 41796
tri 34649 41714 34665 41730 ne
rect 34665 41714 34742 41730
rect 34482 41615 34630 41697
rect 34370 41582 34447 41598
tri 34447 41582 34463 41598 sw
rect 34370 41516 34463 41582
rect 34370 41414 34463 41480
rect 34370 41398 34447 41414
tri 34447 41398 34463 41414 nw
rect 34499 41381 34613 41615
tri 34649 41582 34665 41598 se
rect 34665 41582 34742 41598
rect 34649 41516 34742 41582
rect 34649 41414 34742 41480
tri 34649 41398 34665 41414 ne
rect 34665 41398 34742 41414
rect 34482 41299 34630 41381
rect 34370 41266 34447 41282
tri 34447 41266 34463 41282 sw
rect 34370 41200 34463 41266
rect 34499 41141 34613 41299
tri 34649 41266 34665 41282 se
rect 34665 41266 34742 41282
rect 34649 41200 34742 41266
rect 34370 41065 34742 41141
rect 34370 40940 34463 41006
rect 34370 40924 34447 40940
tri 34447 40924 34463 40940 nw
rect 34499 40907 34613 41065
rect 34649 40940 34742 41006
tri 34649 40924 34665 40940 ne
rect 34665 40924 34742 40940
rect 34482 40825 34630 40907
rect 34370 40792 34447 40808
tri 34447 40792 34463 40808 sw
rect 34370 40726 34463 40792
rect 34370 40624 34463 40690
rect 34370 40608 34447 40624
tri 34447 40608 34463 40624 nw
rect 34499 40591 34613 40825
tri 34649 40792 34665 40808 se
rect 34665 40792 34742 40808
rect 34649 40726 34742 40792
rect 34649 40624 34742 40690
tri 34649 40608 34665 40624 ne
rect 34665 40608 34742 40624
rect 34482 40509 34630 40591
rect 34370 40476 34447 40492
tri 34447 40476 34463 40492 sw
rect 34370 40410 34463 40476
rect 34499 40351 34613 40509
tri 34649 40476 34665 40492 se
rect 34665 40476 34742 40492
rect 34649 40410 34742 40476
rect 34370 40275 34742 40351
rect 34370 40150 34463 40216
rect 34370 40134 34447 40150
tri 34447 40134 34463 40150 nw
rect 34499 40117 34613 40275
rect 34649 40150 34742 40216
tri 34649 40134 34665 40150 ne
rect 34665 40134 34742 40150
rect 34482 40035 34630 40117
rect 34370 40002 34447 40018
tri 34447 40002 34463 40018 sw
rect 34370 39936 34463 40002
rect 34370 39834 34463 39900
rect 34370 39818 34447 39834
tri 34447 39818 34463 39834 nw
rect 34499 39801 34613 40035
tri 34649 40002 34665 40018 se
rect 34665 40002 34742 40018
rect 34649 39936 34742 40002
rect 34649 39834 34742 39900
tri 34649 39818 34665 39834 ne
rect 34665 39818 34742 39834
rect 34482 39719 34630 39801
rect 34370 39686 34447 39702
tri 34447 39686 34463 39702 sw
rect 34370 39620 34463 39686
rect 34499 39561 34613 39719
tri 34649 39686 34665 39702 se
rect 34665 39686 34742 39702
rect 34649 39620 34742 39686
rect 34370 39485 34742 39561
rect 34370 39360 34463 39426
rect 34370 39344 34447 39360
tri 34447 39344 34463 39360 nw
rect 34499 39327 34613 39485
rect 34649 39360 34742 39426
tri 34649 39344 34665 39360 ne
rect 34665 39344 34742 39360
rect 34482 39245 34630 39327
rect 34370 39212 34447 39228
tri 34447 39212 34463 39228 sw
rect 34370 39146 34463 39212
rect 34370 39044 34463 39110
rect 34370 39028 34447 39044
tri 34447 39028 34463 39044 nw
rect 34499 39011 34613 39245
tri 34649 39212 34665 39228 se
rect 34665 39212 34742 39228
rect 34649 39146 34742 39212
rect 34649 39044 34742 39110
tri 34649 39028 34665 39044 ne
rect 34665 39028 34742 39044
rect 34482 38929 34630 39011
rect 34370 38896 34447 38912
tri 34447 38896 34463 38912 sw
rect 34370 38830 34463 38896
rect 34499 38771 34613 38929
tri 34649 38896 34665 38912 se
rect 34665 38896 34742 38912
rect 34649 38830 34742 38896
rect 34370 38695 34742 38771
rect 34370 38570 34463 38636
rect 34370 38554 34447 38570
tri 34447 38554 34463 38570 nw
rect 34499 38537 34613 38695
rect 34649 38570 34742 38636
tri 34649 38554 34665 38570 ne
rect 34665 38554 34742 38570
rect 34482 38455 34630 38537
rect 34370 38422 34447 38438
tri 34447 38422 34463 38438 sw
rect 34370 38356 34463 38422
rect 34370 38254 34463 38320
rect 34370 38238 34447 38254
tri 34447 38238 34463 38254 nw
rect 34499 38221 34613 38455
tri 34649 38422 34665 38438 se
rect 34665 38422 34742 38438
rect 34649 38356 34742 38422
rect 34649 38254 34742 38320
tri 34649 38238 34665 38254 ne
rect 34665 38238 34742 38254
rect 34482 38139 34630 38221
rect 34370 38106 34447 38122
tri 34447 38106 34463 38122 sw
rect 34370 38040 34463 38106
rect 34499 37981 34613 38139
tri 34649 38106 34665 38122 se
rect 34665 38106 34742 38122
rect 34649 38040 34742 38106
rect 34370 37905 34742 37981
rect 34370 37780 34463 37846
rect 34370 37764 34447 37780
tri 34447 37764 34463 37780 nw
rect 34499 37747 34613 37905
rect 34649 37780 34742 37846
tri 34649 37764 34665 37780 ne
rect 34665 37764 34742 37780
rect 34482 37665 34630 37747
rect 34370 37632 34447 37648
tri 34447 37632 34463 37648 sw
rect 34370 37566 34463 37632
rect 34370 37464 34463 37530
rect 34370 37448 34447 37464
tri 34447 37448 34463 37464 nw
rect 34499 37431 34613 37665
tri 34649 37632 34665 37648 se
rect 34665 37632 34742 37648
rect 34649 37566 34742 37632
rect 34649 37464 34742 37530
tri 34649 37448 34665 37464 ne
rect 34665 37448 34742 37464
rect 34482 37349 34630 37431
rect 34370 37316 34447 37332
tri 34447 37316 34463 37332 sw
rect 34370 37250 34463 37316
rect 34499 37191 34613 37349
tri 34649 37316 34665 37332 se
rect 34665 37316 34742 37332
rect 34649 37250 34742 37316
rect 34370 37115 34742 37191
rect 34370 36990 34463 37056
rect 34370 36974 34447 36990
tri 34447 36974 34463 36990 nw
rect 34499 36957 34613 37115
rect 34649 36990 34742 37056
tri 34649 36974 34665 36990 ne
rect 34665 36974 34742 36990
rect 34482 36875 34630 36957
rect 34370 36842 34447 36858
tri 34447 36842 34463 36858 sw
rect 34370 36776 34463 36842
rect 34370 36674 34463 36740
rect 34370 36658 34447 36674
tri 34447 36658 34463 36674 nw
rect 34499 36641 34613 36875
tri 34649 36842 34665 36858 se
rect 34665 36842 34742 36858
rect 34649 36776 34742 36842
rect 34649 36674 34742 36740
tri 34649 36658 34665 36674 ne
rect 34665 36658 34742 36674
rect 34482 36559 34630 36641
rect 34370 36526 34447 36542
tri 34447 36526 34463 36542 sw
rect 34370 36460 34463 36526
rect 34499 36401 34613 36559
tri 34649 36526 34665 36542 se
rect 34665 36526 34742 36542
rect 34649 36460 34742 36526
rect 34370 36325 34742 36401
rect 34370 36200 34463 36266
rect 34370 36184 34447 36200
tri 34447 36184 34463 36200 nw
rect 34499 36167 34613 36325
rect 34649 36200 34742 36266
tri 34649 36184 34665 36200 ne
rect 34665 36184 34742 36200
rect 34482 36085 34630 36167
rect 34370 36052 34447 36068
tri 34447 36052 34463 36068 sw
rect 34370 35986 34463 36052
rect 34370 35884 34463 35950
rect 34370 35868 34447 35884
tri 34447 35868 34463 35884 nw
rect 34499 35851 34613 36085
tri 34649 36052 34665 36068 se
rect 34665 36052 34742 36068
rect 34649 35986 34742 36052
rect 34649 35884 34742 35950
tri 34649 35868 34665 35884 ne
rect 34665 35868 34742 35884
rect 34482 35769 34630 35851
rect 34370 35736 34447 35752
tri 34447 35736 34463 35752 sw
rect 34370 35670 34463 35736
rect 34499 35611 34613 35769
tri 34649 35736 34665 35752 se
rect 34665 35736 34742 35752
rect 34649 35670 34742 35736
rect 34370 35535 34742 35611
rect 34370 35410 34463 35476
rect 34370 35394 34447 35410
tri 34447 35394 34463 35410 nw
rect 34499 35377 34613 35535
rect 34649 35410 34742 35476
tri 34649 35394 34665 35410 ne
rect 34665 35394 34742 35410
rect 34482 35295 34630 35377
rect 34370 35262 34447 35278
tri 34447 35262 34463 35278 sw
rect 34370 35196 34463 35262
rect 34370 35094 34463 35160
rect 34370 35078 34447 35094
tri 34447 35078 34463 35094 nw
rect 34499 35061 34613 35295
tri 34649 35262 34665 35278 se
rect 34665 35262 34742 35278
rect 34649 35196 34742 35262
rect 34649 35094 34742 35160
tri 34649 35078 34665 35094 ne
rect 34665 35078 34742 35094
rect 34482 34979 34630 35061
rect 34370 34946 34447 34962
tri 34447 34946 34463 34962 sw
rect 34370 34880 34463 34946
rect 34499 34821 34613 34979
tri 34649 34946 34665 34962 se
rect 34665 34946 34742 34962
rect 34649 34880 34742 34946
rect 34370 34745 34742 34821
rect 34370 34620 34463 34686
rect 34370 34604 34447 34620
tri 34447 34604 34463 34620 nw
rect 34499 34587 34613 34745
rect 34649 34620 34742 34686
tri 34649 34604 34665 34620 ne
rect 34665 34604 34742 34620
rect 34482 34505 34630 34587
rect 34370 34472 34447 34488
tri 34447 34472 34463 34488 sw
rect 34370 34406 34463 34472
rect 34370 34304 34463 34370
rect 34370 34288 34447 34304
tri 34447 34288 34463 34304 nw
rect 34499 34271 34613 34505
tri 34649 34472 34665 34488 se
rect 34665 34472 34742 34488
rect 34649 34406 34742 34472
rect 34649 34304 34742 34370
tri 34649 34288 34665 34304 ne
rect 34665 34288 34742 34304
rect 34482 34189 34630 34271
rect 34370 34156 34447 34172
tri 34447 34156 34463 34172 sw
rect 34370 34090 34463 34156
rect 34499 34031 34613 34189
tri 34649 34156 34665 34172 se
rect 34665 34156 34742 34172
rect 34649 34090 34742 34156
rect 34370 33955 34742 34031
rect 34370 33830 34463 33896
rect 34370 33814 34447 33830
tri 34447 33814 34463 33830 nw
rect 34499 33797 34613 33955
rect 34649 33830 34742 33896
tri 34649 33814 34665 33830 ne
rect 34665 33814 34742 33830
rect 34482 33715 34630 33797
rect 34370 33682 34447 33698
tri 34447 33682 34463 33698 sw
rect 34370 33616 34463 33682
rect 34370 33514 34463 33580
rect 34370 33498 34447 33514
tri 34447 33498 34463 33514 nw
rect 34499 33481 34613 33715
tri 34649 33682 34665 33698 se
rect 34665 33682 34742 33698
rect 34649 33616 34742 33682
rect 34649 33514 34742 33580
tri 34649 33498 34665 33514 ne
rect 34665 33498 34742 33514
rect 34482 33399 34630 33481
rect 34370 33366 34447 33382
tri 34447 33366 34463 33382 sw
rect 34370 33300 34463 33366
rect 34499 33241 34613 33399
tri 34649 33366 34665 33382 se
rect 34665 33366 34742 33382
rect 34649 33300 34742 33366
rect 34370 33165 34742 33241
rect 34370 33040 34463 33106
rect 34370 33024 34447 33040
tri 34447 33024 34463 33040 nw
rect 34499 33007 34613 33165
rect 34649 33040 34742 33106
tri 34649 33024 34665 33040 ne
rect 34665 33024 34742 33040
rect 34482 32925 34630 33007
rect 34370 32892 34447 32908
tri 34447 32892 34463 32908 sw
rect 34370 32826 34463 32892
rect 34370 32724 34463 32790
rect 34370 32708 34447 32724
tri 34447 32708 34463 32724 nw
rect 34499 32691 34613 32925
tri 34649 32892 34665 32908 se
rect 34665 32892 34742 32908
rect 34649 32826 34742 32892
rect 34649 32724 34742 32790
tri 34649 32708 34665 32724 ne
rect 34665 32708 34742 32724
rect 34482 32609 34630 32691
rect 34370 32576 34447 32592
tri 34447 32576 34463 32592 sw
rect 34370 32510 34463 32576
rect 34499 32451 34613 32609
tri 34649 32576 34665 32592 se
rect 34665 32576 34742 32592
rect 34649 32510 34742 32576
rect 34370 32375 34742 32451
rect 34370 32250 34463 32316
rect 34370 32234 34447 32250
tri 34447 32234 34463 32250 nw
rect 34499 32217 34613 32375
rect 34649 32250 34742 32316
tri 34649 32234 34665 32250 ne
rect 34665 32234 34742 32250
rect 34482 32135 34630 32217
rect 34370 32102 34447 32118
tri 34447 32102 34463 32118 sw
rect 34370 32036 34463 32102
rect 34370 31934 34463 32000
rect 34370 31918 34447 31934
tri 34447 31918 34463 31934 nw
rect 34499 31901 34613 32135
tri 34649 32102 34665 32118 se
rect 34665 32102 34742 32118
rect 34649 32036 34742 32102
rect 34649 31934 34742 32000
tri 34649 31918 34665 31934 ne
rect 34665 31918 34742 31934
rect 34482 31819 34630 31901
rect 34370 31786 34447 31802
tri 34447 31786 34463 31802 sw
rect 34370 31720 34463 31786
rect 34499 31661 34613 31819
tri 34649 31786 34665 31802 se
rect 34665 31786 34742 31802
rect 34649 31720 34742 31786
rect 34370 31585 34742 31661
rect 34370 31460 34463 31526
rect 34370 31444 34447 31460
tri 34447 31444 34463 31460 nw
rect 34499 31427 34613 31585
rect 34649 31460 34742 31526
tri 34649 31444 34665 31460 ne
rect 34665 31444 34742 31460
rect 34482 31345 34630 31427
rect 34370 31312 34447 31328
tri 34447 31312 34463 31328 sw
rect 34370 31246 34463 31312
rect 34370 31144 34463 31210
rect 34370 31128 34447 31144
tri 34447 31128 34463 31144 nw
rect 34499 31111 34613 31345
tri 34649 31312 34665 31328 se
rect 34665 31312 34742 31328
rect 34649 31246 34742 31312
rect 34649 31144 34742 31210
tri 34649 31128 34665 31144 ne
rect 34665 31128 34742 31144
rect 34482 31029 34630 31111
rect 34370 30996 34447 31012
tri 34447 30996 34463 31012 sw
rect 34370 30930 34463 30996
rect 34499 30871 34613 31029
tri 34649 30996 34665 31012 se
rect 34665 30996 34742 31012
rect 34649 30930 34742 30996
rect 34370 30795 34742 30871
rect 34370 30670 34463 30736
rect 34370 30654 34447 30670
tri 34447 30654 34463 30670 nw
rect 34499 30637 34613 30795
rect 34649 30670 34742 30736
tri 34649 30654 34665 30670 ne
rect 34665 30654 34742 30670
rect 34482 30555 34630 30637
rect 34370 30522 34447 30538
tri 34447 30522 34463 30538 sw
rect 34370 30456 34463 30522
rect 34370 30354 34463 30420
rect 34370 30338 34447 30354
tri 34447 30338 34463 30354 nw
rect 34499 30321 34613 30555
tri 34649 30522 34665 30538 se
rect 34665 30522 34742 30538
rect 34649 30456 34742 30522
rect 34649 30354 34742 30420
tri 34649 30338 34665 30354 ne
rect 34665 30338 34742 30354
rect 34482 30239 34630 30321
rect 34370 30206 34447 30222
tri 34447 30206 34463 30222 sw
rect 34370 30140 34463 30206
rect 34499 30081 34613 30239
tri 34649 30206 34665 30222 se
rect 34665 30206 34742 30222
rect 34649 30140 34742 30206
rect 34370 30005 34742 30081
rect 34370 29880 34463 29946
rect 34370 29864 34447 29880
tri 34447 29864 34463 29880 nw
rect 34499 29847 34613 30005
rect 34649 29880 34742 29946
tri 34649 29864 34665 29880 ne
rect 34665 29864 34742 29880
rect 34482 29765 34630 29847
rect 34370 29732 34447 29748
tri 34447 29732 34463 29748 sw
rect 34370 29666 34463 29732
rect 34370 29564 34463 29630
rect 34370 29548 34447 29564
tri 34447 29548 34463 29564 nw
rect 34499 29531 34613 29765
tri 34649 29732 34665 29748 se
rect 34665 29732 34742 29748
rect 34649 29666 34742 29732
rect 34649 29564 34742 29630
tri 34649 29548 34665 29564 ne
rect 34665 29548 34742 29564
rect 34482 29449 34630 29531
rect 34370 29416 34447 29432
tri 34447 29416 34463 29432 sw
rect 34370 29350 34463 29416
rect 34499 29291 34613 29449
tri 34649 29416 34665 29432 se
rect 34665 29416 34742 29432
rect 34649 29350 34742 29416
rect 34370 29215 34742 29291
rect 34370 29090 34463 29156
rect 34370 29074 34447 29090
tri 34447 29074 34463 29090 nw
rect 34499 29057 34613 29215
rect 34649 29090 34742 29156
tri 34649 29074 34665 29090 ne
rect 34665 29074 34742 29090
rect 34482 28975 34630 29057
rect 34370 28942 34447 28958
tri 34447 28942 34463 28958 sw
rect 34370 28876 34463 28942
rect 34499 28833 34613 28975
tri 34649 28942 34665 28958 se
rect 34665 28942 34742 28958
rect 34649 28876 34742 28942
rect 34778 28463 34814 80603
rect 34850 28463 34886 80603
rect 34922 80445 34958 80603
rect 34914 80303 34966 80445
rect 34922 28763 34958 80303
rect 34914 28621 34966 28763
rect 34922 28463 34958 28621
rect 34994 28463 35030 80603
rect 35066 28463 35102 80603
rect 35138 28833 35222 80233
rect 35258 28463 35294 80603
rect 35330 28463 35366 80603
rect 35402 80445 35438 80603
rect 35394 80303 35446 80445
rect 35402 28763 35438 80303
rect 35394 28621 35446 28763
rect 35402 28463 35438 28621
rect 35474 28463 35510 80603
rect 35546 28463 35582 80603
rect 35618 80124 35711 80190
rect 35618 80108 35695 80124
tri 35695 80108 35711 80124 nw
rect 35747 80091 35861 80233
rect 35897 80124 35990 80190
tri 35897 80108 35913 80124 ne
rect 35913 80108 35990 80124
rect 35730 80009 35878 80091
rect 35618 79976 35695 79992
tri 35695 79976 35711 79992 sw
rect 35618 79910 35711 79976
rect 35747 79851 35861 80009
tri 35897 79976 35913 79992 se
rect 35913 79976 35990 79992
rect 35897 79910 35990 79976
rect 35618 79775 35990 79851
rect 35618 79650 35711 79716
rect 35618 79634 35695 79650
tri 35695 79634 35711 79650 nw
rect 35747 79617 35861 79775
rect 35897 79650 35990 79716
tri 35897 79634 35913 79650 ne
rect 35913 79634 35990 79650
rect 35730 79535 35878 79617
rect 35618 79502 35695 79518
tri 35695 79502 35711 79518 sw
rect 35618 79436 35711 79502
rect 35618 79334 35711 79400
rect 35618 79318 35695 79334
tri 35695 79318 35711 79334 nw
rect 35747 79301 35861 79535
tri 35897 79502 35913 79518 se
rect 35913 79502 35990 79518
rect 35897 79436 35990 79502
rect 35897 79334 35990 79400
tri 35897 79318 35913 79334 ne
rect 35913 79318 35990 79334
rect 35730 79219 35878 79301
rect 35618 79186 35695 79202
tri 35695 79186 35711 79202 sw
rect 35618 79120 35711 79186
rect 35747 79061 35861 79219
tri 35897 79186 35913 79202 se
rect 35913 79186 35990 79202
rect 35897 79120 35990 79186
rect 35618 78985 35990 79061
rect 35618 78860 35711 78926
rect 35618 78844 35695 78860
tri 35695 78844 35711 78860 nw
rect 35747 78827 35861 78985
rect 35897 78860 35990 78926
tri 35897 78844 35913 78860 ne
rect 35913 78844 35990 78860
rect 35730 78745 35878 78827
rect 35618 78712 35695 78728
tri 35695 78712 35711 78728 sw
rect 35618 78646 35711 78712
rect 35618 78544 35711 78610
rect 35618 78528 35695 78544
tri 35695 78528 35711 78544 nw
rect 35747 78511 35861 78745
tri 35897 78712 35913 78728 se
rect 35913 78712 35990 78728
rect 35897 78646 35990 78712
rect 35897 78544 35990 78610
tri 35897 78528 35913 78544 ne
rect 35913 78528 35990 78544
rect 35730 78429 35878 78511
rect 35618 78396 35695 78412
tri 35695 78396 35711 78412 sw
rect 35618 78330 35711 78396
rect 35747 78271 35861 78429
tri 35897 78396 35913 78412 se
rect 35913 78396 35990 78412
rect 35897 78330 35990 78396
rect 35618 78195 35990 78271
rect 35618 78070 35711 78136
rect 35618 78054 35695 78070
tri 35695 78054 35711 78070 nw
rect 35747 78037 35861 78195
rect 35897 78070 35990 78136
tri 35897 78054 35913 78070 ne
rect 35913 78054 35990 78070
rect 35730 77955 35878 78037
rect 35618 77922 35695 77938
tri 35695 77922 35711 77938 sw
rect 35618 77856 35711 77922
rect 35618 77754 35711 77820
rect 35618 77738 35695 77754
tri 35695 77738 35711 77754 nw
rect 35747 77721 35861 77955
tri 35897 77922 35913 77938 se
rect 35913 77922 35990 77938
rect 35897 77856 35990 77922
rect 35897 77754 35990 77820
tri 35897 77738 35913 77754 ne
rect 35913 77738 35990 77754
rect 35730 77639 35878 77721
rect 35618 77606 35695 77622
tri 35695 77606 35711 77622 sw
rect 35618 77540 35711 77606
rect 35747 77481 35861 77639
tri 35897 77606 35913 77622 se
rect 35913 77606 35990 77622
rect 35897 77540 35990 77606
rect 35618 77405 35990 77481
rect 35618 77280 35711 77346
rect 35618 77264 35695 77280
tri 35695 77264 35711 77280 nw
rect 35747 77247 35861 77405
rect 35897 77280 35990 77346
tri 35897 77264 35913 77280 ne
rect 35913 77264 35990 77280
rect 35730 77165 35878 77247
rect 35618 77132 35695 77148
tri 35695 77132 35711 77148 sw
rect 35618 77066 35711 77132
rect 35618 76964 35711 77030
rect 35618 76948 35695 76964
tri 35695 76948 35711 76964 nw
rect 35747 76931 35861 77165
tri 35897 77132 35913 77148 se
rect 35913 77132 35990 77148
rect 35897 77066 35990 77132
rect 35897 76964 35990 77030
tri 35897 76948 35913 76964 ne
rect 35913 76948 35990 76964
rect 35730 76849 35878 76931
rect 35618 76816 35695 76832
tri 35695 76816 35711 76832 sw
rect 35618 76750 35711 76816
rect 35747 76691 35861 76849
tri 35897 76816 35913 76832 se
rect 35913 76816 35990 76832
rect 35897 76750 35990 76816
rect 35618 76615 35990 76691
rect 35618 76490 35711 76556
rect 35618 76474 35695 76490
tri 35695 76474 35711 76490 nw
rect 35747 76457 35861 76615
rect 35897 76490 35990 76556
tri 35897 76474 35913 76490 ne
rect 35913 76474 35990 76490
rect 35730 76375 35878 76457
rect 35618 76342 35695 76358
tri 35695 76342 35711 76358 sw
rect 35618 76276 35711 76342
rect 35618 76174 35711 76240
rect 35618 76158 35695 76174
tri 35695 76158 35711 76174 nw
rect 35747 76141 35861 76375
tri 35897 76342 35913 76358 se
rect 35913 76342 35990 76358
rect 35897 76276 35990 76342
rect 35897 76174 35990 76240
tri 35897 76158 35913 76174 ne
rect 35913 76158 35990 76174
rect 35730 76059 35878 76141
rect 35618 76026 35695 76042
tri 35695 76026 35711 76042 sw
rect 35618 75960 35711 76026
rect 35747 75901 35861 76059
tri 35897 76026 35913 76042 se
rect 35913 76026 35990 76042
rect 35897 75960 35990 76026
rect 35618 75825 35990 75901
rect 35618 75700 35711 75766
rect 35618 75684 35695 75700
tri 35695 75684 35711 75700 nw
rect 35747 75667 35861 75825
rect 35897 75700 35990 75766
tri 35897 75684 35913 75700 ne
rect 35913 75684 35990 75700
rect 35730 75585 35878 75667
rect 35618 75552 35695 75568
tri 35695 75552 35711 75568 sw
rect 35618 75486 35711 75552
rect 35618 75384 35711 75450
rect 35618 75368 35695 75384
tri 35695 75368 35711 75384 nw
rect 35747 75351 35861 75585
tri 35897 75552 35913 75568 se
rect 35913 75552 35990 75568
rect 35897 75486 35990 75552
rect 35897 75384 35990 75450
tri 35897 75368 35913 75384 ne
rect 35913 75368 35990 75384
rect 35730 75269 35878 75351
rect 35618 75236 35695 75252
tri 35695 75236 35711 75252 sw
rect 35618 75170 35711 75236
rect 35747 75111 35861 75269
tri 35897 75236 35913 75252 se
rect 35913 75236 35990 75252
rect 35897 75170 35990 75236
rect 35618 75035 35990 75111
rect 35618 74910 35711 74976
rect 35618 74894 35695 74910
tri 35695 74894 35711 74910 nw
rect 35747 74877 35861 75035
rect 35897 74910 35990 74976
tri 35897 74894 35913 74910 ne
rect 35913 74894 35990 74910
rect 35730 74795 35878 74877
rect 35618 74762 35695 74778
tri 35695 74762 35711 74778 sw
rect 35618 74696 35711 74762
rect 35618 74594 35711 74660
rect 35618 74578 35695 74594
tri 35695 74578 35711 74594 nw
rect 35747 74561 35861 74795
tri 35897 74762 35913 74778 se
rect 35913 74762 35990 74778
rect 35897 74696 35990 74762
rect 35897 74594 35990 74660
tri 35897 74578 35913 74594 ne
rect 35913 74578 35990 74594
rect 35730 74479 35878 74561
rect 35618 74446 35695 74462
tri 35695 74446 35711 74462 sw
rect 35618 74380 35711 74446
rect 35747 74321 35861 74479
tri 35897 74446 35913 74462 se
rect 35913 74446 35990 74462
rect 35897 74380 35990 74446
rect 35618 74245 35990 74321
rect 35618 74120 35711 74186
rect 35618 74104 35695 74120
tri 35695 74104 35711 74120 nw
rect 35747 74087 35861 74245
rect 35897 74120 35990 74186
tri 35897 74104 35913 74120 ne
rect 35913 74104 35990 74120
rect 35730 74005 35878 74087
rect 35618 73972 35695 73988
tri 35695 73972 35711 73988 sw
rect 35618 73906 35711 73972
rect 35618 73804 35711 73870
rect 35618 73788 35695 73804
tri 35695 73788 35711 73804 nw
rect 35747 73771 35861 74005
tri 35897 73972 35913 73988 se
rect 35913 73972 35990 73988
rect 35897 73906 35990 73972
rect 35897 73804 35990 73870
tri 35897 73788 35913 73804 ne
rect 35913 73788 35990 73804
rect 35730 73689 35878 73771
rect 35618 73656 35695 73672
tri 35695 73656 35711 73672 sw
rect 35618 73590 35711 73656
rect 35747 73531 35861 73689
tri 35897 73656 35913 73672 se
rect 35913 73656 35990 73672
rect 35897 73590 35990 73656
rect 35618 73455 35990 73531
rect 35618 73330 35711 73396
rect 35618 73314 35695 73330
tri 35695 73314 35711 73330 nw
rect 35747 73297 35861 73455
rect 35897 73330 35990 73396
tri 35897 73314 35913 73330 ne
rect 35913 73314 35990 73330
rect 35730 73215 35878 73297
rect 35618 73182 35695 73198
tri 35695 73182 35711 73198 sw
rect 35618 73116 35711 73182
rect 35618 73014 35711 73080
rect 35618 72998 35695 73014
tri 35695 72998 35711 73014 nw
rect 35747 72981 35861 73215
tri 35897 73182 35913 73198 se
rect 35913 73182 35990 73198
rect 35897 73116 35990 73182
rect 35897 73014 35990 73080
tri 35897 72998 35913 73014 ne
rect 35913 72998 35990 73014
rect 35730 72899 35878 72981
rect 35618 72866 35695 72882
tri 35695 72866 35711 72882 sw
rect 35618 72800 35711 72866
rect 35747 72741 35861 72899
tri 35897 72866 35913 72882 se
rect 35913 72866 35990 72882
rect 35897 72800 35990 72866
rect 35618 72665 35990 72741
rect 35618 72540 35711 72606
rect 35618 72524 35695 72540
tri 35695 72524 35711 72540 nw
rect 35747 72507 35861 72665
rect 35897 72540 35990 72606
tri 35897 72524 35913 72540 ne
rect 35913 72524 35990 72540
rect 35730 72425 35878 72507
rect 35618 72392 35695 72408
tri 35695 72392 35711 72408 sw
rect 35618 72326 35711 72392
rect 35618 72224 35711 72290
rect 35618 72208 35695 72224
tri 35695 72208 35711 72224 nw
rect 35747 72191 35861 72425
tri 35897 72392 35913 72408 se
rect 35913 72392 35990 72408
rect 35897 72326 35990 72392
rect 35897 72224 35990 72290
tri 35897 72208 35913 72224 ne
rect 35913 72208 35990 72224
rect 35730 72109 35878 72191
rect 35618 72076 35695 72092
tri 35695 72076 35711 72092 sw
rect 35618 72010 35711 72076
rect 35747 71951 35861 72109
tri 35897 72076 35913 72092 se
rect 35913 72076 35990 72092
rect 35897 72010 35990 72076
rect 35618 71875 35990 71951
rect 35618 71750 35711 71816
rect 35618 71734 35695 71750
tri 35695 71734 35711 71750 nw
rect 35747 71717 35861 71875
rect 35897 71750 35990 71816
tri 35897 71734 35913 71750 ne
rect 35913 71734 35990 71750
rect 35730 71635 35878 71717
rect 35618 71602 35695 71618
tri 35695 71602 35711 71618 sw
rect 35618 71536 35711 71602
rect 35618 71434 35711 71500
rect 35618 71418 35695 71434
tri 35695 71418 35711 71434 nw
rect 35747 71401 35861 71635
tri 35897 71602 35913 71618 se
rect 35913 71602 35990 71618
rect 35897 71536 35990 71602
rect 35897 71434 35990 71500
tri 35897 71418 35913 71434 ne
rect 35913 71418 35990 71434
rect 35730 71319 35878 71401
rect 35618 71286 35695 71302
tri 35695 71286 35711 71302 sw
rect 35618 71220 35711 71286
rect 35747 71161 35861 71319
tri 35897 71286 35913 71302 se
rect 35913 71286 35990 71302
rect 35897 71220 35990 71286
rect 35618 71085 35990 71161
rect 35618 70960 35711 71026
rect 35618 70944 35695 70960
tri 35695 70944 35711 70960 nw
rect 35747 70927 35861 71085
rect 35897 70960 35990 71026
tri 35897 70944 35913 70960 ne
rect 35913 70944 35990 70960
rect 35730 70845 35878 70927
rect 35618 70812 35695 70828
tri 35695 70812 35711 70828 sw
rect 35618 70746 35711 70812
rect 35618 70644 35711 70710
rect 35618 70628 35695 70644
tri 35695 70628 35711 70644 nw
rect 35747 70611 35861 70845
tri 35897 70812 35913 70828 se
rect 35913 70812 35990 70828
rect 35897 70746 35990 70812
rect 35897 70644 35990 70710
tri 35897 70628 35913 70644 ne
rect 35913 70628 35990 70644
rect 35730 70529 35878 70611
rect 35618 70496 35695 70512
tri 35695 70496 35711 70512 sw
rect 35618 70430 35711 70496
rect 35747 70371 35861 70529
tri 35897 70496 35913 70512 se
rect 35913 70496 35990 70512
rect 35897 70430 35990 70496
rect 35618 70295 35990 70371
rect 35618 70170 35711 70236
rect 35618 70154 35695 70170
tri 35695 70154 35711 70170 nw
rect 35747 70137 35861 70295
rect 35897 70170 35990 70236
tri 35897 70154 35913 70170 ne
rect 35913 70154 35990 70170
rect 35730 70055 35878 70137
rect 35618 70022 35695 70038
tri 35695 70022 35711 70038 sw
rect 35618 69956 35711 70022
rect 35618 69854 35711 69920
rect 35618 69838 35695 69854
tri 35695 69838 35711 69854 nw
rect 35747 69821 35861 70055
tri 35897 70022 35913 70038 se
rect 35913 70022 35990 70038
rect 35897 69956 35990 70022
rect 35897 69854 35990 69920
tri 35897 69838 35913 69854 ne
rect 35913 69838 35990 69854
rect 35730 69739 35878 69821
rect 35618 69706 35695 69722
tri 35695 69706 35711 69722 sw
rect 35618 69640 35711 69706
rect 35747 69581 35861 69739
tri 35897 69706 35913 69722 se
rect 35913 69706 35990 69722
rect 35897 69640 35990 69706
rect 35618 69505 35990 69581
rect 35618 69380 35711 69446
rect 35618 69364 35695 69380
tri 35695 69364 35711 69380 nw
rect 35747 69347 35861 69505
rect 35897 69380 35990 69446
tri 35897 69364 35913 69380 ne
rect 35913 69364 35990 69380
rect 35730 69265 35878 69347
rect 35618 69232 35695 69248
tri 35695 69232 35711 69248 sw
rect 35618 69166 35711 69232
rect 35618 69064 35711 69130
rect 35618 69048 35695 69064
tri 35695 69048 35711 69064 nw
rect 35747 69031 35861 69265
tri 35897 69232 35913 69248 se
rect 35913 69232 35990 69248
rect 35897 69166 35990 69232
rect 35897 69064 35990 69130
tri 35897 69048 35913 69064 ne
rect 35913 69048 35990 69064
rect 35730 68949 35878 69031
rect 35618 68916 35695 68932
tri 35695 68916 35711 68932 sw
rect 35618 68850 35711 68916
rect 35747 68791 35861 68949
tri 35897 68916 35913 68932 se
rect 35913 68916 35990 68932
rect 35897 68850 35990 68916
rect 35618 68715 35990 68791
rect 35618 68590 35711 68656
rect 35618 68574 35695 68590
tri 35695 68574 35711 68590 nw
rect 35747 68557 35861 68715
rect 35897 68590 35990 68656
tri 35897 68574 35913 68590 ne
rect 35913 68574 35990 68590
rect 35730 68475 35878 68557
rect 35618 68442 35695 68458
tri 35695 68442 35711 68458 sw
rect 35618 68376 35711 68442
rect 35618 68274 35711 68340
rect 35618 68258 35695 68274
tri 35695 68258 35711 68274 nw
rect 35747 68241 35861 68475
tri 35897 68442 35913 68458 se
rect 35913 68442 35990 68458
rect 35897 68376 35990 68442
rect 35897 68274 35990 68340
tri 35897 68258 35913 68274 ne
rect 35913 68258 35990 68274
rect 35730 68159 35878 68241
rect 35618 68126 35695 68142
tri 35695 68126 35711 68142 sw
rect 35618 68060 35711 68126
rect 35747 68001 35861 68159
tri 35897 68126 35913 68142 se
rect 35913 68126 35990 68142
rect 35897 68060 35990 68126
rect 35618 67925 35990 68001
rect 35618 67800 35711 67866
rect 35618 67784 35695 67800
tri 35695 67784 35711 67800 nw
rect 35747 67767 35861 67925
rect 35897 67800 35990 67866
tri 35897 67784 35913 67800 ne
rect 35913 67784 35990 67800
rect 35730 67685 35878 67767
rect 35618 67652 35695 67668
tri 35695 67652 35711 67668 sw
rect 35618 67586 35711 67652
rect 35618 67484 35711 67550
rect 35618 67468 35695 67484
tri 35695 67468 35711 67484 nw
rect 35747 67451 35861 67685
tri 35897 67652 35913 67668 se
rect 35913 67652 35990 67668
rect 35897 67586 35990 67652
rect 35897 67484 35990 67550
tri 35897 67468 35913 67484 ne
rect 35913 67468 35990 67484
rect 35730 67369 35878 67451
rect 35618 67336 35695 67352
tri 35695 67336 35711 67352 sw
rect 35618 67270 35711 67336
rect 35747 67211 35861 67369
tri 35897 67336 35913 67352 se
rect 35913 67336 35990 67352
rect 35897 67270 35990 67336
rect 35618 67135 35990 67211
rect 35618 67010 35711 67076
rect 35618 66994 35695 67010
tri 35695 66994 35711 67010 nw
rect 35747 66977 35861 67135
rect 35897 67010 35990 67076
tri 35897 66994 35913 67010 ne
rect 35913 66994 35990 67010
rect 35730 66895 35878 66977
rect 35618 66862 35695 66878
tri 35695 66862 35711 66878 sw
rect 35618 66796 35711 66862
rect 35618 66694 35711 66760
rect 35618 66678 35695 66694
tri 35695 66678 35711 66694 nw
rect 35747 66661 35861 66895
tri 35897 66862 35913 66878 se
rect 35913 66862 35990 66878
rect 35897 66796 35990 66862
rect 35897 66694 35990 66760
tri 35897 66678 35913 66694 ne
rect 35913 66678 35990 66694
rect 35730 66579 35878 66661
rect 35618 66546 35695 66562
tri 35695 66546 35711 66562 sw
rect 35618 66480 35711 66546
rect 35747 66421 35861 66579
tri 35897 66546 35913 66562 se
rect 35913 66546 35990 66562
rect 35897 66480 35990 66546
rect 35618 66345 35990 66421
rect 35618 66220 35711 66286
rect 35618 66204 35695 66220
tri 35695 66204 35711 66220 nw
rect 35747 66187 35861 66345
rect 35897 66220 35990 66286
tri 35897 66204 35913 66220 ne
rect 35913 66204 35990 66220
rect 35730 66105 35878 66187
rect 35618 66072 35695 66088
tri 35695 66072 35711 66088 sw
rect 35618 66006 35711 66072
rect 35618 65904 35711 65970
rect 35618 65888 35695 65904
tri 35695 65888 35711 65904 nw
rect 35747 65871 35861 66105
tri 35897 66072 35913 66088 se
rect 35913 66072 35990 66088
rect 35897 66006 35990 66072
rect 35897 65904 35990 65970
tri 35897 65888 35913 65904 ne
rect 35913 65888 35990 65904
rect 35730 65789 35878 65871
rect 35618 65756 35695 65772
tri 35695 65756 35711 65772 sw
rect 35618 65690 35711 65756
rect 35747 65631 35861 65789
tri 35897 65756 35913 65772 se
rect 35913 65756 35990 65772
rect 35897 65690 35990 65756
rect 35618 65555 35990 65631
rect 35618 65430 35711 65496
rect 35618 65414 35695 65430
tri 35695 65414 35711 65430 nw
rect 35747 65397 35861 65555
rect 35897 65430 35990 65496
tri 35897 65414 35913 65430 ne
rect 35913 65414 35990 65430
rect 35730 65315 35878 65397
rect 35618 65282 35695 65298
tri 35695 65282 35711 65298 sw
rect 35618 65216 35711 65282
rect 35618 65114 35711 65180
rect 35618 65098 35695 65114
tri 35695 65098 35711 65114 nw
rect 35747 65081 35861 65315
tri 35897 65282 35913 65298 se
rect 35913 65282 35990 65298
rect 35897 65216 35990 65282
rect 35897 65114 35990 65180
tri 35897 65098 35913 65114 ne
rect 35913 65098 35990 65114
rect 35730 64999 35878 65081
rect 35618 64966 35695 64982
tri 35695 64966 35711 64982 sw
rect 35618 64900 35711 64966
rect 35747 64841 35861 64999
tri 35897 64966 35913 64982 se
rect 35913 64966 35990 64982
rect 35897 64900 35990 64966
rect 35618 64765 35990 64841
rect 35618 64640 35711 64706
rect 35618 64624 35695 64640
tri 35695 64624 35711 64640 nw
rect 35747 64607 35861 64765
rect 35897 64640 35990 64706
tri 35897 64624 35913 64640 ne
rect 35913 64624 35990 64640
rect 35730 64525 35878 64607
rect 35618 64492 35695 64508
tri 35695 64492 35711 64508 sw
rect 35618 64426 35711 64492
rect 35618 64324 35711 64390
rect 35618 64308 35695 64324
tri 35695 64308 35711 64324 nw
rect 35747 64291 35861 64525
tri 35897 64492 35913 64508 se
rect 35913 64492 35990 64508
rect 35897 64426 35990 64492
rect 35897 64324 35990 64390
tri 35897 64308 35913 64324 ne
rect 35913 64308 35990 64324
rect 35730 64209 35878 64291
rect 35618 64176 35695 64192
tri 35695 64176 35711 64192 sw
rect 35618 64110 35711 64176
rect 35747 64051 35861 64209
tri 35897 64176 35913 64192 se
rect 35913 64176 35990 64192
rect 35897 64110 35990 64176
rect 35618 63975 35990 64051
rect 35618 63850 35711 63916
rect 35618 63834 35695 63850
tri 35695 63834 35711 63850 nw
rect 35747 63817 35861 63975
rect 35897 63850 35990 63916
tri 35897 63834 35913 63850 ne
rect 35913 63834 35990 63850
rect 35730 63735 35878 63817
rect 35618 63702 35695 63718
tri 35695 63702 35711 63718 sw
rect 35618 63636 35711 63702
rect 35618 63534 35711 63600
rect 35618 63518 35695 63534
tri 35695 63518 35711 63534 nw
rect 35747 63501 35861 63735
tri 35897 63702 35913 63718 se
rect 35913 63702 35990 63718
rect 35897 63636 35990 63702
rect 35897 63534 35990 63600
tri 35897 63518 35913 63534 ne
rect 35913 63518 35990 63534
rect 35730 63419 35878 63501
rect 35618 63386 35695 63402
tri 35695 63386 35711 63402 sw
rect 35618 63320 35711 63386
rect 35747 63261 35861 63419
tri 35897 63386 35913 63402 se
rect 35913 63386 35990 63402
rect 35897 63320 35990 63386
rect 35618 63185 35990 63261
rect 35618 63060 35711 63126
rect 35618 63044 35695 63060
tri 35695 63044 35711 63060 nw
rect 35747 63027 35861 63185
rect 35897 63060 35990 63126
tri 35897 63044 35913 63060 ne
rect 35913 63044 35990 63060
rect 35730 62945 35878 63027
rect 35618 62912 35695 62928
tri 35695 62912 35711 62928 sw
rect 35618 62846 35711 62912
rect 35618 62744 35711 62810
rect 35618 62728 35695 62744
tri 35695 62728 35711 62744 nw
rect 35747 62711 35861 62945
tri 35897 62912 35913 62928 se
rect 35913 62912 35990 62928
rect 35897 62846 35990 62912
rect 35897 62744 35990 62810
tri 35897 62728 35913 62744 ne
rect 35913 62728 35990 62744
rect 35730 62629 35878 62711
rect 35618 62596 35695 62612
tri 35695 62596 35711 62612 sw
rect 35618 62530 35711 62596
rect 35747 62471 35861 62629
tri 35897 62596 35913 62612 se
rect 35913 62596 35990 62612
rect 35897 62530 35990 62596
rect 35618 62395 35990 62471
rect 35618 62270 35711 62336
rect 35618 62254 35695 62270
tri 35695 62254 35711 62270 nw
rect 35747 62237 35861 62395
rect 35897 62270 35990 62336
tri 35897 62254 35913 62270 ne
rect 35913 62254 35990 62270
rect 35730 62155 35878 62237
rect 35618 62122 35695 62138
tri 35695 62122 35711 62138 sw
rect 35618 62056 35711 62122
rect 35618 61954 35711 62020
rect 35618 61938 35695 61954
tri 35695 61938 35711 61954 nw
rect 35747 61921 35861 62155
tri 35897 62122 35913 62138 se
rect 35913 62122 35990 62138
rect 35897 62056 35990 62122
rect 35897 61954 35990 62020
tri 35897 61938 35913 61954 ne
rect 35913 61938 35990 61954
rect 35730 61839 35878 61921
rect 35618 61806 35695 61822
tri 35695 61806 35711 61822 sw
rect 35618 61740 35711 61806
rect 35747 61681 35861 61839
tri 35897 61806 35913 61822 se
rect 35913 61806 35990 61822
rect 35897 61740 35990 61806
rect 35618 61605 35990 61681
rect 35618 61480 35711 61546
rect 35618 61464 35695 61480
tri 35695 61464 35711 61480 nw
rect 35747 61447 35861 61605
rect 35897 61480 35990 61546
tri 35897 61464 35913 61480 ne
rect 35913 61464 35990 61480
rect 35730 61365 35878 61447
rect 35618 61332 35695 61348
tri 35695 61332 35711 61348 sw
rect 35618 61266 35711 61332
rect 35618 61164 35711 61230
rect 35618 61148 35695 61164
tri 35695 61148 35711 61164 nw
rect 35747 61131 35861 61365
tri 35897 61332 35913 61348 se
rect 35913 61332 35990 61348
rect 35897 61266 35990 61332
rect 35897 61164 35990 61230
tri 35897 61148 35913 61164 ne
rect 35913 61148 35990 61164
rect 35730 61049 35878 61131
rect 35618 61016 35695 61032
tri 35695 61016 35711 61032 sw
rect 35618 60950 35711 61016
rect 35747 60891 35861 61049
tri 35897 61016 35913 61032 se
rect 35913 61016 35990 61032
rect 35897 60950 35990 61016
rect 35618 60815 35990 60891
rect 35618 60690 35711 60756
rect 35618 60674 35695 60690
tri 35695 60674 35711 60690 nw
rect 35747 60657 35861 60815
rect 35897 60690 35990 60756
tri 35897 60674 35913 60690 ne
rect 35913 60674 35990 60690
rect 35730 60575 35878 60657
rect 35618 60542 35695 60558
tri 35695 60542 35711 60558 sw
rect 35618 60476 35711 60542
rect 35618 60374 35711 60440
rect 35618 60358 35695 60374
tri 35695 60358 35711 60374 nw
rect 35747 60341 35861 60575
tri 35897 60542 35913 60558 se
rect 35913 60542 35990 60558
rect 35897 60476 35990 60542
rect 35897 60374 35990 60440
tri 35897 60358 35913 60374 ne
rect 35913 60358 35990 60374
rect 35730 60259 35878 60341
rect 35618 60226 35695 60242
tri 35695 60226 35711 60242 sw
rect 35618 60160 35711 60226
rect 35747 60101 35861 60259
tri 35897 60226 35913 60242 se
rect 35913 60226 35990 60242
rect 35897 60160 35990 60226
rect 35618 60025 35990 60101
rect 35618 59900 35711 59966
rect 35618 59884 35695 59900
tri 35695 59884 35711 59900 nw
rect 35747 59867 35861 60025
rect 35897 59900 35990 59966
tri 35897 59884 35913 59900 ne
rect 35913 59884 35990 59900
rect 35730 59785 35878 59867
rect 35618 59752 35695 59768
tri 35695 59752 35711 59768 sw
rect 35618 59686 35711 59752
rect 35618 59584 35711 59650
rect 35618 59568 35695 59584
tri 35695 59568 35711 59584 nw
rect 35747 59551 35861 59785
tri 35897 59752 35913 59768 se
rect 35913 59752 35990 59768
rect 35897 59686 35990 59752
rect 35897 59584 35990 59650
tri 35897 59568 35913 59584 ne
rect 35913 59568 35990 59584
rect 35730 59469 35878 59551
rect 35618 59436 35695 59452
tri 35695 59436 35711 59452 sw
rect 35618 59370 35711 59436
rect 35747 59311 35861 59469
tri 35897 59436 35913 59452 se
rect 35913 59436 35990 59452
rect 35897 59370 35990 59436
rect 35618 59235 35990 59311
rect 35618 59110 35711 59176
rect 35618 59094 35695 59110
tri 35695 59094 35711 59110 nw
rect 35747 59077 35861 59235
rect 35897 59110 35990 59176
tri 35897 59094 35913 59110 ne
rect 35913 59094 35990 59110
rect 35730 58995 35878 59077
rect 35618 58962 35695 58978
tri 35695 58962 35711 58978 sw
rect 35618 58896 35711 58962
rect 35618 58794 35711 58860
rect 35618 58778 35695 58794
tri 35695 58778 35711 58794 nw
rect 35747 58761 35861 58995
tri 35897 58962 35913 58978 se
rect 35913 58962 35990 58978
rect 35897 58896 35990 58962
rect 35897 58794 35990 58860
tri 35897 58778 35913 58794 ne
rect 35913 58778 35990 58794
rect 35730 58679 35878 58761
rect 35618 58646 35695 58662
tri 35695 58646 35711 58662 sw
rect 35618 58580 35711 58646
rect 35747 58521 35861 58679
tri 35897 58646 35913 58662 se
rect 35913 58646 35990 58662
rect 35897 58580 35990 58646
rect 35618 58445 35990 58521
rect 35618 58320 35711 58386
rect 35618 58304 35695 58320
tri 35695 58304 35711 58320 nw
rect 35747 58287 35861 58445
rect 35897 58320 35990 58386
tri 35897 58304 35913 58320 ne
rect 35913 58304 35990 58320
rect 35730 58205 35878 58287
rect 35618 58172 35695 58188
tri 35695 58172 35711 58188 sw
rect 35618 58106 35711 58172
rect 35618 58004 35711 58070
rect 35618 57988 35695 58004
tri 35695 57988 35711 58004 nw
rect 35747 57971 35861 58205
tri 35897 58172 35913 58188 se
rect 35913 58172 35990 58188
rect 35897 58106 35990 58172
rect 35897 58004 35990 58070
tri 35897 57988 35913 58004 ne
rect 35913 57988 35990 58004
rect 35730 57889 35878 57971
rect 35618 57856 35695 57872
tri 35695 57856 35711 57872 sw
rect 35618 57790 35711 57856
rect 35747 57731 35861 57889
tri 35897 57856 35913 57872 se
rect 35913 57856 35990 57872
rect 35897 57790 35990 57856
rect 35618 57655 35990 57731
rect 35618 57530 35711 57596
rect 35618 57514 35695 57530
tri 35695 57514 35711 57530 nw
rect 35747 57497 35861 57655
rect 35897 57530 35990 57596
tri 35897 57514 35913 57530 ne
rect 35913 57514 35990 57530
rect 35730 57415 35878 57497
rect 35618 57382 35695 57398
tri 35695 57382 35711 57398 sw
rect 35618 57316 35711 57382
rect 35618 57214 35711 57280
rect 35618 57198 35695 57214
tri 35695 57198 35711 57214 nw
rect 35747 57181 35861 57415
tri 35897 57382 35913 57398 se
rect 35913 57382 35990 57398
rect 35897 57316 35990 57382
rect 35897 57214 35990 57280
tri 35897 57198 35913 57214 ne
rect 35913 57198 35990 57214
rect 35730 57099 35878 57181
rect 35618 57066 35695 57082
tri 35695 57066 35711 57082 sw
rect 35618 57000 35711 57066
rect 35747 56941 35861 57099
tri 35897 57066 35913 57082 se
rect 35913 57066 35990 57082
rect 35897 57000 35990 57066
rect 35618 56865 35990 56941
rect 35618 56740 35711 56806
rect 35618 56724 35695 56740
tri 35695 56724 35711 56740 nw
rect 35747 56707 35861 56865
rect 35897 56740 35990 56806
tri 35897 56724 35913 56740 ne
rect 35913 56724 35990 56740
rect 35730 56625 35878 56707
rect 35618 56592 35695 56608
tri 35695 56592 35711 56608 sw
rect 35618 56526 35711 56592
rect 35618 56424 35711 56490
rect 35618 56408 35695 56424
tri 35695 56408 35711 56424 nw
rect 35747 56391 35861 56625
tri 35897 56592 35913 56608 se
rect 35913 56592 35990 56608
rect 35897 56526 35990 56592
rect 35897 56424 35990 56490
tri 35897 56408 35913 56424 ne
rect 35913 56408 35990 56424
rect 35730 56309 35878 56391
rect 35618 56276 35695 56292
tri 35695 56276 35711 56292 sw
rect 35618 56210 35711 56276
rect 35747 56151 35861 56309
tri 35897 56276 35913 56292 se
rect 35913 56276 35990 56292
rect 35897 56210 35990 56276
rect 35618 56075 35990 56151
rect 35618 55950 35711 56016
rect 35618 55934 35695 55950
tri 35695 55934 35711 55950 nw
rect 35747 55917 35861 56075
rect 35897 55950 35990 56016
tri 35897 55934 35913 55950 ne
rect 35913 55934 35990 55950
rect 35730 55835 35878 55917
rect 35618 55802 35695 55818
tri 35695 55802 35711 55818 sw
rect 35618 55736 35711 55802
rect 35618 55634 35711 55700
rect 35618 55618 35695 55634
tri 35695 55618 35711 55634 nw
rect 35747 55601 35861 55835
tri 35897 55802 35913 55818 se
rect 35913 55802 35990 55818
rect 35897 55736 35990 55802
rect 35897 55634 35990 55700
tri 35897 55618 35913 55634 ne
rect 35913 55618 35990 55634
rect 35730 55519 35878 55601
rect 35618 55486 35695 55502
tri 35695 55486 35711 55502 sw
rect 35618 55420 35711 55486
rect 35747 55361 35861 55519
tri 35897 55486 35913 55502 se
rect 35913 55486 35990 55502
rect 35897 55420 35990 55486
rect 35618 55285 35990 55361
rect 35618 55160 35711 55226
rect 35618 55144 35695 55160
tri 35695 55144 35711 55160 nw
rect 35747 55127 35861 55285
rect 35897 55160 35990 55226
tri 35897 55144 35913 55160 ne
rect 35913 55144 35990 55160
rect 35730 55045 35878 55127
rect 35618 55012 35695 55028
tri 35695 55012 35711 55028 sw
rect 35618 54946 35711 55012
rect 35618 54844 35711 54910
rect 35618 54828 35695 54844
tri 35695 54828 35711 54844 nw
rect 35747 54811 35861 55045
tri 35897 55012 35913 55028 se
rect 35913 55012 35990 55028
rect 35897 54946 35990 55012
rect 35897 54844 35990 54910
tri 35897 54828 35913 54844 ne
rect 35913 54828 35990 54844
rect 35730 54729 35878 54811
rect 35618 54696 35695 54712
tri 35695 54696 35711 54712 sw
rect 35618 54630 35711 54696
rect 35747 54571 35861 54729
tri 35897 54696 35913 54712 se
rect 35913 54696 35990 54712
rect 35897 54630 35990 54696
rect 35618 54495 35990 54571
rect 35618 54370 35711 54436
rect 35618 54354 35695 54370
tri 35695 54354 35711 54370 nw
rect 35747 54337 35861 54495
rect 35897 54370 35990 54436
tri 35897 54354 35913 54370 ne
rect 35913 54354 35990 54370
rect 35730 54255 35878 54337
rect 35618 54222 35695 54238
tri 35695 54222 35711 54238 sw
rect 35618 54156 35711 54222
rect 35618 54054 35711 54120
rect 35618 54038 35695 54054
tri 35695 54038 35711 54054 nw
rect 35747 54021 35861 54255
tri 35897 54222 35913 54238 se
rect 35913 54222 35990 54238
rect 35897 54156 35990 54222
rect 35897 54054 35990 54120
tri 35897 54038 35913 54054 ne
rect 35913 54038 35990 54054
rect 35730 53939 35878 54021
rect 35618 53906 35695 53922
tri 35695 53906 35711 53922 sw
rect 35618 53840 35711 53906
rect 35747 53781 35861 53939
tri 35897 53906 35913 53922 se
rect 35913 53906 35990 53922
rect 35897 53840 35990 53906
rect 35618 53705 35990 53781
rect 35618 53580 35711 53646
rect 35618 53564 35695 53580
tri 35695 53564 35711 53580 nw
rect 35747 53547 35861 53705
rect 35897 53580 35990 53646
tri 35897 53564 35913 53580 ne
rect 35913 53564 35990 53580
rect 35730 53465 35878 53547
rect 35618 53432 35695 53448
tri 35695 53432 35711 53448 sw
rect 35618 53366 35711 53432
rect 35618 53264 35711 53330
rect 35618 53248 35695 53264
tri 35695 53248 35711 53264 nw
rect 35747 53231 35861 53465
tri 35897 53432 35913 53448 se
rect 35913 53432 35990 53448
rect 35897 53366 35990 53432
rect 35897 53264 35990 53330
tri 35897 53248 35913 53264 ne
rect 35913 53248 35990 53264
rect 35730 53149 35878 53231
rect 35618 53116 35695 53132
tri 35695 53116 35711 53132 sw
rect 35618 53050 35711 53116
rect 35747 52991 35861 53149
tri 35897 53116 35913 53132 se
rect 35913 53116 35990 53132
rect 35897 53050 35990 53116
rect 35618 52915 35990 52991
rect 35618 52790 35711 52856
rect 35618 52774 35695 52790
tri 35695 52774 35711 52790 nw
rect 35747 52757 35861 52915
rect 35897 52790 35990 52856
tri 35897 52774 35913 52790 ne
rect 35913 52774 35990 52790
rect 35730 52675 35878 52757
rect 35618 52642 35695 52658
tri 35695 52642 35711 52658 sw
rect 35618 52576 35711 52642
rect 35618 52474 35711 52540
rect 35618 52458 35695 52474
tri 35695 52458 35711 52474 nw
rect 35747 52441 35861 52675
tri 35897 52642 35913 52658 se
rect 35913 52642 35990 52658
rect 35897 52576 35990 52642
rect 35897 52474 35990 52540
tri 35897 52458 35913 52474 ne
rect 35913 52458 35990 52474
rect 35730 52359 35878 52441
rect 35618 52326 35695 52342
tri 35695 52326 35711 52342 sw
rect 35618 52260 35711 52326
rect 35747 52201 35861 52359
tri 35897 52326 35913 52342 se
rect 35913 52326 35990 52342
rect 35897 52260 35990 52326
rect 35618 52125 35990 52201
rect 35618 52000 35711 52066
rect 35618 51984 35695 52000
tri 35695 51984 35711 52000 nw
rect 35747 51967 35861 52125
rect 35897 52000 35990 52066
tri 35897 51984 35913 52000 ne
rect 35913 51984 35990 52000
rect 35730 51885 35878 51967
rect 35618 51852 35695 51868
tri 35695 51852 35711 51868 sw
rect 35618 51786 35711 51852
rect 35618 51684 35711 51750
rect 35618 51668 35695 51684
tri 35695 51668 35711 51684 nw
rect 35747 51651 35861 51885
tri 35897 51852 35913 51868 se
rect 35913 51852 35990 51868
rect 35897 51786 35990 51852
rect 35897 51684 35990 51750
tri 35897 51668 35913 51684 ne
rect 35913 51668 35990 51684
rect 35730 51569 35878 51651
rect 35618 51536 35695 51552
tri 35695 51536 35711 51552 sw
rect 35618 51470 35711 51536
rect 35747 51411 35861 51569
tri 35897 51536 35913 51552 se
rect 35913 51536 35990 51552
rect 35897 51470 35990 51536
rect 35618 51335 35990 51411
rect 35618 51210 35711 51276
rect 35618 51194 35695 51210
tri 35695 51194 35711 51210 nw
rect 35747 51177 35861 51335
rect 35897 51210 35990 51276
tri 35897 51194 35913 51210 ne
rect 35913 51194 35990 51210
rect 35730 51095 35878 51177
rect 35618 51062 35695 51078
tri 35695 51062 35711 51078 sw
rect 35618 50996 35711 51062
rect 35618 50894 35711 50960
rect 35618 50878 35695 50894
tri 35695 50878 35711 50894 nw
rect 35747 50861 35861 51095
tri 35897 51062 35913 51078 se
rect 35913 51062 35990 51078
rect 35897 50996 35990 51062
rect 35897 50894 35990 50960
tri 35897 50878 35913 50894 ne
rect 35913 50878 35990 50894
rect 35730 50779 35878 50861
rect 35618 50746 35695 50762
tri 35695 50746 35711 50762 sw
rect 35618 50680 35711 50746
rect 35747 50621 35861 50779
tri 35897 50746 35913 50762 se
rect 35913 50746 35990 50762
rect 35897 50680 35990 50746
rect 35618 50545 35990 50621
rect 35618 50420 35711 50486
rect 35618 50404 35695 50420
tri 35695 50404 35711 50420 nw
rect 35747 50387 35861 50545
rect 35897 50420 35990 50486
tri 35897 50404 35913 50420 ne
rect 35913 50404 35990 50420
rect 35730 50305 35878 50387
rect 35618 50272 35695 50288
tri 35695 50272 35711 50288 sw
rect 35618 50206 35711 50272
rect 35618 50104 35711 50170
rect 35618 50088 35695 50104
tri 35695 50088 35711 50104 nw
rect 35747 50071 35861 50305
tri 35897 50272 35913 50288 se
rect 35913 50272 35990 50288
rect 35897 50206 35990 50272
rect 35897 50104 35990 50170
tri 35897 50088 35913 50104 ne
rect 35913 50088 35990 50104
rect 35730 49989 35878 50071
rect 35618 49956 35695 49972
tri 35695 49956 35711 49972 sw
rect 35618 49890 35711 49956
rect 35747 49831 35861 49989
tri 35897 49956 35913 49972 se
rect 35913 49956 35990 49972
rect 35897 49890 35990 49956
rect 35618 49755 35990 49831
rect 35618 49630 35711 49696
rect 35618 49614 35695 49630
tri 35695 49614 35711 49630 nw
rect 35747 49597 35861 49755
rect 35897 49630 35990 49696
tri 35897 49614 35913 49630 ne
rect 35913 49614 35990 49630
rect 35730 49515 35878 49597
rect 35618 49482 35695 49498
tri 35695 49482 35711 49498 sw
rect 35618 49416 35711 49482
rect 35618 49314 35711 49380
rect 35618 49298 35695 49314
tri 35695 49298 35711 49314 nw
rect 35747 49281 35861 49515
tri 35897 49482 35913 49498 se
rect 35913 49482 35990 49498
rect 35897 49416 35990 49482
rect 35897 49314 35990 49380
tri 35897 49298 35913 49314 ne
rect 35913 49298 35990 49314
rect 35730 49199 35878 49281
rect 35618 49166 35695 49182
tri 35695 49166 35711 49182 sw
rect 35618 49100 35711 49166
rect 35747 49041 35861 49199
tri 35897 49166 35913 49182 se
rect 35913 49166 35990 49182
rect 35897 49100 35990 49166
rect 35618 48965 35990 49041
rect 35618 48840 35711 48906
rect 35618 48824 35695 48840
tri 35695 48824 35711 48840 nw
rect 35747 48807 35861 48965
rect 35897 48840 35990 48906
tri 35897 48824 35913 48840 ne
rect 35913 48824 35990 48840
rect 35730 48725 35878 48807
rect 35618 48692 35695 48708
tri 35695 48692 35711 48708 sw
rect 35618 48626 35711 48692
rect 35618 48524 35711 48590
rect 35618 48508 35695 48524
tri 35695 48508 35711 48524 nw
rect 35747 48491 35861 48725
tri 35897 48692 35913 48708 se
rect 35913 48692 35990 48708
rect 35897 48626 35990 48692
rect 35897 48524 35990 48590
tri 35897 48508 35913 48524 ne
rect 35913 48508 35990 48524
rect 35730 48409 35878 48491
rect 35618 48376 35695 48392
tri 35695 48376 35711 48392 sw
rect 35618 48310 35711 48376
rect 35747 48251 35861 48409
tri 35897 48376 35913 48392 se
rect 35913 48376 35990 48392
rect 35897 48310 35990 48376
rect 35618 48175 35990 48251
rect 35618 48050 35711 48116
rect 35618 48034 35695 48050
tri 35695 48034 35711 48050 nw
rect 35747 48017 35861 48175
rect 35897 48050 35990 48116
tri 35897 48034 35913 48050 ne
rect 35913 48034 35990 48050
rect 35730 47935 35878 48017
rect 35618 47902 35695 47918
tri 35695 47902 35711 47918 sw
rect 35618 47836 35711 47902
rect 35618 47734 35711 47800
rect 35618 47718 35695 47734
tri 35695 47718 35711 47734 nw
rect 35747 47701 35861 47935
tri 35897 47902 35913 47918 se
rect 35913 47902 35990 47918
rect 35897 47836 35990 47902
rect 35897 47734 35990 47800
tri 35897 47718 35913 47734 ne
rect 35913 47718 35990 47734
rect 35730 47619 35878 47701
rect 35618 47586 35695 47602
tri 35695 47586 35711 47602 sw
rect 35618 47520 35711 47586
rect 35747 47461 35861 47619
tri 35897 47586 35913 47602 se
rect 35913 47586 35990 47602
rect 35897 47520 35990 47586
rect 35618 47385 35990 47461
rect 35618 47260 35711 47326
rect 35618 47244 35695 47260
tri 35695 47244 35711 47260 nw
rect 35747 47227 35861 47385
rect 35897 47260 35990 47326
tri 35897 47244 35913 47260 ne
rect 35913 47244 35990 47260
rect 35730 47145 35878 47227
rect 35618 47112 35695 47128
tri 35695 47112 35711 47128 sw
rect 35618 47046 35711 47112
rect 35618 46944 35711 47010
rect 35618 46928 35695 46944
tri 35695 46928 35711 46944 nw
rect 35747 46911 35861 47145
tri 35897 47112 35913 47128 se
rect 35913 47112 35990 47128
rect 35897 47046 35990 47112
rect 35897 46944 35990 47010
tri 35897 46928 35913 46944 ne
rect 35913 46928 35990 46944
rect 35730 46829 35878 46911
rect 35618 46796 35695 46812
tri 35695 46796 35711 46812 sw
rect 35618 46730 35711 46796
rect 35747 46671 35861 46829
tri 35897 46796 35913 46812 se
rect 35913 46796 35990 46812
rect 35897 46730 35990 46796
rect 35618 46595 35990 46671
rect 35618 46470 35711 46536
rect 35618 46454 35695 46470
tri 35695 46454 35711 46470 nw
rect 35747 46437 35861 46595
rect 35897 46470 35990 46536
tri 35897 46454 35913 46470 ne
rect 35913 46454 35990 46470
rect 35730 46355 35878 46437
rect 35618 46322 35695 46338
tri 35695 46322 35711 46338 sw
rect 35618 46256 35711 46322
rect 35618 46154 35711 46220
rect 35618 46138 35695 46154
tri 35695 46138 35711 46154 nw
rect 35747 46121 35861 46355
tri 35897 46322 35913 46338 se
rect 35913 46322 35990 46338
rect 35897 46256 35990 46322
rect 35897 46154 35990 46220
tri 35897 46138 35913 46154 ne
rect 35913 46138 35990 46154
rect 35730 46039 35878 46121
rect 35618 46006 35695 46022
tri 35695 46006 35711 46022 sw
rect 35618 45940 35711 46006
rect 35747 45881 35861 46039
tri 35897 46006 35913 46022 se
rect 35913 46006 35990 46022
rect 35897 45940 35990 46006
rect 35618 45805 35990 45881
rect 35618 45680 35711 45746
rect 35618 45664 35695 45680
tri 35695 45664 35711 45680 nw
rect 35747 45647 35861 45805
rect 35897 45680 35990 45746
tri 35897 45664 35913 45680 ne
rect 35913 45664 35990 45680
rect 35730 45565 35878 45647
rect 35618 45532 35695 45548
tri 35695 45532 35711 45548 sw
rect 35618 45466 35711 45532
rect 35618 45364 35711 45430
rect 35618 45348 35695 45364
tri 35695 45348 35711 45364 nw
rect 35747 45331 35861 45565
tri 35897 45532 35913 45548 se
rect 35913 45532 35990 45548
rect 35897 45466 35990 45532
rect 35897 45364 35990 45430
tri 35897 45348 35913 45364 ne
rect 35913 45348 35990 45364
rect 35730 45249 35878 45331
rect 35618 45216 35695 45232
tri 35695 45216 35711 45232 sw
rect 35618 45150 35711 45216
rect 35747 45091 35861 45249
tri 35897 45216 35913 45232 se
rect 35913 45216 35990 45232
rect 35897 45150 35990 45216
rect 35618 45015 35990 45091
rect 35618 44890 35711 44956
rect 35618 44874 35695 44890
tri 35695 44874 35711 44890 nw
rect 35747 44857 35861 45015
rect 35897 44890 35990 44956
tri 35897 44874 35913 44890 ne
rect 35913 44874 35990 44890
rect 35730 44775 35878 44857
rect 35618 44742 35695 44758
tri 35695 44742 35711 44758 sw
rect 35618 44676 35711 44742
rect 35618 44574 35711 44640
rect 35618 44558 35695 44574
tri 35695 44558 35711 44574 nw
rect 35747 44541 35861 44775
tri 35897 44742 35913 44758 se
rect 35913 44742 35990 44758
rect 35897 44676 35990 44742
rect 35897 44574 35990 44640
tri 35897 44558 35913 44574 ne
rect 35913 44558 35990 44574
rect 35730 44459 35878 44541
rect 35618 44426 35695 44442
tri 35695 44426 35711 44442 sw
rect 35618 44360 35711 44426
rect 35747 44301 35861 44459
tri 35897 44426 35913 44442 se
rect 35913 44426 35990 44442
rect 35897 44360 35990 44426
rect 35618 44225 35990 44301
rect 35618 44100 35711 44166
rect 35618 44084 35695 44100
tri 35695 44084 35711 44100 nw
rect 35747 44067 35861 44225
rect 35897 44100 35990 44166
tri 35897 44084 35913 44100 ne
rect 35913 44084 35990 44100
rect 35730 43985 35878 44067
rect 35618 43952 35695 43968
tri 35695 43952 35711 43968 sw
rect 35618 43886 35711 43952
rect 35618 43784 35711 43850
rect 35618 43768 35695 43784
tri 35695 43768 35711 43784 nw
rect 35747 43751 35861 43985
tri 35897 43952 35913 43968 se
rect 35913 43952 35990 43968
rect 35897 43886 35990 43952
rect 35897 43784 35990 43850
tri 35897 43768 35913 43784 ne
rect 35913 43768 35990 43784
rect 35730 43669 35878 43751
rect 35618 43636 35695 43652
tri 35695 43636 35711 43652 sw
rect 35618 43570 35711 43636
rect 35747 43511 35861 43669
tri 35897 43636 35913 43652 se
rect 35913 43636 35990 43652
rect 35897 43570 35990 43636
rect 35618 43435 35990 43511
rect 35618 43310 35711 43376
rect 35618 43294 35695 43310
tri 35695 43294 35711 43310 nw
rect 35747 43277 35861 43435
rect 35897 43310 35990 43376
tri 35897 43294 35913 43310 ne
rect 35913 43294 35990 43310
rect 35730 43195 35878 43277
rect 35618 43162 35695 43178
tri 35695 43162 35711 43178 sw
rect 35618 43096 35711 43162
rect 35618 42994 35711 43060
rect 35618 42978 35695 42994
tri 35695 42978 35711 42994 nw
rect 35747 42961 35861 43195
tri 35897 43162 35913 43178 se
rect 35913 43162 35990 43178
rect 35897 43096 35990 43162
rect 35897 42994 35990 43060
tri 35897 42978 35913 42994 ne
rect 35913 42978 35990 42994
rect 35730 42879 35878 42961
rect 35618 42846 35695 42862
tri 35695 42846 35711 42862 sw
rect 35618 42780 35711 42846
rect 35747 42721 35861 42879
tri 35897 42846 35913 42862 se
rect 35913 42846 35990 42862
rect 35897 42780 35990 42846
rect 35618 42645 35990 42721
rect 35618 42520 35711 42586
rect 35618 42504 35695 42520
tri 35695 42504 35711 42520 nw
rect 35747 42487 35861 42645
rect 35897 42520 35990 42586
tri 35897 42504 35913 42520 ne
rect 35913 42504 35990 42520
rect 35730 42405 35878 42487
rect 35618 42372 35695 42388
tri 35695 42372 35711 42388 sw
rect 35618 42306 35711 42372
rect 35618 42204 35711 42270
rect 35618 42188 35695 42204
tri 35695 42188 35711 42204 nw
rect 35747 42171 35861 42405
tri 35897 42372 35913 42388 se
rect 35913 42372 35990 42388
rect 35897 42306 35990 42372
rect 35897 42204 35990 42270
tri 35897 42188 35913 42204 ne
rect 35913 42188 35990 42204
rect 35730 42089 35878 42171
rect 35618 42056 35695 42072
tri 35695 42056 35711 42072 sw
rect 35618 41990 35711 42056
rect 35747 41931 35861 42089
tri 35897 42056 35913 42072 se
rect 35913 42056 35990 42072
rect 35897 41990 35990 42056
rect 35618 41855 35990 41931
rect 35618 41730 35711 41796
rect 35618 41714 35695 41730
tri 35695 41714 35711 41730 nw
rect 35747 41697 35861 41855
rect 35897 41730 35990 41796
tri 35897 41714 35913 41730 ne
rect 35913 41714 35990 41730
rect 35730 41615 35878 41697
rect 35618 41582 35695 41598
tri 35695 41582 35711 41598 sw
rect 35618 41516 35711 41582
rect 35618 41414 35711 41480
rect 35618 41398 35695 41414
tri 35695 41398 35711 41414 nw
rect 35747 41381 35861 41615
tri 35897 41582 35913 41598 se
rect 35913 41582 35990 41598
rect 35897 41516 35990 41582
rect 35897 41414 35990 41480
tri 35897 41398 35913 41414 ne
rect 35913 41398 35990 41414
rect 35730 41299 35878 41381
rect 35618 41266 35695 41282
tri 35695 41266 35711 41282 sw
rect 35618 41200 35711 41266
rect 35747 41141 35861 41299
tri 35897 41266 35913 41282 se
rect 35913 41266 35990 41282
rect 35897 41200 35990 41266
rect 35618 41065 35990 41141
rect 35618 40940 35711 41006
rect 35618 40924 35695 40940
tri 35695 40924 35711 40940 nw
rect 35747 40907 35861 41065
rect 35897 40940 35990 41006
tri 35897 40924 35913 40940 ne
rect 35913 40924 35990 40940
rect 35730 40825 35878 40907
rect 35618 40792 35695 40808
tri 35695 40792 35711 40808 sw
rect 35618 40726 35711 40792
rect 35618 40624 35711 40690
rect 35618 40608 35695 40624
tri 35695 40608 35711 40624 nw
rect 35747 40591 35861 40825
tri 35897 40792 35913 40808 se
rect 35913 40792 35990 40808
rect 35897 40726 35990 40792
rect 35897 40624 35990 40690
tri 35897 40608 35913 40624 ne
rect 35913 40608 35990 40624
rect 35730 40509 35878 40591
rect 35618 40476 35695 40492
tri 35695 40476 35711 40492 sw
rect 35618 40410 35711 40476
rect 35747 40351 35861 40509
tri 35897 40476 35913 40492 se
rect 35913 40476 35990 40492
rect 35897 40410 35990 40476
rect 35618 40275 35990 40351
rect 35618 40150 35711 40216
rect 35618 40134 35695 40150
tri 35695 40134 35711 40150 nw
rect 35747 40117 35861 40275
rect 35897 40150 35990 40216
tri 35897 40134 35913 40150 ne
rect 35913 40134 35990 40150
rect 35730 40035 35878 40117
rect 35618 40002 35695 40018
tri 35695 40002 35711 40018 sw
rect 35618 39936 35711 40002
rect 35618 39834 35711 39900
rect 35618 39818 35695 39834
tri 35695 39818 35711 39834 nw
rect 35747 39801 35861 40035
tri 35897 40002 35913 40018 se
rect 35913 40002 35990 40018
rect 35897 39936 35990 40002
rect 35897 39834 35990 39900
tri 35897 39818 35913 39834 ne
rect 35913 39818 35990 39834
rect 35730 39719 35878 39801
rect 35618 39686 35695 39702
tri 35695 39686 35711 39702 sw
rect 35618 39620 35711 39686
rect 35747 39561 35861 39719
tri 35897 39686 35913 39702 se
rect 35913 39686 35990 39702
rect 35897 39620 35990 39686
rect 35618 39485 35990 39561
rect 35618 39360 35711 39426
rect 35618 39344 35695 39360
tri 35695 39344 35711 39360 nw
rect 35747 39327 35861 39485
rect 35897 39360 35990 39426
tri 35897 39344 35913 39360 ne
rect 35913 39344 35990 39360
rect 35730 39245 35878 39327
rect 35618 39212 35695 39228
tri 35695 39212 35711 39228 sw
rect 35618 39146 35711 39212
rect 35618 39044 35711 39110
rect 35618 39028 35695 39044
tri 35695 39028 35711 39044 nw
rect 35747 39011 35861 39245
tri 35897 39212 35913 39228 se
rect 35913 39212 35990 39228
rect 35897 39146 35990 39212
rect 35897 39044 35990 39110
tri 35897 39028 35913 39044 ne
rect 35913 39028 35990 39044
rect 35730 38929 35878 39011
rect 35618 38896 35695 38912
tri 35695 38896 35711 38912 sw
rect 35618 38830 35711 38896
rect 35747 38771 35861 38929
tri 35897 38896 35913 38912 se
rect 35913 38896 35990 38912
rect 35897 38830 35990 38896
rect 35618 38695 35990 38771
rect 35618 38570 35711 38636
rect 35618 38554 35695 38570
tri 35695 38554 35711 38570 nw
rect 35747 38537 35861 38695
rect 35897 38570 35990 38636
tri 35897 38554 35913 38570 ne
rect 35913 38554 35990 38570
rect 35730 38455 35878 38537
rect 35618 38422 35695 38438
tri 35695 38422 35711 38438 sw
rect 35618 38356 35711 38422
rect 35618 38254 35711 38320
rect 35618 38238 35695 38254
tri 35695 38238 35711 38254 nw
rect 35747 38221 35861 38455
tri 35897 38422 35913 38438 se
rect 35913 38422 35990 38438
rect 35897 38356 35990 38422
rect 35897 38254 35990 38320
tri 35897 38238 35913 38254 ne
rect 35913 38238 35990 38254
rect 35730 38139 35878 38221
rect 35618 38106 35695 38122
tri 35695 38106 35711 38122 sw
rect 35618 38040 35711 38106
rect 35747 37981 35861 38139
tri 35897 38106 35913 38122 se
rect 35913 38106 35990 38122
rect 35897 38040 35990 38106
rect 35618 37905 35990 37981
rect 35618 37780 35711 37846
rect 35618 37764 35695 37780
tri 35695 37764 35711 37780 nw
rect 35747 37747 35861 37905
rect 35897 37780 35990 37846
tri 35897 37764 35913 37780 ne
rect 35913 37764 35990 37780
rect 35730 37665 35878 37747
rect 35618 37632 35695 37648
tri 35695 37632 35711 37648 sw
rect 35618 37566 35711 37632
rect 35618 37464 35711 37530
rect 35618 37448 35695 37464
tri 35695 37448 35711 37464 nw
rect 35747 37431 35861 37665
tri 35897 37632 35913 37648 se
rect 35913 37632 35990 37648
rect 35897 37566 35990 37632
rect 35897 37464 35990 37530
tri 35897 37448 35913 37464 ne
rect 35913 37448 35990 37464
rect 35730 37349 35878 37431
rect 35618 37316 35695 37332
tri 35695 37316 35711 37332 sw
rect 35618 37250 35711 37316
rect 35747 37191 35861 37349
tri 35897 37316 35913 37332 se
rect 35913 37316 35990 37332
rect 35897 37250 35990 37316
rect 35618 37115 35990 37191
rect 35618 36990 35711 37056
rect 35618 36974 35695 36990
tri 35695 36974 35711 36990 nw
rect 35747 36957 35861 37115
rect 35897 36990 35990 37056
tri 35897 36974 35913 36990 ne
rect 35913 36974 35990 36990
rect 35730 36875 35878 36957
rect 35618 36842 35695 36858
tri 35695 36842 35711 36858 sw
rect 35618 36776 35711 36842
rect 35618 36674 35711 36740
rect 35618 36658 35695 36674
tri 35695 36658 35711 36674 nw
rect 35747 36641 35861 36875
tri 35897 36842 35913 36858 se
rect 35913 36842 35990 36858
rect 35897 36776 35990 36842
rect 35897 36674 35990 36740
tri 35897 36658 35913 36674 ne
rect 35913 36658 35990 36674
rect 35730 36559 35878 36641
rect 35618 36526 35695 36542
tri 35695 36526 35711 36542 sw
rect 35618 36460 35711 36526
rect 35747 36401 35861 36559
tri 35897 36526 35913 36542 se
rect 35913 36526 35990 36542
rect 35897 36460 35990 36526
rect 35618 36325 35990 36401
rect 35618 36200 35711 36266
rect 35618 36184 35695 36200
tri 35695 36184 35711 36200 nw
rect 35747 36167 35861 36325
rect 35897 36200 35990 36266
tri 35897 36184 35913 36200 ne
rect 35913 36184 35990 36200
rect 35730 36085 35878 36167
rect 35618 36052 35695 36068
tri 35695 36052 35711 36068 sw
rect 35618 35986 35711 36052
rect 35618 35884 35711 35950
rect 35618 35868 35695 35884
tri 35695 35868 35711 35884 nw
rect 35747 35851 35861 36085
tri 35897 36052 35913 36068 se
rect 35913 36052 35990 36068
rect 35897 35986 35990 36052
rect 35897 35884 35990 35950
tri 35897 35868 35913 35884 ne
rect 35913 35868 35990 35884
rect 35730 35769 35878 35851
rect 35618 35736 35695 35752
tri 35695 35736 35711 35752 sw
rect 35618 35670 35711 35736
rect 35747 35611 35861 35769
tri 35897 35736 35913 35752 se
rect 35913 35736 35990 35752
rect 35897 35670 35990 35736
rect 35618 35535 35990 35611
rect 35618 35410 35711 35476
rect 35618 35394 35695 35410
tri 35695 35394 35711 35410 nw
rect 35747 35377 35861 35535
rect 35897 35410 35990 35476
tri 35897 35394 35913 35410 ne
rect 35913 35394 35990 35410
rect 35730 35295 35878 35377
rect 35618 35262 35695 35278
tri 35695 35262 35711 35278 sw
rect 35618 35196 35711 35262
rect 35618 35094 35711 35160
rect 35618 35078 35695 35094
tri 35695 35078 35711 35094 nw
rect 35747 35061 35861 35295
tri 35897 35262 35913 35278 se
rect 35913 35262 35990 35278
rect 35897 35196 35990 35262
rect 35897 35094 35990 35160
tri 35897 35078 35913 35094 ne
rect 35913 35078 35990 35094
rect 35730 34979 35878 35061
rect 35618 34946 35695 34962
tri 35695 34946 35711 34962 sw
rect 35618 34880 35711 34946
rect 35747 34821 35861 34979
tri 35897 34946 35913 34962 se
rect 35913 34946 35990 34962
rect 35897 34880 35990 34946
rect 35618 34745 35990 34821
rect 35618 34620 35711 34686
rect 35618 34604 35695 34620
tri 35695 34604 35711 34620 nw
rect 35747 34587 35861 34745
rect 35897 34620 35990 34686
tri 35897 34604 35913 34620 ne
rect 35913 34604 35990 34620
rect 35730 34505 35878 34587
rect 35618 34472 35695 34488
tri 35695 34472 35711 34488 sw
rect 35618 34406 35711 34472
rect 35618 34304 35711 34370
rect 35618 34288 35695 34304
tri 35695 34288 35711 34304 nw
rect 35747 34271 35861 34505
tri 35897 34472 35913 34488 se
rect 35913 34472 35990 34488
rect 35897 34406 35990 34472
rect 35897 34304 35990 34370
tri 35897 34288 35913 34304 ne
rect 35913 34288 35990 34304
rect 35730 34189 35878 34271
rect 35618 34156 35695 34172
tri 35695 34156 35711 34172 sw
rect 35618 34090 35711 34156
rect 35747 34031 35861 34189
tri 35897 34156 35913 34172 se
rect 35913 34156 35990 34172
rect 35897 34090 35990 34156
rect 35618 33955 35990 34031
rect 35618 33830 35711 33896
rect 35618 33814 35695 33830
tri 35695 33814 35711 33830 nw
rect 35747 33797 35861 33955
rect 35897 33830 35990 33896
tri 35897 33814 35913 33830 ne
rect 35913 33814 35990 33830
rect 35730 33715 35878 33797
rect 35618 33682 35695 33698
tri 35695 33682 35711 33698 sw
rect 35618 33616 35711 33682
rect 35618 33514 35711 33580
rect 35618 33498 35695 33514
tri 35695 33498 35711 33514 nw
rect 35747 33481 35861 33715
tri 35897 33682 35913 33698 se
rect 35913 33682 35990 33698
rect 35897 33616 35990 33682
rect 35897 33514 35990 33580
tri 35897 33498 35913 33514 ne
rect 35913 33498 35990 33514
rect 35730 33399 35878 33481
rect 35618 33366 35695 33382
tri 35695 33366 35711 33382 sw
rect 35618 33300 35711 33366
rect 35747 33241 35861 33399
tri 35897 33366 35913 33382 se
rect 35913 33366 35990 33382
rect 35897 33300 35990 33366
rect 35618 33165 35990 33241
rect 35618 33040 35711 33106
rect 35618 33024 35695 33040
tri 35695 33024 35711 33040 nw
rect 35747 33007 35861 33165
rect 35897 33040 35990 33106
tri 35897 33024 35913 33040 ne
rect 35913 33024 35990 33040
rect 35730 32925 35878 33007
rect 35618 32892 35695 32908
tri 35695 32892 35711 32908 sw
rect 35618 32826 35711 32892
rect 35618 32724 35711 32790
rect 35618 32708 35695 32724
tri 35695 32708 35711 32724 nw
rect 35747 32691 35861 32925
tri 35897 32892 35913 32908 se
rect 35913 32892 35990 32908
rect 35897 32826 35990 32892
rect 35897 32724 35990 32790
tri 35897 32708 35913 32724 ne
rect 35913 32708 35990 32724
rect 35730 32609 35878 32691
rect 35618 32576 35695 32592
tri 35695 32576 35711 32592 sw
rect 35618 32510 35711 32576
rect 35747 32451 35861 32609
tri 35897 32576 35913 32592 se
rect 35913 32576 35990 32592
rect 35897 32510 35990 32576
rect 35618 32375 35990 32451
rect 35618 32250 35711 32316
rect 35618 32234 35695 32250
tri 35695 32234 35711 32250 nw
rect 35747 32217 35861 32375
rect 35897 32250 35990 32316
tri 35897 32234 35913 32250 ne
rect 35913 32234 35990 32250
rect 35730 32135 35878 32217
rect 35618 32102 35695 32118
tri 35695 32102 35711 32118 sw
rect 35618 32036 35711 32102
rect 35618 31934 35711 32000
rect 35618 31918 35695 31934
tri 35695 31918 35711 31934 nw
rect 35747 31901 35861 32135
tri 35897 32102 35913 32118 se
rect 35913 32102 35990 32118
rect 35897 32036 35990 32102
rect 35897 31934 35990 32000
tri 35897 31918 35913 31934 ne
rect 35913 31918 35990 31934
rect 35730 31819 35878 31901
rect 35618 31786 35695 31802
tri 35695 31786 35711 31802 sw
rect 35618 31720 35711 31786
rect 35747 31661 35861 31819
tri 35897 31786 35913 31802 se
rect 35913 31786 35990 31802
rect 35897 31720 35990 31786
rect 35618 31585 35990 31661
rect 35618 31460 35711 31526
rect 35618 31444 35695 31460
tri 35695 31444 35711 31460 nw
rect 35747 31427 35861 31585
rect 35897 31460 35990 31526
tri 35897 31444 35913 31460 ne
rect 35913 31444 35990 31460
rect 35730 31345 35878 31427
rect 35618 31312 35695 31328
tri 35695 31312 35711 31328 sw
rect 35618 31246 35711 31312
rect 35618 31144 35711 31210
rect 35618 31128 35695 31144
tri 35695 31128 35711 31144 nw
rect 35747 31111 35861 31345
tri 35897 31312 35913 31328 se
rect 35913 31312 35990 31328
rect 35897 31246 35990 31312
rect 35897 31144 35990 31210
tri 35897 31128 35913 31144 ne
rect 35913 31128 35990 31144
rect 35730 31029 35878 31111
rect 35618 30996 35695 31012
tri 35695 30996 35711 31012 sw
rect 35618 30930 35711 30996
rect 35747 30871 35861 31029
tri 35897 30996 35913 31012 se
rect 35913 30996 35990 31012
rect 35897 30930 35990 30996
rect 35618 30795 35990 30871
rect 35618 30670 35711 30736
rect 35618 30654 35695 30670
tri 35695 30654 35711 30670 nw
rect 35747 30637 35861 30795
rect 35897 30670 35990 30736
tri 35897 30654 35913 30670 ne
rect 35913 30654 35990 30670
rect 35730 30555 35878 30637
rect 35618 30522 35695 30538
tri 35695 30522 35711 30538 sw
rect 35618 30456 35711 30522
rect 35618 30354 35711 30420
rect 35618 30338 35695 30354
tri 35695 30338 35711 30354 nw
rect 35747 30321 35861 30555
tri 35897 30522 35913 30538 se
rect 35913 30522 35990 30538
rect 35897 30456 35990 30522
rect 35897 30354 35990 30420
tri 35897 30338 35913 30354 ne
rect 35913 30338 35990 30354
rect 35730 30239 35878 30321
rect 35618 30206 35695 30222
tri 35695 30206 35711 30222 sw
rect 35618 30140 35711 30206
rect 35747 30081 35861 30239
tri 35897 30206 35913 30222 se
rect 35913 30206 35990 30222
rect 35897 30140 35990 30206
rect 35618 30005 35990 30081
rect 35618 29880 35711 29946
rect 35618 29864 35695 29880
tri 35695 29864 35711 29880 nw
rect 35747 29847 35861 30005
rect 35897 29880 35990 29946
tri 35897 29864 35913 29880 ne
rect 35913 29864 35990 29880
rect 35730 29765 35878 29847
rect 35618 29732 35695 29748
tri 35695 29732 35711 29748 sw
rect 35618 29666 35711 29732
rect 35618 29564 35711 29630
rect 35618 29548 35695 29564
tri 35695 29548 35711 29564 nw
rect 35747 29531 35861 29765
tri 35897 29732 35913 29748 se
rect 35913 29732 35990 29748
rect 35897 29666 35990 29732
rect 35897 29564 35990 29630
tri 35897 29548 35913 29564 ne
rect 35913 29548 35990 29564
rect 35730 29449 35878 29531
rect 35618 29416 35695 29432
tri 35695 29416 35711 29432 sw
rect 35618 29350 35711 29416
rect 35747 29291 35861 29449
tri 35897 29416 35913 29432 se
rect 35913 29416 35990 29432
rect 35897 29350 35990 29416
rect 35618 29215 35990 29291
rect 35618 29090 35711 29156
rect 35618 29074 35695 29090
tri 35695 29074 35711 29090 nw
rect 35747 29057 35861 29215
rect 35897 29090 35990 29156
tri 35897 29074 35913 29090 ne
rect 35913 29074 35990 29090
rect 35730 28975 35878 29057
rect 35618 28942 35695 28958
tri 35695 28942 35711 28958 sw
rect 35618 28876 35711 28942
rect 35747 28833 35861 28975
tri 35897 28942 35913 28958 se
rect 35913 28942 35990 28958
rect 35897 28876 35990 28942
rect 36026 28463 36062 80603
rect 36098 28463 36134 80603
rect 36170 80445 36206 80603
rect 36162 80303 36214 80445
rect 36170 28763 36206 80303
rect 36162 28621 36214 28763
rect 36170 28463 36206 28621
rect 36242 28463 36278 80603
rect 36314 28463 36350 80603
rect 36386 28833 36470 80233
rect 36506 28463 36542 80603
rect 36578 28463 36614 80603
rect 36650 80445 36686 80603
rect 36642 80303 36694 80445
rect 36650 28763 36686 80303
rect 36642 28621 36694 28763
rect 36650 28463 36686 28621
rect 36722 28463 36758 80603
rect 36794 28463 36830 80603
rect 36866 80124 36959 80190
rect 36866 80108 36943 80124
tri 36943 80108 36959 80124 nw
rect 36995 80091 37109 80233
rect 37145 80124 37238 80190
tri 37145 80108 37161 80124 ne
rect 37161 80108 37238 80124
rect 36978 80009 37126 80091
rect 36866 79976 36943 79992
tri 36943 79976 36959 79992 sw
rect 36866 79910 36959 79976
rect 36995 79851 37109 80009
tri 37145 79976 37161 79992 se
rect 37161 79976 37238 79992
rect 37145 79910 37238 79976
rect 36866 79775 37238 79851
rect 36866 79650 36959 79716
rect 36866 79634 36943 79650
tri 36943 79634 36959 79650 nw
rect 36995 79617 37109 79775
rect 37145 79650 37238 79716
tri 37145 79634 37161 79650 ne
rect 37161 79634 37238 79650
rect 36978 79535 37126 79617
rect 36866 79502 36943 79518
tri 36943 79502 36959 79518 sw
rect 36866 79436 36959 79502
rect 36866 79334 36959 79400
rect 36866 79318 36943 79334
tri 36943 79318 36959 79334 nw
rect 36995 79301 37109 79535
tri 37145 79502 37161 79518 se
rect 37161 79502 37238 79518
rect 37145 79436 37238 79502
rect 37145 79334 37238 79400
tri 37145 79318 37161 79334 ne
rect 37161 79318 37238 79334
rect 36978 79219 37126 79301
rect 36866 79186 36943 79202
tri 36943 79186 36959 79202 sw
rect 36866 79120 36959 79186
rect 36995 79061 37109 79219
tri 37145 79186 37161 79202 se
rect 37161 79186 37238 79202
rect 37145 79120 37238 79186
rect 36866 78985 37238 79061
rect 36866 78860 36959 78926
rect 36866 78844 36943 78860
tri 36943 78844 36959 78860 nw
rect 36995 78827 37109 78985
rect 37145 78860 37238 78926
tri 37145 78844 37161 78860 ne
rect 37161 78844 37238 78860
rect 36978 78745 37126 78827
rect 36866 78712 36943 78728
tri 36943 78712 36959 78728 sw
rect 36866 78646 36959 78712
rect 36866 78544 36959 78610
rect 36866 78528 36943 78544
tri 36943 78528 36959 78544 nw
rect 36995 78511 37109 78745
tri 37145 78712 37161 78728 se
rect 37161 78712 37238 78728
rect 37145 78646 37238 78712
rect 37145 78544 37238 78610
tri 37145 78528 37161 78544 ne
rect 37161 78528 37238 78544
rect 36978 78429 37126 78511
rect 36866 78396 36943 78412
tri 36943 78396 36959 78412 sw
rect 36866 78330 36959 78396
rect 36995 78271 37109 78429
tri 37145 78396 37161 78412 se
rect 37161 78396 37238 78412
rect 37145 78330 37238 78396
rect 36866 78195 37238 78271
rect 36866 78070 36959 78136
rect 36866 78054 36943 78070
tri 36943 78054 36959 78070 nw
rect 36995 78037 37109 78195
rect 37145 78070 37238 78136
tri 37145 78054 37161 78070 ne
rect 37161 78054 37238 78070
rect 36978 77955 37126 78037
rect 36866 77922 36943 77938
tri 36943 77922 36959 77938 sw
rect 36866 77856 36959 77922
rect 36866 77754 36959 77820
rect 36866 77738 36943 77754
tri 36943 77738 36959 77754 nw
rect 36995 77721 37109 77955
tri 37145 77922 37161 77938 se
rect 37161 77922 37238 77938
rect 37145 77856 37238 77922
rect 37145 77754 37238 77820
tri 37145 77738 37161 77754 ne
rect 37161 77738 37238 77754
rect 36978 77639 37126 77721
rect 36866 77606 36943 77622
tri 36943 77606 36959 77622 sw
rect 36866 77540 36959 77606
rect 36995 77481 37109 77639
tri 37145 77606 37161 77622 se
rect 37161 77606 37238 77622
rect 37145 77540 37238 77606
rect 36866 77405 37238 77481
rect 36866 77280 36959 77346
rect 36866 77264 36943 77280
tri 36943 77264 36959 77280 nw
rect 36995 77247 37109 77405
rect 37145 77280 37238 77346
tri 37145 77264 37161 77280 ne
rect 37161 77264 37238 77280
rect 36978 77165 37126 77247
rect 36866 77132 36943 77148
tri 36943 77132 36959 77148 sw
rect 36866 77066 36959 77132
rect 36866 76964 36959 77030
rect 36866 76948 36943 76964
tri 36943 76948 36959 76964 nw
rect 36995 76931 37109 77165
tri 37145 77132 37161 77148 se
rect 37161 77132 37238 77148
rect 37145 77066 37238 77132
rect 37145 76964 37238 77030
tri 37145 76948 37161 76964 ne
rect 37161 76948 37238 76964
rect 36978 76849 37126 76931
rect 36866 76816 36943 76832
tri 36943 76816 36959 76832 sw
rect 36866 76750 36959 76816
rect 36995 76691 37109 76849
tri 37145 76816 37161 76832 se
rect 37161 76816 37238 76832
rect 37145 76750 37238 76816
rect 36866 76615 37238 76691
rect 36866 76490 36959 76556
rect 36866 76474 36943 76490
tri 36943 76474 36959 76490 nw
rect 36995 76457 37109 76615
rect 37145 76490 37238 76556
tri 37145 76474 37161 76490 ne
rect 37161 76474 37238 76490
rect 36978 76375 37126 76457
rect 36866 76342 36943 76358
tri 36943 76342 36959 76358 sw
rect 36866 76276 36959 76342
rect 36866 76174 36959 76240
rect 36866 76158 36943 76174
tri 36943 76158 36959 76174 nw
rect 36995 76141 37109 76375
tri 37145 76342 37161 76358 se
rect 37161 76342 37238 76358
rect 37145 76276 37238 76342
rect 37145 76174 37238 76240
tri 37145 76158 37161 76174 ne
rect 37161 76158 37238 76174
rect 36978 76059 37126 76141
rect 36866 76026 36943 76042
tri 36943 76026 36959 76042 sw
rect 36866 75960 36959 76026
rect 36995 75901 37109 76059
tri 37145 76026 37161 76042 se
rect 37161 76026 37238 76042
rect 37145 75960 37238 76026
rect 36866 75825 37238 75901
rect 36866 75700 36959 75766
rect 36866 75684 36943 75700
tri 36943 75684 36959 75700 nw
rect 36995 75667 37109 75825
rect 37145 75700 37238 75766
tri 37145 75684 37161 75700 ne
rect 37161 75684 37238 75700
rect 36978 75585 37126 75667
rect 36866 75552 36943 75568
tri 36943 75552 36959 75568 sw
rect 36866 75486 36959 75552
rect 36866 75384 36959 75450
rect 36866 75368 36943 75384
tri 36943 75368 36959 75384 nw
rect 36995 75351 37109 75585
tri 37145 75552 37161 75568 se
rect 37161 75552 37238 75568
rect 37145 75486 37238 75552
rect 37145 75384 37238 75450
tri 37145 75368 37161 75384 ne
rect 37161 75368 37238 75384
rect 36978 75269 37126 75351
rect 36866 75236 36943 75252
tri 36943 75236 36959 75252 sw
rect 36866 75170 36959 75236
rect 36995 75111 37109 75269
tri 37145 75236 37161 75252 se
rect 37161 75236 37238 75252
rect 37145 75170 37238 75236
rect 36866 75035 37238 75111
rect 36866 74910 36959 74976
rect 36866 74894 36943 74910
tri 36943 74894 36959 74910 nw
rect 36995 74877 37109 75035
rect 37145 74910 37238 74976
tri 37145 74894 37161 74910 ne
rect 37161 74894 37238 74910
rect 36978 74795 37126 74877
rect 36866 74762 36943 74778
tri 36943 74762 36959 74778 sw
rect 36866 74696 36959 74762
rect 36866 74594 36959 74660
rect 36866 74578 36943 74594
tri 36943 74578 36959 74594 nw
rect 36995 74561 37109 74795
tri 37145 74762 37161 74778 se
rect 37161 74762 37238 74778
rect 37145 74696 37238 74762
rect 37145 74594 37238 74660
tri 37145 74578 37161 74594 ne
rect 37161 74578 37238 74594
rect 36978 74479 37126 74561
rect 36866 74446 36943 74462
tri 36943 74446 36959 74462 sw
rect 36866 74380 36959 74446
rect 36995 74321 37109 74479
tri 37145 74446 37161 74462 se
rect 37161 74446 37238 74462
rect 37145 74380 37238 74446
rect 36866 74245 37238 74321
rect 36866 74120 36959 74186
rect 36866 74104 36943 74120
tri 36943 74104 36959 74120 nw
rect 36995 74087 37109 74245
rect 37145 74120 37238 74186
tri 37145 74104 37161 74120 ne
rect 37161 74104 37238 74120
rect 36978 74005 37126 74087
rect 36866 73972 36943 73988
tri 36943 73972 36959 73988 sw
rect 36866 73906 36959 73972
rect 36866 73804 36959 73870
rect 36866 73788 36943 73804
tri 36943 73788 36959 73804 nw
rect 36995 73771 37109 74005
tri 37145 73972 37161 73988 se
rect 37161 73972 37238 73988
rect 37145 73906 37238 73972
rect 37145 73804 37238 73870
tri 37145 73788 37161 73804 ne
rect 37161 73788 37238 73804
rect 36978 73689 37126 73771
rect 36866 73656 36943 73672
tri 36943 73656 36959 73672 sw
rect 36866 73590 36959 73656
rect 36995 73531 37109 73689
tri 37145 73656 37161 73672 se
rect 37161 73656 37238 73672
rect 37145 73590 37238 73656
rect 36866 73455 37238 73531
rect 36866 73330 36959 73396
rect 36866 73314 36943 73330
tri 36943 73314 36959 73330 nw
rect 36995 73297 37109 73455
rect 37145 73330 37238 73396
tri 37145 73314 37161 73330 ne
rect 37161 73314 37238 73330
rect 36978 73215 37126 73297
rect 36866 73182 36943 73198
tri 36943 73182 36959 73198 sw
rect 36866 73116 36959 73182
rect 36866 73014 36959 73080
rect 36866 72998 36943 73014
tri 36943 72998 36959 73014 nw
rect 36995 72981 37109 73215
tri 37145 73182 37161 73198 se
rect 37161 73182 37238 73198
rect 37145 73116 37238 73182
rect 37145 73014 37238 73080
tri 37145 72998 37161 73014 ne
rect 37161 72998 37238 73014
rect 36978 72899 37126 72981
rect 36866 72866 36943 72882
tri 36943 72866 36959 72882 sw
rect 36866 72800 36959 72866
rect 36995 72741 37109 72899
tri 37145 72866 37161 72882 se
rect 37161 72866 37238 72882
rect 37145 72800 37238 72866
rect 36866 72665 37238 72741
rect 36866 72540 36959 72606
rect 36866 72524 36943 72540
tri 36943 72524 36959 72540 nw
rect 36995 72507 37109 72665
rect 37145 72540 37238 72606
tri 37145 72524 37161 72540 ne
rect 37161 72524 37238 72540
rect 36978 72425 37126 72507
rect 36866 72392 36943 72408
tri 36943 72392 36959 72408 sw
rect 36866 72326 36959 72392
rect 36866 72224 36959 72290
rect 36866 72208 36943 72224
tri 36943 72208 36959 72224 nw
rect 36995 72191 37109 72425
tri 37145 72392 37161 72408 se
rect 37161 72392 37238 72408
rect 37145 72326 37238 72392
rect 37145 72224 37238 72290
tri 37145 72208 37161 72224 ne
rect 37161 72208 37238 72224
rect 36978 72109 37126 72191
rect 36866 72076 36943 72092
tri 36943 72076 36959 72092 sw
rect 36866 72010 36959 72076
rect 36995 71951 37109 72109
tri 37145 72076 37161 72092 se
rect 37161 72076 37238 72092
rect 37145 72010 37238 72076
rect 36866 71875 37238 71951
rect 36866 71750 36959 71816
rect 36866 71734 36943 71750
tri 36943 71734 36959 71750 nw
rect 36995 71717 37109 71875
rect 37145 71750 37238 71816
tri 37145 71734 37161 71750 ne
rect 37161 71734 37238 71750
rect 36978 71635 37126 71717
rect 36866 71602 36943 71618
tri 36943 71602 36959 71618 sw
rect 36866 71536 36959 71602
rect 36866 71434 36959 71500
rect 36866 71418 36943 71434
tri 36943 71418 36959 71434 nw
rect 36995 71401 37109 71635
tri 37145 71602 37161 71618 se
rect 37161 71602 37238 71618
rect 37145 71536 37238 71602
rect 37145 71434 37238 71500
tri 37145 71418 37161 71434 ne
rect 37161 71418 37238 71434
rect 36978 71319 37126 71401
rect 36866 71286 36943 71302
tri 36943 71286 36959 71302 sw
rect 36866 71220 36959 71286
rect 36995 71161 37109 71319
tri 37145 71286 37161 71302 se
rect 37161 71286 37238 71302
rect 37145 71220 37238 71286
rect 36866 71085 37238 71161
rect 36866 70960 36959 71026
rect 36866 70944 36943 70960
tri 36943 70944 36959 70960 nw
rect 36995 70927 37109 71085
rect 37145 70960 37238 71026
tri 37145 70944 37161 70960 ne
rect 37161 70944 37238 70960
rect 36978 70845 37126 70927
rect 36866 70812 36943 70828
tri 36943 70812 36959 70828 sw
rect 36866 70746 36959 70812
rect 36866 70644 36959 70710
rect 36866 70628 36943 70644
tri 36943 70628 36959 70644 nw
rect 36995 70611 37109 70845
tri 37145 70812 37161 70828 se
rect 37161 70812 37238 70828
rect 37145 70746 37238 70812
rect 37145 70644 37238 70710
tri 37145 70628 37161 70644 ne
rect 37161 70628 37238 70644
rect 36978 70529 37126 70611
rect 36866 70496 36943 70512
tri 36943 70496 36959 70512 sw
rect 36866 70430 36959 70496
rect 36995 70371 37109 70529
tri 37145 70496 37161 70512 se
rect 37161 70496 37238 70512
rect 37145 70430 37238 70496
rect 36866 70295 37238 70371
rect 36866 70170 36959 70236
rect 36866 70154 36943 70170
tri 36943 70154 36959 70170 nw
rect 36995 70137 37109 70295
rect 37145 70170 37238 70236
tri 37145 70154 37161 70170 ne
rect 37161 70154 37238 70170
rect 36978 70055 37126 70137
rect 36866 70022 36943 70038
tri 36943 70022 36959 70038 sw
rect 36866 69956 36959 70022
rect 36866 69854 36959 69920
rect 36866 69838 36943 69854
tri 36943 69838 36959 69854 nw
rect 36995 69821 37109 70055
tri 37145 70022 37161 70038 se
rect 37161 70022 37238 70038
rect 37145 69956 37238 70022
rect 37145 69854 37238 69920
tri 37145 69838 37161 69854 ne
rect 37161 69838 37238 69854
rect 36978 69739 37126 69821
rect 36866 69706 36943 69722
tri 36943 69706 36959 69722 sw
rect 36866 69640 36959 69706
rect 36995 69581 37109 69739
tri 37145 69706 37161 69722 se
rect 37161 69706 37238 69722
rect 37145 69640 37238 69706
rect 36866 69505 37238 69581
rect 36866 69380 36959 69446
rect 36866 69364 36943 69380
tri 36943 69364 36959 69380 nw
rect 36995 69347 37109 69505
rect 37145 69380 37238 69446
tri 37145 69364 37161 69380 ne
rect 37161 69364 37238 69380
rect 36978 69265 37126 69347
rect 36866 69232 36943 69248
tri 36943 69232 36959 69248 sw
rect 36866 69166 36959 69232
rect 36866 69064 36959 69130
rect 36866 69048 36943 69064
tri 36943 69048 36959 69064 nw
rect 36995 69031 37109 69265
tri 37145 69232 37161 69248 se
rect 37161 69232 37238 69248
rect 37145 69166 37238 69232
rect 37145 69064 37238 69130
tri 37145 69048 37161 69064 ne
rect 37161 69048 37238 69064
rect 36978 68949 37126 69031
rect 36866 68916 36943 68932
tri 36943 68916 36959 68932 sw
rect 36866 68850 36959 68916
rect 36995 68791 37109 68949
tri 37145 68916 37161 68932 se
rect 37161 68916 37238 68932
rect 37145 68850 37238 68916
rect 36866 68715 37238 68791
rect 36866 68590 36959 68656
rect 36866 68574 36943 68590
tri 36943 68574 36959 68590 nw
rect 36995 68557 37109 68715
rect 37145 68590 37238 68656
tri 37145 68574 37161 68590 ne
rect 37161 68574 37238 68590
rect 36978 68475 37126 68557
rect 36866 68442 36943 68458
tri 36943 68442 36959 68458 sw
rect 36866 68376 36959 68442
rect 36866 68274 36959 68340
rect 36866 68258 36943 68274
tri 36943 68258 36959 68274 nw
rect 36995 68241 37109 68475
tri 37145 68442 37161 68458 se
rect 37161 68442 37238 68458
rect 37145 68376 37238 68442
rect 37145 68274 37238 68340
tri 37145 68258 37161 68274 ne
rect 37161 68258 37238 68274
rect 36978 68159 37126 68241
rect 36866 68126 36943 68142
tri 36943 68126 36959 68142 sw
rect 36866 68060 36959 68126
rect 36995 68001 37109 68159
tri 37145 68126 37161 68142 se
rect 37161 68126 37238 68142
rect 37145 68060 37238 68126
rect 36866 67925 37238 68001
rect 36866 67800 36959 67866
rect 36866 67784 36943 67800
tri 36943 67784 36959 67800 nw
rect 36995 67767 37109 67925
rect 37145 67800 37238 67866
tri 37145 67784 37161 67800 ne
rect 37161 67784 37238 67800
rect 36978 67685 37126 67767
rect 36866 67652 36943 67668
tri 36943 67652 36959 67668 sw
rect 36866 67586 36959 67652
rect 36866 67484 36959 67550
rect 36866 67468 36943 67484
tri 36943 67468 36959 67484 nw
rect 36995 67451 37109 67685
tri 37145 67652 37161 67668 se
rect 37161 67652 37238 67668
rect 37145 67586 37238 67652
rect 37145 67484 37238 67550
tri 37145 67468 37161 67484 ne
rect 37161 67468 37238 67484
rect 36978 67369 37126 67451
rect 36866 67336 36943 67352
tri 36943 67336 36959 67352 sw
rect 36866 67270 36959 67336
rect 36995 67211 37109 67369
tri 37145 67336 37161 67352 se
rect 37161 67336 37238 67352
rect 37145 67270 37238 67336
rect 36866 67135 37238 67211
rect 36866 67010 36959 67076
rect 36866 66994 36943 67010
tri 36943 66994 36959 67010 nw
rect 36995 66977 37109 67135
rect 37145 67010 37238 67076
tri 37145 66994 37161 67010 ne
rect 37161 66994 37238 67010
rect 36978 66895 37126 66977
rect 36866 66862 36943 66878
tri 36943 66862 36959 66878 sw
rect 36866 66796 36959 66862
rect 36866 66694 36959 66760
rect 36866 66678 36943 66694
tri 36943 66678 36959 66694 nw
rect 36995 66661 37109 66895
tri 37145 66862 37161 66878 se
rect 37161 66862 37238 66878
rect 37145 66796 37238 66862
rect 37145 66694 37238 66760
tri 37145 66678 37161 66694 ne
rect 37161 66678 37238 66694
rect 36978 66579 37126 66661
rect 36866 66546 36943 66562
tri 36943 66546 36959 66562 sw
rect 36866 66480 36959 66546
rect 36995 66421 37109 66579
tri 37145 66546 37161 66562 se
rect 37161 66546 37238 66562
rect 37145 66480 37238 66546
rect 36866 66345 37238 66421
rect 36866 66220 36959 66286
rect 36866 66204 36943 66220
tri 36943 66204 36959 66220 nw
rect 36995 66187 37109 66345
rect 37145 66220 37238 66286
tri 37145 66204 37161 66220 ne
rect 37161 66204 37238 66220
rect 36978 66105 37126 66187
rect 36866 66072 36943 66088
tri 36943 66072 36959 66088 sw
rect 36866 66006 36959 66072
rect 36866 65904 36959 65970
rect 36866 65888 36943 65904
tri 36943 65888 36959 65904 nw
rect 36995 65871 37109 66105
tri 37145 66072 37161 66088 se
rect 37161 66072 37238 66088
rect 37145 66006 37238 66072
rect 37145 65904 37238 65970
tri 37145 65888 37161 65904 ne
rect 37161 65888 37238 65904
rect 36978 65789 37126 65871
rect 36866 65756 36943 65772
tri 36943 65756 36959 65772 sw
rect 36866 65690 36959 65756
rect 36995 65631 37109 65789
tri 37145 65756 37161 65772 se
rect 37161 65756 37238 65772
rect 37145 65690 37238 65756
rect 36866 65555 37238 65631
rect 36866 65430 36959 65496
rect 36866 65414 36943 65430
tri 36943 65414 36959 65430 nw
rect 36995 65397 37109 65555
rect 37145 65430 37238 65496
tri 37145 65414 37161 65430 ne
rect 37161 65414 37238 65430
rect 36978 65315 37126 65397
rect 36866 65282 36943 65298
tri 36943 65282 36959 65298 sw
rect 36866 65216 36959 65282
rect 36866 65114 36959 65180
rect 36866 65098 36943 65114
tri 36943 65098 36959 65114 nw
rect 36995 65081 37109 65315
tri 37145 65282 37161 65298 se
rect 37161 65282 37238 65298
rect 37145 65216 37238 65282
rect 37145 65114 37238 65180
tri 37145 65098 37161 65114 ne
rect 37161 65098 37238 65114
rect 36978 64999 37126 65081
rect 36866 64966 36943 64982
tri 36943 64966 36959 64982 sw
rect 36866 64900 36959 64966
rect 36995 64841 37109 64999
tri 37145 64966 37161 64982 se
rect 37161 64966 37238 64982
rect 37145 64900 37238 64966
rect 36866 64765 37238 64841
rect 36866 64640 36959 64706
rect 36866 64624 36943 64640
tri 36943 64624 36959 64640 nw
rect 36995 64607 37109 64765
rect 37145 64640 37238 64706
tri 37145 64624 37161 64640 ne
rect 37161 64624 37238 64640
rect 36978 64525 37126 64607
rect 36866 64492 36943 64508
tri 36943 64492 36959 64508 sw
rect 36866 64426 36959 64492
rect 36866 64324 36959 64390
rect 36866 64308 36943 64324
tri 36943 64308 36959 64324 nw
rect 36995 64291 37109 64525
tri 37145 64492 37161 64508 se
rect 37161 64492 37238 64508
rect 37145 64426 37238 64492
rect 37145 64324 37238 64390
tri 37145 64308 37161 64324 ne
rect 37161 64308 37238 64324
rect 36978 64209 37126 64291
rect 36866 64176 36943 64192
tri 36943 64176 36959 64192 sw
rect 36866 64110 36959 64176
rect 36995 64051 37109 64209
tri 37145 64176 37161 64192 se
rect 37161 64176 37238 64192
rect 37145 64110 37238 64176
rect 36866 63975 37238 64051
rect 36866 63850 36959 63916
rect 36866 63834 36943 63850
tri 36943 63834 36959 63850 nw
rect 36995 63817 37109 63975
rect 37145 63850 37238 63916
tri 37145 63834 37161 63850 ne
rect 37161 63834 37238 63850
rect 36978 63735 37126 63817
rect 36866 63702 36943 63718
tri 36943 63702 36959 63718 sw
rect 36866 63636 36959 63702
rect 36866 63534 36959 63600
rect 36866 63518 36943 63534
tri 36943 63518 36959 63534 nw
rect 36995 63501 37109 63735
tri 37145 63702 37161 63718 se
rect 37161 63702 37238 63718
rect 37145 63636 37238 63702
rect 37145 63534 37238 63600
tri 37145 63518 37161 63534 ne
rect 37161 63518 37238 63534
rect 36978 63419 37126 63501
rect 36866 63386 36943 63402
tri 36943 63386 36959 63402 sw
rect 36866 63320 36959 63386
rect 36995 63261 37109 63419
tri 37145 63386 37161 63402 se
rect 37161 63386 37238 63402
rect 37145 63320 37238 63386
rect 36866 63185 37238 63261
rect 36866 63060 36959 63126
rect 36866 63044 36943 63060
tri 36943 63044 36959 63060 nw
rect 36995 63027 37109 63185
rect 37145 63060 37238 63126
tri 37145 63044 37161 63060 ne
rect 37161 63044 37238 63060
rect 36978 62945 37126 63027
rect 36866 62912 36943 62928
tri 36943 62912 36959 62928 sw
rect 36866 62846 36959 62912
rect 36866 62744 36959 62810
rect 36866 62728 36943 62744
tri 36943 62728 36959 62744 nw
rect 36995 62711 37109 62945
tri 37145 62912 37161 62928 se
rect 37161 62912 37238 62928
rect 37145 62846 37238 62912
rect 37145 62744 37238 62810
tri 37145 62728 37161 62744 ne
rect 37161 62728 37238 62744
rect 36978 62629 37126 62711
rect 36866 62596 36943 62612
tri 36943 62596 36959 62612 sw
rect 36866 62530 36959 62596
rect 36995 62471 37109 62629
tri 37145 62596 37161 62612 se
rect 37161 62596 37238 62612
rect 37145 62530 37238 62596
rect 36866 62395 37238 62471
rect 36866 62270 36959 62336
rect 36866 62254 36943 62270
tri 36943 62254 36959 62270 nw
rect 36995 62237 37109 62395
rect 37145 62270 37238 62336
tri 37145 62254 37161 62270 ne
rect 37161 62254 37238 62270
rect 36978 62155 37126 62237
rect 36866 62122 36943 62138
tri 36943 62122 36959 62138 sw
rect 36866 62056 36959 62122
rect 36866 61954 36959 62020
rect 36866 61938 36943 61954
tri 36943 61938 36959 61954 nw
rect 36995 61921 37109 62155
tri 37145 62122 37161 62138 se
rect 37161 62122 37238 62138
rect 37145 62056 37238 62122
rect 37145 61954 37238 62020
tri 37145 61938 37161 61954 ne
rect 37161 61938 37238 61954
rect 36978 61839 37126 61921
rect 36866 61806 36943 61822
tri 36943 61806 36959 61822 sw
rect 36866 61740 36959 61806
rect 36995 61681 37109 61839
tri 37145 61806 37161 61822 se
rect 37161 61806 37238 61822
rect 37145 61740 37238 61806
rect 36866 61605 37238 61681
rect 36866 61480 36959 61546
rect 36866 61464 36943 61480
tri 36943 61464 36959 61480 nw
rect 36995 61447 37109 61605
rect 37145 61480 37238 61546
tri 37145 61464 37161 61480 ne
rect 37161 61464 37238 61480
rect 36978 61365 37126 61447
rect 36866 61332 36943 61348
tri 36943 61332 36959 61348 sw
rect 36866 61266 36959 61332
rect 36866 61164 36959 61230
rect 36866 61148 36943 61164
tri 36943 61148 36959 61164 nw
rect 36995 61131 37109 61365
tri 37145 61332 37161 61348 se
rect 37161 61332 37238 61348
rect 37145 61266 37238 61332
rect 37145 61164 37238 61230
tri 37145 61148 37161 61164 ne
rect 37161 61148 37238 61164
rect 36978 61049 37126 61131
rect 36866 61016 36943 61032
tri 36943 61016 36959 61032 sw
rect 36866 60950 36959 61016
rect 36995 60891 37109 61049
tri 37145 61016 37161 61032 se
rect 37161 61016 37238 61032
rect 37145 60950 37238 61016
rect 36866 60815 37238 60891
rect 36866 60690 36959 60756
rect 36866 60674 36943 60690
tri 36943 60674 36959 60690 nw
rect 36995 60657 37109 60815
rect 37145 60690 37238 60756
tri 37145 60674 37161 60690 ne
rect 37161 60674 37238 60690
rect 36978 60575 37126 60657
rect 36866 60542 36943 60558
tri 36943 60542 36959 60558 sw
rect 36866 60476 36959 60542
rect 36866 60374 36959 60440
rect 36866 60358 36943 60374
tri 36943 60358 36959 60374 nw
rect 36995 60341 37109 60575
tri 37145 60542 37161 60558 se
rect 37161 60542 37238 60558
rect 37145 60476 37238 60542
rect 37145 60374 37238 60440
tri 37145 60358 37161 60374 ne
rect 37161 60358 37238 60374
rect 36978 60259 37126 60341
rect 36866 60226 36943 60242
tri 36943 60226 36959 60242 sw
rect 36866 60160 36959 60226
rect 36995 60101 37109 60259
tri 37145 60226 37161 60242 se
rect 37161 60226 37238 60242
rect 37145 60160 37238 60226
rect 36866 60025 37238 60101
rect 36866 59900 36959 59966
rect 36866 59884 36943 59900
tri 36943 59884 36959 59900 nw
rect 36995 59867 37109 60025
rect 37145 59900 37238 59966
tri 37145 59884 37161 59900 ne
rect 37161 59884 37238 59900
rect 36978 59785 37126 59867
rect 36866 59752 36943 59768
tri 36943 59752 36959 59768 sw
rect 36866 59686 36959 59752
rect 36866 59584 36959 59650
rect 36866 59568 36943 59584
tri 36943 59568 36959 59584 nw
rect 36995 59551 37109 59785
tri 37145 59752 37161 59768 se
rect 37161 59752 37238 59768
rect 37145 59686 37238 59752
rect 37145 59584 37238 59650
tri 37145 59568 37161 59584 ne
rect 37161 59568 37238 59584
rect 36978 59469 37126 59551
rect 36866 59436 36943 59452
tri 36943 59436 36959 59452 sw
rect 36866 59370 36959 59436
rect 36995 59311 37109 59469
tri 37145 59436 37161 59452 se
rect 37161 59436 37238 59452
rect 37145 59370 37238 59436
rect 36866 59235 37238 59311
rect 36866 59110 36959 59176
rect 36866 59094 36943 59110
tri 36943 59094 36959 59110 nw
rect 36995 59077 37109 59235
rect 37145 59110 37238 59176
tri 37145 59094 37161 59110 ne
rect 37161 59094 37238 59110
rect 36978 58995 37126 59077
rect 36866 58962 36943 58978
tri 36943 58962 36959 58978 sw
rect 36866 58896 36959 58962
rect 36866 58794 36959 58860
rect 36866 58778 36943 58794
tri 36943 58778 36959 58794 nw
rect 36995 58761 37109 58995
tri 37145 58962 37161 58978 se
rect 37161 58962 37238 58978
rect 37145 58896 37238 58962
rect 37145 58794 37238 58860
tri 37145 58778 37161 58794 ne
rect 37161 58778 37238 58794
rect 36978 58679 37126 58761
rect 36866 58646 36943 58662
tri 36943 58646 36959 58662 sw
rect 36866 58580 36959 58646
rect 36995 58521 37109 58679
tri 37145 58646 37161 58662 se
rect 37161 58646 37238 58662
rect 37145 58580 37238 58646
rect 36866 58445 37238 58521
rect 36866 58320 36959 58386
rect 36866 58304 36943 58320
tri 36943 58304 36959 58320 nw
rect 36995 58287 37109 58445
rect 37145 58320 37238 58386
tri 37145 58304 37161 58320 ne
rect 37161 58304 37238 58320
rect 36978 58205 37126 58287
rect 36866 58172 36943 58188
tri 36943 58172 36959 58188 sw
rect 36866 58106 36959 58172
rect 36866 58004 36959 58070
rect 36866 57988 36943 58004
tri 36943 57988 36959 58004 nw
rect 36995 57971 37109 58205
tri 37145 58172 37161 58188 se
rect 37161 58172 37238 58188
rect 37145 58106 37238 58172
rect 37145 58004 37238 58070
tri 37145 57988 37161 58004 ne
rect 37161 57988 37238 58004
rect 36978 57889 37126 57971
rect 36866 57856 36943 57872
tri 36943 57856 36959 57872 sw
rect 36866 57790 36959 57856
rect 36995 57731 37109 57889
tri 37145 57856 37161 57872 se
rect 37161 57856 37238 57872
rect 37145 57790 37238 57856
rect 36866 57655 37238 57731
rect 36866 57530 36959 57596
rect 36866 57514 36943 57530
tri 36943 57514 36959 57530 nw
rect 36995 57497 37109 57655
rect 37145 57530 37238 57596
tri 37145 57514 37161 57530 ne
rect 37161 57514 37238 57530
rect 36978 57415 37126 57497
rect 36866 57382 36943 57398
tri 36943 57382 36959 57398 sw
rect 36866 57316 36959 57382
rect 36866 57214 36959 57280
rect 36866 57198 36943 57214
tri 36943 57198 36959 57214 nw
rect 36995 57181 37109 57415
tri 37145 57382 37161 57398 se
rect 37161 57382 37238 57398
rect 37145 57316 37238 57382
rect 37145 57214 37238 57280
tri 37145 57198 37161 57214 ne
rect 37161 57198 37238 57214
rect 36978 57099 37126 57181
rect 36866 57066 36943 57082
tri 36943 57066 36959 57082 sw
rect 36866 57000 36959 57066
rect 36995 56941 37109 57099
tri 37145 57066 37161 57082 se
rect 37161 57066 37238 57082
rect 37145 57000 37238 57066
rect 36866 56865 37238 56941
rect 36866 56740 36959 56806
rect 36866 56724 36943 56740
tri 36943 56724 36959 56740 nw
rect 36995 56707 37109 56865
rect 37145 56740 37238 56806
tri 37145 56724 37161 56740 ne
rect 37161 56724 37238 56740
rect 36978 56625 37126 56707
rect 36866 56592 36943 56608
tri 36943 56592 36959 56608 sw
rect 36866 56526 36959 56592
rect 36866 56424 36959 56490
rect 36866 56408 36943 56424
tri 36943 56408 36959 56424 nw
rect 36995 56391 37109 56625
tri 37145 56592 37161 56608 se
rect 37161 56592 37238 56608
rect 37145 56526 37238 56592
rect 37145 56424 37238 56490
tri 37145 56408 37161 56424 ne
rect 37161 56408 37238 56424
rect 36978 56309 37126 56391
rect 36866 56276 36943 56292
tri 36943 56276 36959 56292 sw
rect 36866 56210 36959 56276
rect 36995 56151 37109 56309
tri 37145 56276 37161 56292 se
rect 37161 56276 37238 56292
rect 37145 56210 37238 56276
rect 36866 56075 37238 56151
rect 36866 55950 36959 56016
rect 36866 55934 36943 55950
tri 36943 55934 36959 55950 nw
rect 36995 55917 37109 56075
rect 37145 55950 37238 56016
tri 37145 55934 37161 55950 ne
rect 37161 55934 37238 55950
rect 36978 55835 37126 55917
rect 36866 55802 36943 55818
tri 36943 55802 36959 55818 sw
rect 36866 55736 36959 55802
rect 36866 55634 36959 55700
rect 36866 55618 36943 55634
tri 36943 55618 36959 55634 nw
rect 36995 55601 37109 55835
tri 37145 55802 37161 55818 se
rect 37161 55802 37238 55818
rect 37145 55736 37238 55802
rect 37145 55634 37238 55700
tri 37145 55618 37161 55634 ne
rect 37161 55618 37238 55634
rect 36978 55519 37126 55601
rect 36866 55486 36943 55502
tri 36943 55486 36959 55502 sw
rect 36866 55420 36959 55486
rect 36995 55361 37109 55519
tri 37145 55486 37161 55502 se
rect 37161 55486 37238 55502
rect 37145 55420 37238 55486
rect 36866 55285 37238 55361
rect 36866 55160 36959 55226
rect 36866 55144 36943 55160
tri 36943 55144 36959 55160 nw
rect 36995 55127 37109 55285
rect 37145 55160 37238 55226
tri 37145 55144 37161 55160 ne
rect 37161 55144 37238 55160
rect 36978 55045 37126 55127
rect 36866 55012 36943 55028
tri 36943 55012 36959 55028 sw
rect 36866 54946 36959 55012
rect 36866 54844 36959 54910
rect 36866 54828 36943 54844
tri 36943 54828 36959 54844 nw
rect 36995 54811 37109 55045
tri 37145 55012 37161 55028 se
rect 37161 55012 37238 55028
rect 37145 54946 37238 55012
rect 37145 54844 37238 54910
tri 37145 54828 37161 54844 ne
rect 37161 54828 37238 54844
rect 36978 54729 37126 54811
rect 36866 54696 36943 54712
tri 36943 54696 36959 54712 sw
rect 36866 54630 36959 54696
rect 36995 54571 37109 54729
tri 37145 54696 37161 54712 se
rect 37161 54696 37238 54712
rect 37145 54630 37238 54696
rect 36866 54495 37238 54571
rect 36866 54370 36959 54436
rect 36866 54354 36943 54370
tri 36943 54354 36959 54370 nw
rect 36995 54337 37109 54495
rect 37145 54370 37238 54436
tri 37145 54354 37161 54370 ne
rect 37161 54354 37238 54370
rect 36978 54255 37126 54337
rect 36866 54222 36943 54238
tri 36943 54222 36959 54238 sw
rect 36866 54156 36959 54222
rect 36866 54054 36959 54120
rect 36866 54038 36943 54054
tri 36943 54038 36959 54054 nw
rect 36995 54021 37109 54255
tri 37145 54222 37161 54238 se
rect 37161 54222 37238 54238
rect 37145 54156 37238 54222
rect 37145 54054 37238 54120
tri 37145 54038 37161 54054 ne
rect 37161 54038 37238 54054
rect 36978 53939 37126 54021
rect 36866 53906 36943 53922
tri 36943 53906 36959 53922 sw
rect 36866 53840 36959 53906
rect 36995 53781 37109 53939
tri 37145 53906 37161 53922 se
rect 37161 53906 37238 53922
rect 37145 53840 37238 53906
rect 36866 53705 37238 53781
rect 36866 53580 36959 53646
rect 36866 53564 36943 53580
tri 36943 53564 36959 53580 nw
rect 36995 53547 37109 53705
rect 37145 53580 37238 53646
tri 37145 53564 37161 53580 ne
rect 37161 53564 37238 53580
rect 36978 53465 37126 53547
rect 36866 53432 36943 53448
tri 36943 53432 36959 53448 sw
rect 36866 53366 36959 53432
rect 36866 53264 36959 53330
rect 36866 53248 36943 53264
tri 36943 53248 36959 53264 nw
rect 36995 53231 37109 53465
tri 37145 53432 37161 53448 se
rect 37161 53432 37238 53448
rect 37145 53366 37238 53432
rect 37145 53264 37238 53330
tri 37145 53248 37161 53264 ne
rect 37161 53248 37238 53264
rect 36978 53149 37126 53231
rect 36866 53116 36943 53132
tri 36943 53116 36959 53132 sw
rect 36866 53050 36959 53116
rect 36995 52991 37109 53149
tri 37145 53116 37161 53132 se
rect 37161 53116 37238 53132
rect 37145 53050 37238 53116
rect 36866 52915 37238 52991
rect 36866 52790 36959 52856
rect 36866 52774 36943 52790
tri 36943 52774 36959 52790 nw
rect 36995 52757 37109 52915
rect 37145 52790 37238 52856
tri 37145 52774 37161 52790 ne
rect 37161 52774 37238 52790
rect 36978 52675 37126 52757
rect 36866 52642 36943 52658
tri 36943 52642 36959 52658 sw
rect 36866 52576 36959 52642
rect 36866 52474 36959 52540
rect 36866 52458 36943 52474
tri 36943 52458 36959 52474 nw
rect 36995 52441 37109 52675
tri 37145 52642 37161 52658 se
rect 37161 52642 37238 52658
rect 37145 52576 37238 52642
rect 37145 52474 37238 52540
tri 37145 52458 37161 52474 ne
rect 37161 52458 37238 52474
rect 36978 52359 37126 52441
rect 36866 52326 36943 52342
tri 36943 52326 36959 52342 sw
rect 36866 52260 36959 52326
rect 36995 52201 37109 52359
tri 37145 52326 37161 52342 se
rect 37161 52326 37238 52342
rect 37145 52260 37238 52326
rect 36866 52125 37238 52201
rect 36866 52000 36959 52066
rect 36866 51984 36943 52000
tri 36943 51984 36959 52000 nw
rect 36995 51967 37109 52125
rect 37145 52000 37238 52066
tri 37145 51984 37161 52000 ne
rect 37161 51984 37238 52000
rect 36978 51885 37126 51967
rect 36866 51852 36943 51868
tri 36943 51852 36959 51868 sw
rect 36866 51786 36959 51852
rect 36866 51684 36959 51750
rect 36866 51668 36943 51684
tri 36943 51668 36959 51684 nw
rect 36995 51651 37109 51885
tri 37145 51852 37161 51868 se
rect 37161 51852 37238 51868
rect 37145 51786 37238 51852
rect 37145 51684 37238 51750
tri 37145 51668 37161 51684 ne
rect 37161 51668 37238 51684
rect 36978 51569 37126 51651
rect 36866 51536 36943 51552
tri 36943 51536 36959 51552 sw
rect 36866 51470 36959 51536
rect 36995 51411 37109 51569
tri 37145 51536 37161 51552 se
rect 37161 51536 37238 51552
rect 37145 51470 37238 51536
rect 36866 51335 37238 51411
rect 36866 51210 36959 51276
rect 36866 51194 36943 51210
tri 36943 51194 36959 51210 nw
rect 36995 51177 37109 51335
rect 37145 51210 37238 51276
tri 37145 51194 37161 51210 ne
rect 37161 51194 37238 51210
rect 36978 51095 37126 51177
rect 36866 51062 36943 51078
tri 36943 51062 36959 51078 sw
rect 36866 50996 36959 51062
rect 36866 50894 36959 50960
rect 36866 50878 36943 50894
tri 36943 50878 36959 50894 nw
rect 36995 50861 37109 51095
tri 37145 51062 37161 51078 se
rect 37161 51062 37238 51078
rect 37145 50996 37238 51062
rect 37145 50894 37238 50960
tri 37145 50878 37161 50894 ne
rect 37161 50878 37238 50894
rect 36978 50779 37126 50861
rect 36866 50746 36943 50762
tri 36943 50746 36959 50762 sw
rect 36866 50680 36959 50746
rect 36995 50621 37109 50779
tri 37145 50746 37161 50762 se
rect 37161 50746 37238 50762
rect 37145 50680 37238 50746
rect 36866 50545 37238 50621
rect 36866 50420 36959 50486
rect 36866 50404 36943 50420
tri 36943 50404 36959 50420 nw
rect 36995 50387 37109 50545
rect 37145 50420 37238 50486
tri 37145 50404 37161 50420 ne
rect 37161 50404 37238 50420
rect 36978 50305 37126 50387
rect 36866 50272 36943 50288
tri 36943 50272 36959 50288 sw
rect 36866 50206 36959 50272
rect 36866 50104 36959 50170
rect 36866 50088 36943 50104
tri 36943 50088 36959 50104 nw
rect 36995 50071 37109 50305
tri 37145 50272 37161 50288 se
rect 37161 50272 37238 50288
rect 37145 50206 37238 50272
rect 37145 50104 37238 50170
tri 37145 50088 37161 50104 ne
rect 37161 50088 37238 50104
rect 36978 49989 37126 50071
rect 36866 49956 36943 49972
tri 36943 49956 36959 49972 sw
rect 36866 49890 36959 49956
rect 36995 49831 37109 49989
tri 37145 49956 37161 49972 se
rect 37161 49956 37238 49972
rect 37145 49890 37238 49956
rect 36866 49755 37238 49831
rect 36866 49630 36959 49696
rect 36866 49614 36943 49630
tri 36943 49614 36959 49630 nw
rect 36995 49597 37109 49755
rect 37145 49630 37238 49696
tri 37145 49614 37161 49630 ne
rect 37161 49614 37238 49630
rect 36978 49515 37126 49597
rect 36866 49482 36943 49498
tri 36943 49482 36959 49498 sw
rect 36866 49416 36959 49482
rect 36866 49314 36959 49380
rect 36866 49298 36943 49314
tri 36943 49298 36959 49314 nw
rect 36995 49281 37109 49515
tri 37145 49482 37161 49498 se
rect 37161 49482 37238 49498
rect 37145 49416 37238 49482
rect 37145 49314 37238 49380
tri 37145 49298 37161 49314 ne
rect 37161 49298 37238 49314
rect 36978 49199 37126 49281
rect 36866 49166 36943 49182
tri 36943 49166 36959 49182 sw
rect 36866 49100 36959 49166
rect 36995 49041 37109 49199
tri 37145 49166 37161 49182 se
rect 37161 49166 37238 49182
rect 37145 49100 37238 49166
rect 36866 48965 37238 49041
rect 36866 48840 36959 48906
rect 36866 48824 36943 48840
tri 36943 48824 36959 48840 nw
rect 36995 48807 37109 48965
rect 37145 48840 37238 48906
tri 37145 48824 37161 48840 ne
rect 37161 48824 37238 48840
rect 36978 48725 37126 48807
rect 36866 48692 36943 48708
tri 36943 48692 36959 48708 sw
rect 36866 48626 36959 48692
rect 36866 48524 36959 48590
rect 36866 48508 36943 48524
tri 36943 48508 36959 48524 nw
rect 36995 48491 37109 48725
tri 37145 48692 37161 48708 se
rect 37161 48692 37238 48708
rect 37145 48626 37238 48692
rect 37145 48524 37238 48590
tri 37145 48508 37161 48524 ne
rect 37161 48508 37238 48524
rect 36978 48409 37126 48491
rect 36866 48376 36943 48392
tri 36943 48376 36959 48392 sw
rect 36866 48310 36959 48376
rect 36995 48251 37109 48409
tri 37145 48376 37161 48392 se
rect 37161 48376 37238 48392
rect 37145 48310 37238 48376
rect 36866 48175 37238 48251
rect 36866 48050 36959 48116
rect 36866 48034 36943 48050
tri 36943 48034 36959 48050 nw
rect 36995 48017 37109 48175
rect 37145 48050 37238 48116
tri 37145 48034 37161 48050 ne
rect 37161 48034 37238 48050
rect 36978 47935 37126 48017
rect 36866 47902 36943 47918
tri 36943 47902 36959 47918 sw
rect 36866 47836 36959 47902
rect 36866 47734 36959 47800
rect 36866 47718 36943 47734
tri 36943 47718 36959 47734 nw
rect 36995 47701 37109 47935
tri 37145 47902 37161 47918 se
rect 37161 47902 37238 47918
rect 37145 47836 37238 47902
rect 37145 47734 37238 47800
tri 37145 47718 37161 47734 ne
rect 37161 47718 37238 47734
rect 36978 47619 37126 47701
rect 36866 47586 36943 47602
tri 36943 47586 36959 47602 sw
rect 36866 47520 36959 47586
rect 36995 47461 37109 47619
tri 37145 47586 37161 47602 se
rect 37161 47586 37238 47602
rect 37145 47520 37238 47586
rect 36866 47385 37238 47461
rect 36866 47260 36959 47326
rect 36866 47244 36943 47260
tri 36943 47244 36959 47260 nw
rect 36995 47227 37109 47385
rect 37145 47260 37238 47326
tri 37145 47244 37161 47260 ne
rect 37161 47244 37238 47260
rect 36978 47145 37126 47227
rect 36866 47112 36943 47128
tri 36943 47112 36959 47128 sw
rect 36866 47046 36959 47112
rect 36866 46944 36959 47010
rect 36866 46928 36943 46944
tri 36943 46928 36959 46944 nw
rect 36995 46911 37109 47145
tri 37145 47112 37161 47128 se
rect 37161 47112 37238 47128
rect 37145 47046 37238 47112
rect 37145 46944 37238 47010
tri 37145 46928 37161 46944 ne
rect 37161 46928 37238 46944
rect 36978 46829 37126 46911
rect 36866 46796 36943 46812
tri 36943 46796 36959 46812 sw
rect 36866 46730 36959 46796
rect 36995 46671 37109 46829
tri 37145 46796 37161 46812 se
rect 37161 46796 37238 46812
rect 37145 46730 37238 46796
rect 36866 46595 37238 46671
rect 36866 46470 36959 46536
rect 36866 46454 36943 46470
tri 36943 46454 36959 46470 nw
rect 36995 46437 37109 46595
rect 37145 46470 37238 46536
tri 37145 46454 37161 46470 ne
rect 37161 46454 37238 46470
rect 36978 46355 37126 46437
rect 36866 46322 36943 46338
tri 36943 46322 36959 46338 sw
rect 36866 46256 36959 46322
rect 36866 46154 36959 46220
rect 36866 46138 36943 46154
tri 36943 46138 36959 46154 nw
rect 36995 46121 37109 46355
tri 37145 46322 37161 46338 se
rect 37161 46322 37238 46338
rect 37145 46256 37238 46322
rect 37145 46154 37238 46220
tri 37145 46138 37161 46154 ne
rect 37161 46138 37238 46154
rect 36978 46039 37126 46121
rect 36866 46006 36943 46022
tri 36943 46006 36959 46022 sw
rect 36866 45940 36959 46006
rect 36995 45881 37109 46039
tri 37145 46006 37161 46022 se
rect 37161 46006 37238 46022
rect 37145 45940 37238 46006
rect 36866 45805 37238 45881
rect 36866 45680 36959 45746
rect 36866 45664 36943 45680
tri 36943 45664 36959 45680 nw
rect 36995 45647 37109 45805
rect 37145 45680 37238 45746
tri 37145 45664 37161 45680 ne
rect 37161 45664 37238 45680
rect 36978 45565 37126 45647
rect 36866 45532 36943 45548
tri 36943 45532 36959 45548 sw
rect 36866 45466 36959 45532
rect 36866 45364 36959 45430
rect 36866 45348 36943 45364
tri 36943 45348 36959 45364 nw
rect 36995 45331 37109 45565
tri 37145 45532 37161 45548 se
rect 37161 45532 37238 45548
rect 37145 45466 37238 45532
rect 37145 45364 37238 45430
tri 37145 45348 37161 45364 ne
rect 37161 45348 37238 45364
rect 36978 45249 37126 45331
rect 36866 45216 36943 45232
tri 36943 45216 36959 45232 sw
rect 36866 45150 36959 45216
rect 36995 45091 37109 45249
tri 37145 45216 37161 45232 se
rect 37161 45216 37238 45232
rect 37145 45150 37238 45216
rect 36866 45015 37238 45091
rect 36866 44890 36959 44956
rect 36866 44874 36943 44890
tri 36943 44874 36959 44890 nw
rect 36995 44857 37109 45015
rect 37145 44890 37238 44956
tri 37145 44874 37161 44890 ne
rect 37161 44874 37238 44890
rect 36978 44775 37126 44857
rect 36866 44742 36943 44758
tri 36943 44742 36959 44758 sw
rect 36866 44676 36959 44742
rect 36866 44574 36959 44640
rect 36866 44558 36943 44574
tri 36943 44558 36959 44574 nw
rect 36995 44541 37109 44775
tri 37145 44742 37161 44758 se
rect 37161 44742 37238 44758
rect 37145 44676 37238 44742
rect 37145 44574 37238 44640
tri 37145 44558 37161 44574 ne
rect 37161 44558 37238 44574
rect 36978 44459 37126 44541
rect 36866 44426 36943 44442
tri 36943 44426 36959 44442 sw
rect 36866 44360 36959 44426
rect 36995 44301 37109 44459
tri 37145 44426 37161 44442 se
rect 37161 44426 37238 44442
rect 37145 44360 37238 44426
rect 36866 44225 37238 44301
rect 36866 44100 36959 44166
rect 36866 44084 36943 44100
tri 36943 44084 36959 44100 nw
rect 36995 44067 37109 44225
rect 37145 44100 37238 44166
tri 37145 44084 37161 44100 ne
rect 37161 44084 37238 44100
rect 36978 43985 37126 44067
rect 36866 43952 36943 43968
tri 36943 43952 36959 43968 sw
rect 36866 43886 36959 43952
rect 36866 43784 36959 43850
rect 36866 43768 36943 43784
tri 36943 43768 36959 43784 nw
rect 36995 43751 37109 43985
tri 37145 43952 37161 43968 se
rect 37161 43952 37238 43968
rect 37145 43886 37238 43952
rect 37145 43784 37238 43850
tri 37145 43768 37161 43784 ne
rect 37161 43768 37238 43784
rect 36978 43669 37126 43751
rect 36866 43636 36943 43652
tri 36943 43636 36959 43652 sw
rect 36866 43570 36959 43636
rect 36995 43511 37109 43669
tri 37145 43636 37161 43652 se
rect 37161 43636 37238 43652
rect 37145 43570 37238 43636
rect 36866 43435 37238 43511
rect 36866 43310 36959 43376
rect 36866 43294 36943 43310
tri 36943 43294 36959 43310 nw
rect 36995 43277 37109 43435
rect 37145 43310 37238 43376
tri 37145 43294 37161 43310 ne
rect 37161 43294 37238 43310
rect 36978 43195 37126 43277
rect 36866 43162 36943 43178
tri 36943 43162 36959 43178 sw
rect 36866 43096 36959 43162
rect 36866 42994 36959 43060
rect 36866 42978 36943 42994
tri 36943 42978 36959 42994 nw
rect 36995 42961 37109 43195
tri 37145 43162 37161 43178 se
rect 37161 43162 37238 43178
rect 37145 43096 37238 43162
rect 37145 42994 37238 43060
tri 37145 42978 37161 42994 ne
rect 37161 42978 37238 42994
rect 36978 42879 37126 42961
rect 36866 42846 36943 42862
tri 36943 42846 36959 42862 sw
rect 36866 42780 36959 42846
rect 36995 42721 37109 42879
tri 37145 42846 37161 42862 se
rect 37161 42846 37238 42862
rect 37145 42780 37238 42846
rect 36866 42645 37238 42721
rect 36866 42520 36959 42586
rect 36866 42504 36943 42520
tri 36943 42504 36959 42520 nw
rect 36995 42487 37109 42645
rect 37145 42520 37238 42586
tri 37145 42504 37161 42520 ne
rect 37161 42504 37238 42520
rect 36978 42405 37126 42487
rect 36866 42372 36943 42388
tri 36943 42372 36959 42388 sw
rect 36866 42306 36959 42372
rect 36866 42204 36959 42270
rect 36866 42188 36943 42204
tri 36943 42188 36959 42204 nw
rect 36995 42171 37109 42405
tri 37145 42372 37161 42388 se
rect 37161 42372 37238 42388
rect 37145 42306 37238 42372
rect 37145 42204 37238 42270
tri 37145 42188 37161 42204 ne
rect 37161 42188 37238 42204
rect 36978 42089 37126 42171
rect 36866 42056 36943 42072
tri 36943 42056 36959 42072 sw
rect 36866 41990 36959 42056
rect 36995 41931 37109 42089
tri 37145 42056 37161 42072 se
rect 37161 42056 37238 42072
rect 37145 41990 37238 42056
rect 36866 41855 37238 41931
rect 36866 41730 36959 41796
rect 36866 41714 36943 41730
tri 36943 41714 36959 41730 nw
rect 36995 41697 37109 41855
rect 37145 41730 37238 41796
tri 37145 41714 37161 41730 ne
rect 37161 41714 37238 41730
rect 36978 41615 37126 41697
rect 36866 41582 36943 41598
tri 36943 41582 36959 41598 sw
rect 36866 41516 36959 41582
rect 36866 41414 36959 41480
rect 36866 41398 36943 41414
tri 36943 41398 36959 41414 nw
rect 36995 41381 37109 41615
tri 37145 41582 37161 41598 se
rect 37161 41582 37238 41598
rect 37145 41516 37238 41582
rect 37145 41414 37238 41480
tri 37145 41398 37161 41414 ne
rect 37161 41398 37238 41414
rect 36978 41299 37126 41381
rect 36866 41266 36943 41282
tri 36943 41266 36959 41282 sw
rect 36866 41200 36959 41266
rect 36995 41141 37109 41299
tri 37145 41266 37161 41282 se
rect 37161 41266 37238 41282
rect 37145 41200 37238 41266
rect 36866 41065 37238 41141
rect 36866 40940 36959 41006
rect 36866 40924 36943 40940
tri 36943 40924 36959 40940 nw
rect 36995 40907 37109 41065
rect 37145 40940 37238 41006
tri 37145 40924 37161 40940 ne
rect 37161 40924 37238 40940
rect 36978 40825 37126 40907
rect 36866 40792 36943 40808
tri 36943 40792 36959 40808 sw
rect 36866 40726 36959 40792
rect 36866 40624 36959 40690
rect 36866 40608 36943 40624
tri 36943 40608 36959 40624 nw
rect 36995 40591 37109 40825
tri 37145 40792 37161 40808 se
rect 37161 40792 37238 40808
rect 37145 40726 37238 40792
rect 37145 40624 37238 40690
tri 37145 40608 37161 40624 ne
rect 37161 40608 37238 40624
rect 36978 40509 37126 40591
rect 36866 40476 36943 40492
tri 36943 40476 36959 40492 sw
rect 36866 40410 36959 40476
rect 36995 40351 37109 40509
tri 37145 40476 37161 40492 se
rect 37161 40476 37238 40492
rect 37145 40410 37238 40476
rect 36866 40275 37238 40351
rect 36866 40150 36959 40216
rect 36866 40134 36943 40150
tri 36943 40134 36959 40150 nw
rect 36995 40117 37109 40275
rect 37145 40150 37238 40216
tri 37145 40134 37161 40150 ne
rect 37161 40134 37238 40150
rect 36978 40035 37126 40117
rect 36866 40002 36943 40018
tri 36943 40002 36959 40018 sw
rect 36866 39936 36959 40002
rect 36866 39834 36959 39900
rect 36866 39818 36943 39834
tri 36943 39818 36959 39834 nw
rect 36995 39801 37109 40035
tri 37145 40002 37161 40018 se
rect 37161 40002 37238 40018
rect 37145 39936 37238 40002
rect 37145 39834 37238 39900
tri 37145 39818 37161 39834 ne
rect 37161 39818 37238 39834
rect 36978 39719 37126 39801
rect 36866 39686 36943 39702
tri 36943 39686 36959 39702 sw
rect 36866 39620 36959 39686
rect 36995 39561 37109 39719
tri 37145 39686 37161 39702 se
rect 37161 39686 37238 39702
rect 37145 39620 37238 39686
rect 36866 39485 37238 39561
rect 36866 39360 36959 39426
rect 36866 39344 36943 39360
tri 36943 39344 36959 39360 nw
rect 36995 39327 37109 39485
rect 37145 39360 37238 39426
tri 37145 39344 37161 39360 ne
rect 37161 39344 37238 39360
rect 36978 39245 37126 39327
rect 36866 39212 36943 39228
tri 36943 39212 36959 39228 sw
rect 36866 39146 36959 39212
rect 36866 39044 36959 39110
rect 36866 39028 36943 39044
tri 36943 39028 36959 39044 nw
rect 36995 39011 37109 39245
tri 37145 39212 37161 39228 se
rect 37161 39212 37238 39228
rect 37145 39146 37238 39212
rect 37145 39044 37238 39110
tri 37145 39028 37161 39044 ne
rect 37161 39028 37238 39044
rect 36978 38929 37126 39011
rect 36866 38896 36943 38912
tri 36943 38896 36959 38912 sw
rect 36866 38830 36959 38896
rect 36995 38771 37109 38929
tri 37145 38896 37161 38912 se
rect 37161 38896 37238 38912
rect 37145 38830 37238 38896
rect 36866 38695 37238 38771
rect 36866 38570 36959 38636
rect 36866 38554 36943 38570
tri 36943 38554 36959 38570 nw
rect 36995 38537 37109 38695
rect 37145 38570 37238 38636
tri 37145 38554 37161 38570 ne
rect 37161 38554 37238 38570
rect 36978 38455 37126 38537
rect 36866 38422 36943 38438
tri 36943 38422 36959 38438 sw
rect 36866 38356 36959 38422
rect 36866 38254 36959 38320
rect 36866 38238 36943 38254
tri 36943 38238 36959 38254 nw
rect 36995 38221 37109 38455
tri 37145 38422 37161 38438 se
rect 37161 38422 37238 38438
rect 37145 38356 37238 38422
rect 37145 38254 37238 38320
tri 37145 38238 37161 38254 ne
rect 37161 38238 37238 38254
rect 36978 38139 37126 38221
rect 36866 38106 36943 38122
tri 36943 38106 36959 38122 sw
rect 36866 38040 36959 38106
rect 36995 37981 37109 38139
tri 37145 38106 37161 38122 se
rect 37161 38106 37238 38122
rect 37145 38040 37238 38106
rect 36866 37905 37238 37981
rect 36866 37780 36959 37846
rect 36866 37764 36943 37780
tri 36943 37764 36959 37780 nw
rect 36995 37747 37109 37905
rect 37145 37780 37238 37846
tri 37145 37764 37161 37780 ne
rect 37161 37764 37238 37780
rect 36978 37665 37126 37747
rect 36866 37632 36943 37648
tri 36943 37632 36959 37648 sw
rect 36866 37566 36959 37632
rect 36866 37464 36959 37530
rect 36866 37448 36943 37464
tri 36943 37448 36959 37464 nw
rect 36995 37431 37109 37665
tri 37145 37632 37161 37648 se
rect 37161 37632 37238 37648
rect 37145 37566 37238 37632
rect 37145 37464 37238 37530
tri 37145 37448 37161 37464 ne
rect 37161 37448 37238 37464
rect 36978 37349 37126 37431
rect 36866 37316 36943 37332
tri 36943 37316 36959 37332 sw
rect 36866 37250 36959 37316
rect 36995 37191 37109 37349
tri 37145 37316 37161 37332 se
rect 37161 37316 37238 37332
rect 37145 37250 37238 37316
rect 36866 37115 37238 37191
rect 36866 36990 36959 37056
rect 36866 36974 36943 36990
tri 36943 36974 36959 36990 nw
rect 36995 36957 37109 37115
rect 37145 36990 37238 37056
tri 37145 36974 37161 36990 ne
rect 37161 36974 37238 36990
rect 36978 36875 37126 36957
rect 36866 36842 36943 36858
tri 36943 36842 36959 36858 sw
rect 36866 36776 36959 36842
rect 36866 36674 36959 36740
rect 36866 36658 36943 36674
tri 36943 36658 36959 36674 nw
rect 36995 36641 37109 36875
tri 37145 36842 37161 36858 se
rect 37161 36842 37238 36858
rect 37145 36776 37238 36842
rect 37145 36674 37238 36740
tri 37145 36658 37161 36674 ne
rect 37161 36658 37238 36674
rect 36978 36559 37126 36641
rect 36866 36526 36943 36542
tri 36943 36526 36959 36542 sw
rect 36866 36460 36959 36526
rect 36995 36401 37109 36559
tri 37145 36526 37161 36542 se
rect 37161 36526 37238 36542
rect 37145 36460 37238 36526
rect 36866 36325 37238 36401
rect 36866 36200 36959 36266
rect 36866 36184 36943 36200
tri 36943 36184 36959 36200 nw
rect 36995 36167 37109 36325
rect 37145 36200 37238 36266
tri 37145 36184 37161 36200 ne
rect 37161 36184 37238 36200
rect 36978 36085 37126 36167
rect 36866 36052 36943 36068
tri 36943 36052 36959 36068 sw
rect 36866 35986 36959 36052
rect 36866 35884 36959 35950
rect 36866 35868 36943 35884
tri 36943 35868 36959 35884 nw
rect 36995 35851 37109 36085
tri 37145 36052 37161 36068 se
rect 37161 36052 37238 36068
rect 37145 35986 37238 36052
rect 37145 35884 37238 35950
tri 37145 35868 37161 35884 ne
rect 37161 35868 37238 35884
rect 36978 35769 37126 35851
rect 36866 35736 36943 35752
tri 36943 35736 36959 35752 sw
rect 36866 35670 36959 35736
rect 36995 35611 37109 35769
tri 37145 35736 37161 35752 se
rect 37161 35736 37238 35752
rect 37145 35670 37238 35736
rect 36866 35535 37238 35611
rect 36866 35410 36959 35476
rect 36866 35394 36943 35410
tri 36943 35394 36959 35410 nw
rect 36995 35377 37109 35535
rect 37145 35410 37238 35476
tri 37145 35394 37161 35410 ne
rect 37161 35394 37238 35410
rect 36978 35295 37126 35377
rect 36866 35262 36943 35278
tri 36943 35262 36959 35278 sw
rect 36866 35196 36959 35262
rect 36866 35094 36959 35160
rect 36866 35078 36943 35094
tri 36943 35078 36959 35094 nw
rect 36995 35061 37109 35295
tri 37145 35262 37161 35278 se
rect 37161 35262 37238 35278
rect 37145 35196 37238 35262
rect 37145 35094 37238 35160
tri 37145 35078 37161 35094 ne
rect 37161 35078 37238 35094
rect 36978 34979 37126 35061
rect 36866 34946 36943 34962
tri 36943 34946 36959 34962 sw
rect 36866 34880 36959 34946
rect 36995 34821 37109 34979
tri 37145 34946 37161 34962 se
rect 37161 34946 37238 34962
rect 37145 34880 37238 34946
rect 36866 34745 37238 34821
rect 36866 34620 36959 34686
rect 36866 34604 36943 34620
tri 36943 34604 36959 34620 nw
rect 36995 34587 37109 34745
rect 37145 34620 37238 34686
tri 37145 34604 37161 34620 ne
rect 37161 34604 37238 34620
rect 36978 34505 37126 34587
rect 36866 34472 36943 34488
tri 36943 34472 36959 34488 sw
rect 36866 34406 36959 34472
rect 36866 34304 36959 34370
rect 36866 34288 36943 34304
tri 36943 34288 36959 34304 nw
rect 36995 34271 37109 34505
tri 37145 34472 37161 34488 se
rect 37161 34472 37238 34488
rect 37145 34406 37238 34472
rect 37145 34304 37238 34370
tri 37145 34288 37161 34304 ne
rect 37161 34288 37238 34304
rect 36978 34189 37126 34271
rect 36866 34156 36943 34172
tri 36943 34156 36959 34172 sw
rect 36866 34090 36959 34156
rect 36995 34031 37109 34189
tri 37145 34156 37161 34172 se
rect 37161 34156 37238 34172
rect 37145 34090 37238 34156
rect 36866 33955 37238 34031
rect 36866 33830 36959 33896
rect 36866 33814 36943 33830
tri 36943 33814 36959 33830 nw
rect 36995 33797 37109 33955
rect 37145 33830 37238 33896
tri 37145 33814 37161 33830 ne
rect 37161 33814 37238 33830
rect 36978 33715 37126 33797
rect 36866 33682 36943 33698
tri 36943 33682 36959 33698 sw
rect 36866 33616 36959 33682
rect 36866 33514 36959 33580
rect 36866 33498 36943 33514
tri 36943 33498 36959 33514 nw
rect 36995 33481 37109 33715
tri 37145 33682 37161 33698 se
rect 37161 33682 37238 33698
rect 37145 33616 37238 33682
rect 37145 33514 37238 33580
tri 37145 33498 37161 33514 ne
rect 37161 33498 37238 33514
rect 36978 33399 37126 33481
rect 36866 33366 36943 33382
tri 36943 33366 36959 33382 sw
rect 36866 33300 36959 33366
rect 36995 33241 37109 33399
tri 37145 33366 37161 33382 se
rect 37161 33366 37238 33382
rect 37145 33300 37238 33366
rect 36866 33165 37238 33241
rect 36866 33040 36959 33106
rect 36866 33024 36943 33040
tri 36943 33024 36959 33040 nw
rect 36995 33007 37109 33165
rect 37145 33040 37238 33106
tri 37145 33024 37161 33040 ne
rect 37161 33024 37238 33040
rect 36978 32925 37126 33007
rect 36866 32892 36943 32908
tri 36943 32892 36959 32908 sw
rect 36866 32826 36959 32892
rect 36866 32724 36959 32790
rect 36866 32708 36943 32724
tri 36943 32708 36959 32724 nw
rect 36995 32691 37109 32925
tri 37145 32892 37161 32908 se
rect 37161 32892 37238 32908
rect 37145 32826 37238 32892
rect 37145 32724 37238 32790
tri 37145 32708 37161 32724 ne
rect 37161 32708 37238 32724
rect 36978 32609 37126 32691
rect 36866 32576 36943 32592
tri 36943 32576 36959 32592 sw
rect 36866 32510 36959 32576
rect 36995 32451 37109 32609
tri 37145 32576 37161 32592 se
rect 37161 32576 37238 32592
rect 37145 32510 37238 32576
rect 36866 32375 37238 32451
rect 36866 32250 36959 32316
rect 36866 32234 36943 32250
tri 36943 32234 36959 32250 nw
rect 36995 32217 37109 32375
rect 37145 32250 37238 32316
tri 37145 32234 37161 32250 ne
rect 37161 32234 37238 32250
rect 36978 32135 37126 32217
rect 36866 32102 36943 32118
tri 36943 32102 36959 32118 sw
rect 36866 32036 36959 32102
rect 36866 31934 36959 32000
rect 36866 31918 36943 31934
tri 36943 31918 36959 31934 nw
rect 36995 31901 37109 32135
tri 37145 32102 37161 32118 se
rect 37161 32102 37238 32118
rect 37145 32036 37238 32102
rect 37145 31934 37238 32000
tri 37145 31918 37161 31934 ne
rect 37161 31918 37238 31934
rect 36978 31819 37126 31901
rect 36866 31786 36943 31802
tri 36943 31786 36959 31802 sw
rect 36866 31720 36959 31786
rect 36995 31661 37109 31819
tri 37145 31786 37161 31802 se
rect 37161 31786 37238 31802
rect 37145 31720 37238 31786
rect 36866 31585 37238 31661
rect 36866 31460 36959 31526
rect 36866 31444 36943 31460
tri 36943 31444 36959 31460 nw
rect 36995 31427 37109 31585
rect 37145 31460 37238 31526
tri 37145 31444 37161 31460 ne
rect 37161 31444 37238 31460
rect 36978 31345 37126 31427
rect 36866 31312 36943 31328
tri 36943 31312 36959 31328 sw
rect 36866 31246 36959 31312
rect 36866 31144 36959 31210
rect 36866 31128 36943 31144
tri 36943 31128 36959 31144 nw
rect 36995 31111 37109 31345
tri 37145 31312 37161 31328 se
rect 37161 31312 37238 31328
rect 37145 31246 37238 31312
rect 37145 31144 37238 31210
tri 37145 31128 37161 31144 ne
rect 37161 31128 37238 31144
rect 36978 31029 37126 31111
rect 36866 30996 36943 31012
tri 36943 30996 36959 31012 sw
rect 36866 30930 36959 30996
rect 36995 30871 37109 31029
tri 37145 30996 37161 31012 se
rect 37161 30996 37238 31012
rect 37145 30930 37238 30996
rect 36866 30795 37238 30871
rect 36866 30670 36959 30736
rect 36866 30654 36943 30670
tri 36943 30654 36959 30670 nw
rect 36995 30637 37109 30795
rect 37145 30670 37238 30736
tri 37145 30654 37161 30670 ne
rect 37161 30654 37238 30670
rect 36978 30555 37126 30637
rect 36866 30522 36943 30538
tri 36943 30522 36959 30538 sw
rect 36866 30456 36959 30522
rect 36866 30354 36959 30420
rect 36866 30338 36943 30354
tri 36943 30338 36959 30354 nw
rect 36995 30321 37109 30555
tri 37145 30522 37161 30538 se
rect 37161 30522 37238 30538
rect 37145 30456 37238 30522
rect 37145 30354 37238 30420
tri 37145 30338 37161 30354 ne
rect 37161 30338 37238 30354
rect 36978 30239 37126 30321
rect 36866 30206 36943 30222
tri 36943 30206 36959 30222 sw
rect 36866 30140 36959 30206
rect 36995 30081 37109 30239
tri 37145 30206 37161 30222 se
rect 37161 30206 37238 30222
rect 37145 30140 37238 30206
rect 36866 30005 37238 30081
rect 36866 29880 36959 29946
rect 36866 29864 36943 29880
tri 36943 29864 36959 29880 nw
rect 36995 29847 37109 30005
rect 37145 29880 37238 29946
tri 37145 29864 37161 29880 ne
rect 37161 29864 37238 29880
rect 36978 29765 37126 29847
rect 36866 29732 36943 29748
tri 36943 29732 36959 29748 sw
rect 36866 29666 36959 29732
rect 36866 29564 36959 29630
rect 36866 29548 36943 29564
tri 36943 29548 36959 29564 nw
rect 36995 29531 37109 29765
tri 37145 29732 37161 29748 se
rect 37161 29732 37238 29748
rect 37145 29666 37238 29732
rect 37145 29564 37238 29630
tri 37145 29548 37161 29564 ne
rect 37161 29548 37238 29564
rect 36978 29449 37126 29531
rect 36866 29416 36943 29432
tri 36943 29416 36959 29432 sw
rect 36866 29350 36959 29416
rect 36995 29291 37109 29449
tri 37145 29416 37161 29432 se
rect 37161 29416 37238 29432
rect 37145 29350 37238 29416
rect 36866 29215 37238 29291
rect 36866 29090 36959 29156
rect 36866 29074 36943 29090
tri 36943 29074 36959 29090 nw
rect 36995 29057 37109 29215
rect 37145 29090 37238 29156
tri 37145 29074 37161 29090 ne
rect 37161 29074 37238 29090
rect 36978 28975 37126 29057
rect 36866 28942 36943 28958
tri 36943 28942 36959 28958 sw
rect 36866 28876 36959 28942
rect 36995 28833 37109 28975
tri 37145 28942 37161 28958 se
rect 37161 28942 37238 28958
rect 37145 28876 37238 28942
rect 37274 28463 37310 80603
rect 37346 28463 37382 80603
rect 37418 80445 37454 80603
rect 37410 80303 37462 80445
rect 37418 28763 37454 80303
rect 37410 28621 37462 28763
rect 37418 28463 37454 28621
rect 37490 28463 37526 80603
rect 37562 28463 37598 80603
rect 37634 28833 37718 80233
rect 37754 28463 37790 80603
rect 37826 28463 37862 80603
rect 37898 80445 37934 80603
rect 37890 80303 37942 80445
rect 37898 28763 37934 80303
rect 37890 28621 37942 28763
rect 37898 28463 37934 28621
rect 37970 28463 38006 80603
rect 38042 28463 38078 80603
rect 38114 80124 38207 80190
rect 38114 80108 38191 80124
tri 38191 80108 38207 80124 nw
rect 38243 80091 38357 80233
rect 38393 80124 38486 80190
tri 38393 80108 38409 80124 ne
rect 38409 80108 38486 80124
rect 38226 80009 38374 80091
rect 38114 79976 38191 79992
tri 38191 79976 38207 79992 sw
rect 38114 79910 38207 79976
rect 38243 79851 38357 80009
tri 38393 79976 38409 79992 se
rect 38409 79976 38486 79992
rect 38393 79910 38486 79976
rect 38114 79775 38486 79851
rect 38114 79650 38207 79716
rect 38114 79634 38191 79650
tri 38191 79634 38207 79650 nw
rect 38243 79617 38357 79775
rect 38393 79650 38486 79716
tri 38393 79634 38409 79650 ne
rect 38409 79634 38486 79650
rect 38226 79535 38374 79617
rect 38114 79502 38191 79518
tri 38191 79502 38207 79518 sw
rect 38114 79436 38207 79502
rect 38114 79334 38207 79400
rect 38114 79318 38191 79334
tri 38191 79318 38207 79334 nw
rect 38243 79301 38357 79535
tri 38393 79502 38409 79518 se
rect 38409 79502 38486 79518
rect 38393 79436 38486 79502
rect 38393 79334 38486 79400
tri 38393 79318 38409 79334 ne
rect 38409 79318 38486 79334
rect 38226 79219 38374 79301
rect 38114 79186 38191 79202
tri 38191 79186 38207 79202 sw
rect 38114 79120 38207 79186
rect 38243 79061 38357 79219
tri 38393 79186 38409 79202 se
rect 38409 79186 38486 79202
rect 38393 79120 38486 79186
rect 38114 78985 38486 79061
rect 38114 78860 38207 78926
rect 38114 78844 38191 78860
tri 38191 78844 38207 78860 nw
rect 38243 78827 38357 78985
rect 38393 78860 38486 78926
tri 38393 78844 38409 78860 ne
rect 38409 78844 38486 78860
rect 38226 78745 38374 78827
rect 38114 78712 38191 78728
tri 38191 78712 38207 78728 sw
rect 38114 78646 38207 78712
rect 38114 78544 38207 78610
rect 38114 78528 38191 78544
tri 38191 78528 38207 78544 nw
rect 38243 78511 38357 78745
tri 38393 78712 38409 78728 se
rect 38409 78712 38486 78728
rect 38393 78646 38486 78712
rect 38393 78544 38486 78610
tri 38393 78528 38409 78544 ne
rect 38409 78528 38486 78544
rect 38226 78429 38374 78511
rect 38114 78396 38191 78412
tri 38191 78396 38207 78412 sw
rect 38114 78330 38207 78396
rect 38243 78271 38357 78429
tri 38393 78396 38409 78412 se
rect 38409 78396 38486 78412
rect 38393 78330 38486 78396
rect 38114 78195 38486 78271
rect 38114 78070 38207 78136
rect 38114 78054 38191 78070
tri 38191 78054 38207 78070 nw
rect 38243 78037 38357 78195
rect 38393 78070 38486 78136
tri 38393 78054 38409 78070 ne
rect 38409 78054 38486 78070
rect 38226 77955 38374 78037
rect 38114 77922 38191 77938
tri 38191 77922 38207 77938 sw
rect 38114 77856 38207 77922
rect 38114 77754 38207 77820
rect 38114 77738 38191 77754
tri 38191 77738 38207 77754 nw
rect 38243 77721 38357 77955
tri 38393 77922 38409 77938 se
rect 38409 77922 38486 77938
rect 38393 77856 38486 77922
rect 38393 77754 38486 77820
tri 38393 77738 38409 77754 ne
rect 38409 77738 38486 77754
rect 38226 77639 38374 77721
rect 38114 77606 38191 77622
tri 38191 77606 38207 77622 sw
rect 38114 77540 38207 77606
rect 38243 77481 38357 77639
tri 38393 77606 38409 77622 se
rect 38409 77606 38486 77622
rect 38393 77540 38486 77606
rect 38114 77405 38486 77481
rect 38114 77280 38207 77346
rect 38114 77264 38191 77280
tri 38191 77264 38207 77280 nw
rect 38243 77247 38357 77405
rect 38393 77280 38486 77346
tri 38393 77264 38409 77280 ne
rect 38409 77264 38486 77280
rect 38226 77165 38374 77247
rect 38114 77132 38191 77148
tri 38191 77132 38207 77148 sw
rect 38114 77066 38207 77132
rect 38114 76964 38207 77030
rect 38114 76948 38191 76964
tri 38191 76948 38207 76964 nw
rect 38243 76931 38357 77165
tri 38393 77132 38409 77148 se
rect 38409 77132 38486 77148
rect 38393 77066 38486 77132
rect 38393 76964 38486 77030
tri 38393 76948 38409 76964 ne
rect 38409 76948 38486 76964
rect 38226 76849 38374 76931
rect 38114 76816 38191 76832
tri 38191 76816 38207 76832 sw
rect 38114 76750 38207 76816
rect 38243 76691 38357 76849
tri 38393 76816 38409 76832 se
rect 38409 76816 38486 76832
rect 38393 76750 38486 76816
rect 38114 76615 38486 76691
rect 38114 76490 38207 76556
rect 38114 76474 38191 76490
tri 38191 76474 38207 76490 nw
rect 38243 76457 38357 76615
rect 38393 76490 38486 76556
tri 38393 76474 38409 76490 ne
rect 38409 76474 38486 76490
rect 38226 76375 38374 76457
rect 38114 76342 38191 76358
tri 38191 76342 38207 76358 sw
rect 38114 76276 38207 76342
rect 38114 76174 38207 76240
rect 38114 76158 38191 76174
tri 38191 76158 38207 76174 nw
rect 38243 76141 38357 76375
tri 38393 76342 38409 76358 se
rect 38409 76342 38486 76358
rect 38393 76276 38486 76342
rect 38393 76174 38486 76240
tri 38393 76158 38409 76174 ne
rect 38409 76158 38486 76174
rect 38226 76059 38374 76141
rect 38114 76026 38191 76042
tri 38191 76026 38207 76042 sw
rect 38114 75960 38207 76026
rect 38243 75901 38357 76059
tri 38393 76026 38409 76042 se
rect 38409 76026 38486 76042
rect 38393 75960 38486 76026
rect 38114 75825 38486 75901
rect 38114 75700 38207 75766
rect 38114 75684 38191 75700
tri 38191 75684 38207 75700 nw
rect 38243 75667 38357 75825
rect 38393 75700 38486 75766
tri 38393 75684 38409 75700 ne
rect 38409 75684 38486 75700
rect 38226 75585 38374 75667
rect 38114 75552 38191 75568
tri 38191 75552 38207 75568 sw
rect 38114 75486 38207 75552
rect 38114 75384 38207 75450
rect 38114 75368 38191 75384
tri 38191 75368 38207 75384 nw
rect 38243 75351 38357 75585
tri 38393 75552 38409 75568 se
rect 38409 75552 38486 75568
rect 38393 75486 38486 75552
rect 38393 75384 38486 75450
tri 38393 75368 38409 75384 ne
rect 38409 75368 38486 75384
rect 38226 75269 38374 75351
rect 38114 75236 38191 75252
tri 38191 75236 38207 75252 sw
rect 38114 75170 38207 75236
rect 38243 75111 38357 75269
tri 38393 75236 38409 75252 se
rect 38409 75236 38486 75252
rect 38393 75170 38486 75236
rect 38114 75035 38486 75111
rect 38114 74910 38207 74976
rect 38114 74894 38191 74910
tri 38191 74894 38207 74910 nw
rect 38243 74877 38357 75035
rect 38393 74910 38486 74976
tri 38393 74894 38409 74910 ne
rect 38409 74894 38486 74910
rect 38226 74795 38374 74877
rect 38114 74762 38191 74778
tri 38191 74762 38207 74778 sw
rect 38114 74696 38207 74762
rect 38114 74594 38207 74660
rect 38114 74578 38191 74594
tri 38191 74578 38207 74594 nw
rect 38243 74561 38357 74795
tri 38393 74762 38409 74778 se
rect 38409 74762 38486 74778
rect 38393 74696 38486 74762
rect 38393 74594 38486 74660
tri 38393 74578 38409 74594 ne
rect 38409 74578 38486 74594
rect 38226 74479 38374 74561
rect 38114 74446 38191 74462
tri 38191 74446 38207 74462 sw
rect 38114 74380 38207 74446
rect 38243 74321 38357 74479
tri 38393 74446 38409 74462 se
rect 38409 74446 38486 74462
rect 38393 74380 38486 74446
rect 38114 74245 38486 74321
rect 38114 74120 38207 74186
rect 38114 74104 38191 74120
tri 38191 74104 38207 74120 nw
rect 38243 74087 38357 74245
rect 38393 74120 38486 74186
tri 38393 74104 38409 74120 ne
rect 38409 74104 38486 74120
rect 38226 74005 38374 74087
rect 38114 73972 38191 73988
tri 38191 73972 38207 73988 sw
rect 38114 73906 38207 73972
rect 38114 73804 38207 73870
rect 38114 73788 38191 73804
tri 38191 73788 38207 73804 nw
rect 38243 73771 38357 74005
tri 38393 73972 38409 73988 se
rect 38409 73972 38486 73988
rect 38393 73906 38486 73972
rect 38393 73804 38486 73870
tri 38393 73788 38409 73804 ne
rect 38409 73788 38486 73804
rect 38226 73689 38374 73771
rect 38114 73656 38191 73672
tri 38191 73656 38207 73672 sw
rect 38114 73590 38207 73656
rect 38243 73531 38357 73689
tri 38393 73656 38409 73672 se
rect 38409 73656 38486 73672
rect 38393 73590 38486 73656
rect 38114 73455 38486 73531
rect 38114 73330 38207 73396
rect 38114 73314 38191 73330
tri 38191 73314 38207 73330 nw
rect 38243 73297 38357 73455
rect 38393 73330 38486 73396
tri 38393 73314 38409 73330 ne
rect 38409 73314 38486 73330
rect 38226 73215 38374 73297
rect 38114 73182 38191 73198
tri 38191 73182 38207 73198 sw
rect 38114 73116 38207 73182
rect 38114 73014 38207 73080
rect 38114 72998 38191 73014
tri 38191 72998 38207 73014 nw
rect 38243 72981 38357 73215
tri 38393 73182 38409 73198 se
rect 38409 73182 38486 73198
rect 38393 73116 38486 73182
rect 38393 73014 38486 73080
tri 38393 72998 38409 73014 ne
rect 38409 72998 38486 73014
rect 38226 72899 38374 72981
rect 38114 72866 38191 72882
tri 38191 72866 38207 72882 sw
rect 38114 72800 38207 72866
rect 38243 72741 38357 72899
tri 38393 72866 38409 72882 se
rect 38409 72866 38486 72882
rect 38393 72800 38486 72866
rect 38114 72665 38486 72741
rect 38114 72540 38207 72606
rect 38114 72524 38191 72540
tri 38191 72524 38207 72540 nw
rect 38243 72507 38357 72665
rect 38393 72540 38486 72606
tri 38393 72524 38409 72540 ne
rect 38409 72524 38486 72540
rect 38226 72425 38374 72507
rect 38114 72392 38191 72408
tri 38191 72392 38207 72408 sw
rect 38114 72326 38207 72392
rect 38114 72224 38207 72290
rect 38114 72208 38191 72224
tri 38191 72208 38207 72224 nw
rect 38243 72191 38357 72425
tri 38393 72392 38409 72408 se
rect 38409 72392 38486 72408
rect 38393 72326 38486 72392
rect 38393 72224 38486 72290
tri 38393 72208 38409 72224 ne
rect 38409 72208 38486 72224
rect 38226 72109 38374 72191
rect 38114 72076 38191 72092
tri 38191 72076 38207 72092 sw
rect 38114 72010 38207 72076
rect 38243 71951 38357 72109
tri 38393 72076 38409 72092 se
rect 38409 72076 38486 72092
rect 38393 72010 38486 72076
rect 38114 71875 38486 71951
rect 38114 71750 38207 71816
rect 38114 71734 38191 71750
tri 38191 71734 38207 71750 nw
rect 38243 71717 38357 71875
rect 38393 71750 38486 71816
tri 38393 71734 38409 71750 ne
rect 38409 71734 38486 71750
rect 38226 71635 38374 71717
rect 38114 71602 38191 71618
tri 38191 71602 38207 71618 sw
rect 38114 71536 38207 71602
rect 38114 71434 38207 71500
rect 38114 71418 38191 71434
tri 38191 71418 38207 71434 nw
rect 38243 71401 38357 71635
tri 38393 71602 38409 71618 se
rect 38409 71602 38486 71618
rect 38393 71536 38486 71602
rect 38393 71434 38486 71500
tri 38393 71418 38409 71434 ne
rect 38409 71418 38486 71434
rect 38226 71319 38374 71401
rect 38114 71286 38191 71302
tri 38191 71286 38207 71302 sw
rect 38114 71220 38207 71286
rect 38243 71161 38357 71319
tri 38393 71286 38409 71302 se
rect 38409 71286 38486 71302
rect 38393 71220 38486 71286
rect 38114 71085 38486 71161
rect 38114 70960 38207 71026
rect 38114 70944 38191 70960
tri 38191 70944 38207 70960 nw
rect 38243 70927 38357 71085
rect 38393 70960 38486 71026
tri 38393 70944 38409 70960 ne
rect 38409 70944 38486 70960
rect 38226 70845 38374 70927
rect 38114 70812 38191 70828
tri 38191 70812 38207 70828 sw
rect 38114 70746 38207 70812
rect 38114 70644 38207 70710
rect 38114 70628 38191 70644
tri 38191 70628 38207 70644 nw
rect 38243 70611 38357 70845
tri 38393 70812 38409 70828 se
rect 38409 70812 38486 70828
rect 38393 70746 38486 70812
rect 38393 70644 38486 70710
tri 38393 70628 38409 70644 ne
rect 38409 70628 38486 70644
rect 38226 70529 38374 70611
rect 38114 70496 38191 70512
tri 38191 70496 38207 70512 sw
rect 38114 70430 38207 70496
rect 38243 70371 38357 70529
tri 38393 70496 38409 70512 se
rect 38409 70496 38486 70512
rect 38393 70430 38486 70496
rect 38114 70295 38486 70371
rect 38114 70170 38207 70236
rect 38114 70154 38191 70170
tri 38191 70154 38207 70170 nw
rect 38243 70137 38357 70295
rect 38393 70170 38486 70236
tri 38393 70154 38409 70170 ne
rect 38409 70154 38486 70170
rect 38226 70055 38374 70137
rect 38114 70022 38191 70038
tri 38191 70022 38207 70038 sw
rect 38114 69956 38207 70022
rect 38114 69854 38207 69920
rect 38114 69838 38191 69854
tri 38191 69838 38207 69854 nw
rect 38243 69821 38357 70055
tri 38393 70022 38409 70038 se
rect 38409 70022 38486 70038
rect 38393 69956 38486 70022
rect 38393 69854 38486 69920
tri 38393 69838 38409 69854 ne
rect 38409 69838 38486 69854
rect 38226 69739 38374 69821
rect 38114 69706 38191 69722
tri 38191 69706 38207 69722 sw
rect 38114 69640 38207 69706
rect 38243 69581 38357 69739
tri 38393 69706 38409 69722 se
rect 38409 69706 38486 69722
rect 38393 69640 38486 69706
rect 38114 69505 38486 69581
rect 38114 69380 38207 69446
rect 38114 69364 38191 69380
tri 38191 69364 38207 69380 nw
rect 38243 69347 38357 69505
rect 38393 69380 38486 69446
tri 38393 69364 38409 69380 ne
rect 38409 69364 38486 69380
rect 38226 69265 38374 69347
rect 38114 69232 38191 69248
tri 38191 69232 38207 69248 sw
rect 38114 69166 38207 69232
rect 38114 69064 38207 69130
rect 38114 69048 38191 69064
tri 38191 69048 38207 69064 nw
rect 38243 69031 38357 69265
tri 38393 69232 38409 69248 se
rect 38409 69232 38486 69248
rect 38393 69166 38486 69232
rect 38393 69064 38486 69130
tri 38393 69048 38409 69064 ne
rect 38409 69048 38486 69064
rect 38226 68949 38374 69031
rect 38114 68916 38191 68932
tri 38191 68916 38207 68932 sw
rect 38114 68850 38207 68916
rect 38243 68791 38357 68949
tri 38393 68916 38409 68932 se
rect 38409 68916 38486 68932
rect 38393 68850 38486 68916
rect 38114 68715 38486 68791
rect 38114 68590 38207 68656
rect 38114 68574 38191 68590
tri 38191 68574 38207 68590 nw
rect 38243 68557 38357 68715
rect 38393 68590 38486 68656
tri 38393 68574 38409 68590 ne
rect 38409 68574 38486 68590
rect 38226 68475 38374 68557
rect 38114 68442 38191 68458
tri 38191 68442 38207 68458 sw
rect 38114 68376 38207 68442
rect 38114 68274 38207 68340
rect 38114 68258 38191 68274
tri 38191 68258 38207 68274 nw
rect 38243 68241 38357 68475
tri 38393 68442 38409 68458 se
rect 38409 68442 38486 68458
rect 38393 68376 38486 68442
rect 38393 68274 38486 68340
tri 38393 68258 38409 68274 ne
rect 38409 68258 38486 68274
rect 38226 68159 38374 68241
rect 38114 68126 38191 68142
tri 38191 68126 38207 68142 sw
rect 38114 68060 38207 68126
rect 38243 68001 38357 68159
tri 38393 68126 38409 68142 se
rect 38409 68126 38486 68142
rect 38393 68060 38486 68126
rect 38114 67925 38486 68001
rect 38114 67800 38207 67866
rect 38114 67784 38191 67800
tri 38191 67784 38207 67800 nw
rect 38243 67767 38357 67925
rect 38393 67800 38486 67866
tri 38393 67784 38409 67800 ne
rect 38409 67784 38486 67800
rect 38226 67685 38374 67767
rect 38114 67652 38191 67668
tri 38191 67652 38207 67668 sw
rect 38114 67586 38207 67652
rect 38114 67484 38207 67550
rect 38114 67468 38191 67484
tri 38191 67468 38207 67484 nw
rect 38243 67451 38357 67685
tri 38393 67652 38409 67668 se
rect 38409 67652 38486 67668
rect 38393 67586 38486 67652
rect 38393 67484 38486 67550
tri 38393 67468 38409 67484 ne
rect 38409 67468 38486 67484
rect 38226 67369 38374 67451
rect 38114 67336 38191 67352
tri 38191 67336 38207 67352 sw
rect 38114 67270 38207 67336
rect 38243 67211 38357 67369
tri 38393 67336 38409 67352 se
rect 38409 67336 38486 67352
rect 38393 67270 38486 67336
rect 38114 67135 38486 67211
rect 38114 67010 38207 67076
rect 38114 66994 38191 67010
tri 38191 66994 38207 67010 nw
rect 38243 66977 38357 67135
rect 38393 67010 38486 67076
tri 38393 66994 38409 67010 ne
rect 38409 66994 38486 67010
rect 38226 66895 38374 66977
rect 38114 66862 38191 66878
tri 38191 66862 38207 66878 sw
rect 38114 66796 38207 66862
rect 38114 66694 38207 66760
rect 38114 66678 38191 66694
tri 38191 66678 38207 66694 nw
rect 38243 66661 38357 66895
tri 38393 66862 38409 66878 se
rect 38409 66862 38486 66878
rect 38393 66796 38486 66862
rect 38393 66694 38486 66760
tri 38393 66678 38409 66694 ne
rect 38409 66678 38486 66694
rect 38226 66579 38374 66661
rect 38114 66546 38191 66562
tri 38191 66546 38207 66562 sw
rect 38114 66480 38207 66546
rect 38243 66421 38357 66579
tri 38393 66546 38409 66562 se
rect 38409 66546 38486 66562
rect 38393 66480 38486 66546
rect 38114 66345 38486 66421
rect 38114 66220 38207 66286
rect 38114 66204 38191 66220
tri 38191 66204 38207 66220 nw
rect 38243 66187 38357 66345
rect 38393 66220 38486 66286
tri 38393 66204 38409 66220 ne
rect 38409 66204 38486 66220
rect 38226 66105 38374 66187
rect 38114 66072 38191 66088
tri 38191 66072 38207 66088 sw
rect 38114 66006 38207 66072
rect 38114 65904 38207 65970
rect 38114 65888 38191 65904
tri 38191 65888 38207 65904 nw
rect 38243 65871 38357 66105
tri 38393 66072 38409 66088 se
rect 38409 66072 38486 66088
rect 38393 66006 38486 66072
rect 38393 65904 38486 65970
tri 38393 65888 38409 65904 ne
rect 38409 65888 38486 65904
rect 38226 65789 38374 65871
rect 38114 65756 38191 65772
tri 38191 65756 38207 65772 sw
rect 38114 65690 38207 65756
rect 38243 65631 38357 65789
tri 38393 65756 38409 65772 se
rect 38409 65756 38486 65772
rect 38393 65690 38486 65756
rect 38114 65555 38486 65631
rect 38114 65430 38207 65496
rect 38114 65414 38191 65430
tri 38191 65414 38207 65430 nw
rect 38243 65397 38357 65555
rect 38393 65430 38486 65496
tri 38393 65414 38409 65430 ne
rect 38409 65414 38486 65430
rect 38226 65315 38374 65397
rect 38114 65282 38191 65298
tri 38191 65282 38207 65298 sw
rect 38114 65216 38207 65282
rect 38114 65114 38207 65180
rect 38114 65098 38191 65114
tri 38191 65098 38207 65114 nw
rect 38243 65081 38357 65315
tri 38393 65282 38409 65298 se
rect 38409 65282 38486 65298
rect 38393 65216 38486 65282
rect 38393 65114 38486 65180
tri 38393 65098 38409 65114 ne
rect 38409 65098 38486 65114
rect 38226 64999 38374 65081
rect 38114 64966 38191 64982
tri 38191 64966 38207 64982 sw
rect 38114 64900 38207 64966
rect 38243 64841 38357 64999
tri 38393 64966 38409 64982 se
rect 38409 64966 38486 64982
rect 38393 64900 38486 64966
rect 38114 64765 38486 64841
rect 38114 64640 38207 64706
rect 38114 64624 38191 64640
tri 38191 64624 38207 64640 nw
rect 38243 64607 38357 64765
rect 38393 64640 38486 64706
tri 38393 64624 38409 64640 ne
rect 38409 64624 38486 64640
rect 38226 64525 38374 64607
rect 38114 64492 38191 64508
tri 38191 64492 38207 64508 sw
rect 38114 64426 38207 64492
rect 38114 64324 38207 64390
rect 38114 64308 38191 64324
tri 38191 64308 38207 64324 nw
rect 38243 64291 38357 64525
tri 38393 64492 38409 64508 se
rect 38409 64492 38486 64508
rect 38393 64426 38486 64492
rect 38393 64324 38486 64390
tri 38393 64308 38409 64324 ne
rect 38409 64308 38486 64324
rect 38226 64209 38374 64291
rect 38114 64176 38191 64192
tri 38191 64176 38207 64192 sw
rect 38114 64110 38207 64176
rect 38243 64051 38357 64209
tri 38393 64176 38409 64192 se
rect 38409 64176 38486 64192
rect 38393 64110 38486 64176
rect 38114 63975 38486 64051
rect 38114 63850 38207 63916
rect 38114 63834 38191 63850
tri 38191 63834 38207 63850 nw
rect 38243 63817 38357 63975
rect 38393 63850 38486 63916
tri 38393 63834 38409 63850 ne
rect 38409 63834 38486 63850
rect 38226 63735 38374 63817
rect 38114 63702 38191 63718
tri 38191 63702 38207 63718 sw
rect 38114 63636 38207 63702
rect 38114 63534 38207 63600
rect 38114 63518 38191 63534
tri 38191 63518 38207 63534 nw
rect 38243 63501 38357 63735
tri 38393 63702 38409 63718 se
rect 38409 63702 38486 63718
rect 38393 63636 38486 63702
rect 38393 63534 38486 63600
tri 38393 63518 38409 63534 ne
rect 38409 63518 38486 63534
rect 38226 63419 38374 63501
rect 38114 63386 38191 63402
tri 38191 63386 38207 63402 sw
rect 38114 63320 38207 63386
rect 38243 63261 38357 63419
tri 38393 63386 38409 63402 se
rect 38409 63386 38486 63402
rect 38393 63320 38486 63386
rect 38114 63185 38486 63261
rect 38114 63060 38207 63126
rect 38114 63044 38191 63060
tri 38191 63044 38207 63060 nw
rect 38243 63027 38357 63185
rect 38393 63060 38486 63126
tri 38393 63044 38409 63060 ne
rect 38409 63044 38486 63060
rect 38226 62945 38374 63027
rect 38114 62912 38191 62928
tri 38191 62912 38207 62928 sw
rect 38114 62846 38207 62912
rect 38114 62744 38207 62810
rect 38114 62728 38191 62744
tri 38191 62728 38207 62744 nw
rect 38243 62711 38357 62945
tri 38393 62912 38409 62928 se
rect 38409 62912 38486 62928
rect 38393 62846 38486 62912
rect 38393 62744 38486 62810
tri 38393 62728 38409 62744 ne
rect 38409 62728 38486 62744
rect 38226 62629 38374 62711
rect 38114 62596 38191 62612
tri 38191 62596 38207 62612 sw
rect 38114 62530 38207 62596
rect 38243 62471 38357 62629
tri 38393 62596 38409 62612 se
rect 38409 62596 38486 62612
rect 38393 62530 38486 62596
rect 38114 62395 38486 62471
rect 38114 62270 38207 62336
rect 38114 62254 38191 62270
tri 38191 62254 38207 62270 nw
rect 38243 62237 38357 62395
rect 38393 62270 38486 62336
tri 38393 62254 38409 62270 ne
rect 38409 62254 38486 62270
rect 38226 62155 38374 62237
rect 38114 62122 38191 62138
tri 38191 62122 38207 62138 sw
rect 38114 62056 38207 62122
rect 38114 61954 38207 62020
rect 38114 61938 38191 61954
tri 38191 61938 38207 61954 nw
rect 38243 61921 38357 62155
tri 38393 62122 38409 62138 se
rect 38409 62122 38486 62138
rect 38393 62056 38486 62122
rect 38393 61954 38486 62020
tri 38393 61938 38409 61954 ne
rect 38409 61938 38486 61954
rect 38226 61839 38374 61921
rect 38114 61806 38191 61822
tri 38191 61806 38207 61822 sw
rect 38114 61740 38207 61806
rect 38243 61681 38357 61839
tri 38393 61806 38409 61822 se
rect 38409 61806 38486 61822
rect 38393 61740 38486 61806
rect 38114 61605 38486 61681
rect 38114 61480 38207 61546
rect 38114 61464 38191 61480
tri 38191 61464 38207 61480 nw
rect 38243 61447 38357 61605
rect 38393 61480 38486 61546
tri 38393 61464 38409 61480 ne
rect 38409 61464 38486 61480
rect 38226 61365 38374 61447
rect 38114 61332 38191 61348
tri 38191 61332 38207 61348 sw
rect 38114 61266 38207 61332
rect 38114 61164 38207 61230
rect 38114 61148 38191 61164
tri 38191 61148 38207 61164 nw
rect 38243 61131 38357 61365
tri 38393 61332 38409 61348 se
rect 38409 61332 38486 61348
rect 38393 61266 38486 61332
rect 38393 61164 38486 61230
tri 38393 61148 38409 61164 ne
rect 38409 61148 38486 61164
rect 38226 61049 38374 61131
rect 38114 61016 38191 61032
tri 38191 61016 38207 61032 sw
rect 38114 60950 38207 61016
rect 38243 60891 38357 61049
tri 38393 61016 38409 61032 se
rect 38409 61016 38486 61032
rect 38393 60950 38486 61016
rect 38114 60815 38486 60891
rect 38114 60690 38207 60756
rect 38114 60674 38191 60690
tri 38191 60674 38207 60690 nw
rect 38243 60657 38357 60815
rect 38393 60690 38486 60756
tri 38393 60674 38409 60690 ne
rect 38409 60674 38486 60690
rect 38226 60575 38374 60657
rect 38114 60542 38191 60558
tri 38191 60542 38207 60558 sw
rect 38114 60476 38207 60542
rect 38114 60374 38207 60440
rect 38114 60358 38191 60374
tri 38191 60358 38207 60374 nw
rect 38243 60341 38357 60575
tri 38393 60542 38409 60558 se
rect 38409 60542 38486 60558
rect 38393 60476 38486 60542
rect 38393 60374 38486 60440
tri 38393 60358 38409 60374 ne
rect 38409 60358 38486 60374
rect 38226 60259 38374 60341
rect 38114 60226 38191 60242
tri 38191 60226 38207 60242 sw
rect 38114 60160 38207 60226
rect 38243 60101 38357 60259
tri 38393 60226 38409 60242 se
rect 38409 60226 38486 60242
rect 38393 60160 38486 60226
rect 38114 60025 38486 60101
rect 38114 59900 38207 59966
rect 38114 59884 38191 59900
tri 38191 59884 38207 59900 nw
rect 38243 59867 38357 60025
rect 38393 59900 38486 59966
tri 38393 59884 38409 59900 ne
rect 38409 59884 38486 59900
rect 38226 59785 38374 59867
rect 38114 59752 38191 59768
tri 38191 59752 38207 59768 sw
rect 38114 59686 38207 59752
rect 38114 59584 38207 59650
rect 38114 59568 38191 59584
tri 38191 59568 38207 59584 nw
rect 38243 59551 38357 59785
tri 38393 59752 38409 59768 se
rect 38409 59752 38486 59768
rect 38393 59686 38486 59752
rect 38393 59584 38486 59650
tri 38393 59568 38409 59584 ne
rect 38409 59568 38486 59584
rect 38226 59469 38374 59551
rect 38114 59436 38191 59452
tri 38191 59436 38207 59452 sw
rect 38114 59370 38207 59436
rect 38243 59311 38357 59469
tri 38393 59436 38409 59452 se
rect 38409 59436 38486 59452
rect 38393 59370 38486 59436
rect 38114 59235 38486 59311
rect 38114 59110 38207 59176
rect 38114 59094 38191 59110
tri 38191 59094 38207 59110 nw
rect 38243 59077 38357 59235
rect 38393 59110 38486 59176
tri 38393 59094 38409 59110 ne
rect 38409 59094 38486 59110
rect 38226 58995 38374 59077
rect 38114 58962 38191 58978
tri 38191 58962 38207 58978 sw
rect 38114 58896 38207 58962
rect 38114 58794 38207 58860
rect 38114 58778 38191 58794
tri 38191 58778 38207 58794 nw
rect 38243 58761 38357 58995
tri 38393 58962 38409 58978 se
rect 38409 58962 38486 58978
rect 38393 58896 38486 58962
rect 38393 58794 38486 58860
tri 38393 58778 38409 58794 ne
rect 38409 58778 38486 58794
rect 38226 58679 38374 58761
rect 38114 58646 38191 58662
tri 38191 58646 38207 58662 sw
rect 38114 58580 38207 58646
rect 38243 58521 38357 58679
tri 38393 58646 38409 58662 se
rect 38409 58646 38486 58662
rect 38393 58580 38486 58646
rect 38114 58445 38486 58521
rect 38114 58320 38207 58386
rect 38114 58304 38191 58320
tri 38191 58304 38207 58320 nw
rect 38243 58287 38357 58445
rect 38393 58320 38486 58386
tri 38393 58304 38409 58320 ne
rect 38409 58304 38486 58320
rect 38226 58205 38374 58287
rect 38114 58172 38191 58188
tri 38191 58172 38207 58188 sw
rect 38114 58106 38207 58172
rect 38114 58004 38207 58070
rect 38114 57988 38191 58004
tri 38191 57988 38207 58004 nw
rect 38243 57971 38357 58205
tri 38393 58172 38409 58188 se
rect 38409 58172 38486 58188
rect 38393 58106 38486 58172
rect 38393 58004 38486 58070
tri 38393 57988 38409 58004 ne
rect 38409 57988 38486 58004
rect 38226 57889 38374 57971
rect 38114 57856 38191 57872
tri 38191 57856 38207 57872 sw
rect 38114 57790 38207 57856
rect 38243 57731 38357 57889
tri 38393 57856 38409 57872 se
rect 38409 57856 38486 57872
rect 38393 57790 38486 57856
rect 38114 57655 38486 57731
rect 38114 57530 38207 57596
rect 38114 57514 38191 57530
tri 38191 57514 38207 57530 nw
rect 38243 57497 38357 57655
rect 38393 57530 38486 57596
tri 38393 57514 38409 57530 ne
rect 38409 57514 38486 57530
rect 38226 57415 38374 57497
rect 38114 57382 38191 57398
tri 38191 57382 38207 57398 sw
rect 38114 57316 38207 57382
rect 38114 57214 38207 57280
rect 38114 57198 38191 57214
tri 38191 57198 38207 57214 nw
rect 38243 57181 38357 57415
tri 38393 57382 38409 57398 se
rect 38409 57382 38486 57398
rect 38393 57316 38486 57382
rect 38393 57214 38486 57280
tri 38393 57198 38409 57214 ne
rect 38409 57198 38486 57214
rect 38226 57099 38374 57181
rect 38114 57066 38191 57082
tri 38191 57066 38207 57082 sw
rect 38114 57000 38207 57066
rect 38243 56941 38357 57099
tri 38393 57066 38409 57082 se
rect 38409 57066 38486 57082
rect 38393 57000 38486 57066
rect 38114 56865 38486 56941
rect 38114 56740 38207 56806
rect 38114 56724 38191 56740
tri 38191 56724 38207 56740 nw
rect 38243 56707 38357 56865
rect 38393 56740 38486 56806
tri 38393 56724 38409 56740 ne
rect 38409 56724 38486 56740
rect 38226 56625 38374 56707
rect 38114 56592 38191 56608
tri 38191 56592 38207 56608 sw
rect 38114 56526 38207 56592
rect 38114 56424 38207 56490
rect 38114 56408 38191 56424
tri 38191 56408 38207 56424 nw
rect 38243 56391 38357 56625
tri 38393 56592 38409 56608 se
rect 38409 56592 38486 56608
rect 38393 56526 38486 56592
rect 38393 56424 38486 56490
tri 38393 56408 38409 56424 ne
rect 38409 56408 38486 56424
rect 38226 56309 38374 56391
rect 38114 56276 38191 56292
tri 38191 56276 38207 56292 sw
rect 38114 56210 38207 56276
rect 38243 56151 38357 56309
tri 38393 56276 38409 56292 se
rect 38409 56276 38486 56292
rect 38393 56210 38486 56276
rect 38114 56075 38486 56151
rect 38114 55950 38207 56016
rect 38114 55934 38191 55950
tri 38191 55934 38207 55950 nw
rect 38243 55917 38357 56075
rect 38393 55950 38486 56016
tri 38393 55934 38409 55950 ne
rect 38409 55934 38486 55950
rect 38226 55835 38374 55917
rect 38114 55802 38191 55818
tri 38191 55802 38207 55818 sw
rect 38114 55736 38207 55802
rect 38114 55634 38207 55700
rect 38114 55618 38191 55634
tri 38191 55618 38207 55634 nw
rect 38243 55601 38357 55835
tri 38393 55802 38409 55818 se
rect 38409 55802 38486 55818
rect 38393 55736 38486 55802
rect 38393 55634 38486 55700
tri 38393 55618 38409 55634 ne
rect 38409 55618 38486 55634
rect 38226 55519 38374 55601
rect 38114 55486 38191 55502
tri 38191 55486 38207 55502 sw
rect 38114 55420 38207 55486
rect 38243 55361 38357 55519
tri 38393 55486 38409 55502 se
rect 38409 55486 38486 55502
rect 38393 55420 38486 55486
rect 38114 55285 38486 55361
rect 38114 55160 38207 55226
rect 38114 55144 38191 55160
tri 38191 55144 38207 55160 nw
rect 38243 55127 38357 55285
rect 38393 55160 38486 55226
tri 38393 55144 38409 55160 ne
rect 38409 55144 38486 55160
rect 38226 55045 38374 55127
rect 38114 55012 38191 55028
tri 38191 55012 38207 55028 sw
rect 38114 54946 38207 55012
rect 38114 54844 38207 54910
rect 38114 54828 38191 54844
tri 38191 54828 38207 54844 nw
rect 38243 54811 38357 55045
tri 38393 55012 38409 55028 se
rect 38409 55012 38486 55028
rect 38393 54946 38486 55012
rect 38393 54844 38486 54910
tri 38393 54828 38409 54844 ne
rect 38409 54828 38486 54844
rect 38226 54729 38374 54811
rect 38114 54696 38191 54712
tri 38191 54696 38207 54712 sw
rect 38114 54630 38207 54696
rect 38243 54571 38357 54729
tri 38393 54696 38409 54712 se
rect 38409 54696 38486 54712
rect 38393 54630 38486 54696
rect 38114 54495 38486 54571
rect 38114 54370 38207 54436
rect 38114 54354 38191 54370
tri 38191 54354 38207 54370 nw
rect 38243 54337 38357 54495
rect 38393 54370 38486 54436
tri 38393 54354 38409 54370 ne
rect 38409 54354 38486 54370
rect 38226 54255 38374 54337
rect 38114 54222 38191 54238
tri 38191 54222 38207 54238 sw
rect 38114 54156 38207 54222
rect 38114 54054 38207 54120
rect 38114 54038 38191 54054
tri 38191 54038 38207 54054 nw
rect 38243 54021 38357 54255
tri 38393 54222 38409 54238 se
rect 38409 54222 38486 54238
rect 38393 54156 38486 54222
rect 38393 54054 38486 54120
tri 38393 54038 38409 54054 ne
rect 38409 54038 38486 54054
rect 38226 53939 38374 54021
rect 38114 53906 38191 53922
tri 38191 53906 38207 53922 sw
rect 38114 53840 38207 53906
rect 38243 53781 38357 53939
tri 38393 53906 38409 53922 se
rect 38409 53906 38486 53922
rect 38393 53840 38486 53906
rect 38114 53705 38486 53781
rect 38114 53580 38207 53646
rect 38114 53564 38191 53580
tri 38191 53564 38207 53580 nw
rect 38243 53547 38357 53705
rect 38393 53580 38486 53646
tri 38393 53564 38409 53580 ne
rect 38409 53564 38486 53580
rect 38226 53465 38374 53547
rect 38114 53432 38191 53448
tri 38191 53432 38207 53448 sw
rect 38114 53366 38207 53432
rect 38114 53264 38207 53330
rect 38114 53248 38191 53264
tri 38191 53248 38207 53264 nw
rect 38243 53231 38357 53465
tri 38393 53432 38409 53448 se
rect 38409 53432 38486 53448
rect 38393 53366 38486 53432
rect 38393 53264 38486 53330
tri 38393 53248 38409 53264 ne
rect 38409 53248 38486 53264
rect 38226 53149 38374 53231
rect 38114 53116 38191 53132
tri 38191 53116 38207 53132 sw
rect 38114 53050 38207 53116
rect 38243 52991 38357 53149
tri 38393 53116 38409 53132 se
rect 38409 53116 38486 53132
rect 38393 53050 38486 53116
rect 38114 52915 38486 52991
rect 38114 52790 38207 52856
rect 38114 52774 38191 52790
tri 38191 52774 38207 52790 nw
rect 38243 52757 38357 52915
rect 38393 52790 38486 52856
tri 38393 52774 38409 52790 ne
rect 38409 52774 38486 52790
rect 38226 52675 38374 52757
rect 38114 52642 38191 52658
tri 38191 52642 38207 52658 sw
rect 38114 52576 38207 52642
rect 38114 52474 38207 52540
rect 38114 52458 38191 52474
tri 38191 52458 38207 52474 nw
rect 38243 52441 38357 52675
tri 38393 52642 38409 52658 se
rect 38409 52642 38486 52658
rect 38393 52576 38486 52642
rect 38393 52474 38486 52540
tri 38393 52458 38409 52474 ne
rect 38409 52458 38486 52474
rect 38226 52359 38374 52441
rect 38114 52326 38191 52342
tri 38191 52326 38207 52342 sw
rect 38114 52260 38207 52326
rect 38243 52201 38357 52359
tri 38393 52326 38409 52342 se
rect 38409 52326 38486 52342
rect 38393 52260 38486 52326
rect 38114 52125 38486 52201
rect 38114 52000 38207 52066
rect 38114 51984 38191 52000
tri 38191 51984 38207 52000 nw
rect 38243 51967 38357 52125
rect 38393 52000 38486 52066
tri 38393 51984 38409 52000 ne
rect 38409 51984 38486 52000
rect 38226 51885 38374 51967
rect 38114 51852 38191 51868
tri 38191 51852 38207 51868 sw
rect 38114 51786 38207 51852
rect 38114 51684 38207 51750
rect 38114 51668 38191 51684
tri 38191 51668 38207 51684 nw
rect 38243 51651 38357 51885
tri 38393 51852 38409 51868 se
rect 38409 51852 38486 51868
rect 38393 51786 38486 51852
rect 38393 51684 38486 51750
tri 38393 51668 38409 51684 ne
rect 38409 51668 38486 51684
rect 38226 51569 38374 51651
rect 38114 51536 38191 51552
tri 38191 51536 38207 51552 sw
rect 38114 51470 38207 51536
rect 38243 51411 38357 51569
tri 38393 51536 38409 51552 se
rect 38409 51536 38486 51552
rect 38393 51470 38486 51536
rect 38114 51335 38486 51411
rect 38114 51210 38207 51276
rect 38114 51194 38191 51210
tri 38191 51194 38207 51210 nw
rect 38243 51177 38357 51335
rect 38393 51210 38486 51276
tri 38393 51194 38409 51210 ne
rect 38409 51194 38486 51210
rect 38226 51095 38374 51177
rect 38114 51062 38191 51078
tri 38191 51062 38207 51078 sw
rect 38114 50996 38207 51062
rect 38114 50894 38207 50960
rect 38114 50878 38191 50894
tri 38191 50878 38207 50894 nw
rect 38243 50861 38357 51095
tri 38393 51062 38409 51078 se
rect 38409 51062 38486 51078
rect 38393 50996 38486 51062
rect 38393 50894 38486 50960
tri 38393 50878 38409 50894 ne
rect 38409 50878 38486 50894
rect 38226 50779 38374 50861
rect 38114 50746 38191 50762
tri 38191 50746 38207 50762 sw
rect 38114 50680 38207 50746
rect 38243 50621 38357 50779
tri 38393 50746 38409 50762 se
rect 38409 50746 38486 50762
rect 38393 50680 38486 50746
rect 38114 50545 38486 50621
rect 38114 50420 38207 50486
rect 38114 50404 38191 50420
tri 38191 50404 38207 50420 nw
rect 38243 50387 38357 50545
rect 38393 50420 38486 50486
tri 38393 50404 38409 50420 ne
rect 38409 50404 38486 50420
rect 38226 50305 38374 50387
rect 38114 50272 38191 50288
tri 38191 50272 38207 50288 sw
rect 38114 50206 38207 50272
rect 38114 50104 38207 50170
rect 38114 50088 38191 50104
tri 38191 50088 38207 50104 nw
rect 38243 50071 38357 50305
tri 38393 50272 38409 50288 se
rect 38409 50272 38486 50288
rect 38393 50206 38486 50272
rect 38393 50104 38486 50170
tri 38393 50088 38409 50104 ne
rect 38409 50088 38486 50104
rect 38226 49989 38374 50071
rect 38114 49956 38191 49972
tri 38191 49956 38207 49972 sw
rect 38114 49890 38207 49956
rect 38243 49831 38357 49989
tri 38393 49956 38409 49972 se
rect 38409 49956 38486 49972
rect 38393 49890 38486 49956
rect 38114 49755 38486 49831
rect 38114 49630 38207 49696
rect 38114 49614 38191 49630
tri 38191 49614 38207 49630 nw
rect 38243 49597 38357 49755
rect 38393 49630 38486 49696
tri 38393 49614 38409 49630 ne
rect 38409 49614 38486 49630
rect 38226 49515 38374 49597
rect 38114 49482 38191 49498
tri 38191 49482 38207 49498 sw
rect 38114 49416 38207 49482
rect 38114 49314 38207 49380
rect 38114 49298 38191 49314
tri 38191 49298 38207 49314 nw
rect 38243 49281 38357 49515
tri 38393 49482 38409 49498 se
rect 38409 49482 38486 49498
rect 38393 49416 38486 49482
rect 38393 49314 38486 49380
tri 38393 49298 38409 49314 ne
rect 38409 49298 38486 49314
rect 38226 49199 38374 49281
rect 38114 49166 38191 49182
tri 38191 49166 38207 49182 sw
rect 38114 49100 38207 49166
rect 38243 49041 38357 49199
tri 38393 49166 38409 49182 se
rect 38409 49166 38486 49182
rect 38393 49100 38486 49166
rect 38114 48965 38486 49041
rect 38114 48840 38207 48906
rect 38114 48824 38191 48840
tri 38191 48824 38207 48840 nw
rect 38243 48807 38357 48965
rect 38393 48840 38486 48906
tri 38393 48824 38409 48840 ne
rect 38409 48824 38486 48840
rect 38226 48725 38374 48807
rect 38114 48692 38191 48708
tri 38191 48692 38207 48708 sw
rect 38114 48626 38207 48692
rect 38114 48524 38207 48590
rect 38114 48508 38191 48524
tri 38191 48508 38207 48524 nw
rect 38243 48491 38357 48725
tri 38393 48692 38409 48708 se
rect 38409 48692 38486 48708
rect 38393 48626 38486 48692
rect 38393 48524 38486 48590
tri 38393 48508 38409 48524 ne
rect 38409 48508 38486 48524
rect 38226 48409 38374 48491
rect 38114 48376 38191 48392
tri 38191 48376 38207 48392 sw
rect 38114 48310 38207 48376
rect 38243 48251 38357 48409
tri 38393 48376 38409 48392 se
rect 38409 48376 38486 48392
rect 38393 48310 38486 48376
rect 38114 48175 38486 48251
rect 38114 48050 38207 48116
rect 38114 48034 38191 48050
tri 38191 48034 38207 48050 nw
rect 38243 48017 38357 48175
rect 38393 48050 38486 48116
tri 38393 48034 38409 48050 ne
rect 38409 48034 38486 48050
rect 38226 47935 38374 48017
rect 38114 47902 38191 47918
tri 38191 47902 38207 47918 sw
rect 38114 47836 38207 47902
rect 38114 47734 38207 47800
rect 38114 47718 38191 47734
tri 38191 47718 38207 47734 nw
rect 38243 47701 38357 47935
tri 38393 47902 38409 47918 se
rect 38409 47902 38486 47918
rect 38393 47836 38486 47902
rect 38393 47734 38486 47800
tri 38393 47718 38409 47734 ne
rect 38409 47718 38486 47734
rect 38226 47619 38374 47701
rect 38114 47586 38191 47602
tri 38191 47586 38207 47602 sw
rect 38114 47520 38207 47586
rect 38243 47461 38357 47619
tri 38393 47586 38409 47602 se
rect 38409 47586 38486 47602
rect 38393 47520 38486 47586
rect 38114 47385 38486 47461
rect 38114 47260 38207 47326
rect 38114 47244 38191 47260
tri 38191 47244 38207 47260 nw
rect 38243 47227 38357 47385
rect 38393 47260 38486 47326
tri 38393 47244 38409 47260 ne
rect 38409 47244 38486 47260
rect 38226 47145 38374 47227
rect 38114 47112 38191 47128
tri 38191 47112 38207 47128 sw
rect 38114 47046 38207 47112
rect 38114 46944 38207 47010
rect 38114 46928 38191 46944
tri 38191 46928 38207 46944 nw
rect 38243 46911 38357 47145
tri 38393 47112 38409 47128 se
rect 38409 47112 38486 47128
rect 38393 47046 38486 47112
rect 38393 46944 38486 47010
tri 38393 46928 38409 46944 ne
rect 38409 46928 38486 46944
rect 38226 46829 38374 46911
rect 38114 46796 38191 46812
tri 38191 46796 38207 46812 sw
rect 38114 46730 38207 46796
rect 38243 46671 38357 46829
tri 38393 46796 38409 46812 se
rect 38409 46796 38486 46812
rect 38393 46730 38486 46796
rect 38114 46595 38486 46671
rect 38114 46470 38207 46536
rect 38114 46454 38191 46470
tri 38191 46454 38207 46470 nw
rect 38243 46437 38357 46595
rect 38393 46470 38486 46536
tri 38393 46454 38409 46470 ne
rect 38409 46454 38486 46470
rect 38226 46355 38374 46437
rect 38114 46322 38191 46338
tri 38191 46322 38207 46338 sw
rect 38114 46256 38207 46322
rect 38114 46154 38207 46220
rect 38114 46138 38191 46154
tri 38191 46138 38207 46154 nw
rect 38243 46121 38357 46355
tri 38393 46322 38409 46338 se
rect 38409 46322 38486 46338
rect 38393 46256 38486 46322
rect 38393 46154 38486 46220
tri 38393 46138 38409 46154 ne
rect 38409 46138 38486 46154
rect 38226 46039 38374 46121
rect 38114 46006 38191 46022
tri 38191 46006 38207 46022 sw
rect 38114 45940 38207 46006
rect 38243 45881 38357 46039
tri 38393 46006 38409 46022 se
rect 38409 46006 38486 46022
rect 38393 45940 38486 46006
rect 38114 45805 38486 45881
rect 38114 45680 38207 45746
rect 38114 45664 38191 45680
tri 38191 45664 38207 45680 nw
rect 38243 45647 38357 45805
rect 38393 45680 38486 45746
tri 38393 45664 38409 45680 ne
rect 38409 45664 38486 45680
rect 38226 45565 38374 45647
rect 38114 45532 38191 45548
tri 38191 45532 38207 45548 sw
rect 38114 45466 38207 45532
rect 38114 45364 38207 45430
rect 38114 45348 38191 45364
tri 38191 45348 38207 45364 nw
rect 38243 45331 38357 45565
tri 38393 45532 38409 45548 se
rect 38409 45532 38486 45548
rect 38393 45466 38486 45532
rect 38393 45364 38486 45430
tri 38393 45348 38409 45364 ne
rect 38409 45348 38486 45364
rect 38226 45249 38374 45331
rect 38114 45216 38191 45232
tri 38191 45216 38207 45232 sw
rect 38114 45150 38207 45216
rect 38243 45091 38357 45249
tri 38393 45216 38409 45232 se
rect 38409 45216 38486 45232
rect 38393 45150 38486 45216
rect 38114 45015 38486 45091
rect 38114 44890 38207 44956
rect 38114 44874 38191 44890
tri 38191 44874 38207 44890 nw
rect 38243 44857 38357 45015
rect 38393 44890 38486 44956
tri 38393 44874 38409 44890 ne
rect 38409 44874 38486 44890
rect 38226 44775 38374 44857
rect 38114 44742 38191 44758
tri 38191 44742 38207 44758 sw
rect 38114 44676 38207 44742
rect 38114 44574 38207 44640
rect 38114 44558 38191 44574
tri 38191 44558 38207 44574 nw
rect 38243 44541 38357 44775
tri 38393 44742 38409 44758 se
rect 38409 44742 38486 44758
rect 38393 44676 38486 44742
rect 38393 44574 38486 44640
tri 38393 44558 38409 44574 ne
rect 38409 44558 38486 44574
rect 38226 44459 38374 44541
rect 38114 44426 38191 44442
tri 38191 44426 38207 44442 sw
rect 38114 44360 38207 44426
rect 38243 44301 38357 44459
tri 38393 44426 38409 44442 se
rect 38409 44426 38486 44442
rect 38393 44360 38486 44426
rect 38114 44225 38486 44301
rect 38114 44100 38207 44166
rect 38114 44084 38191 44100
tri 38191 44084 38207 44100 nw
rect 38243 44067 38357 44225
rect 38393 44100 38486 44166
tri 38393 44084 38409 44100 ne
rect 38409 44084 38486 44100
rect 38226 43985 38374 44067
rect 38114 43952 38191 43968
tri 38191 43952 38207 43968 sw
rect 38114 43886 38207 43952
rect 38114 43784 38207 43850
rect 38114 43768 38191 43784
tri 38191 43768 38207 43784 nw
rect 38243 43751 38357 43985
tri 38393 43952 38409 43968 se
rect 38409 43952 38486 43968
rect 38393 43886 38486 43952
rect 38393 43784 38486 43850
tri 38393 43768 38409 43784 ne
rect 38409 43768 38486 43784
rect 38226 43669 38374 43751
rect 38114 43636 38191 43652
tri 38191 43636 38207 43652 sw
rect 38114 43570 38207 43636
rect 38243 43511 38357 43669
tri 38393 43636 38409 43652 se
rect 38409 43636 38486 43652
rect 38393 43570 38486 43636
rect 38114 43435 38486 43511
rect 38114 43310 38207 43376
rect 38114 43294 38191 43310
tri 38191 43294 38207 43310 nw
rect 38243 43277 38357 43435
rect 38393 43310 38486 43376
tri 38393 43294 38409 43310 ne
rect 38409 43294 38486 43310
rect 38226 43195 38374 43277
rect 38114 43162 38191 43178
tri 38191 43162 38207 43178 sw
rect 38114 43096 38207 43162
rect 38114 42994 38207 43060
rect 38114 42978 38191 42994
tri 38191 42978 38207 42994 nw
rect 38243 42961 38357 43195
tri 38393 43162 38409 43178 se
rect 38409 43162 38486 43178
rect 38393 43096 38486 43162
rect 38393 42994 38486 43060
tri 38393 42978 38409 42994 ne
rect 38409 42978 38486 42994
rect 38226 42879 38374 42961
rect 38114 42846 38191 42862
tri 38191 42846 38207 42862 sw
rect 38114 42780 38207 42846
rect 38243 42721 38357 42879
tri 38393 42846 38409 42862 se
rect 38409 42846 38486 42862
rect 38393 42780 38486 42846
rect 38114 42645 38486 42721
rect 38114 42520 38207 42586
rect 38114 42504 38191 42520
tri 38191 42504 38207 42520 nw
rect 38243 42487 38357 42645
rect 38393 42520 38486 42586
tri 38393 42504 38409 42520 ne
rect 38409 42504 38486 42520
rect 38226 42405 38374 42487
rect 38114 42372 38191 42388
tri 38191 42372 38207 42388 sw
rect 38114 42306 38207 42372
rect 38114 42204 38207 42270
rect 38114 42188 38191 42204
tri 38191 42188 38207 42204 nw
rect 38243 42171 38357 42405
tri 38393 42372 38409 42388 se
rect 38409 42372 38486 42388
rect 38393 42306 38486 42372
rect 38393 42204 38486 42270
tri 38393 42188 38409 42204 ne
rect 38409 42188 38486 42204
rect 38226 42089 38374 42171
rect 38114 42056 38191 42072
tri 38191 42056 38207 42072 sw
rect 38114 41990 38207 42056
rect 38243 41931 38357 42089
tri 38393 42056 38409 42072 se
rect 38409 42056 38486 42072
rect 38393 41990 38486 42056
rect 38114 41855 38486 41931
rect 38114 41730 38207 41796
rect 38114 41714 38191 41730
tri 38191 41714 38207 41730 nw
rect 38243 41697 38357 41855
rect 38393 41730 38486 41796
tri 38393 41714 38409 41730 ne
rect 38409 41714 38486 41730
rect 38226 41615 38374 41697
rect 38114 41582 38191 41598
tri 38191 41582 38207 41598 sw
rect 38114 41516 38207 41582
rect 38114 41414 38207 41480
rect 38114 41398 38191 41414
tri 38191 41398 38207 41414 nw
rect 38243 41381 38357 41615
tri 38393 41582 38409 41598 se
rect 38409 41582 38486 41598
rect 38393 41516 38486 41582
rect 38393 41414 38486 41480
tri 38393 41398 38409 41414 ne
rect 38409 41398 38486 41414
rect 38226 41299 38374 41381
rect 38114 41266 38191 41282
tri 38191 41266 38207 41282 sw
rect 38114 41200 38207 41266
rect 38243 41141 38357 41299
tri 38393 41266 38409 41282 se
rect 38409 41266 38486 41282
rect 38393 41200 38486 41266
rect 38114 41065 38486 41141
rect 38114 40940 38207 41006
rect 38114 40924 38191 40940
tri 38191 40924 38207 40940 nw
rect 38243 40907 38357 41065
rect 38393 40940 38486 41006
tri 38393 40924 38409 40940 ne
rect 38409 40924 38486 40940
rect 38226 40825 38374 40907
rect 38114 40792 38191 40808
tri 38191 40792 38207 40808 sw
rect 38114 40726 38207 40792
rect 38114 40624 38207 40690
rect 38114 40608 38191 40624
tri 38191 40608 38207 40624 nw
rect 38243 40591 38357 40825
tri 38393 40792 38409 40808 se
rect 38409 40792 38486 40808
rect 38393 40726 38486 40792
rect 38393 40624 38486 40690
tri 38393 40608 38409 40624 ne
rect 38409 40608 38486 40624
rect 38226 40509 38374 40591
rect 38114 40476 38191 40492
tri 38191 40476 38207 40492 sw
rect 38114 40410 38207 40476
rect 38243 40351 38357 40509
tri 38393 40476 38409 40492 se
rect 38409 40476 38486 40492
rect 38393 40410 38486 40476
rect 38114 40275 38486 40351
rect 38114 40150 38207 40216
rect 38114 40134 38191 40150
tri 38191 40134 38207 40150 nw
rect 38243 40117 38357 40275
rect 38393 40150 38486 40216
tri 38393 40134 38409 40150 ne
rect 38409 40134 38486 40150
rect 38226 40035 38374 40117
rect 38114 40002 38191 40018
tri 38191 40002 38207 40018 sw
rect 38114 39936 38207 40002
rect 38114 39834 38207 39900
rect 38114 39818 38191 39834
tri 38191 39818 38207 39834 nw
rect 38243 39801 38357 40035
tri 38393 40002 38409 40018 se
rect 38409 40002 38486 40018
rect 38393 39936 38486 40002
rect 38393 39834 38486 39900
tri 38393 39818 38409 39834 ne
rect 38409 39818 38486 39834
rect 38226 39719 38374 39801
rect 38114 39686 38191 39702
tri 38191 39686 38207 39702 sw
rect 38114 39620 38207 39686
rect 38243 39561 38357 39719
tri 38393 39686 38409 39702 se
rect 38409 39686 38486 39702
rect 38393 39620 38486 39686
rect 38114 39485 38486 39561
rect 38114 39360 38207 39426
rect 38114 39344 38191 39360
tri 38191 39344 38207 39360 nw
rect 38243 39327 38357 39485
rect 38393 39360 38486 39426
tri 38393 39344 38409 39360 ne
rect 38409 39344 38486 39360
rect 38226 39245 38374 39327
rect 38114 39212 38191 39228
tri 38191 39212 38207 39228 sw
rect 38114 39146 38207 39212
rect 38114 39044 38207 39110
rect 38114 39028 38191 39044
tri 38191 39028 38207 39044 nw
rect 38243 39011 38357 39245
tri 38393 39212 38409 39228 se
rect 38409 39212 38486 39228
rect 38393 39146 38486 39212
rect 38393 39044 38486 39110
tri 38393 39028 38409 39044 ne
rect 38409 39028 38486 39044
rect 38226 38929 38374 39011
rect 38114 38896 38191 38912
tri 38191 38896 38207 38912 sw
rect 38114 38830 38207 38896
rect 38243 38771 38357 38929
tri 38393 38896 38409 38912 se
rect 38409 38896 38486 38912
rect 38393 38830 38486 38896
rect 38114 38695 38486 38771
rect 38114 38570 38207 38636
rect 38114 38554 38191 38570
tri 38191 38554 38207 38570 nw
rect 38243 38537 38357 38695
rect 38393 38570 38486 38636
tri 38393 38554 38409 38570 ne
rect 38409 38554 38486 38570
rect 38226 38455 38374 38537
rect 38114 38422 38191 38438
tri 38191 38422 38207 38438 sw
rect 38114 38356 38207 38422
rect 38114 38254 38207 38320
rect 38114 38238 38191 38254
tri 38191 38238 38207 38254 nw
rect 38243 38221 38357 38455
tri 38393 38422 38409 38438 se
rect 38409 38422 38486 38438
rect 38393 38356 38486 38422
rect 38393 38254 38486 38320
tri 38393 38238 38409 38254 ne
rect 38409 38238 38486 38254
rect 38226 38139 38374 38221
rect 38114 38106 38191 38122
tri 38191 38106 38207 38122 sw
rect 38114 38040 38207 38106
rect 38243 37981 38357 38139
tri 38393 38106 38409 38122 se
rect 38409 38106 38486 38122
rect 38393 38040 38486 38106
rect 38114 37905 38486 37981
rect 38114 37780 38207 37846
rect 38114 37764 38191 37780
tri 38191 37764 38207 37780 nw
rect 38243 37747 38357 37905
rect 38393 37780 38486 37846
tri 38393 37764 38409 37780 ne
rect 38409 37764 38486 37780
rect 38226 37665 38374 37747
rect 38114 37632 38191 37648
tri 38191 37632 38207 37648 sw
rect 38114 37566 38207 37632
rect 38114 37464 38207 37530
rect 38114 37448 38191 37464
tri 38191 37448 38207 37464 nw
rect 38243 37431 38357 37665
tri 38393 37632 38409 37648 se
rect 38409 37632 38486 37648
rect 38393 37566 38486 37632
rect 38393 37464 38486 37530
tri 38393 37448 38409 37464 ne
rect 38409 37448 38486 37464
rect 38226 37349 38374 37431
rect 38114 37316 38191 37332
tri 38191 37316 38207 37332 sw
rect 38114 37250 38207 37316
rect 38243 37191 38357 37349
tri 38393 37316 38409 37332 se
rect 38409 37316 38486 37332
rect 38393 37250 38486 37316
rect 38114 37115 38486 37191
rect 38114 36990 38207 37056
rect 38114 36974 38191 36990
tri 38191 36974 38207 36990 nw
rect 38243 36957 38357 37115
rect 38393 36990 38486 37056
tri 38393 36974 38409 36990 ne
rect 38409 36974 38486 36990
rect 38226 36875 38374 36957
rect 38114 36842 38191 36858
tri 38191 36842 38207 36858 sw
rect 38114 36776 38207 36842
rect 38114 36674 38207 36740
rect 38114 36658 38191 36674
tri 38191 36658 38207 36674 nw
rect 38243 36641 38357 36875
tri 38393 36842 38409 36858 se
rect 38409 36842 38486 36858
rect 38393 36776 38486 36842
rect 38393 36674 38486 36740
tri 38393 36658 38409 36674 ne
rect 38409 36658 38486 36674
rect 38226 36559 38374 36641
rect 38114 36526 38191 36542
tri 38191 36526 38207 36542 sw
rect 38114 36460 38207 36526
rect 38243 36401 38357 36559
tri 38393 36526 38409 36542 se
rect 38409 36526 38486 36542
rect 38393 36460 38486 36526
rect 38114 36325 38486 36401
rect 38114 36200 38207 36266
rect 38114 36184 38191 36200
tri 38191 36184 38207 36200 nw
rect 38243 36167 38357 36325
rect 38393 36200 38486 36266
tri 38393 36184 38409 36200 ne
rect 38409 36184 38486 36200
rect 38226 36085 38374 36167
rect 38114 36052 38191 36068
tri 38191 36052 38207 36068 sw
rect 38114 35986 38207 36052
rect 38114 35884 38207 35950
rect 38114 35868 38191 35884
tri 38191 35868 38207 35884 nw
rect 38243 35851 38357 36085
tri 38393 36052 38409 36068 se
rect 38409 36052 38486 36068
rect 38393 35986 38486 36052
rect 38393 35884 38486 35950
tri 38393 35868 38409 35884 ne
rect 38409 35868 38486 35884
rect 38226 35769 38374 35851
rect 38114 35736 38191 35752
tri 38191 35736 38207 35752 sw
rect 38114 35670 38207 35736
rect 38243 35611 38357 35769
tri 38393 35736 38409 35752 se
rect 38409 35736 38486 35752
rect 38393 35670 38486 35736
rect 38114 35535 38486 35611
rect 38114 35410 38207 35476
rect 38114 35394 38191 35410
tri 38191 35394 38207 35410 nw
rect 38243 35377 38357 35535
rect 38393 35410 38486 35476
tri 38393 35394 38409 35410 ne
rect 38409 35394 38486 35410
rect 38226 35295 38374 35377
rect 38114 35262 38191 35278
tri 38191 35262 38207 35278 sw
rect 38114 35196 38207 35262
rect 38114 35094 38207 35160
rect 38114 35078 38191 35094
tri 38191 35078 38207 35094 nw
rect 38243 35061 38357 35295
tri 38393 35262 38409 35278 se
rect 38409 35262 38486 35278
rect 38393 35196 38486 35262
rect 38393 35094 38486 35160
tri 38393 35078 38409 35094 ne
rect 38409 35078 38486 35094
rect 38226 34979 38374 35061
rect 38114 34946 38191 34962
tri 38191 34946 38207 34962 sw
rect 38114 34880 38207 34946
rect 38243 34821 38357 34979
tri 38393 34946 38409 34962 se
rect 38409 34946 38486 34962
rect 38393 34880 38486 34946
rect 38114 34745 38486 34821
rect 38114 34620 38207 34686
rect 38114 34604 38191 34620
tri 38191 34604 38207 34620 nw
rect 38243 34587 38357 34745
rect 38393 34620 38486 34686
tri 38393 34604 38409 34620 ne
rect 38409 34604 38486 34620
rect 38226 34505 38374 34587
rect 38114 34472 38191 34488
tri 38191 34472 38207 34488 sw
rect 38114 34406 38207 34472
rect 38114 34304 38207 34370
rect 38114 34288 38191 34304
tri 38191 34288 38207 34304 nw
rect 38243 34271 38357 34505
tri 38393 34472 38409 34488 se
rect 38409 34472 38486 34488
rect 38393 34406 38486 34472
rect 38393 34304 38486 34370
tri 38393 34288 38409 34304 ne
rect 38409 34288 38486 34304
rect 38226 34189 38374 34271
rect 38114 34156 38191 34172
tri 38191 34156 38207 34172 sw
rect 38114 34090 38207 34156
rect 38243 34031 38357 34189
tri 38393 34156 38409 34172 se
rect 38409 34156 38486 34172
rect 38393 34090 38486 34156
rect 38114 33955 38486 34031
rect 38114 33830 38207 33896
rect 38114 33814 38191 33830
tri 38191 33814 38207 33830 nw
rect 38243 33797 38357 33955
rect 38393 33830 38486 33896
tri 38393 33814 38409 33830 ne
rect 38409 33814 38486 33830
rect 38226 33715 38374 33797
rect 38114 33682 38191 33698
tri 38191 33682 38207 33698 sw
rect 38114 33616 38207 33682
rect 38114 33514 38207 33580
rect 38114 33498 38191 33514
tri 38191 33498 38207 33514 nw
rect 38243 33481 38357 33715
tri 38393 33682 38409 33698 se
rect 38409 33682 38486 33698
rect 38393 33616 38486 33682
rect 38393 33514 38486 33580
tri 38393 33498 38409 33514 ne
rect 38409 33498 38486 33514
rect 38226 33399 38374 33481
rect 38114 33366 38191 33382
tri 38191 33366 38207 33382 sw
rect 38114 33300 38207 33366
rect 38243 33241 38357 33399
tri 38393 33366 38409 33382 se
rect 38409 33366 38486 33382
rect 38393 33300 38486 33366
rect 38114 33165 38486 33241
rect 38114 33040 38207 33106
rect 38114 33024 38191 33040
tri 38191 33024 38207 33040 nw
rect 38243 33007 38357 33165
rect 38393 33040 38486 33106
tri 38393 33024 38409 33040 ne
rect 38409 33024 38486 33040
rect 38226 32925 38374 33007
rect 38114 32892 38191 32908
tri 38191 32892 38207 32908 sw
rect 38114 32826 38207 32892
rect 38114 32724 38207 32790
rect 38114 32708 38191 32724
tri 38191 32708 38207 32724 nw
rect 38243 32691 38357 32925
tri 38393 32892 38409 32908 se
rect 38409 32892 38486 32908
rect 38393 32826 38486 32892
rect 38393 32724 38486 32790
tri 38393 32708 38409 32724 ne
rect 38409 32708 38486 32724
rect 38226 32609 38374 32691
rect 38114 32576 38191 32592
tri 38191 32576 38207 32592 sw
rect 38114 32510 38207 32576
rect 38243 32451 38357 32609
tri 38393 32576 38409 32592 se
rect 38409 32576 38486 32592
rect 38393 32510 38486 32576
rect 38114 32375 38486 32451
rect 38114 32250 38207 32316
rect 38114 32234 38191 32250
tri 38191 32234 38207 32250 nw
rect 38243 32217 38357 32375
rect 38393 32250 38486 32316
tri 38393 32234 38409 32250 ne
rect 38409 32234 38486 32250
rect 38226 32135 38374 32217
rect 38114 32102 38191 32118
tri 38191 32102 38207 32118 sw
rect 38114 32036 38207 32102
rect 38114 31934 38207 32000
rect 38114 31918 38191 31934
tri 38191 31918 38207 31934 nw
rect 38243 31901 38357 32135
tri 38393 32102 38409 32118 se
rect 38409 32102 38486 32118
rect 38393 32036 38486 32102
rect 38393 31934 38486 32000
tri 38393 31918 38409 31934 ne
rect 38409 31918 38486 31934
rect 38226 31819 38374 31901
rect 38114 31786 38191 31802
tri 38191 31786 38207 31802 sw
rect 38114 31720 38207 31786
rect 38243 31661 38357 31819
tri 38393 31786 38409 31802 se
rect 38409 31786 38486 31802
rect 38393 31720 38486 31786
rect 38114 31585 38486 31661
rect 38114 31460 38207 31526
rect 38114 31444 38191 31460
tri 38191 31444 38207 31460 nw
rect 38243 31427 38357 31585
rect 38393 31460 38486 31526
tri 38393 31444 38409 31460 ne
rect 38409 31444 38486 31460
rect 38226 31345 38374 31427
rect 38114 31312 38191 31328
tri 38191 31312 38207 31328 sw
rect 38114 31246 38207 31312
rect 38114 31144 38207 31210
rect 38114 31128 38191 31144
tri 38191 31128 38207 31144 nw
rect 38243 31111 38357 31345
tri 38393 31312 38409 31328 se
rect 38409 31312 38486 31328
rect 38393 31246 38486 31312
rect 38393 31144 38486 31210
tri 38393 31128 38409 31144 ne
rect 38409 31128 38486 31144
rect 38226 31029 38374 31111
rect 38114 30996 38191 31012
tri 38191 30996 38207 31012 sw
rect 38114 30930 38207 30996
rect 38243 30871 38357 31029
tri 38393 30996 38409 31012 se
rect 38409 30996 38486 31012
rect 38393 30930 38486 30996
rect 38114 30795 38486 30871
rect 38114 30670 38207 30736
rect 38114 30654 38191 30670
tri 38191 30654 38207 30670 nw
rect 38243 30637 38357 30795
rect 38393 30670 38486 30736
tri 38393 30654 38409 30670 ne
rect 38409 30654 38486 30670
rect 38226 30555 38374 30637
rect 38114 30522 38191 30538
tri 38191 30522 38207 30538 sw
rect 38114 30456 38207 30522
rect 38114 30354 38207 30420
rect 38114 30338 38191 30354
tri 38191 30338 38207 30354 nw
rect 38243 30321 38357 30555
tri 38393 30522 38409 30538 se
rect 38409 30522 38486 30538
rect 38393 30456 38486 30522
rect 38393 30354 38486 30420
tri 38393 30338 38409 30354 ne
rect 38409 30338 38486 30354
rect 38226 30239 38374 30321
rect 38114 30206 38191 30222
tri 38191 30206 38207 30222 sw
rect 38114 30140 38207 30206
rect 38243 30081 38357 30239
tri 38393 30206 38409 30222 se
rect 38409 30206 38486 30222
rect 38393 30140 38486 30206
rect 38114 30005 38486 30081
rect 38114 29880 38207 29946
rect 38114 29864 38191 29880
tri 38191 29864 38207 29880 nw
rect 38243 29847 38357 30005
rect 38393 29880 38486 29946
tri 38393 29864 38409 29880 ne
rect 38409 29864 38486 29880
rect 38226 29765 38374 29847
rect 38114 29732 38191 29748
tri 38191 29732 38207 29748 sw
rect 38114 29666 38207 29732
rect 38114 29564 38207 29630
rect 38114 29548 38191 29564
tri 38191 29548 38207 29564 nw
rect 38243 29531 38357 29765
tri 38393 29732 38409 29748 se
rect 38409 29732 38486 29748
rect 38393 29666 38486 29732
rect 38393 29564 38486 29630
tri 38393 29548 38409 29564 ne
rect 38409 29548 38486 29564
rect 38226 29449 38374 29531
rect 38114 29416 38191 29432
tri 38191 29416 38207 29432 sw
rect 38114 29350 38207 29416
rect 38243 29291 38357 29449
tri 38393 29416 38409 29432 se
rect 38409 29416 38486 29432
rect 38393 29350 38486 29416
rect 38114 29215 38486 29291
rect 38114 29090 38207 29156
rect 38114 29074 38191 29090
tri 38191 29074 38207 29090 nw
rect 38243 29057 38357 29215
rect 38393 29090 38486 29156
tri 38393 29074 38409 29090 ne
rect 38409 29074 38486 29090
rect 38226 28975 38374 29057
rect 38114 28942 38191 28958
tri 38191 28942 38207 28958 sw
rect 38114 28876 38207 28942
rect 38243 28833 38357 28975
tri 38393 28942 38409 28958 se
rect 38409 28942 38486 28958
rect 38393 28876 38486 28942
rect 38522 28463 38558 80603
rect 38594 28463 38630 80603
rect 38666 80445 38702 80603
rect 38658 80303 38710 80445
rect 38666 28763 38702 80303
rect 38658 28621 38710 28763
rect 38666 28463 38702 28621
rect 38738 28463 38774 80603
rect 38810 28463 38846 80603
rect 38882 28833 38966 80233
rect 39002 28463 39038 80603
rect 39074 28463 39110 80603
rect 39146 80445 39182 80603
rect 39138 80303 39190 80445
rect 39146 28763 39182 80303
rect 39138 28621 39190 28763
rect 39146 28463 39182 28621
rect 39218 28463 39254 80603
rect 39290 28463 39326 80603
rect 39362 80124 39455 80190
rect 39362 80108 39439 80124
tri 39439 80108 39455 80124 nw
rect 39491 80091 39605 80233
rect 39641 80124 39734 80190
tri 39641 80108 39657 80124 ne
rect 39657 80108 39734 80124
rect 39474 80009 39622 80091
rect 39362 79976 39439 79992
tri 39439 79976 39455 79992 sw
rect 39362 79910 39455 79976
rect 39491 79851 39605 80009
tri 39641 79976 39657 79992 se
rect 39657 79976 39734 79992
rect 39641 79910 39734 79976
rect 39362 79775 39734 79851
rect 39362 79650 39455 79716
rect 39362 79634 39439 79650
tri 39439 79634 39455 79650 nw
rect 39491 79617 39605 79775
rect 39641 79650 39734 79716
tri 39641 79634 39657 79650 ne
rect 39657 79634 39734 79650
rect 39474 79535 39622 79617
rect 39362 79502 39439 79518
tri 39439 79502 39455 79518 sw
rect 39362 79436 39455 79502
rect 39362 79334 39455 79400
rect 39362 79318 39439 79334
tri 39439 79318 39455 79334 nw
rect 39491 79301 39605 79535
tri 39641 79502 39657 79518 se
rect 39657 79502 39734 79518
rect 39641 79436 39734 79502
rect 39641 79334 39734 79400
tri 39641 79318 39657 79334 ne
rect 39657 79318 39734 79334
rect 39474 79219 39622 79301
rect 39362 79186 39439 79202
tri 39439 79186 39455 79202 sw
rect 39362 79120 39455 79186
rect 39491 79061 39605 79219
tri 39641 79186 39657 79202 se
rect 39657 79186 39734 79202
rect 39641 79120 39734 79186
rect 39362 78985 39734 79061
rect 39362 78860 39455 78926
rect 39362 78844 39439 78860
tri 39439 78844 39455 78860 nw
rect 39491 78827 39605 78985
rect 39641 78860 39734 78926
tri 39641 78844 39657 78860 ne
rect 39657 78844 39734 78860
rect 39474 78745 39622 78827
rect 39362 78712 39439 78728
tri 39439 78712 39455 78728 sw
rect 39362 78646 39455 78712
rect 39362 78544 39455 78610
rect 39362 78528 39439 78544
tri 39439 78528 39455 78544 nw
rect 39491 78511 39605 78745
tri 39641 78712 39657 78728 se
rect 39657 78712 39734 78728
rect 39641 78646 39734 78712
rect 39641 78544 39734 78610
tri 39641 78528 39657 78544 ne
rect 39657 78528 39734 78544
rect 39474 78429 39622 78511
rect 39362 78396 39439 78412
tri 39439 78396 39455 78412 sw
rect 39362 78330 39455 78396
rect 39491 78271 39605 78429
tri 39641 78396 39657 78412 se
rect 39657 78396 39734 78412
rect 39641 78330 39734 78396
rect 39362 78195 39734 78271
rect 39362 78070 39455 78136
rect 39362 78054 39439 78070
tri 39439 78054 39455 78070 nw
rect 39491 78037 39605 78195
rect 39641 78070 39734 78136
tri 39641 78054 39657 78070 ne
rect 39657 78054 39734 78070
rect 39474 77955 39622 78037
rect 39362 77922 39439 77938
tri 39439 77922 39455 77938 sw
rect 39362 77856 39455 77922
rect 39362 77754 39455 77820
rect 39362 77738 39439 77754
tri 39439 77738 39455 77754 nw
rect 39491 77721 39605 77955
tri 39641 77922 39657 77938 se
rect 39657 77922 39734 77938
rect 39641 77856 39734 77922
rect 39641 77754 39734 77820
tri 39641 77738 39657 77754 ne
rect 39657 77738 39734 77754
rect 39474 77639 39622 77721
rect 39362 77606 39439 77622
tri 39439 77606 39455 77622 sw
rect 39362 77540 39455 77606
rect 39491 77481 39605 77639
tri 39641 77606 39657 77622 se
rect 39657 77606 39734 77622
rect 39641 77540 39734 77606
rect 39362 77405 39734 77481
rect 39362 77280 39455 77346
rect 39362 77264 39439 77280
tri 39439 77264 39455 77280 nw
rect 39491 77247 39605 77405
rect 39641 77280 39734 77346
tri 39641 77264 39657 77280 ne
rect 39657 77264 39734 77280
rect 39474 77165 39622 77247
rect 39362 77132 39439 77148
tri 39439 77132 39455 77148 sw
rect 39362 77066 39455 77132
rect 39362 76964 39455 77030
rect 39362 76948 39439 76964
tri 39439 76948 39455 76964 nw
rect 39491 76931 39605 77165
tri 39641 77132 39657 77148 se
rect 39657 77132 39734 77148
rect 39641 77066 39734 77132
rect 39641 76964 39734 77030
tri 39641 76948 39657 76964 ne
rect 39657 76948 39734 76964
rect 39474 76849 39622 76931
rect 39362 76816 39439 76832
tri 39439 76816 39455 76832 sw
rect 39362 76750 39455 76816
rect 39491 76691 39605 76849
tri 39641 76816 39657 76832 se
rect 39657 76816 39734 76832
rect 39641 76750 39734 76816
rect 39362 76615 39734 76691
rect 39362 76490 39455 76556
rect 39362 76474 39439 76490
tri 39439 76474 39455 76490 nw
rect 39491 76457 39605 76615
rect 39641 76490 39734 76556
tri 39641 76474 39657 76490 ne
rect 39657 76474 39734 76490
rect 39474 76375 39622 76457
rect 39362 76342 39439 76358
tri 39439 76342 39455 76358 sw
rect 39362 76276 39455 76342
rect 39362 76174 39455 76240
rect 39362 76158 39439 76174
tri 39439 76158 39455 76174 nw
rect 39491 76141 39605 76375
tri 39641 76342 39657 76358 se
rect 39657 76342 39734 76358
rect 39641 76276 39734 76342
rect 39641 76174 39734 76240
tri 39641 76158 39657 76174 ne
rect 39657 76158 39734 76174
rect 39474 76059 39622 76141
rect 39362 76026 39439 76042
tri 39439 76026 39455 76042 sw
rect 39362 75960 39455 76026
rect 39491 75901 39605 76059
tri 39641 76026 39657 76042 se
rect 39657 76026 39734 76042
rect 39641 75960 39734 76026
rect 39362 75825 39734 75901
rect 39362 75700 39455 75766
rect 39362 75684 39439 75700
tri 39439 75684 39455 75700 nw
rect 39491 75667 39605 75825
rect 39641 75700 39734 75766
tri 39641 75684 39657 75700 ne
rect 39657 75684 39734 75700
rect 39474 75585 39622 75667
rect 39362 75552 39439 75568
tri 39439 75552 39455 75568 sw
rect 39362 75486 39455 75552
rect 39362 75384 39455 75450
rect 39362 75368 39439 75384
tri 39439 75368 39455 75384 nw
rect 39491 75351 39605 75585
tri 39641 75552 39657 75568 se
rect 39657 75552 39734 75568
rect 39641 75486 39734 75552
rect 39641 75384 39734 75450
tri 39641 75368 39657 75384 ne
rect 39657 75368 39734 75384
rect 39474 75269 39622 75351
rect 39362 75236 39439 75252
tri 39439 75236 39455 75252 sw
rect 39362 75170 39455 75236
rect 39491 75111 39605 75269
tri 39641 75236 39657 75252 se
rect 39657 75236 39734 75252
rect 39641 75170 39734 75236
rect 39362 75035 39734 75111
rect 39362 74910 39455 74976
rect 39362 74894 39439 74910
tri 39439 74894 39455 74910 nw
rect 39491 74877 39605 75035
rect 39641 74910 39734 74976
tri 39641 74894 39657 74910 ne
rect 39657 74894 39734 74910
rect 39474 74795 39622 74877
rect 39362 74762 39439 74778
tri 39439 74762 39455 74778 sw
rect 39362 74696 39455 74762
rect 39362 74594 39455 74660
rect 39362 74578 39439 74594
tri 39439 74578 39455 74594 nw
rect 39491 74561 39605 74795
tri 39641 74762 39657 74778 se
rect 39657 74762 39734 74778
rect 39641 74696 39734 74762
rect 39641 74594 39734 74660
tri 39641 74578 39657 74594 ne
rect 39657 74578 39734 74594
rect 39474 74479 39622 74561
rect 39362 74446 39439 74462
tri 39439 74446 39455 74462 sw
rect 39362 74380 39455 74446
rect 39491 74321 39605 74479
tri 39641 74446 39657 74462 se
rect 39657 74446 39734 74462
rect 39641 74380 39734 74446
rect 39362 74245 39734 74321
rect 39362 74120 39455 74186
rect 39362 74104 39439 74120
tri 39439 74104 39455 74120 nw
rect 39491 74087 39605 74245
rect 39641 74120 39734 74186
tri 39641 74104 39657 74120 ne
rect 39657 74104 39734 74120
rect 39474 74005 39622 74087
rect 39362 73972 39439 73988
tri 39439 73972 39455 73988 sw
rect 39362 73906 39455 73972
rect 39362 73804 39455 73870
rect 39362 73788 39439 73804
tri 39439 73788 39455 73804 nw
rect 39491 73771 39605 74005
tri 39641 73972 39657 73988 se
rect 39657 73972 39734 73988
rect 39641 73906 39734 73972
rect 39641 73804 39734 73870
tri 39641 73788 39657 73804 ne
rect 39657 73788 39734 73804
rect 39474 73689 39622 73771
rect 39362 73656 39439 73672
tri 39439 73656 39455 73672 sw
rect 39362 73590 39455 73656
rect 39491 73531 39605 73689
tri 39641 73656 39657 73672 se
rect 39657 73656 39734 73672
rect 39641 73590 39734 73656
rect 39362 73455 39734 73531
rect 39362 73330 39455 73396
rect 39362 73314 39439 73330
tri 39439 73314 39455 73330 nw
rect 39491 73297 39605 73455
rect 39641 73330 39734 73396
tri 39641 73314 39657 73330 ne
rect 39657 73314 39734 73330
rect 39474 73215 39622 73297
rect 39362 73182 39439 73198
tri 39439 73182 39455 73198 sw
rect 39362 73116 39455 73182
rect 39362 73014 39455 73080
rect 39362 72998 39439 73014
tri 39439 72998 39455 73014 nw
rect 39491 72981 39605 73215
tri 39641 73182 39657 73198 se
rect 39657 73182 39734 73198
rect 39641 73116 39734 73182
rect 39641 73014 39734 73080
tri 39641 72998 39657 73014 ne
rect 39657 72998 39734 73014
rect 39474 72899 39622 72981
rect 39362 72866 39439 72882
tri 39439 72866 39455 72882 sw
rect 39362 72800 39455 72866
rect 39491 72741 39605 72899
tri 39641 72866 39657 72882 se
rect 39657 72866 39734 72882
rect 39641 72800 39734 72866
rect 39362 72665 39734 72741
rect 39362 72540 39455 72606
rect 39362 72524 39439 72540
tri 39439 72524 39455 72540 nw
rect 39491 72507 39605 72665
rect 39641 72540 39734 72606
tri 39641 72524 39657 72540 ne
rect 39657 72524 39734 72540
rect 39474 72425 39622 72507
rect 39362 72392 39439 72408
tri 39439 72392 39455 72408 sw
rect 39362 72326 39455 72392
rect 39362 72224 39455 72290
rect 39362 72208 39439 72224
tri 39439 72208 39455 72224 nw
rect 39491 72191 39605 72425
tri 39641 72392 39657 72408 se
rect 39657 72392 39734 72408
rect 39641 72326 39734 72392
rect 39641 72224 39734 72290
tri 39641 72208 39657 72224 ne
rect 39657 72208 39734 72224
rect 39474 72109 39622 72191
rect 39362 72076 39439 72092
tri 39439 72076 39455 72092 sw
rect 39362 72010 39455 72076
rect 39491 71951 39605 72109
tri 39641 72076 39657 72092 se
rect 39657 72076 39734 72092
rect 39641 72010 39734 72076
rect 39362 71875 39734 71951
rect 39362 71750 39455 71816
rect 39362 71734 39439 71750
tri 39439 71734 39455 71750 nw
rect 39491 71717 39605 71875
rect 39641 71750 39734 71816
tri 39641 71734 39657 71750 ne
rect 39657 71734 39734 71750
rect 39474 71635 39622 71717
rect 39362 71602 39439 71618
tri 39439 71602 39455 71618 sw
rect 39362 71536 39455 71602
rect 39362 71434 39455 71500
rect 39362 71418 39439 71434
tri 39439 71418 39455 71434 nw
rect 39491 71401 39605 71635
tri 39641 71602 39657 71618 se
rect 39657 71602 39734 71618
rect 39641 71536 39734 71602
rect 39641 71434 39734 71500
tri 39641 71418 39657 71434 ne
rect 39657 71418 39734 71434
rect 39474 71319 39622 71401
rect 39362 71286 39439 71302
tri 39439 71286 39455 71302 sw
rect 39362 71220 39455 71286
rect 39491 71161 39605 71319
tri 39641 71286 39657 71302 se
rect 39657 71286 39734 71302
rect 39641 71220 39734 71286
rect 39362 71085 39734 71161
rect 39362 70960 39455 71026
rect 39362 70944 39439 70960
tri 39439 70944 39455 70960 nw
rect 39491 70927 39605 71085
rect 39641 70960 39734 71026
tri 39641 70944 39657 70960 ne
rect 39657 70944 39734 70960
rect 39474 70845 39622 70927
rect 39362 70812 39439 70828
tri 39439 70812 39455 70828 sw
rect 39362 70746 39455 70812
rect 39362 70644 39455 70710
rect 39362 70628 39439 70644
tri 39439 70628 39455 70644 nw
rect 39491 70611 39605 70845
tri 39641 70812 39657 70828 se
rect 39657 70812 39734 70828
rect 39641 70746 39734 70812
rect 39641 70644 39734 70710
tri 39641 70628 39657 70644 ne
rect 39657 70628 39734 70644
rect 39474 70529 39622 70611
rect 39362 70496 39439 70512
tri 39439 70496 39455 70512 sw
rect 39362 70430 39455 70496
rect 39491 70371 39605 70529
tri 39641 70496 39657 70512 se
rect 39657 70496 39734 70512
rect 39641 70430 39734 70496
rect 39362 70295 39734 70371
rect 39362 70170 39455 70236
rect 39362 70154 39439 70170
tri 39439 70154 39455 70170 nw
rect 39491 70137 39605 70295
rect 39641 70170 39734 70236
tri 39641 70154 39657 70170 ne
rect 39657 70154 39734 70170
rect 39474 70055 39622 70137
rect 39362 70022 39439 70038
tri 39439 70022 39455 70038 sw
rect 39362 69956 39455 70022
rect 39362 69854 39455 69920
rect 39362 69838 39439 69854
tri 39439 69838 39455 69854 nw
rect 39491 69821 39605 70055
tri 39641 70022 39657 70038 se
rect 39657 70022 39734 70038
rect 39641 69956 39734 70022
rect 39641 69854 39734 69920
tri 39641 69838 39657 69854 ne
rect 39657 69838 39734 69854
rect 39474 69739 39622 69821
rect 39362 69706 39439 69722
tri 39439 69706 39455 69722 sw
rect 39362 69640 39455 69706
rect 39491 69581 39605 69739
tri 39641 69706 39657 69722 se
rect 39657 69706 39734 69722
rect 39641 69640 39734 69706
rect 39362 69505 39734 69581
rect 39362 69380 39455 69446
rect 39362 69364 39439 69380
tri 39439 69364 39455 69380 nw
rect 39491 69347 39605 69505
rect 39641 69380 39734 69446
tri 39641 69364 39657 69380 ne
rect 39657 69364 39734 69380
rect 39474 69265 39622 69347
rect 39362 69232 39439 69248
tri 39439 69232 39455 69248 sw
rect 39362 69166 39455 69232
rect 39362 69064 39455 69130
rect 39362 69048 39439 69064
tri 39439 69048 39455 69064 nw
rect 39491 69031 39605 69265
tri 39641 69232 39657 69248 se
rect 39657 69232 39734 69248
rect 39641 69166 39734 69232
rect 39641 69064 39734 69130
tri 39641 69048 39657 69064 ne
rect 39657 69048 39734 69064
rect 39474 68949 39622 69031
rect 39362 68916 39439 68932
tri 39439 68916 39455 68932 sw
rect 39362 68850 39455 68916
rect 39491 68791 39605 68949
tri 39641 68916 39657 68932 se
rect 39657 68916 39734 68932
rect 39641 68850 39734 68916
rect 39362 68715 39734 68791
rect 39362 68590 39455 68656
rect 39362 68574 39439 68590
tri 39439 68574 39455 68590 nw
rect 39491 68557 39605 68715
rect 39641 68590 39734 68656
tri 39641 68574 39657 68590 ne
rect 39657 68574 39734 68590
rect 39474 68475 39622 68557
rect 39362 68442 39439 68458
tri 39439 68442 39455 68458 sw
rect 39362 68376 39455 68442
rect 39362 68274 39455 68340
rect 39362 68258 39439 68274
tri 39439 68258 39455 68274 nw
rect 39491 68241 39605 68475
tri 39641 68442 39657 68458 se
rect 39657 68442 39734 68458
rect 39641 68376 39734 68442
rect 39641 68274 39734 68340
tri 39641 68258 39657 68274 ne
rect 39657 68258 39734 68274
rect 39474 68159 39622 68241
rect 39362 68126 39439 68142
tri 39439 68126 39455 68142 sw
rect 39362 68060 39455 68126
rect 39491 68001 39605 68159
tri 39641 68126 39657 68142 se
rect 39657 68126 39734 68142
rect 39641 68060 39734 68126
rect 39362 67925 39734 68001
rect 39362 67800 39455 67866
rect 39362 67784 39439 67800
tri 39439 67784 39455 67800 nw
rect 39491 67767 39605 67925
rect 39641 67800 39734 67866
tri 39641 67784 39657 67800 ne
rect 39657 67784 39734 67800
rect 39474 67685 39622 67767
rect 39362 67652 39439 67668
tri 39439 67652 39455 67668 sw
rect 39362 67586 39455 67652
rect 39362 67484 39455 67550
rect 39362 67468 39439 67484
tri 39439 67468 39455 67484 nw
rect 39491 67451 39605 67685
tri 39641 67652 39657 67668 se
rect 39657 67652 39734 67668
rect 39641 67586 39734 67652
rect 39641 67484 39734 67550
tri 39641 67468 39657 67484 ne
rect 39657 67468 39734 67484
rect 39474 67369 39622 67451
rect 39362 67336 39439 67352
tri 39439 67336 39455 67352 sw
rect 39362 67270 39455 67336
rect 39491 67211 39605 67369
tri 39641 67336 39657 67352 se
rect 39657 67336 39734 67352
rect 39641 67270 39734 67336
rect 39362 67135 39734 67211
rect 39362 67010 39455 67076
rect 39362 66994 39439 67010
tri 39439 66994 39455 67010 nw
rect 39491 66977 39605 67135
rect 39641 67010 39734 67076
tri 39641 66994 39657 67010 ne
rect 39657 66994 39734 67010
rect 39474 66895 39622 66977
rect 39362 66862 39439 66878
tri 39439 66862 39455 66878 sw
rect 39362 66796 39455 66862
rect 39362 66694 39455 66760
rect 39362 66678 39439 66694
tri 39439 66678 39455 66694 nw
rect 39491 66661 39605 66895
tri 39641 66862 39657 66878 se
rect 39657 66862 39734 66878
rect 39641 66796 39734 66862
rect 39641 66694 39734 66760
tri 39641 66678 39657 66694 ne
rect 39657 66678 39734 66694
rect 39474 66579 39622 66661
rect 39362 66546 39439 66562
tri 39439 66546 39455 66562 sw
rect 39362 66480 39455 66546
rect 39491 66421 39605 66579
tri 39641 66546 39657 66562 se
rect 39657 66546 39734 66562
rect 39641 66480 39734 66546
rect 39362 66345 39734 66421
rect 39362 66220 39455 66286
rect 39362 66204 39439 66220
tri 39439 66204 39455 66220 nw
rect 39491 66187 39605 66345
rect 39641 66220 39734 66286
tri 39641 66204 39657 66220 ne
rect 39657 66204 39734 66220
rect 39474 66105 39622 66187
rect 39362 66072 39439 66088
tri 39439 66072 39455 66088 sw
rect 39362 66006 39455 66072
rect 39362 65904 39455 65970
rect 39362 65888 39439 65904
tri 39439 65888 39455 65904 nw
rect 39491 65871 39605 66105
tri 39641 66072 39657 66088 se
rect 39657 66072 39734 66088
rect 39641 66006 39734 66072
rect 39641 65904 39734 65970
tri 39641 65888 39657 65904 ne
rect 39657 65888 39734 65904
rect 39474 65789 39622 65871
rect 39362 65756 39439 65772
tri 39439 65756 39455 65772 sw
rect 39362 65690 39455 65756
rect 39491 65631 39605 65789
tri 39641 65756 39657 65772 se
rect 39657 65756 39734 65772
rect 39641 65690 39734 65756
rect 39362 65555 39734 65631
rect 39362 65430 39455 65496
rect 39362 65414 39439 65430
tri 39439 65414 39455 65430 nw
rect 39491 65397 39605 65555
rect 39641 65430 39734 65496
tri 39641 65414 39657 65430 ne
rect 39657 65414 39734 65430
rect 39474 65315 39622 65397
rect 39362 65282 39439 65298
tri 39439 65282 39455 65298 sw
rect 39362 65216 39455 65282
rect 39362 65114 39455 65180
rect 39362 65098 39439 65114
tri 39439 65098 39455 65114 nw
rect 39491 65081 39605 65315
tri 39641 65282 39657 65298 se
rect 39657 65282 39734 65298
rect 39641 65216 39734 65282
rect 39641 65114 39734 65180
tri 39641 65098 39657 65114 ne
rect 39657 65098 39734 65114
rect 39474 64999 39622 65081
rect 39362 64966 39439 64982
tri 39439 64966 39455 64982 sw
rect 39362 64900 39455 64966
rect 39491 64841 39605 64999
tri 39641 64966 39657 64982 se
rect 39657 64966 39734 64982
rect 39641 64900 39734 64966
rect 39362 64765 39734 64841
rect 39362 64640 39455 64706
rect 39362 64624 39439 64640
tri 39439 64624 39455 64640 nw
rect 39491 64607 39605 64765
rect 39641 64640 39734 64706
tri 39641 64624 39657 64640 ne
rect 39657 64624 39734 64640
rect 39474 64525 39622 64607
rect 39362 64492 39439 64508
tri 39439 64492 39455 64508 sw
rect 39362 64426 39455 64492
rect 39362 64324 39455 64390
rect 39362 64308 39439 64324
tri 39439 64308 39455 64324 nw
rect 39491 64291 39605 64525
tri 39641 64492 39657 64508 se
rect 39657 64492 39734 64508
rect 39641 64426 39734 64492
rect 39641 64324 39734 64390
tri 39641 64308 39657 64324 ne
rect 39657 64308 39734 64324
rect 39474 64209 39622 64291
rect 39362 64176 39439 64192
tri 39439 64176 39455 64192 sw
rect 39362 64110 39455 64176
rect 39491 64051 39605 64209
tri 39641 64176 39657 64192 se
rect 39657 64176 39734 64192
rect 39641 64110 39734 64176
rect 39362 63975 39734 64051
rect 39362 63850 39455 63916
rect 39362 63834 39439 63850
tri 39439 63834 39455 63850 nw
rect 39491 63817 39605 63975
rect 39641 63850 39734 63916
tri 39641 63834 39657 63850 ne
rect 39657 63834 39734 63850
rect 39474 63735 39622 63817
rect 39362 63702 39439 63718
tri 39439 63702 39455 63718 sw
rect 39362 63636 39455 63702
rect 39362 63534 39455 63600
rect 39362 63518 39439 63534
tri 39439 63518 39455 63534 nw
rect 39491 63501 39605 63735
tri 39641 63702 39657 63718 se
rect 39657 63702 39734 63718
rect 39641 63636 39734 63702
rect 39641 63534 39734 63600
tri 39641 63518 39657 63534 ne
rect 39657 63518 39734 63534
rect 39474 63419 39622 63501
rect 39362 63386 39439 63402
tri 39439 63386 39455 63402 sw
rect 39362 63320 39455 63386
rect 39491 63261 39605 63419
tri 39641 63386 39657 63402 se
rect 39657 63386 39734 63402
rect 39641 63320 39734 63386
rect 39362 63185 39734 63261
rect 39362 63060 39455 63126
rect 39362 63044 39439 63060
tri 39439 63044 39455 63060 nw
rect 39491 63027 39605 63185
rect 39641 63060 39734 63126
tri 39641 63044 39657 63060 ne
rect 39657 63044 39734 63060
rect 39474 62945 39622 63027
rect 39362 62912 39439 62928
tri 39439 62912 39455 62928 sw
rect 39362 62846 39455 62912
rect 39362 62744 39455 62810
rect 39362 62728 39439 62744
tri 39439 62728 39455 62744 nw
rect 39491 62711 39605 62945
tri 39641 62912 39657 62928 se
rect 39657 62912 39734 62928
rect 39641 62846 39734 62912
rect 39641 62744 39734 62810
tri 39641 62728 39657 62744 ne
rect 39657 62728 39734 62744
rect 39474 62629 39622 62711
rect 39362 62596 39439 62612
tri 39439 62596 39455 62612 sw
rect 39362 62530 39455 62596
rect 39491 62471 39605 62629
tri 39641 62596 39657 62612 se
rect 39657 62596 39734 62612
rect 39641 62530 39734 62596
rect 39362 62395 39734 62471
rect 39362 62270 39455 62336
rect 39362 62254 39439 62270
tri 39439 62254 39455 62270 nw
rect 39491 62237 39605 62395
rect 39641 62270 39734 62336
tri 39641 62254 39657 62270 ne
rect 39657 62254 39734 62270
rect 39474 62155 39622 62237
rect 39362 62122 39439 62138
tri 39439 62122 39455 62138 sw
rect 39362 62056 39455 62122
rect 39362 61954 39455 62020
rect 39362 61938 39439 61954
tri 39439 61938 39455 61954 nw
rect 39491 61921 39605 62155
tri 39641 62122 39657 62138 se
rect 39657 62122 39734 62138
rect 39641 62056 39734 62122
rect 39641 61954 39734 62020
tri 39641 61938 39657 61954 ne
rect 39657 61938 39734 61954
rect 39474 61839 39622 61921
rect 39362 61806 39439 61822
tri 39439 61806 39455 61822 sw
rect 39362 61740 39455 61806
rect 39491 61681 39605 61839
tri 39641 61806 39657 61822 se
rect 39657 61806 39734 61822
rect 39641 61740 39734 61806
rect 39362 61605 39734 61681
rect 39362 61480 39455 61546
rect 39362 61464 39439 61480
tri 39439 61464 39455 61480 nw
rect 39491 61447 39605 61605
rect 39641 61480 39734 61546
tri 39641 61464 39657 61480 ne
rect 39657 61464 39734 61480
rect 39474 61365 39622 61447
rect 39362 61332 39439 61348
tri 39439 61332 39455 61348 sw
rect 39362 61266 39455 61332
rect 39362 61164 39455 61230
rect 39362 61148 39439 61164
tri 39439 61148 39455 61164 nw
rect 39491 61131 39605 61365
tri 39641 61332 39657 61348 se
rect 39657 61332 39734 61348
rect 39641 61266 39734 61332
rect 39641 61164 39734 61230
tri 39641 61148 39657 61164 ne
rect 39657 61148 39734 61164
rect 39474 61049 39622 61131
rect 39362 61016 39439 61032
tri 39439 61016 39455 61032 sw
rect 39362 60950 39455 61016
rect 39491 60891 39605 61049
tri 39641 61016 39657 61032 se
rect 39657 61016 39734 61032
rect 39641 60950 39734 61016
rect 39362 60815 39734 60891
rect 39362 60690 39455 60756
rect 39362 60674 39439 60690
tri 39439 60674 39455 60690 nw
rect 39491 60657 39605 60815
rect 39641 60690 39734 60756
tri 39641 60674 39657 60690 ne
rect 39657 60674 39734 60690
rect 39474 60575 39622 60657
rect 39362 60542 39439 60558
tri 39439 60542 39455 60558 sw
rect 39362 60476 39455 60542
rect 39362 60374 39455 60440
rect 39362 60358 39439 60374
tri 39439 60358 39455 60374 nw
rect 39491 60341 39605 60575
tri 39641 60542 39657 60558 se
rect 39657 60542 39734 60558
rect 39641 60476 39734 60542
rect 39641 60374 39734 60440
tri 39641 60358 39657 60374 ne
rect 39657 60358 39734 60374
rect 39474 60259 39622 60341
rect 39362 60226 39439 60242
tri 39439 60226 39455 60242 sw
rect 39362 60160 39455 60226
rect 39491 60101 39605 60259
tri 39641 60226 39657 60242 se
rect 39657 60226 39734 60242
rect 39641 60160 39734 60226
rect 39362 60025 39734 60101
rect 39362 59900 39455 59966
rect 39362 59884 39439 59900
tri 39439 59884 39455 59900 nw
rect 39491 59867 39605 60025
rect 39641 59900 39734 59966
tri 39641 59884 39657 59900 ne
rect 39657 59884 39734 59900
rect 39474 59785 39622 59867
rect 39362 59752 39439 59768
tri 39439 59752 39455 59768 sw
rect 39362 59686 39455 59752
rect 39362 59584 39455 59650
rect 39362 59568 39439 59584
tri 39439 59568 39455 59584 nw
rect 39491 59551 39605 59785
tri 39641 59752 39657 59768 se
rect 39657 59752 39734 59768
rect 39641 59686 39734 59752
rect 39641 59584 39734 59650
tri 39641 59568 39657 59584 ne
rect 39657 59568 39734 59584
rect 39474 59469 39622 59551
rect 39362 59436 39439 59452
tri 39439 59436 39455 59452 sw
rect 39362 59370 39455 59436
rect 39491 59311 39605 59469
tri 39641 59436 39657 59452 se
rect 39657 59436 39734 59452
rect 39641 59370 39734 59436
rect 39362 59235 39734 59311
rect 39362 59110 39455 59176
rect 39362 59094 39439 59110
tri 39439 59094 39455 59110 nw
rect 39491 59077 39605 59235
rect 39641 59110 39734 59176
tri 39641 59094 39657 59110 ne
rect 39657 59094 39734 59110
rect 39474 58995 39622 59077
rect 39362 58962 39439 58978
tri 39439 58962 39455 58978 sw
rect 39362 58896 39455 58962
rect 39362 58794 39455 58860
rect 39362 58778 39439 58794
tri 39439 58778 39455 58794 nw
rect 39491 58761 39605 58995
tri 39641 58962 39657 58978 se
rect 39657 58962 39734 58978
rect 39641 58896 39734 58962
rect 39641 58794 39734 58860
tri 39641 58778 39657 58794 ne
rect 39657 58778 39734 58794
rect 39474 58679 39622 58761
rect 39362 58646 39439 58662
tri 39439 58646 39455 58662 sw
rect 39362 58580 39455 58646
rect 39491 58521 39605 58679
tri 39641 58646 39657 58662 se
rect 39657 58646 39734 58662
rect 39641 58580 39734 58646
rect 39362 58445 39734 58521
rect 39362 58320 39455 58386
rect 39362 58304 39439 58320
tri 39439 58304 39455 58320 nw
rect 39491 58287 39605 58445
rect 39641 58320 39734 58386
tri 39641 58304 39657 58320 ne
rect 39657 58304 39734 58320
rect 39474 58205 39622 58287
rect 39362 58172 39439 58188
tri 39439 58172 39455 58188 sw
rect 39362 58106 39455 58172
rect 39362 58004 39455 58070
rect 39362 57988 39439 58004
tri 39439 57988 39455 58004 nw
rect 39491 57971 39605 58205
tri 39641 58172 39657 58188 se
rect 39657 58172 39734 58188
rect 39641 58106 39734 58172
rect 39641 58004 39734 58070
tri 39641 57988 39657 58004 ne
rect 39657 57988 39734 58004
rect 39474 57889 39622 57971
rect 39362 57856 39439 57872
tri 39439 57856 39455 57872 sw
rect 39362 57790 39455 57856
rect 39491 57731 39605 57889
tri 39641 57856 39657 57872 se
rect 39657 57856 39734 57872
rect 39641 57790 39734 57856
rect 39362 57655 39734 57731
rect 39362 57530 39455 57596
rect 39362 57514 39439 57530
tri 39439 57514 39455 57530 nw
rect 39491 57497 39605 57655
rect 39641 57530 39734 57596
tri 39641 57514 39657 57530 ne
rect 39657 57514 39734 57530
rect 39474 57415 39622 57497
rect 39362 57382 39439 57398
tri 39439 57382 39455 57398 sw
rect 39362 57316 39455 57382
rect 39362 57214 39455 57280
rect 39362 57198 39439 57214
tri 39439 57198 39455 57214 nw
rect 39491 57181 39605 57415
tri 39641 57382 39657 57398 se
rect 39657 57382 39734 57398
rect 39641 57316 39734 57382
rect 39641 57214 39734 57280
tri 39641 57198 39657 57214 ne
rect 39657 57198 39734 57214
rect 39474 57099 39622 57181
rect 39362 57066 39439 57082
tri 39439 57066 39455 57082 sw
rect 39362 57000 39455 57066
rect 39491 56941 39605 57099
tri 39641 57066 39657 57082 se
rect 39657 57066 39734 57082
rect 39641 57000 39734 57066
rect 39362 56865 39734 56941
rect 39362 56740 39455 56806
rect 39362 56724 39439 56740
tri 39439 56724 39455 56740 nw
rect 39491 56707 39605 56865
rect 39641 56740 39734 56806
tri 39641 56724 39657 56740 ne
rect 39657 56724 39734 56740
rect 39474 56625 39622 56707
rect 39362 56592 39439 56608
tri 39439 56592 39455 56608 sw
rect 39362 56526 39455 56592
rect 39362 56424 39455 56490
rect 39362 56408 39439 56424
tri 39439 56408 39455 56424 nw
rect 39491 56391 39605 56625
tri 39641 56592 39657 56608 se
rect 39657 56592 39734 56608
rect 39641 56526 39734 56592
rect 39641 56424 39734 56490
tri 39641 56408 39657 56424 ne
rect 39657 56408 39734 56424
rect 39474 56309 39622 56391
rect 39362 56276 39439 56292
tri 39439 56276 39455 56292 sw
rect 39362 56210 39455 56276
rect 39491 56151 39605 56309
tri 39641 56276 39657 56292 se
rect 39657 56276 39734 56292
rect 39641 56210 39734 56276
rect 39362 56075 39734 56151
rect 39362 55950 39455 56016
rect 39362 55934 39439 55950
tri 39439 55934 39455 55950 nw
rect 39491 55917 39605 56075
rect 39641 55950 39734 56016
tri 39641 55934 39657 55950 ne
rect 39657 55934 39734 55950
rect 39474 55835 39622 55917
rect 39362 55802 39439 55818
tri 39439 55802 39455 55818 sw
rect 39362 55736 39455 55802
rect 39362 55634 39455 55700
rect 39362 55618 39439 55634
tri 39439 55618 39455 55634 nw
rect 39491 55601 39605 55835
tri 39641 55802 39657 55818 se
rect 39657 55802 39734 55818
rect 39641 55736 39734 55802
rect 39641 55634 39734 55700
tri 39641 55618 39657 55634 ne
rect 39657 55618 39734 55634
rect 39474 55519 39622 55601
rect 39362 55486 39439 55502
tri 39439 55486 39455 55502 sw
rect 39362 55420 39455 55486
rect 39491 55361 39605 55519
tri 39641 55486 39657 55502 se
rect 39657 55486 39734 55502
rect 39641 55420 39734 55486
rect 39362 55285 39734 55361
rect 39362 55160 39455 55226
rect 39362 55144 39439 55160
tri 39439 55144 39455 55160 nw
rect 39491 55127 39605 55285
rect 39641 55160 39734 55226
tri 39641 55144 39657 55160 ne
rect 39657 55144 39734 55160
rect 39474 55045 39622 55127
rect 39362 55012 39439 55028
tri 39439 55012 39455 55028 sw
rect 39362 54946 39455 55012
rect 39362 54844 39455 54910
rect 39362 54828 39439 54844
tri 39439 54828 39455 54844 nw
rect 39491 54811 39605 55045
tri 39641 55012 39657 55028 se
rect 39657 55012 39734 55028
rect 39641 54946 39734 55012
rect 39641 54844 39734 54910
tri 39641 54828 39657 54844 ne
rect 39657 54828 39734 54844
rect 39474 54729 39622 54811
rect 39362 54696 39439 54712
tri 39439 54696 39455 54712 sw
rect 39362 54630 39455 54696
rect 39491 54571 39605 54729
tri 39641 54696 39657 54712 se
rect 39657 54696 39734 54712
rect 39641 54630 39734 54696
rect 39362 54495 39734 54571
rect 39362 54370 39455 54436
rect 39362 54354 39439 54370
tri 39439 54354 39455 54370 nw
rect 39491 54337 39605 54495
rect 39641 54370 39734 54436
tri 39641 54354 39657 54370 ne
rect 39657 54354 39734 54370
rect 39474 54255 39622 54337
rect 39362 54222 39439 54238
tri 39439 54222 39455 54238 sw
rect 39362 54156 39455 54222
rect 39362 54054 39455 54120
rect 39362 54038 39439 54054
tri 39439 54038 39455 54054 nw
rect 39491 54021 39605 54255
tri 39641 54222 39657 54238 se
rect 39657 54222 39734 54238
rect 39641 54156 39734 54222
rect 39641 54054 39734 54120
tri 39641 54038 39657 54054 ne
rect 39657 54038 39734 54054
rect 39474 53939 39622 54021
rect 39362 53906 39439 53922
tri 39439 53906 39455 53922 sw
rect 39362 53840 39455 53906
rect 39491 53781 39605 53939
tri 39641 53906 39657 53922 se
rect 39657 53906 39734 53922
rect 39641 53840 39734 53906
rect 39362 53705 39734 53781
rect 39362 53580 39455 53646
rect 39362 53564 39439 53580
tri 39439 53564 39455 53580 nw
rect 39491 53547 39605 53705
rect 39641 53580 39734 53646
tri 39641 53564 39657 53580 ne
rect 39657 53564 39734 53580
rect 39474 53465 39622 53547
rect 39362 53432 39439 53448
tri 39439 53432 39455 53448 sw
rect 39362 53366 39455 53432
rect 39362 53264 39455 53330
rect 39362 53248 39439 53264
tri 39439 53248 39455 53264 nw
rect 39491 53231 39605 53465
tri 39641 53432 39657 53448 se
rect 39657 53432 39734 53448
rect 39641 53366 39734 53432
rect 39641 53264 39734 53330
tri 39641 53248 39657 53264 ne
rect 39657 53248 39734 53264
rect 39474 53149 39622 53231
rect 39362 53116 39439 53132
tri 39439 53116 39455 53132 sw
rect 39362 53050 39455 53116
rect 39491 52991 39605 53149
tri 39641 53116 39657 53132 se
rect 39657 53116 39734 53132
rect 39641 53050 39734 53116
rect 39362 52915 39734 52991
rect 39362 52790 39455 52856
rect 39362 52774 39439 52790
tri 39439 52774 39455 52790 nw
rect 39491 52757 39605 52915
rect 39641 52790 39734 52856
tri 39641 52774 39657 52790 ne
rect 39657 52774 39734 52790
rect 39474 52675 39622 52757
rect 39362 52642 39439 52658
tri 39439 52642 39455 52658 sw
rect 39362 52576 39455 52642
rect 39362 52474 39455 52540
rect 39362 52458 39439 52474
tri 39439 52458 39455 52474 nw
rect 39491 52441 39605 52675
tri 39641 52642 39657 52658 se
rect 39657 52642 39734 52658
rect 39641 52576 39734 52642
rect 39641 52474 39734 52540
tri 39641 52458 39657 52474 ne
rect 39657 52458 39734 52474
rect 39474 52359 39622 52441
rect 39362 52326 39439 52342
tri 39439 52326 39455 52342 sw
rect 39362 52260 39455 52326
rect 39491 52201 39605 52359
tri 39641 52326 39657 52342 se
rect 39657 52326 39734 52342
rect 39641 52260 39734 52326
rect 39362 52125 39734 52201
rect 39362 52000 39455 52066
rect 39362 51984 39439 52000
tri 39439 51984 39455 52000 nw
rect 39491 51967 39605 52125
rect 39641 52000 39734 52066
tri 39641 51984 39657 52000 ne
rect 39657 51984 39734 52000
rect 39474 51885 39622 51967
rect 39362 51852 39439 51868
tri 39439 51852 39455 51868 sw
rect 39362 51786 39455 51852
rect 39362 51684 39455 51750
rect 39362 51668 39439 51684
tri 39439 51668 39455 51684 nw
rect 39491 51651 39605 51885
tri 39641 51852 39657 51868 se
rect 39657 51852 39734 51868
rect 39641 51786 39734 51852
rect 39641 51684 39734 51750
tri 39641 51668 39657 51684 ne
rect 39657 51668 39734 51684
rect 39474 51569 39622 51651
rect 39362 51536 39439 51552
tri 39439 51536 39455 51552 sw
rect 39362 51470 39455 51536
rect 39491 51411 39605 51569
tri 39641 51536 39657 51552 se
rect 39657 51536 39734 51552
rect 39641 51470 39734 51536
rect 39362 51335 39734 51411
rect 39362 51210 39455 51276
rect 39362 51194 39439 51210
tri 39439 51194 39455 51210 nw
rect 39491 51177 39605 51335
rect 39641 51210 39734 51276
tri 39641 51194 39657 51210 ne
rect 39657 51194 39734 51210
rect 39474 51095 39622 51177
rect 39362 51062 39439 51078
tri 39439 51062 39455 51078 sw
rect 39362 50996 39455 51062
rect 39362 50894 39455 50960
rect 39362 50878 39439 50894
tri 39439 50878 39455 50894 nw
rect 39491 50861 39605 51095
tri 39641 51062 39657 51078 se
rect 39657 51062 39734 51078
rect 39641 50996 39734 51062
rect 39641 50894 39734 50960
tri 39641 50878 39657 50894 ne
rect 39657 50878 39734 50894
rect 39474 50779 39622 50861
rect 39362 50746 39439 50762
tri 39439 50746 39455 50762 sw
rect 39362 50680 39455 50746
rect 39491 50621 39605 50779
tri 39641 50746 39657 50762 se
rect 39657 50746 39734 50762
rect 39641 50680 39734 50746
rect 39362 50545 39734 50621
rect 39362 50420 39455 50486
rect 39362 50404 39439 50420
tri 39439 50404 39455 50420 nw
rect 39491 50387 39605 50545
rect 39641 50420 39734 50486
tri 39641 50404 39657 50420 ne
rect 39657 50404 39734 50420
rect 39474 50305 39622 50387
rect 39362 50272 39439 50288
tri 39439 50272 39455 50288 sw
rect 39362 50206 39455 50272
rect 39362 50104 39455 50170
rect 39362 50088 39439 50104
tri 39439 50088 39455 50104 nw
rect 39491 50071 39605 50305
tri 39641 50272 39657 50288 se
rect 39657 50272 39734 50288
rect 39641 50206 39734 50272
rect 39641 50104 39734 50170
tri 39641 50088 39657 50104 ne
rect 39657 50088 39734 50104
rect 39474 49989 39622 50071
rect 39362 49956 39439 49972
tri 39439 49956 39455 49972 sw
rect 39362 49890 39455 49956
rect 39491 49831 39605 49989
tri 39641 49956 39657 49972 se
rect 39657 49956 39734 49972
rect 39641 49890 39734 49956
rect 39362 49755 39734 49831
rect 39362 49630 39455 49696
rect 39362 49614 39439 49630
tri 39439 49614 39455 49630 nw
rect 39491 49597 39605 49755
rect 39641 49630 39734 49696
tri 39641 49614 39657 49630 ne
rect 39657 49614 39734 49630
rect 39474 49515 39622 49597
rect 39362 49482 39439 49498
tri 39439 49482 39455 49498 sw
rect 39362 49416 39455 49482
rect 39362 49314 39455 49380
rect 39362 49298 39439 49314
tri 39439 49298 39455 49314 nw
rect 39491 49281 39605 49515
tri 39641 49482 39657 49498 se
rect 39657 49482 39734 49498
rect 39641 49416 39734 49482
rect 39641 49314 39734 49380
tri 39641 49298 39657 49314 ne
rect 39657 49298 39734 49314
rect 39474 49199 39622 49281
rect 39362 49166 39439 49182
tri 39439 49166 39455 49182 sw
rect 39362 49100 39455 49166
rect 39491 49041 39605 49199
tri 39641 49166 39657 49182 se
rect 39657 49166 39734 49182
rect 39641 49100 39734 49166
rect 39362 48965 39734 49041
rect 39362 48840 39455 48906
rect 39362 48824 39439 48840
tri 39439 48824 39455 48840 nw
rect 39491 48807 39605 48965
rect 39641 48840 39734 48906
tri 39641 48824 39657 48840 ne
rect 39657 48824 39734 48840
rect 39474 48725 39622 48807
rect 39362 48692 39439 48708
tri 39439 48692 39455 48708 sw
rect 39362 48626 39455 48692
rect 39362 48524 39455 48590
rect 39362 48508 39439 48524
tri 39439 48508 39455 48524 nw
rect 39491 48491 39605 48725
tri 39641 48692 39657 48708 se
rect 39657 48692 39734 48708
rect 39641 48626 39734 48692
rect 39641 48524 39734 48590
tri 39641 48508 39657 48524 ne
rect 39657 48508 39734 48524
rect 39474 48409 39622 48491
rect 39362 48376 39439 48392
tri 39439 48376 39455 48392 sw
rect 39362 48310 39455 48376
rect 39491 48251 39605 48409
tri 39641 48376 39657 48392 se
rect 39657 48376 39734 48392
rect 39641 48310 39734 48376
rect 39362 48175 39734 48251
rect 39362 48050 39455 48116
rect 39362 48034 39439 48050
tri 39439 48034 39455 48050 nw
rect 39491 48017 39605 48175
rect 39641 48050 39734 48116
tri 39641 48034 39657 48050 ne
rect 39657 48034 39734 48050
rect 39474 47935 39622 48017
rect 39362 47902 39439 47918
tri 39439 47902 39455 47918 sw
rect 39362 47836 39455 47902
rect 39362 47734 39455 47800
rect 39362 47718 39439 47734
tri 39439 47718 39455 47734 nw
rect 39491 47701 39605 47935
tri 39641 47902 39657 47918 se
rect 39657 47902 39734 47918
rect 39641 47836 39734 47902
rect 39641 47734 39734 47800
tri 39641 47718 39657 47734 ne
rect 39657 47718 39734 47734
rect 39474 47619 39622 47701
rect 39362 47586 39439 47602
tri 39439 47586 39455 47602 sw
rect 39362 47520 39455 47586
rect 39491 47461 39605 47619
tri 39641 47586 39657 47602 se
rect 39657 47586 39734 47602
rect 39641 47520 39734 47586
rect 39362 47385 39734 47461
rect 39362 47260 39455 47326
rect 39362 47244 39439 47260
tri 39439 47244 39455 47260 nw
rect 39491 47227 39605 47385
rect 39641 47260 39734 47326
tri 39641 47244 39657 47260 ne
rect 39657 47244 39734 47260
rect 39474 47145 39622 47227
rect 39362 47112 39439 47128
tri 39439 47112 39455 47128 sw
rect 39362 47046 39455 47112
rect 39362 46944 39455 47010
rect 39362 46928 39439 46944
tri 39439 46928 39455 46944 nw
rect 39491 46911 39605 47145
tri 39641 47112 39657 47128 se
rect 39657 47112 39734 47128
rect 39641 47046 39734 47112
rect 39641 46944 39734 47010
tri 39641 46928 39657 46944 ne
rect 39657 46928 39734 46944
rect 39474 46829 39622 46911
rect 39362 46796 39439 46812
tri 39439 46796 39455 46812 sw
rect 39362 46730 39455 46796
rect 39491 46671 39605 46829
tri 39641 46796 39657 46812 se
rect 39657 46796 39734 46812
rect 39641 46730 39734 46796
rect 39362 46595 39734 46671
rect 39362 46470 39455 46536
rect 39362 46454 39439 46470
tri 39439 46454 39455 46470 nw
rect 39491 46437 39605 46595
rect 39641 46470 39734 46536
tri 39641 46454 39657 46470 ne
rect 39657 46454 39734 46470
rect 39474 46355 39622 46437
rect 39362 46322 39439 46338
tri 39439 46322 39455 46338 sw
rect 39362 46256 39455 46322
rect 39362 46154 39455 46220
rect 39362 46138 39439 46154
tri 39439 46138 39455 46154 nw
rect 39491 46121 39605 46355
tri 39641 46322 39657 46338 se
rect 39657 46322 39734 46338
rect 39641 46256 39734 46322
rect 39641 46154 39734 46220
tri 39641 46138 39657 46154 ne
rect 39657 46138 39734 46154
rect 39474 46039 39622 46121
rect 39362 46006 39439 46022
tri 39439 46006 39455 46022 sw
rect 39362 45940 39455 46006
rect 39491 45881 39605 46039
tri 39641 46006 39657 46022 se
rect 39657 46006 39734 46022
rect 39641 45940 39734 46006
rect 39362 45805 39734 45881
rect 39362 45680 39455 45746
rect 39362 45664 39439 45680
tri 39439 45664 39455 45680 nw
rect 39491 45647 39605 45805
rect 39641 45680 39734 45746
tri 39641 45664 39657 45680 ne
rect 39657 45664 39734 45680
rect 39474 45565 39622 45647
rect 39362 45532 39439 45548
tri 39439 45532 39455 45548 sw
rect 39362 45466 39455 45532
rect 39362 45364 39455 45430
rect 39362 45348 39439 45364
tri 39439 45348 39455 45364 nw
rect 39491 45331 39605 45565
tri 39641 45532 39657 45548 se
rect 39657 45532 39734 45548
rect 39641 45466 39734 45532
rect 39641 45364 39734 45430
tri 39641 45348 39657 45364 ne
rect 39657 45348 39734 45364
rect 39474 45249 39622 45331
rect 39362 45216 39439 45232
tri 39439 45216 39455 45232 sw
rect 39362 45150 39455 45216
rect 39491 45091 39605 45249
tri 39641 45216 39657 45232 se
rect 39657 45216 39734 45232
rect 39641 45150 39734 45216
rect 39362 45015 39734 45091
rect 39362 44890 39455 44956
rect 39362 44874 39439 44890
tri 39439 44874 39455 44890 nw
rect 39491 44857 39605 45015
rect 39641 44890 39734 44956
tri 39641 44874 39657 44890 ne
rect 39657 44874 39734 44890
rect 39474 44775 39622 44857
rect 39362 44742 39439 44758
tri 39439 44742 39455 44758 sw
rect 39362 44676 39455 44742
rect 39362 44574 39455 44640
rect 39362 44558 39439 44574
tri 39439 44558 39455 44574 nw
rect 39491 44541 39605 44775
tri 39641 44742 39657 44758 se
rect 39657 44742 39734 44758
rect 39641 44676 39734 44742
rect 39641 44574 39734 44640
tri 39641 44558 39657 44574 ne
rect 39657 44558 39734 44574
rect 39474 44459 39622 44541
rect 39362 44426 39439 44442
tri 39439 44426 39455 44442 sw
rect 39362 44360 39455 44426
rect 39491 44301 39605 44459
tri 39641 44426 39657 44442 se
rect 39657 44426 39734 44442
rect 39641 44360 39734 44426
rect 39362 44225 39734 44301
rect 39362 44100 39455 44166
rect 39362 44084 39439 44100
tri 39439 44084 39455 44100 nw
rect 39491 44067 39605 44225
rect 39641 44100 39734 44166
tri 39641 44084 39657 44100 ne
rect 39657 44084 39734 44100
rect 39474 43985 39622 44067
rect 39362 43952 39439 43968
tri 39439 43952 39455 43968 sw
rect 39362 43886 39455 43952
rect 39362 43784 39455 43850
rect 39362 43768 39439 43784
tri 39439 43768 39455 43784 nw
rect 39491 43751 39605 43985
tri 39641 43952 39657 43968 se
rect 39657 43952 39734 43968
rect 39641 43886 39734 43952
rect 39641 43784 39734 43850
tri 39641 43768 39657 43784 ne
rect 39657 43768 39734 43784
rect 39474 43669 39622 43751
rect 39362 43636 39439 43652
tri 39439 43636 39455 43652 sw
rect 39362 43570 39455 43636
rect 39491 43511 39605 43669
tri 39641 43636 39657 43652 se
rect 39657 43636 39734 43652
rect 39641 43570 39734 43636
rect 39362 43435 39734 43511
rect 39362 43310 39455 43376
rect 39362 43294 39439 43310
tri 39439 43294 39455 43310 nw
rect 39491 43277 39605 43435
rect 39641 43310 39734 43376
tri 39641 43294 39657 43310 ne
rect 39657 43294 39734 43310
rect 39474 43195 39622 43277
rect 39362 43162 39439 43178
tri 39439 43162 39455 43178 sw
rect 39362 43096 39455 43162
rect 39362 42994 39455 43060
rect 39362 42978 39439 42994
tri 39439 42978 39455 42994 nw
rect 39491 42961 39605 43195
tri 39641 43162 39657 43178 se
rect 39657 43162 39734 43178
rect 39641 43096 39734 43162
rect 39641 42994 39734 43060
tri 39641 42978 39657 42994 ne
rect 39657 42978 39734 42994
rect 39474 42879 39622 42961
rect 39362 42846 39439 42862
tri 39439 42846 39455 42862 sw
rect 39362 42780 39455 42846
rect 39491 42721 39605 42879
tri 39641 42846 39657 42862 se
rect 39657 42846 39734 42862
rect 39641 42780 39734 42846
rect 39362 42645 39734 42721
rect 39362 42520 39455 42586
rect 39362 42504 39439 42520
tri 39439 42504 39455 42520 nw
rect 39491 42487 39605 42645
rect 39641 42520 39734 42586
tri 39641 42504 39657 42520 ne
rect 39657 42504 39734 42520
rect 39474 42405 39622 42487
rect 39362 42372 39439 42388
tri 39439 42372 39455 42388 sw
rect 39362 42306 39455 42372
rect 39362 42204 39455 42270
rect 39362 42188 39439 42204
tri 39439 42188 39455 42204 nw
rect 39491 42171 39605 42405
tri 39641 42372 39657 42388 se
rect 39657 42372 39734 42388
rect 39641 42306 39734 42372
rect 39641 42204 39734 42270
tri 39641 42188 39657 42204 ne
rect 39657 42188 39734 42204
rect 39474 42089 39622 42171
rect 39362 42056 39439 42072
tri 39439 42056 39455 42072 sw
rect 39362 41990 39455 42056
rect 39491 41931 39605 42089
tri 39641 42056 39657 42072 se
rect 39657 42056 39734 42072
rect 39641 41990 39734 42056
rect 39362 41855 39734 41931
rect 39362 41730 39455 41796
rect 39362 41714 39439 41730
tri 39439 41714 39455 41730 nw
rect 39491 41697 39605 41855
rect 39641 41730 39734 41796
tri 39641 41714 39657 41730 ne
rect 39657 41714 39734 41730
rect 39474 41615 39622 41697
rect 39362 41582 39439 41598
tri 39439 41582 39455 41598 sw
rect 39362 41516 39455 41582
rect 39362 41414 39455 41480
rect 39362 41398 39439 41414
tri 39439 41398 39455 41414 nw
rect 39491 41381 39605 41615
tri 39641 41582 39657 41598 se
rect 39657 41582 39734 41598
rect 39641 41516 39734 41582
rect 39641 41414 39734 41480
tri 39641 41398 39657 41414 ne
rect 39657 41398 39734 41414
rect 39474 41299 39622 41381
rect 39362 41266 39439 41282
tri 39439 41266 39455 41282 sw
rect 39362 41200 39455 41266
rect 39491 41141 39605 41299
tri 39641 41266 39657 41282 se
rect 39657 41266 39734 41282
rect 39641 41200 39734 41266
rect 39362 41065 39734 41141
rect 39362 40940 39455 41006
rect 39362 40924 39439 40940
tri 39439 40924 39455 40940 nw
rect 39491 40907 39605 41065
rect 39641 40940 39734 41006
tri 39641 40924 39657 40940 ne
rect 39657 40924 39734 40940
rect 39474 40825 39622 40907
rect 39362 40792 39439 40808
tri 39439 40792 39455 40808 sw
rect 39362 40726 39455 40792
rect 39362 40624 39455 40690
rect 39362 40608 39439 40624
tri 39439 40608 39455 40624 nw
rect 39491 40591 39605 40825
tri 39641 40792 39657 40808 se
rect 39657 40792 39734 40808
rect 39641 40726 39734 40792
rect 39641 40624 39734 40690
tri 39641 40608 39657 40624 ne
rect 39657 40608 39734 40624
rect 39474 40509 39622 40591
rect 39362 40476 39439 40492
tri 39439 40476 39455 40492 sw
rect 39362 40410 39455 40476
rect 39491 40351 39605 40509
tri 39641 40476 39657 40492 se
rect 39657 40476 39734 40492
rect 39641 40410 39734 40476
rect 39362 40275 39734 40351
rect 39362 40150 39455 40216
rect 39362 40134 39439 40150
tri 39439 40134 39455 40150 nw
rect 39491 40117 39605 40275
rect 39641 40150 39734 40216
tri 39641 40134 39657 40150 ne
rect 39657 40134 39734 40150
rect 39474 40035 39622 40117
rect 39362 40002 39439 40018
tri 39439 40002 39455 40018 sw
rect 39362 39936 39455 40002
rect 39362 39834 39455 39900
rect 39362 39818 39439 39834
tri 39439 39818 39455 39834 nw
rect 39491 39801 39605 40035
tri 39641 40002 39657 40018 se
rect 39657 40002 39734 40018
rect 39641 39936 39734 40002
rect 39641 39834 39734 39900
tri 39641 39818 39657 39834 ne
rect 39657 39818 39734 39834
rect 39474 39719 39622 39801
rect 39362 39686 39439 39702
tri 39439 39686 39455 39702 sw
rect 39362 39620 39455 39686
rect 39491 39561 39605 39719
tri 39641 39686 39657 39702 se
rect 39657 39686 39734 39702
rect 39641 39620 39734 39686
rect 39362 39485 39734 39561
rect 39362 39360 39455 39426
rect 39362 39344 39439 39360
tri 39439 39344 39455 39360 nw
rect 39491 39327 39605 39485
rect 39641 39360 39734 39426
tri 39641 39344 39657 39360 ne
rect 39657 39344 39734 39360
rect 39474 39245 39622 39327
rect 39362 39212 39439 39228
tri 39439 39212 39455 39228 sw
rect 39362 39146 39455 39212
rect 39362 39044 39455 39110
rect 39362 39028 39439 39044
tri 39439 39028 39455 39044 nw
rect 39491 39011 39605 39245
tri 39641 39212 39657 39228 se
rect 39657 39212 39734 39228
rect 39641 39146 39734 39212
rect 39641 39044 39734 39110
tri 39641 39028 39657 39044 ne
rect 39657 39028 39734 39044
rect 39474 38929 39622 39011
rect 39362 38896 39439 38912
tri 39439 38896 39455 38912 sw
rect 39362 38830 39455 38896
rect 39491 38771 39605 38929
tri 39641 38896 39657 38912 se
rect 39657 38896 39734 38912
rect 39641 38830 39734 38896
rect 39362 38695 39734 38771
rect 39362 38570 39455 38636
rect 39362 38554 39439 38570
tri 39439 38554 39455 38570 nw
rect 39491 38537 39605 38695
rect 39641 38570 39734 38636
tri 39641 38554 39657 38570 ne
rect 39657 38554 39734 38570
rect 39474 38455 39622 38537
rect 39362 38422 39439 38438
tri 39439 38422 39455 38438 sw
rect 39362 38356 39455 38422
rect 39362 38254 39455 38320
rect 39362 38238 39439 38254
tri 39439 38238 39455 38254 nw
rect 39491 38221 39605 38455
tri 39641 38422 39657 38438 se
rect 39657 38422 39734 38438
rect 39641 38356 39734 38422
rect 39641 38254 39734 38320
tri 39641 38238 39657 38254 ne
rect 39657 38238 39734 38254
rect 39474 38139 39622 38221
rect 39362 38106 39439 38122
tri 39439 38106 39455 38122 sw
rect 39362 38040 39455 38106
rect 39491 37981 39605 38139
tri 39641 38106 39657 38122 se
rect 39657 38106 39734 38122
rect 39641 38040 39734 38106
rect 39362 37905 39734 37981
rect 39362 37780 39455 37846
rect 39362 37764 39439 37780
tri 39439 37764 39455 37780 nw
rect 39491 37747 39605 37905
rect 39641 37780 39734 37846
tri 39641 37764 39657 37780 ne
rect 39657 37764 39734 37780
rect 39474 37665 39622 37747
rect 39362 37632 39439 37648
tri 39439 37632 39455 37648 sw
rect 39362 37566 39455 37632
rect 39362 37464 39455 37530
rect 39362 37448 39439 37464
tri 39439 37448 39455 37464 nw
rect 39491 37431 39605 37665
tri 39641 37632 39657 37648 se
rect 39657 37632 39734 37648
rect 39641 37566 39734 37632
rect 39641 37464 39734 37530
tri 39641 37448 39657 37464 ne
rect 39657 37448 39734 37464
rect 39474 37349 39622 37431
rect 39362 37316 39439 37332
tri 39439 37316 39455 37332 sw
rect 39362 37250 39455 37316
rect 39491 37191 39605 37349
tri 39641 37316 39657 37332 se
rect 39657 37316 39734 37332
rect 39641 37250 39734 37316
rect 39362 37115 39734 37191
rect 39362 36990 39455 37056
rect 39362 36974 39439 36990
tri 39439 36974 39455 36990 nw
rect 39491 36957 39605 37115
rect 39641 36990 39734 37056
tri 39641 36974 39657 36990 ne
rect 39657 36974 39734 36990
rect 39474 36875 39622 36957
rect 39362 36842 39439 36858
tri 39439 36842 39455 36858 sw
rect 39362 36776 39455 36842
rect 39362 36674 39455 36740
rect 39362 36658 39439 36674
tri 39439 36658 39455 36674 nw
rect 39491 36641 39605 36875
tri 39641 36842 39657 36858 se
rect 39657 36842 39734 36858
rect 39641 36776 39734 36842
rect 39641 36674 39734 36740
tri 39641 36658 39657 36674 ne
rect 39657 36658 39734 36674
rect 39474 36559 39622 36641
rect 39362 36526 39439 36542
tri 39439 36526 39455 36542 sw
rect 39362 36460 39455 36526
rect 39491 36401 39605 36559
tri 39641 36526 39657 36542 se
rect 39657 36526 39734 36542
rect 39641 36460 39734 36526
rect 39362 36325 39734 36401
rect 39362 36200 39455 36266
rect 39362 36184 39439 36200
tri 39439 36184 39455 36200 nw
rect 39491 36167 39605 36325
rect 39641 36200 39734 36266
tri 39641 36184 39657 36200 ne
rect 39657 36184 39734 36200
rect 39474 36085 39622 36167
rect 39362 36052 39439 36068
tri 39439 36052 39455 36068 sw
rect 39362 35986 39455 36052
rect 39362 35884 39455 35950
rect 39362 35868 39439 35884
tri 39439 35868 39455 35884 nw
rect 39491 35851 39605 36085
tri 39641 36052 39657 36068 se
rect 39657 36052 39734 36068
rect 39641 35986 39734 36052
rect 39641 35884 39734 35950
tri 39641 35868 39657 35884 ne
rect 39657 35868 39734 35884
rect 39474 35769 39622 35851
rect 39362 35736 39439 35752
tri 39439 35736 39455 35752 sw
rect 39362 35670 39455 35736
rect 39491 35611 39605 35769
tri 39641 35736 39657 35752 se
rect 39657 35736 39734 35752
rect 39641 35670 39734 35736
rect 39362 35535 39734 35611
rect 39362 35410 39455 35476
rect 39362 35394 39439 35410
tri 39439 35394 39455 35410 nw
rect 39491 35377 39605 35535
rect 39641 35410 39734 35476
tri 39641 35394 39657 35410 ne
rect 39657 35394 39734 35410
rect 39474 35295 39622 35377
rect 39362 35262 39439 35278
tri 39439 35262 39455 35278 sw
rect 39362 35196 39455 35262
rect 39362 35094 39455 35160
rect 39362 35078 39439 35094
tri 39439 35078 39455 35094 nw
rect 39491 35061 39605 35295
tri 39641 35262 39657 35278 se
rect 39657 35262 39734 35278
rect 39641 35196 39734 35262
rect 39641 35094 39734 35160
tri 39641 35078 39657 35094 ne
rect 39657 35078 39734 35094
rect 39474 34979 39622 35061
rect 39362 34946 39439 34962
tri 39439 34946 39455 34962 sw
rect 39362 34880 39455 34946
rect 39491 34821 39605 34979
tri 39641 34946 39657 34962 se
rect 39657 34946 39734 34962
rect 39641 34880 39734 34946
rect 39362 34745 39734 34821
rect 39362 34620 39455 34686
rect 39362 34604 39439 34620
tri 39439 34604 39455 34620 nw
rect 39491 34587 39605 34745
rect 39641 34620 39734 34686
tri 39641 34604 39657 34620 ne
rect 39657 34604 39734 34620
rect 39474 34505 39622 34587
rect 39362 34472 39439 34488
tri 39439 34472 39455 34488 sw
rect 39362 34406 39455 34472
rect 39362 34304 39455 34370
rect 39362 34288 39439 34304
tri 39439 34288 39455 34304 nw
rect 39491 34271 39605 34505
tri 39641 34472 39657 34488 se
rect 39657 34472 39734 34488
rect 39641 34406 39734 34472
rect 39641 34304 39734 34370
tri 39641 34288 39657 34304 ne
rect 39657 34288 39734 34304
rect 39474 34189 39622 34271
rect 39362 34156 39439 34172
tri 39439 34156 39455 34172 sw
rect 39362 34090 39455 34156
rect 39491 34031 39605 34189
tri 39641 34156 39657 34172 se
rect 39657 34156 39734 34172
rect 39641 34090 39734 34156
rect 39362 33955 39734 34031
rect 39362 33830 39455 33896
rect 39362 33814 39439 33830
tri 39439 33814 39455 33830 nw
rect 39491 33797 39605 33955
rect 39641 33830 39734 33896
tri 39641 33814 39657 33830 ne
rect 39657 33814 39734 33830
rect 39474 33715 39622 33797
rect 39362 33682 39439 33698
tri 39439 33682 39455 33698 sw
rect 39362 33616 39455 33682
rect 39362 33514 39455 33580
rect 39362 33498 39439 33514
tri 39439 33498 39455 33514 nw
rect 39491 33481 39605 33715
tri 39641 33682 39657 33698 se
rect 39657 33682 39734 33698
rect 39641 33616 39734 33682
rect 39641 33514 39734 33580
tri 39641 33498 39657 33514 ne
rect 39657 33498 39734 33514
rect 39474 33399 39622 33481
rect 39362 33366 39439 33382
tri 39439 33366 39455 33382 sw
rect 39362 33300 39455 33366
rect 39491 33241 39605 33399
tri 39641 33366 39657 33382 se
rect 39657 33366 39734 33382
rect 39641 33300 39734 33366
rect 39362 33165 39734 33241
rect 39362 33040 39455 33106
rect 39362 33024 39439 33040
tri 39439 33024 39455 33040 nw
rect 39491 33007 39605 33165
rect 39641 33040 39734 33106
tri 39641 33024 39657 33040 ne
rect 39657 33024 39734 33040
rect 39474 32925 39622 33007
rect 39362 32892 39439 32908
tri 39439 32892 39455 32908 sw
rect 39362 32826 39455 32892
rect 39362 32724 39455 32790
rect 39362 32708 39439 32724
tri 39439 32708 39455 32724 nw
rect 39491 32691 39605 32925
tri 39641 32892 39657 32908 se
rect 39657 32892 39734 32908
rect 39641 32826 39734 32892
rect 39641 32724 39734 32790
tri 39641 32708 39657 32724 ne
rect 39657 32708 39734 32724
rect 39474 32609 39622 32691
rect 39362 32576 39439 32592
tri 39439 32576 39455 32592 sw
rect 39362 32510 39455 32576
rect 39491 32451 39605 32609
tri 39641 32576 39657 32592 se
rect 39657 32576 39734 32592
rect 39641 32510 39734 32576
rect 39362 32375 39734 32451
rect 39362 32250 39455 32316
rect 39362 32234 39439 32250
tri 39439 32234 39455 32250 nw
rect 39491 32217 39605 32375
rect 39641 32250 39734 32316
tri 39641 32234 39657 32250 ne
rect 39657 32234 39734 32250
rect 39474 32135 39622 32217
rect 39362 32102 39439 32118
tri 39439 32102 39455 32118 sw
rect 39362 32036 39455 32102
rect 39362 31934 39455 32000
rect 39362 31918 39439 31934
tri 39439 31918 39455 31934 nw
rect 39491 31901 39605 32135
tri 39641 32102 39657 32118 se
rect 39657 32102 39734 32118
rect 39641 32036 39734 32102
rect 39641 31934 39734 32000
tri 39641 31918 39657 31934 ne
rect 39657 31918 39734 31934
rect 39474 31819 39622 31901
rect 39362 31786 39439 31802
tri 39439 31786 39455 31802 sw
rect 39362 31720 39455 31786
rect 39491 31661 39605 31819
tri 39641 31786 39657 31802 se
rect 39657 31786 39734 31802
rect 39641 31720 39734 31786
rect 39362 31585 39734 31661
rect 39362 31460 39455 31526
rect 39362 31444 39439 31460
tri 39439 31444 39455 31460 nw
rect 39491 31427 39605 31585
rect 39641 31460 39734 31526
tri 39641 31444 39657 31460 ne
rect 39657 31444 39734 31460
rect 39474 31345 39622 31427
rect 39362 31312 39439 31328
tri 39439 31312 39455 31328 sw
rect 39362 31246 39455 31312
rect 39362 31144 39455 31210
rect 39362 31128 39439 31144
tri 39439 31128 39455 31144 nw
rect 39491 31111 39605 31345
tri 39641 31312 39657 31328 se
rect 39657 31312 39734 31328
rect 39641 31246 39734 31312
rect 39641 31144 39734 31210
tri 39641 31128 39657 31144 ne
rect 39657 31128 39734 31144
rect 39474 31029 39622 31111
rect 39362 30996 39439 31012
tri 39439 30996 39455 31012 sw
rect 39362 30930 39455 30996
rect 39491 30871 39605 31029
tri 39641 30996 39657 31012 se
rect 39657 30996 39734 31012
rect 39641 30930 39734 30996
rect 39362 30795 39734 30871
rect 39362 30670 39455 30736
rect 39362 30654 39439 30670
tri 39439 30654 39455 30670 nw
rect 39491 30637 39605 30795
rect 39641 30670 39734 30736
tri 39641 30654 39657 30670 ne
rect 39657 30654 39734 30670
rect 39474 30555 39622 30637
rect 39362 30522 39439 30538
tri 39439 30522 39455 30538 sw
rect 39362 30456 39455 30522
rect 39362 30354 39455 30420
rect 39362 30338 39439 30354
tri 39439 30338 39455 30354 nw
rect 39491 30321 39605 30555
tri 39641 30522 39657 30538 se
rect 39657 30522 39734 30538
rect 39641 30456 39734 30522
rect 39641 30354 39734 30420
tri 39641 30338 39657 30354 ne
rect 39657 30338 39734 30354
rect 39474 30239 39622 30321
rect 39362 30206 39439 30222
tri 39439 30206 39455 30222 sw
rect 39362 30140 39455 30206
rect 39491 30081 39605 30239
tri 39641 30206 39657 30222 se
rect 39657 30206 39734 30222
rect 39641 30140 39734 30206
rect 39362 30005 39734 30081
rect 39362 29880 39455 29946
rect 39362 29864 39439 29880
tri 39439 29864 39455 29880 nw
rect 39491 29847 39605 30005
rect 39641 29880 39734 29946
tri 39641 29864 39657 29880 ne
rect 39657 29864 39734 29880
rect 39474 29765 39622 29847
rect 39362 29732 39439 29748
tri 39439 29732 39455 29748 sw
rect 39362 29666 39455 29732
rect 39362 29564 39455 29630
rect 39362 29548 39439 29564
tri 39439 29548 39455 29564 nw
rect 39491 29531 39605 29765
tri 39641 29732 39657 29748 se
rect 39657 29732 39734 29748
rect 39641 29666 39734 29732
rect 39641 29564 39734 29630
tri 39641 29548 39657 29564 ne
rect 39657 29548 39734 29564
rect 39474 29449 39622 29531
rect 39362 29416 39439 29432
tri 39439 29416 39455 29432 sw
rect 39362 29350 39455 29416
rect 39491 29291 39605 29449
tri 39641 29416 39657 29432 se
rect 39657 29416 39734 29432
rect 39641 29350 39734 29416
rect 39362 29215 39734 29291
rect 39362 29090 39455 29156
rect 39362 29074 39439 29090
tri 39439 29074 39455 29090 nw
rect 39491 29057 39605 29215
rect 39641 29090 39734 29156
tri 39641 29074 39657 29090 ne
rect 39657 29074 39734 29090
rect 39474 28975 39622 29057
rect 39362 28942 39439 28958
tri 39439 28942 39455 28958 sw
rect 39362 28876 39455 28942
rect 39491 28833 39605 28975
tri 39641 28942 39657 28958 se
rect 39657 28942 39734 28958
rect 39641 28876 39734 28942
rect 39770 28463 39806 80603
rect 39842 28463 39878 80603
rect 39914 80445 39950 80603
rect 39906 80303 39958 80445
rect 39914 28763 39950 80303
rect 39906 28621 39958 28763
rect 39914 28463 39950 28621
rect 39986 28463 40022 80603
rect 40058 28463 40094 80603
rect 40130 28833 40214 80233
rect 40250 28463 40286 80603
rect 40322 28463 40358 80603
rect 40394 80445 40430 80603
rect 40386 80303 40438 80445
rect 40394 28763 40430 80303
rect 40386 28621 40438 28763
rect 40394 28463 40430 28621
rect 40466 28463 40502 80603
rect 40538 28463 40574 80603
rect 40610 80124 40703 80190
rect 40610 80108 40687 80124
tri 40687 80108 40703 80124 nw
rect 40739 80091 40853 80233
rect 40889 80124 40982 80190
tri 40889 80108 40905 80124 ne
rect 40905 80108 40982 80124
rect 40722 80009 40870 80091
rect 40610 79976 40687 79992
tri 40687 79976 40703 79992 sw
rect 40610 79910 40703 79976
rect 40739 79851 40853 80009
tri 40889 79976 40905 79992 se
rect 40905 79976 40982 79992
rect 40889 79910 40982 79976
rect 40610 79775 40982 79851
rect 40610 79650 40703 79716
rect 40610 79634 40687 79650
tri 40687 79634 40703 79650 nw
rect 40739 79617 40853 79775
rect 40889 79650 40982 79716
tri 40889 79634 40905 79650 ne
rect 40905 79634 40982 79650
rect 40722 79535 40870 79617
rect 40610 79502 40687 79518
tri 40687 79502 40703 79518 sw
rect 40610 79436 40703 79502
rect 40610 79334 40703 79400
rect 40610 79318 40687 79334
tri 40687 79318 40703 79334 nw
rect 40739 79301 40853 79535
tri 40889 79502 40905 79518 se
rect 40905 79502 40982 79518
rect 40889 79436 40982 79502
rect 40889 79334 40982 79400
tri 40889 79318 40905 79334 ne
rect 40905 79318 40982 79334
rect 40722 79219 40870 79301
rect 40610 79186 40687 79202
tri 40687 79186 40703 79202 sw
rect 40610 79120 40703 79186
rect 40739 79061 40853 79219
tri 40889 79186 40905 79202 se
rect 40905 79186 40982 79202
rect 40889 79120 40982 79186
rect 40610 78985 40982 79061
rect 40610 78860 40703 78926
rect 40610 78844 40687 78860
tri 40687 78844 40703 78860 nw
rect 40739 78827 40853 78985
rect 40889 78860 40982 78926
tri 40889 78844 40905 78860 ne
rect 40905 78844 40982 78860
rect 40722 78745 40870 78827
rect 40610 78712 40687 78728
tri 40687 78712 40703 78728 sw
rect 40610 78646 40703 78712
rect 40610 78544 40703 78610
rect 40610 78528 40687 78544
tri 40687 78528 40703 78544 nw
rect 40739 78511 40853 78745
tri 40889 78712 40905 78728 se
rect 40905 78712 40982 78728
rect 40889 78646 40982 78712
rect 40889 78544 40982 78610
tri 40889 78528 40905 78544 ne
rect 40905 78528 40982 78544
rect 40722 78429 40870 78511
rect 40610 78396 40687 78412
tri 40687 78396 40703 78412 sw
rect 40610 78330 40703 78396
rect 40739 78271 40853 78429
tri 40889 78396 40905 78412 se
rect 40905 78396 40982 78412
rect 40889 78330 40982 78396
rect 40610 78195 40982 78271
rect 40610 78070 40703 78136
rect 40610 78054 40687 78070
tri 40687 78054 40703 78070 nw
rect 40739 78037 40853 78195
rect 40889 78070 40982 78136
tri 40889 78054 40905 78070 ne
rect 40905 78054 40982 78070
rect 40722 77955 40870 78037
rect 40610 77922 40687 77938
tri 40687 77922 40703 77938 sw
rect 40610 77856 40703 77922
rect 40610 77754 40703 77820
rect 40610 77738 40687 77754
tri 40687 77738 40703 77754 nw
rect 40739 77721 40853 77955
tri 40889 77922 40905 77938 se
rect 40905 77922 40982 77938
rect 40889 77856 40982 77922
rect 40889 77754 40982 77820
tri 40889 77738 40905 77754 ne
rect 40905 77738 40982 77754
rect 40722 77639 40870 77721
rect 40610 77606 40687 77622
tri 40687 77606 40703 77622 sw
rect 40610 77540 40703 77606
rect 40739 77481 40853 77639
tri 40889 77606 40905 77622 se
rect 40905 77606 40982 77622
rect 40889 77540 40982 77606
rect 40610 77405 40982 77481
rect 40610 77280 40703 77346
rect 40610 77264 40687 77280
tri 40687 77264 40703 77280 nw
rect 40739 77247 40853 77405
rect 40889 77280 40982 77346
tri 40889 77264 40905 77280 ne
rect 40905 77264 40982 77280
rect 40722 77165 40870 77247
rect 40610 77132 40687 77148
tri 40687 77132 40703 77148 sw
rect 40610 77066 40703 77132
rect 40610 76964 40703 77030
rect 40610 76948 40687 76964
tri 40687 76948 40703 76964 nw
rect 40739 76931 40853 77165
tri 40889 77132 40905 77148 se
rect 40905 77132 40982 77148
rect 40889 77066 40982 77132
rect 40889 76964 40982 77030
tri 40889 76948 40905 76964 ne
rect 40905 76948 40982 76964
rect 40722 76849 40870 76931
rect 40610 76816 40687 76832
tri 40687 76816 40703 76832 sw
rect 40610 76750 40703 76816
rect 40739 76691 40853 76849
tri 40889 76816 40905 76832 se
rect 40905 76816 40982 76832
rect 40889 76750 40982 76816
rect 40610 76615 40982 76691
rect 40610 76490 40703 76556
rect 40610 76474 40687 76490
tri 40687 76474 40703 76490 nw
rect 40739 76457 40853 76615
rect 40889 76490 40982 76556
tri 40889 76474 40905 76490 ne
rect 40905 76474 40982 76490
rect 40722 76375 40870 76457
rect 40610 76342 40687 76358
tri 40687 76342 40703 76358 sw
rect 40610 76276 40703 76342
rect 40610 76174 40703 76240
rect 40610 76158 40687 76174
tri 40687 76158 40703 76174 nw
rect 40739 76141 40853 76375
tri 40889 76342 40905 76358 se
rect 40905 76342 40982 76358
rect 40889 76276 40982 76342
rect 40889 76174 40982 76240
tri 40889 76158 40905 76174 ne
rect 40905 76158 40982 76174
rect 40722 76059 40870 76141
rect 40610 76026 40687 76042
tri 40687 76026 40703 76042 sw
rect 40610 75960 40703 76026
rect 40739 75901 40853 76059
tri 40889 76026 40905 76042 se
rect 40905 76026 40982 76042
rect 40889 75960 40982 76026
rect 40610 75825 40982 75901
rect 40610 75700 40703 75766
rect 40610 75684 40687 75700
tri 40687 75684 40703 75700 nw
rect 40739 75667 40853 75825
rect 40889 75700 40982 75766
tri 40889 75684 40905 75700 ne
rect 40905 75684 40982 75700
rect 40722 75585 40870 75667
rect 40610 75552 40687 75568
tri 40687 75552 40703 75568 sw
rect 40610 75486 40703 75552
rect 40610 75384 40703 75450
rect 40610 75368 40687 75384
tri 40687 75368 40703 75384 nw
rect 40739 75351 40853 75585
tri 40889 75552 40905 75568 se
rect 40905 75552 40982 75568
rect 40889 75486 40982 75552
rect 40889 75384 40982 75450
tri 40889 75368 40905 75384 ne
rect 40905 75368 40982 75384
rect 40722 75269 40870 75351
rect 40610 75236 40687 75252
tri 40687 75236 40703 75252 sw
rect 40610 75170 40703 75236
rect 40739 75111 40853 75269
tri 40889 75236 40905 75252 se
rect 40905 75236 40982 75252
rect 40889 75170 40982 75236
rect 40610 75035 40982 75111
rect 40610 74910 40703 74976
rect 40610 74894 40687 74910
tri 40687 74894 40703 74910 nw
rect 40739 74877 40853 75035
rect 40889 74910 40982 74976
tri 40889 74894 40905 74910 ne
rect 40905 74894 40982 74910
rect 40722 74795 40870 74877
rect 40610 74762 40687 74778
tri 40687 74762 40703 74778 sw
rect 40610 74696 40703 74762
rect 40610 74594 40703 74660
rect 40610 74578 40687 74594
tri 40687 74578 40703 74594 nw
rect 40739 74561 40853 74795
tri 40889 74762 40905 74778 se
rect 40905 74762 40982 74778
rect 40889 74696 40982 74762
rect 40889 74594 40982 74660
tri 40889 74578 40905 74594 ne
rect 40905 74578 40982 74594
rect 40722 74479 40870 74561
rect 40610 74446 40687 74462
tri 40687 74446 40703 74462 sw
rect 40610 74380 40703 74446
rect 40739 74321 40853 74479
tri 40889 74446 40905 74462 se
rect 40905 74446 40982 74462
rect 40889 74380 40982 74446
rect 40610 74245 40982 74321
rect 40610 74120 40703 74186
rect 40610 74104 40687 74120
tri 40687 74104 40703 74120 nw
rect 40739 74087 40853 74245
rect 40889 74120 40982 74186
tri 40889 74104 40905 74120 ne
rect 40905 74104 40982 74120
rect 40722 74005 40870 74087
rect 40610 73972 40687 73988
tri 40687 73972 40703 73988 sw
rect 40610 73906 40703 73972
rect 40610 73804 40703 73870
rect 40610 73788 40687 73804
tri 40687 73788 40703 73804 nw
rect 40739 73771 40853 74005
tri 40889 73972 40905 73988 se
rect 40905 73972 40982 73988
rect 40889 73906 40982 73972
rect 40889 73804 40982 73870
tri 40889 73788 40905 73804 ne
rect 40905 73788 40982 73804
rect 40722 73689 40870 73771
rect 40610 73656 40687 73672
tri 40687 73656 40703 73672 sw
rect 40610 73590 40703 73656
rect 40739 73531 40853 73689
tri 40889 73656 40905 73672 se
rect 40905 73656 40982 73672
rect 40889 73590 40982 73656
rect 40610 73455 40982 73531
rect 40610 73330 40703 73396
rect 40610 73314 40687 73330
tri 40687 73314 40703 73330 nw
rect 40739 73297 40853 73455
rect 40889 73330 40982 73396
tri 40889 73314 40905 73330 ne
rect 40905 73314 40982 73330
rect 40722 73215 40870 73297
rect 40610 73182 40687 73198
tri 40687 73182 40703 73198 sw
rect 40610 73116 40703 73182
rect 40610 73014 40703 73080
rect 40610 72998 40687 73014
tri 40687 72998 40703 73014 nw
rect 40739 72981 40853 73215
tri 40889 73182 40905 73198 se
rect 40905 73182 40982 73198
rect 40889 73116 40982 73182
rect 40889 73014 40982 73080
tri 40889 72998 40905 73014 ne
rect 40905 72998 40982 73014
rect 40722 72899 40870 72981
rect 40610 72866 40687 72882
tri 40687 72866 40703 72882 sw
rect 40610 72800 40703 72866
rect 40739 72741 40853 72899
tri 40889 72866 40905 72882 se
rect 40905 72866 40982 72882
rect 40889 72800 40982 72866
rect 40610 72665 40982 72741
rect 40610 72540 40703 72606
rect 40610 72524 40687 72540
tri 40687 72524 40703 72540 nw
rect 40739 72507 40853 72665
rect 40889 72540 40982 72606
tri 40889 72524 40905 72540 ne
rect 40905 72524 40982 72540
rect 40722 72425 40870 72507
rect 40610 72392 40687 72408
tri 40687 72392 40703 72408 sw
rect 40610 72326 40703 72392
rect 40610 72224 40703 72290
rect 40610 72208 40687 72224
tri 40687 72208 40703 72224 nw
rect 40739 72191 40853 72425
tri 40889 72392 40905 72408 se
rect 40905 72392 40982 72408
rect 40889 72326 40982 72392
rect 40889 72224 40982 72290
tri 40889 72208 40905 72224 ne
rect 40905 72208 40982 72224
rect 40722 72109 40870 72191
rect 40610 72076 40687 72092
tri 40687 72076 40703 72092 sw
rect 40610 72010 40703 72076
rect 40739 71951 40853 72109
tri 40889 72076 40905 72092 se
rect 40905 72076 40982 72092
rect 40889 72010 40982 72076
rect 40610 71875 40982 71951
rect 40610 71750 40703 71816
rect 40610 71734 40687 71750
tri 40687 71734 40703 71750 nw
rect 40739 71717 40853 71875
rect 40889 71750 40982 71816
tri 40889 71734 40905 71750 ne
rect 40905 71734 40982 71750
rect 40722 71635 40870 71717
rect 40610 71602 40687 71618
tri 40687 71602 40703 71618 sw
rect 40610 71536 40703 71602
rect 40610 71434 40703 71500
rect 40610 71418 40687 71434
tri 40687 71418 40703 71434 nw
rect 40739 71401 40853 71635
tri 40889 71602 40905 71618 se
rect 40905 71602 40982 71618
rect 40889 71536 40982 71602
rect 40889 71434 40982 71500
tri 40889 71418 40905 71434 ne
rect 40905 71418 40982 71434
rect 40722 71319 40870 71401
rect 40610 71286 40687 71302
tri 40687 71286 40703 71302 sw
rect 40610 71220 40703 71286
rect 40739 71161 40853 71319
tri 40889 71286 40905 71302 se
rect 40905 71286 40982 71302
rect 40889 71220 40982 71286
rect 40610 71085 40982 71161
rect 40610 70960 40703 71026
rect 40610 70944 40687 70960
tri 40687 70944 40703 70960 nw
rect 40739 70927 40853 71085
rect 40889 70960 40982 71026
tri 40889 70944 40905 70960 ne
rect 40905 70944 40982 70960
rect 40722 70845 40870 70927
rect 40610 70812 40687 70828
tri 40687 70812 40703 70828 sw
rect 40610 70746 40703 70812
rect 40610 70644 40703 70710
rect 40610 70628 40687 70644
tri 40687 70628 40703 70644 nw
rect 40739 70611 40853 70845
tri 40889 70812 40905 70828 se
rect 40905 70812 40982 70828
rect 40889 70746 40982 70812
rect 40889 70644 40982 70710
tri 40889 70628 40905 70644 ne
rect 40905 70628 40982 70644
rect 40722 70529 40870 70611
rect 40610 70496 40687 70512
tri 40687 70496 40703 70512 sw
rect 40610 70430 40703 70496
rect 40739 70371 40853 70529
tri 40889 70496 40905 70512 se
rect 40905 70496 40982 70512
rect 40889 70430 40982 70496
rect 40610 70295 40982 70371
rect 40610 70170 40703 70236
rect 40610 70154 40687 70170
tri 40687 70154 40703 70170 nw
rect 40739 70137 40853 70295
rect 40889 70170 40982 70236
tri 40889 70154 40905 70170 ne
rect 40905 70154 40982 70170
rect 40722 70055 40870 70137
rect 40610 70022 40687 70038
tri 40687 70022 40703 70038 sw
rect 40610 69956 40703 70022
rect 40610 69854 40703 69920
rect 40610 69838 40687 69854
tri 40687 69838 40703 69854 nw
rect 40739 69821 40853 70055
tri 40889 70022 40905 70038 se
rect 40905 70022 40982 70038
rect 40889 69956 40982 70022
rect 40889 69854 40982 69920
tri 40889 69838 40905 69854 ne
rect 40905 69838 40982 69854
rect 40722 69739 40870 69821
rect 40610 69706 40687 69722
tri 40687 69706 40703 69722 sw
rect 40610 69640 40703 69706
rect 40739 69581 40853 69739
tri 40889 69706 40905 69722 se
rect 40905 69706 40982 69722
rect 40889 69640 40982 69706
rect 40610 69505 40982 69581
rect 40610 69380 40703 69446
rect 40610 69364 40687 69380
tri 40687 69364 40703 69380 nw
rect 40739 69347 40853 69505
rect 40889 69380 40982 69446
tri 40889 69364 40905 69380 ne
rect 40905 69364 40982 69380
rect 40722 69265 40870 69347
rect 40610 69232 40687 69248
tri 40687 69232 40703 69248 sw
rect 40610 69166 40703 69232
rect 40610 69064 40703 69130
rect 40610 69048 40687 69064
tri 40687 69048 40703 69064 nw
rect 40739 69031 40853 69265
tri 40889 69232 40905 69248 se
rect 40905 69232 40982 69248
rect 40889 69166 40982 69232
rect 40889 69064 40982 69130
tri 40889 69048 40905 69064 ne
rect 40905 69048 40982 69064
rect 40722 68949 40870 69031
rect 40610 68916 40687 68932
tri 40687 68916 40703 68932 sw
rect 40610 68850 40703 68916
rect 40739 68791 40853 68949
tri 40889 68916 40905 68932 se
rect 40905 68916 40982 68932
rect 40889 68850 40982 68916
rect 40610 68715 40982 68791
rect 40610 68590 40703 68656
rect 40610 68574 40687 68590
tri 40687 68574 40703 68590 nw
rect 40739 68557 40853 68715
rect 40889 68590 40982 68656
tri 40889 68574 40905 68590 ne
rect 40905 68574 40982 68590
rect 40722 68475 40870 68557
rect 40610 68442 40687 68458
tri 40687 68442 40703 68458 sw
rect 40610 68376 40703 68442
rect 40610 68274 40703 68340
rect 40610 68258 40687 68274
tri 40687 68258 40703 68274 nw
rect 40739 68241 40853 68475
tri 40889 68442 40905 68458 se
rect 40905 68442 40982 68458
rect 40889 68376 40982 68442
rect 40889 68274 40982 68340
tri 40889 68258 40905 68274 ne
rect 40905 68258 40982 68274
rect 40722 68159 40870 68241
rect 40610 68126 40687 68142
tri 40687 68126 40703 68142 sw
rect 40610 68060 40703 68126
rect 40739 68001 40853 68159
tri 40889 68126 40905 68142 se
rect 40905 68126 40982 68142
rect 40889 68060 40982 68126
rect 40610 67925 40982 68001
rect 40610 67800 40703 67866
rect 40610 67784 40687 67800
tri 40687 67784 40703 67800 nw
rect 40739 67767 40853 67925
rect 40889 67800 40982 67866
tri 40889 67784 40905 67800 ne
rect 40905 67784 40982 67800
rect 40722 67685 40870 67767
rect 40610 67652 40687 67668
tri 40687 67652 40703 67668 sw
rect 40610 67586 40703 67652
rect 40610 67484 40703 67550
rect 40610 67468 40687 67484
tri 40687 67468 40703 67484 nw
rect 40739 67451 40853 67685
tri 40889 67652 40905 67668 se
rect 40905 67652 40982 67668
rect 40889 67586 40982 67652
rect 40889 67484 40982 67550
tri 40889 67468 40905 67484 ne
rect 40905 67468 40982 67484
rect 40722 67369 40870 67451
rect 40610 67336 40687 67352
tri 40687 67336 40703 67352 sw
rect 40610 67270 40703 67336
rect 40739 67211 40853 67369
tri 40889 67336 40905 67352 se
rect 40905 67336 40982 67352
rect 40889 67270 40982 67336
rect 40610 67135 40982 67211
rect 40610 67010 40703 67076
rect 40610 66994 40687 67010
tri 40687 66994 40703 67010 nw
rect 40739 66977 40853 67135
rect 40889 67010 40982 67076
tri 40889 66994 40905 67010 ne
rect 40905 66994 40982 67010
rect 40722 66895 40870 66977
rect 40610 66862 40687 66878
tri 40687 66862 40703 66878 sw
rect 40610 66796 40703 66862
rect 40610 66694 40703 66760
rect 40610 66678 40687 66694
tri 40687 66678 40703 66694 nw
rect 40739 66661 40853 66895
tri 40889 66862 40905 66878 se
rect 40905 66862 40982 66878
rect 40889 66796 40982 66862
rect 40889 66694 40982 66760
tri 40889 66678 40905 66694 ne
rect 40905 66678 40982 66694
rect 40722 66579 40870 66661
rect 40610 66546 40687 66562
tri 40687 66546 40703 66562 sw
rect 40610 66480 40703 66546
rect 40739 66421 40853 66579
tri 40889 66546 40905 66562 se
rect 40905 66546 40982 66562
rect 40889 66480 40982 66546
rect 40610 66345 40982 66421
rect 40610 66220 40703 66286
rect 40610 66204 40687 66220
tri 40687 66204 40703 66220 nw
rect 40739 66187 40853 66345
rect 40889 66220 40982 66286
tri 40889 66204 40905 66220 ne
rect 40905 66204 40982 66220
rect 40722 66105 40870 66187
rect 40610 66072 40687 66088
tri 40687 66072 40703 66088 sw
rect 40610 66006 40703 66072
rect 40610 65904 40703 65970
rect 40610 65888 40687 65904
tri 40687 65888 40703 65904 nw
rect 40739 65871 40853 66105
tri 40889 66072 40905 66088 se
rect 40905 66072 40982 66088
rect 40889 66006 40982 66072
rect 40889 65904 40982 65970
tri 40889 65888 40905 65904 ne
rect 40905 65888 40982 65904
rect 40722 65789 40870 65871
rect 40610 65756 40687 65772
tri 40687 65756 40703 65772 sw
rect 40610 65690 40703 65756
rect 40739 65631 40853 65789
tri 40889 65756 40905 65772 se
rect 40905 65756 40982 65772
rect 40889 65690 40982 65756
rect 40610 65555 40982 65631
rect 40610 65430 40703 65496
rect 40610 65414 40687 65430
tri 40687 65414 40703 65430 nw
rect 40739 65397 40853 65555
rect 40889 65430 40982 65496
tri 40889 65414 40905 65430 ne
rect 40905 65414 40982 65430
rect 40722 65315 40870 65397
rect 40610 65282 40687 65298
tri 40687 65282 40703 65298 sw
rect 40610 65216 40703 65282
rect 40610 65114 40703 65180
rect 40610 65098 40687 65114
tri 40687 65098 40703 65114 nw
rect 40739 65081 40853 65315
tri 40889 65282 40905 65298 se
rect 40905 65282 40982 65298
rect 40889 65216 40982 65282
rect 40889 65114 40982 65180
tri 40889 65098 40905 65114 ne
rect 40905 65098 40982 65114
rect 40722 64999 40870 65081
rect 40610 64966 40687 64982
tri 40687 64966 40703 64982 sw
rect 40610 64900 40703 64966
rect 40739 64841 40853 64999
tri 40889 64966 40905 64982 se
rect 40905 64966 40982 64982
rect 40889 64900 40982 64966
rect 40610 64765 40982 64841
rect 40610 64640 40703 64706
rect 40610 64624 40687 64640
tri 40687 64624 40703 64640 nw
rect 40739 64607 40853 64765
rect 40889 64640 40982 64706
tri 40889 64624 40905 64640 ne
rect 40905 64624 40982 64640
rect 40722 64525 40870 64607
rect 40610 64492 40687 64508
tri 40687 64492 40703 64508 sw
rect 40610 64426 40703 64492
rect 40610 64324 40703 64390
rect 40610 64308 40687 64324
tri 40687 64308 40703 64324 nw
rect 40739 64291 40853 64525
tri 40889 64492 40905 64508 se
rect 40905 64492 40982 64508
rect 40889 64426 40982 64492
rect 40889 64324 40982 64390
tri 40889 64308 40905 64324 ne
rect 40905 64308 40982 64324
rect 40722 64209 40870 64291
rect 40610 64176 40687 64192
tri 40687 64176 40703 64192 sw
rect 40610 64110 40703 64176
rect 40739 64051 40853 64209
tri 40889 64176 40905 64192 se
rect 40905 64176 40982 64192
rect 40889 64110 40982 64176
rect 40610 63975 40982 64051
rect 40610 63850 40703 63916
rect 40610 63834 40687 63850
tri 40687 63834 40703 63850 nw
rect 40739 63817 40853 63975
rect 40889 63850 40982 63916
tri 40889 63834 40905 63850 ne
rect 40905 63834 40982 63850
rect 40722 63735 40870 63817
rect 40610 63702 40687 63718
tri 40687 63702 40703 63718 sw
rect 40610 63636 40703 63702
rect 40610 63534 40703 63600
rect 40610 63518 40687 63534
tri 40687 63518 40703 63534 nw
rect 40739 63501 40853 63735
tri 40889 63702 40905 63718 se
rect 40905 63702 40982 63718
rect 40889 63636 40982 63702
rect 40889 63534 40982 63600
tri 40889 63518 40905 63534 ne
rect 40905 63518 40982 63534
rect 40722 63419 40870 63501
rect 40610 63386 40687 63402
tri 40687 63386 40703 63402 sw
rect 40610 63320 40703 63386
rect 40739 63261 40853 63419
tri 40889 63386 40905 63402 se
rect 40905 63386 40982 63402
rect 40889 63320 40982 63386
rect 40610 63185 40982 63261
rect 40610 63060 40703 63126
rect 40610 63044 40687 63060
tri 40687 63044 40703 63060 nw
rect 40739 63027 40853 63185
rect 40889 63060 40982 63126
tri 40889 63044 40905 63060 ne
rect 40905 63044 40982 63060
rect 40722 62945 40870 63027
rect 40610 62912 40687 62928
tri 40687 62912 40703 62928 sw
rect 40610 62846 40703 62912
rect 40610 62744 40703 62810
rect 40610 62728 40687 62744
tri 40687 62728 40703 62744 nw
rect 40739 62711 40853 62945
tri 40889 62912 40905 62928 se
rect 40905 62912 40982 62928
rect 40889 62846 40982 62912
rect 40889 62744 40982 62810
tri 40889 62728 40905 62744 ne
rect 40905 62728 40982 62744
rect 40722 62629 40870 62711
rect 40610 62596 40687 62612
tri 40687 62596 40703 62612 sw
rect 40610 62530 40703 62596
rect 40739 62471 40853 62629
tri 40889 62596 40905 62612 se
rect 40905 62596 40982 62612
rect 40889 62530 40982 62596
rect 40610 62395 40982 62471
rect 40610 62270 40703 62336
rect 40610 62254 40687 62270
tri 40687 62254 40703 62270 nw
rect 40739 62237 40853 62395
rect 40889 62270 40982 62336
tri 40889 62254 40905 62270 ne
rect 40905 62254 40982 62270
rect 40722 62155 40870 62237
rect 40610 62122 40687 62138
tri 40687 62122 40703 62138 sw
rect 40610 62056 40703 62122
rect 40610 61954 40703 62020
rect 40610 61938 40687 61954
tri 40687 61938 40703 61954 nw
rect 40739 61921 40853 62155
tri 40889 62122 40905 62138 se
rect 40905 62122 40982 62138
rect 40889 62056 40982 62122
rect 40889 61954 40982 62020
tri 40889 61938 40905 61954 ne
rect 40905 61938 40982 61954
rect 40722 61839 40870 61921
rect 40610 61806 40687 61822
tri 40687 61806 40703 61822 sw
rect 40610 61740 40703 61806
rect 40739 61681 40853 61839
tri 40889 61806 40905 61822 se
rect 40905 61806 40982 61822
rect 40889 61740 40982 61806
rect 40610 61605 40982 61681
rect 40610 61480 40703 61546
rect 40610 61464 40687 61480
tri 40687 61464 40703 61480 nw
rect 40739 61447 40853 61605
rect 40889 61480 40982 61546
tri 40889 61464 40905 61480 ne
rect 40905 61464 40982 61480
rect 40722 61365 40870 61447
rect 40610 61332 40687 61348
tri 40687 61332 40703 61348 sw
rect 40610 61266 40703 61332
rect 40610 61164 40703 61230
rect 40610 61148 40687 61164
tri 40687 61148 40703 61164 nw
rect 40739 61131 40853 61365
tri 40889 61332 40905 61348 se
rect 40905 61332 40982 61348
rect 40889 61266 40982 61332
rect 40889 61164 40982 61230
tri 40889 61148 40905 61164 ne
rect 40905 61148 40982 61164
rect 40722 61049 40870 61131
rect 40610 61016 40687 61032
tri 40687 61016 40703 61032 sw
rect 40610 60950 40703 61016
rect 40739 60891 40853 61049
tri 40889 61016 40905 61032 se
rect 40905 61016 40982 61032
rect 40889 60950 40982 61016
rect 40610 60815 40982 60891
rect 40610 60690 40703 60756
rect 40610 60674 40687 60690
tri 40687 60674 40703 60690 nw
rect 40739 60657 40853 60815
rect 40889 60690 40982 60756
tri 40889 60674 40905 60690 ne
rect 40905 60674 40982 60690
rect 40722 60575 40870 60657
rect 40610 60542 40687 60558
tri 40687 60542 40703 60558 sw
rect 40610 60476 40703 60542
rect 40610 60374 40703 60440
rect 40610 60358 40687 60374
tri 40687 60358 40703 60374 nw
rect 40739 60341 40853 60575
tri 40889 60542 40905 60558 se
rect 40905 60542 40982 60558
rect 40889 60476 40982 60542
rect 40889 60374 40982 60440
tri 40889 60358 40905 60374 ne
rect 40905 60358 40982 60374
rect 40722 60259 40870 60341
rect 40610 60226 40687 60242
tri 40687 60226 40703 60242 sw
rect 40610 60160 40703 60226
rect 40739 60101 40853 60259
tri 40889 60226 40905 60242 se
rect 40905 60226 40982 60242
rect 40889 60160 40982 60226
rect 40610 60025 40982 60101
rect 40610 59900 40703 59966
rect 40610 59884 40687 59900
tri 40687 59884 40703 59900 nw
rect 40739 59867 40853 60025
rect 40889 59900 40982 59966
tri 40889 59884 40905 59900 ne
rect 40905 59884 40982 59900
rect 40722 59785 40870 59867
rect 40610 59752 40687 59768
tri 40687 59752 40703 59768 sw
rect 40610 59686 40703 59752
rect 40610 59584 40703 59650
rect 40610 59568 40687 59584
tri 40687 59568 40703 59584 nw
rect 40739 59551 40853 59785
tri 40889 59752 40905 59768 se
rect 40905 59752 40982 59768
rect 40889 59686 40982 59752
rect 40889 59584 40982 59650
tri 40889 59568 40905 59584 ne
rect 40905 59568 40982 59584
rect 40722 59469 40870 59551
rect 40610 59436 40687 59452
tri 40687 59436 40703 59452 sw
rect 40610 59370 40703 59436
rect 40739 59311 40853 59469
tri 40889 59436 40905 59452 se
rect 40905 59436 40982 59452
rect 40889 59370 40982 59436
rect 40610 59235 40982 59311
rect 40610 59110 40703 59176
rect 40610 59094 40687 59110
tri 40687 59094 40703 59110 nw
rect 40739 59077 40853 59235
rect 40889 59110 40982 59176
tri 40889 59094 40905 59110 ne
rect 40905 59094 40982 59110
rect 40722 58995 40870 59077
rect 40610 58962 40687 58978
tri 40687 58962 40703 58978 sw
rect 40610 58896 40703 58962
rect 40610 58794 40703 58860
rect 40610 58778 40687 58794
tri 40687 58778 40703 58794 nw
rect 40739 58761 40853 58995
tri 40889 58962 40905 58978 se
rect 40905 58962 40982 58978
rect 40889 58896 40982 58962
rect 40889 58794 40982 58860
tri 40889 58778 40905 58794 ne
rect 40905 58778 40982 58794
rect 40722 58679 40870 58761
rect 40610 58646 40687 58662
tri 40687 58646 40703 58662 sw
rect 40610 58580 40703 58646
rect 40739 58521 40853 58679
tri 40889 58646 40905 58662 se
rect 40905 58646 40982 58662
rect 40889 58580 40982 58646
rect 40610 58445 40982 58521
rect 40610 58320 40703 58386
rect 40610 58304 40687 58320
tri 40687 58304 40703 58320 nw
rect 40739 58287 40853 58445
rect 40889 58320 40982 58386
tri 40889 58304 40905 58320 ne
rect 40905 58304 40982 58320
rect 40722 58205 40870 58287
rect 40610 58172 40687 58188
tri 40687 58172 40703 58188 sw
rect 40610 58106 40703 58172
rect 40610 58004 40703 58070
rect 40610 57988 40687 58004
tri 40687 57988 40703 58004 nw
rect 40739 57971 40853 58205
tri 40889 58172 40905 58188 se
rect 40905 58172 40982 58188
rect 40889 58106 40982 58172
rect 40889 58004 40982 58070
tri 40889 57988 40905 58004 ne
rect 40905 57988 40982 58004
rect 40722 57889 40870 57971
rect 40610 57856 40687 57872
tri 40687 57856 40703 57872 sw
rect 40610 57790 40703 57856
rect 40739 57731 40853 57889
tri 40889 57856 40905 57872 se
rect 40905 57856 40982 57872
rect 40889 57790 40982 57856
rect 40610 57655 40982 57731
rect 40610 57530 40703 57596
rect 40610 57514 40687 57530
tri 40687 57514 40703 57530 nw
rect 40739 57497 40853 57655
rect 40889 57530 40982 57596
tri 40889 57514 40905 57530 ne
rect 40905 57514 40982 57530
rect 40722 57415 40870 57497
rect 40610 57382 40687 57398
tri 40687 57382 40703 57398 sw
rect 40610 57316 40703 57382
rect 40610 57214 40703 57280
rect 40610 57198 40687 57214
tri 40687 57198 40703 57214 nw
rect 40739 57181 40853 57415
tri 40889 57382 40905 57398 se
rect 40905 57382 40982 57398
rect 40889 57316 40982 57382
rect 40889 57214 40982 57280
tri 40889 57198 40905 57214 ne
rect 40905 57198 40982 57214
rect 40722 57099 40870 57181
rect 40610 57066 40687 57082
tri 40687 57066 40703 57082 sw
rect 40610 57000 40703 57066
rect 40739 56941 40853 57099
tri 40889 57066 40905 57082 se
rect 40905 57066 40982 57082
rect 40889 57000 40982 57066
rect 40610 56865 40982 56941
rect 40610 56740 40703 56806
rect 40610 56724 40687 56740
tri 40687 56724 40703 56740 nw
rect 40739 56707 40853 56865
rect 40889 56740 40982 56806
tri 40889 56724 40905 56740 ne
rect 40905 56724 40982 56740
rect 40722 56625 40870 56707
rect 40610 56592 40687 56608
tri 40687 56592 40703 56608 sw
rect 40610 56526 40703 56592
rect 40610 56424 40703 56490
rect 40610 56408 40687 56424
tri 40687 56408 40703 56424 nw
rect 40739 56391 40853 56625
tri 40889 56592 40905 56608 se
rect 40905 56592 40982 56608
rect 40889 56526 40982 56592
rect 40889 56424 40982 56490
tri 40889 56408 40905 56424 ne
rect 40905 56408 40982 56424
rect 40722 56309 40870 56391
rect 40610 56276 40687 56292
tri 40687 56276 40703 56292 sw
rect 40610 56210 40703 56276
rect 40739 56151 40853 56309
tri 40889 56276 40905 56292 se
rect 40905 56276 40982 56292
rect 40889 56210 40982 56276
rect 40610 56075 40982 56151
rect 40610 55950 40703 56016
rect 40610 55934 40687 55950
tri 40687 55934 40703 55950 nw
rect 40739 55917 40853 56075
rect 40889 55950 40982 56016
tri 40889 55934 40905 55950 ne
rect 40905 55934 40982 55950
rect 40722 55835 40870 55917
rect 40610 55802 40687 55818
tri 40687 55802 40703 55818 sw
rect 40610 55736 40703 55802
rect 40610 55634 40703 55700
rect 40610 55618 40687 55634
tri 40687 55618 40703 55634 nw
rect 40739 55601 40853 55835
tri 40889 55802 40905 55818 se
rect 40905 55802 40982 55818
rect 40889 55736 40982 55802
rect 40889 55634 40982 55700
tri 40889 55618 40905 55634 ne
rect 40905 55618 40982 55634
rect 40722 55519 40870 55601
rect 40610 55486 40687 55502
tri 40687 55486 40703 55502 sw
rect 40610 55420 40703 55486
rect 40739 55361 40853 55519
tri 40889 55486 40905 55502 se
rect 40905 55486 40982 55502
rect 40889 55420 40982 55486
rect 40610 55285 40982 55361
rect 40610 55160 40703 55226
rect 40610 55144 40687 55160
tri 40687 55144 40703 55160 nw
rect 40739 55127 40853 55285
rect 40889 55160 40982 55226
tri 40889 55144 40905 55160 ne
rect 40905 55144 40982 55160
rect 40722 55045 40870 55127
rect 40610 55012 40687 55028
tri 40687 55012 40703 55028 sw
rect 40610 54946 40703 55012
rect 40610 54844 40703 54910
rect 40610 54828 40687 54844
tri 40687 54828 40703 54844 nw
rect 40739 54811 40853 55045
tri 40889 55012 40905 55028 se
rect 40905 55012 40982 55028
rect 40889 54946 40982 55012
rect 40889 54844 40982 54910
tri 40889 54828 40905 54844 ne
rect 40905 54828 40982 54844
rect 40722 54729 40870 54811
rect 40610 54696 40687 54712
tri 40687 54696 40703 54712 sw
rect 40610 54630 40703 54696
rect 40739 54571 40853 54729
tri 40889 54696 40905 54712 se
rect 40905 54696 40982 54712
rect 40889 54630 40982 54696
rect 40610 54495 40982 54571
rect 40610 54370 40703 54436
rect 40610 54354 40687 54370
tri 40687 54354 40703 54370 nw
rect 40739 54337 40853 54495
rect 40889 54370 40982 54436
tri 40889 54354 40905 54370 ne
rect 40905 54354 40982 54370
rect 40722 54255 40870 54337
rect 40610 54222 40687 54238
tri 40687 54222 40703 54238 sw
rect 40610 54156 40703 54222
rect 40610 54054 40703 54120
rect 40610 54038 40687 54054
tri 40687 54038 40703 54054 nw
rect 40739 54021 40853 54255
tri 40889 54222 40905 54238 se
rect 40905 54222 40982 54238
rect 40889 54156 40982 54222
rect 40889 54054 40982 54120
tri 40889 54038 40905 54054 ne
rect 40905 54038 40982 54054
rect 40722 53939 40870 54021
rect 40610 53906 40687 53922
tri 40687 53906 40703 53922 sw
rect 40610 53840 40703 53906
rect 40739 53781 40853 53939
tri 40889 53906 40905 53922 se
rect 40905 53906 40982 53922
rect 40889 53840 40982 53906
rect 40610 53705 40982 53781
rect 40610 53580 40703 53646
rect 40610 53564 40687 53580
tri 40687 53564 40703 53580 nw
rect 40739 53547 40853 53705
rect 40889 53580 40982 53646
tri 40889 53564 40905 53580 ne
rect 40905 53564 40982 53580
rect 40722 53465 40870 53547
rect 40610 53432 40687 53448
tri 40687 53432 40703 53448 sw
rect 40610 53366 40703 53432
rect 40610 53264 40703 53330
rect 40610 53248 40687 53264
tri 40687 53248 40703 53264 nw
rect 40739 53231 40853 53465
tri 40889 53432 40905 53448 se
rect 40905 53432 40982 53448
rect 40889 53366 40982 53432
rect 40889 53264 40982 53330
tri 40889 53248 40905 53264 ne
rect 40905 53248 40982 53264
rect 40722 53149 40870 53231
rect 40610 53116 40687 53132
tri 40687 53116 40703 53132 sw
rect 40610 53050 40703 53116
rect 40739 52991 40853 53149
tri 40889 53116 40905 53132 se
rect 40905 53116 40982 53132
rect 40889 53050 40982 53116
rect 40610 52915 40982 52991
rect 40610 52790 40703 52856
rect 40610 52774 40687 52790
tri 40687 52774 40703 52790 nw
rect 40739 52757 40853 52915
rect 40889 52790 40982 52856
tri 40889 52774 40905 52790 ne
rect 40905 52774 40982 52790
rect 40722 52675 40870 52757
rect 40610 52642 40687 52658
tri 40687 52642 40703 52658 sw
rect 40610 52576 40703 52642
rect 40610 52474 40703 52540
rect 40610 52458 40687 52474
tri 40687 52458 40703 52474 nw
rect 40739 52441 40853 52675
tri 40889 52642 40905 52658 se
rect 40905 52642 40982 52658
rect 40889 52576 40982 52642
rect 40889 52474 40982 52540
tri 40889 52458 40905 52474 ne
rect 40905 52458 40982 52474
rect 40722 52359 40870 52441
rect 40610 52326 40687 52342
tri 40687 52326 40703 52342 sw
rect 40610 52260 40703 52326
rect 40739 52201 40853 52359
tri 40889 52326 40905 52342 se
rect 40905 52326 40982 52342
rect 40889 52260 40982 52326
rect 40610 52125 40982 52201
rect 40610 52000 40703 52066
rect 40610 51984 40687 52000
tri 40687 51984 40703 52000 nw
rect 40739 51967 40853 52125
rect 40889 52000 40982 52066
tri 40889 51984 40905 52000 ne
rect 40905 51984 40982 52000
rect 40722 51885 40870 51967
rect 40610 51852 40687 51868
tri 40687 51852 40703 51868 sw
rect 40610 51786 40703 51852
rect 40610 51684 40703 51750
rect 40610 51668 40687 51684
tri 40687 51668 40703 51684 nw
rect 40739 51651 40853 51885
tri 40889 51852 40905 51868 se
rect 40905 51852 40982 51868
rect 40889 51786 40982 51852
rect 40889 51684 40982 51750
tri 40889 51668 40905 51684 ne
rect 40905 51668 40982 51684
rect 40722 51569 40870 51651
rect 40610 51536 40687 51552
tri 40687 51536 40703 51552 sw
rect 40610 51470 40703 51536
rect 40739 51411 40853 51569
tri 40889 51536 40905 51552 se
rect 40905 51536 40982 51552
rect 40889 51470 40982 51536
rect 40610 51335 40982 51411
rect 40610 51210 40703 51276
rect 40610 51194 40687 51210
tri 40687 51194 40703 51210 nw
rect 40739 51177 40853 51335
rect 40889 51210 40982 51276
tri 40889 51194 40905 51210 ne
rect 40905 51194 40982 51210
rect 40722 51095 40870 51177
rect 40610 51062 40687 51078
tri 40687 51062 40703 51078 sw
rect 40610 50996 40703 51062
rect 40610 50894 40703 50960
rect 40610 50878 40687 50894
tri 40687 50878 40703 50894 nw
rect 40739 50861 40853 51095
tri 40889 51062 40905 51078 se
rect 40905 51062 40982 51078
rect 40889 50996 40982 51062
rect 40889 50894 40982 50960
tri 40889 50878 40905 50894 ne
rect 40905 50878 40982 50894
rect 40722 50779 40870 50861
rect 40610 50746 40687 50762
tri 40687 50746 40703 50762 sw
rect 40610 50680 40703 50746
rect 40739 50621 40853 50779
tri 40889 50746 40905 50762 se
rect 40905 50746 40982 50762
rect 40889 50680 40982 50746
rect 40610 50545 40982 50621
rect 40610 50420 40703 50486
rect 40610 50404 40687 50420
tri 40687 50404 40703 50420 nw
rect 40739 50387 40853 50545
rect 40889 50420 40982 50486
tri 40889 50404 40905 50420 ne
rect 40905 50404 40982 50420
rect 40722 50305 40870 50387
rect 40610 50272 40687 50288
tri 40687 50272 40703 50288 sw
rect 40610 50206 40703 50272
rect 40610 50104 40703 50170
rect 40610 50088 40687 50104
tri 40687 50088 40703 50104 nw
rect 40739 50071 40853 50305
tri 40889 50272 40905 50288 se
rect 40905 50272 40982 50288
rect 40889 50206 40982 50272
rect 40889 50104 40982 50170
tri 40889 50088 40905 50104 ne
rect 40905 50088 40982 50104
rect 40722 49989 40870 50071
rect 40610 49956 40687 49972
tri 40687 49956 40703 49972 sw
rect 40610 49890 40703 49956
rect 40739 49831 40853 49989
tri 40889 49956 40905 49972 se
rect 40905 49956 40982 49972
rect 40889 49890 40982 49956
rect 40610 49755 40982 49831
rect 40610 49630 40703 49696
rect 40610 49614 40687 49630
tri 40687 49614 40703 49630 nw
rect 40739 49597 40853 49755
rect 40889 49630 40982 49696
tri 40889 49614 40905 49630 ne
rect 40905 49614 40982 49630
rect 40722 49515 40870 49597
rect 40610 49482 40687 49498
tri 40687 49482 40703 49498 sw
rect 40610 49416 40703 49482
rect 40610 49314 40703 49380
rect 40610 49298 40687 49314
tri 40687 49298 40703 49314 nw
rect 40739 49281 40853 49515
tri 40889 49482 40905 49498 se
rect 40905 49482 40982 49498
rect 40889 49416 40982 49482
rect 40889 49314 40982 49380
tri 40889 49298 40905 49314 ne
rect 40905 49298 40982 49314
rect 40722 49199 40870 49281
rect 40610 49166 40687 49182
tri 40687 49166 40703 49182 sw
rect 40610 49100 40703 49166
rect 40739 49041 40853 49199
tri 40889 49166 40905 49182 se
rect 40905 49166 40982 49182
rect 40889 49100 40982 49166
rect 40610 48965 40982 49041
rect 40610 48840 40703 48906
rect 40610 48824 40687 48840
tri 40687 48824 40703 48840 nw
rect 40739 48807 40853 48965
rect 40889 48840 40982 48906
tri 40889 48824 40905 48840 ne
rect 40905 48824 40982 48840
rect 40722 48725 40870 48807
rect 40610 48692 40687 48708
tri 40687 48692 40703 48708 sw
rect 40610 48626 40703 48692
rect 40610 48524 40703 48590
rect 40610 48508 40687 48524
tri 40687 48508 40703 48524 nw
rect 40739 48491 40853 48725
tri 40889 48692 40905 48708 se
rect 40905 48692 40982 48708
rect 40889 48626 40982 48692
rect 40889 48524 40982 48590
tri 40889 48508 40905 48524 ne
rect 40905 48508 40982 48524
rect 40722 48409 40870 48491
rect 40610 48376 40687 48392
tri 40687 48376 40703 48392 sw
rect 40610 48310 40703 48376
rect 40739 48251 40853 48409
tri 40889 48376 40905 48392 se
rect 40905 48376 40982 48392
rect 40889 48310 40982 48376
rect 40610 48175 40982 48251
rect 40610 48050 40703 48116
rect 40610 48034 40687 48050
tri 40687 48034 40703 48050 nw
rect 40739 48017 40853 48175
rect 40889 48050 40982 48116
tri 40889 48034 40905 48050 ne
rect 40905 48034 40982 48050
rect 40722 47935 40870 48017
rect 40610 47902 40687 47918
tri 40687 47902 40703 47918 sw
rect 40610 47836 40703 47902
rect 40610 47734 40703 47800
rect 40610 47718 40687 47734
tri 40687 47718 40703 47734 nw
rect 40739 47701 40853 47935
tri 40889 47902 40905 47918 se
rect 40905 47902 40982 47918
rect 40889 47836 40982 47902
rect 40889 47734 40982 47800
tri 40889 47718 40905 47734 ne
rect 40905 47718 40982 47734
rect 40722 47619 40870 47701
rect 40610 47586 40687 47602
tri 40687 47586 40703 47602 sw
rect 40610 47520 40703 47586
rect 40739 47461 40853 47619
tri 40889 47586 40905 47602 se
rect 40905 47586 40982 47602
rect 40889 47520 40982 47586
rect 40610 47385 40982 47461
rect 40610 47260 40703 47326
rect 40610 47244 40687 47260
tri 40687 47244 40703 47260 nw
rect 40739 47227 40853 47385
rect 40889 47260 40982 47326
tri 40889 47244 40905 47260 ne
rect 40905 47244 40982 47260
rect 40722 47145 40870 47227
rect 40610 47112 40687 47128
tri 40687 47112 40703 47128 sw
rect 40610 47046 40703 47112
rect 40610 46944 40703 47010
rect 40610 46928 40687 46944
tri 40687 46928 40703 46944 nw
rect 40739 46911 40853 47145
tri 40889 47112 40905 47128 se
rect 40905 47112 40982 47128
rect 40889 47046 40982 47112
rect 40889 46944 40982 47010
tri 40889 46928 40905 46944 ne
rect 40905 46928 40982 46944
rect 40722 46829 40870 46911
rect 40610 46796 40687 46812
tri 40687 46796 40703 46812 sw
rect 40610 46730 40703 46796
rect 40739 46671 40853 46829
tri 40889 46796 40905 46812 se
rect 40905 46796 40982 46812
rect 40889 46730 40982 46796
rect 40610 46595 40982 46671
rect 40610 46470 40703 46536
rect 40610 46454 40687 46470
tri 40687 46454 40703 46470 nw
rect 40739 46437 40853 46595
rect 40889 46470 40982 46536
tri 40889 46454 40905 46470 ne
rect 40905 46454 40982 46470
rect 40722 46355 40870 46437
rect 40610 46322 40687 46338
tri 40687 46322 40703 46338 sw
rect 40610 46256 40703 46322
rect 40610 46154 40703 46220
rect 40610 46138 40687 46154
tri 40687 46138 40703 46154 nw
rect 40739 46121 40853 46355
tri 40889 46322 40905 46338 se
rect 40905 46322 40982 46338
rect 40889 46256 40982 46322
rect 40889 46154 40982 46220
tri 40889 46138 40905 46154 ne
rect 40905 46138 40982 46154
rect 40722 46039 40870 46121
rect 40610 46006 40687 46022
tri 40687 46006 40703 46022 sw
rect 40610 45940 40703 46006
rect 40739 45881 40853 46039
tri 40889 46006 40905 46022 se
rect 40905 46006 40982 46022
rect 40889 45940 40982 46006
rect 40610 45805 40982 45881
rect 40610 45680 40703 45746
rect 40610 45664 40687 45680
tri 40687 45664 40703 45680 nw
rect 40739 45647 40853 45805
rect 40889 45680 40982 45746
tri 40889 45664 40905 45680 ne
rect 40905 45664 40982 45680
rect 40722 45565 40870 45647
rect 40610 45532 40687 45548
tri 40687 45532 40703 45548 sw
rect 40610 45466 40703 45532
rect 40610 45364 40703 45430
rect 40610 45348 40687 45364
tri 40687 45348 40703 45364 nw
rect 40739 45331 40853 45565
tri 40889 45532 40905 45548 se
rect 40905 45532 40982 45548
rect 40889 45466 40982 45532
rect 40889 45364 40982 45430
tri 40889 45348 40905 45364 ne
rect 40905 45348 40982 45364
rect 40722 45249 40870 45331
rect 40610 45216 40687 45232
tri 40687 45216 40703 45232 sw
rect 40610 45150 40703 45216
rect 40739 45091 40853 45249
tri 40889 45216 40905 45232 se
rect 40905 45216 40982 45232
rect 40889 45150 40982 45216
rect 40610 45015 40982 45091
rect 40610 44890 40703 44956
rect 40610 44874 40687 44890
tri 40687 44874 40703 44890 nw
rect 40739 44857 40853 45015
rect 40889 44890 40982 44956
tri 40889 44874 40905 44890 ne
rect 40905 44874 40982 44890
rect 40722 44775 40870 44857
rect 40610 44742 40687 44758
tri 40687 44742 40703 44758 sw
rect 40610 44676 40703 44742
rect 40610 44574 40703 44640
rect 40610 44558 40687 44574
tri 40687 44558 40703 44574 nw
rect 40739 44541 40853 44775
tri 40889 44742 40905 44758 se
rect 40905 44742 40982 44758
rect 40889 44676 40982 44742
rect 40889 44574 40982 44640
tri 40889 44558 40905 44574 ne
rect 40905 44558 40982 44574
rect 40722 44459 40870 44541
rect 40610 44426 40687 44442
tri 40687 44426 40703 44442 sw
rect 40610 44360 40703 44426
rect 40739 44301 40853 44459
tri 40889 44426 40905 44442 se
rect 40905 44426 40982 44442
rect 40889 44360 40982 44426
rect 40610 44225 40982 44301
rect 40610 44100 40703 44166
rect 40610 44084 40687 44100
tri 40687 44084 40703 44100 nw
rect 40739 44067 40853 44225
rect 40889 44100 40982 44166
tri 40889 44084 40905 44100 ne
rect 40905 44084 40982 44100
rect 40722 43985 40870 44067
rect 40610 43952 40687 43968
tri 40687 43952 40703 43968 sw
rect 40610 43886 40703 43952
rect 40610 43784 40703 43850
rect 40610 43768 40687 43784
tri 40687 43768 40703 43784 nw
rect 40739 43751 40853 43985
tri 40889 43952 40905 43968 se
rect 40905 43952 40982 43968
rect 40889 43886 40982 43952
rect 40889 43784 40982 43850
tri 40889 43768 40905 43784 ne
rect 40905 43768 40982 43784
rect 40722 43669 40870 43751
rect 40610 43636 40687 43652
tri 40687 43636 40703 43652 sw
rect 40610 43570 40703 43636
rect 40739 43511 40853 43669
tri 40889 43636 40905 43652 se
rect 40905 43636 40982 43652
rect 40889 43570 40982 43636
rect 40610 43435 40982 43511
rect 40610 43310 40703 43376
rect 40610 43294 40687 43310
tri 40687 43294 40703 43310 nw
rect 40739 43277 40853 43435
rect 40889 43310 40982 43376
tri 40889 43294 40905 43310 ne
rect 40905 43294 40982 43310
rect 40722 43195 40870 43277
rect 40610 43162 40687 43178
tri 40687 43162 40703 43178 sw
rect 40610 43096 40703 43162
rect 40610 42994 40703 43060
rect 40610 42978 40687 42994
tri 40687 42978 40703 42994 nw
rect 40739 42961 40853 43195
tri 40889 43162 40905 43178 se
rect 40905 43162 40982 43178
rect 40889 43096 40982 43162
rect 40889 42994 40982 43060
tri 40889 42978 40905 42994 ne
rect 40905 42978 40982 42994
rect 40722 42879 40870 42961
rect 40610 42846 40687 42862
tri 40687 42846 40703 42862 sw
rect 40610 42780 40703 42846
rect 40739 42721 40853 42879
tri 40889 42846 40905 42862 se
rect 40905 42846 40982 42862
rect 40889 42780 40982 42846
rect 40610 42645 40982 42721
rect 40610 42520 40703 42586
rect 40610 42504 40687 42520
tri 40687 42504 40703 42520 nw
rect 40739 42487 40853 42645
rect 40889 42520 40982 42586
tri 40889 42504 40905 42520 ne
rect 40905 42504 40982 42520
rect 40722 42405 40870 42487
rect 40610 42372 40687 42388
tri 40687 42372 40703 42388 sw
rect 40610 42306 40703 42372
rect 40610 42204 40703 42270
rect 40610 42188 40687 42204
tri 40687 42188 40703 42204 nw
rect 40739 42171 40853 42405
tri 40889 42372 40905 42388 se
rect 40905 42372 40982 42388
rect 40889 42306 40982 42372
rect 40889 42204 40982 42270
tri 40889 42188 40905 42204 ne
rect 40905 42188 40982 42204
rect 40722 42089 40870 42171
rect 40610 42056 40687 42072
tri 40687 42056 40703 42072 sw
rect 40610 41990 40703 42056
rect 40739 41931 40853 42089
tri 40889 42056 40905 42072 se
rect 40905 42056 40982 42072
rect 40889 41990 40982 42056
rect 40610 41855 40982 41931
rect 40610 41730 40703 41796
rect 40610 41714 40687 41730
tri 40687 41714 40703 41730 nw
rect 40739 41697 40853 41855
rect 40889 41730 40982 41796
tri 40889 41714 40905 41730 ne
rect 40905 41714 40982 41730
rect 40722 41615 40870 41697
rect 40610 41582 40687 41598
tri 40687 41582 40703 41598 sw
rect 40610 41516 40703 41582
rect 40610 41414 40703 41480
rect 40610 41398 40687 41414
tri 40687 41398 40703 41414 nw
rect 40739 41381 40853 41615
tri 40889 41582 40905 41598 se
rect 40905 41582 40982 41598
rect 40889 41516 40982 41582
rect 40889 41414 40982 41480
tri 40889 41398 40905 41414 ne
rect 40905 41398 40982 41414
rect 40722 41299 40870 41381
rect 40610 41266 40687 41282
tri 40687 41266 40703 41282 sw
rect 40610 41200 40703 41266
rect 40739 41141 40853 41299
tri 40889 41266 40905 41282 se
rect 40905 41266 40982 41282
rect 40889 41200 40982 41266
rect 40610 41065 40982 41141
rect 40610 40940 40703 41006
rect 40610 40924 40687 40940
tri 40687 40924 40703 40940 nw
rect 40739 40907 40853 41065
rect 40889 40940 40982 41006
tri 40889 40924 40905 40940 ne
rect 40905 40924 40982 40940
rect 40722 40825 40870 40907
rect 40610 40792 40687 40808
tri 40687 40792 40703 40808 sw
rect 40610 40726 40703 40792
rect 40610 40624 40703 40690
rect 40610 40608 40687 40624
tri 40687 40608 40703 40624 nw
rect 40739 40591 40853 40825
tri 40889 40792 40905 40808 se
rect 40905 40792 40982 40808
rect 40889 40726 40982 40792
rect 40889 40624 40982 40690
tri 40889 40608 40905 40624 ne
rect 40905 40608 40982 40624
rect 40722 40509 40870 40591
rect 40610 40476 40687 40492
tri 40687 40476 40703 40492 sw
rect 40610 40410 40703 40476
rect 40739 40351 40853 40509
tri 40889 40476 40905 40492 se
rect 40905 40476 40982 40492
rect 40889 40410 40982 40476
rect 40610 40275 40982 40351
rect 40610 40150 40703 40216
rect 40610 40134 40687 40150
tri 40687 40134 40703 40150 nw
rect 40739 40117 40853 40275
rect 40889 40150 40982 40216
tri 40889 40134 40905 40150 ne
rect 40905 40134 40982 40150
rect 40722 40035 40870 40117
rect 40610 40002 40687 40018
tri 40687 40002 40703 40018 sw
rect 40610 39936 40703 40002
rect 40610 39834 40703 39900
rect 40610 39818 40687 39834
tri 40687 39818 40703 39834 nw
rect 40739 39801 40853 40035
tri 40889 40002 40905 40018 se
rect 40905 40002 40982 40018
rect 40889 39936 40982 40002
rect 40889 39834 40982 39900
tri 40889 39818 40905 39834 ne
rect 40905 39818 40982 39834
rect 40722 39719 40870 39801
rect 40610 39686 40687 39702
tri 40687 39686 40703 39702 sw
rect 40610 39620 40703 39686
rect 40739 39561 40853 39719
tri 40889 39686 40905 39702 se
rect 40905 39686 40982 39702
rect 40889 39620 40982 39686
rect 40610 39485 40982 39561
rect 40610 39360 40703 39426
rect 40610 39344 40687 39360
tri 40687 39344 40703 39360 nw
rect 40739 39327 40853 39485
rect 40889 39360 40982 39426
tri 40889 39344 40905 39360 ne
rect 40905 39344 40982 39360
rect 40722 39245 40870 39327
rect 40610 39212 40687 39228
tri 40687 39212 40703 39228 sw
rect 40610 39146 40703 39212
rect 40610 39044 40703 39110
rect 40610 39028 40687 39044
tri 40687 39028 40703 39044 nw
rect 40739 39011 40853 39245
tri 40889 39212 40905 39228 se
rect 40905 39212 40982 39228
rect 40889 39146 40982 39212
rect 40889 39044 40982 39110
tri 40889 39028 40905 39044 ne
rect 40905 39028 40982 39044
rect 40722 38929 40870 39011
rect 40610 38896 40687 38912
tri 40687 38896 40703 38912 sw
rect 40610 38830 40703 38896
rect 40739 38771 40853 38929
tri 40889 38896 40905 38912 se
rect 40905 38896 40982 38912
rect 40889 38830 40982 38896
rect 40610 38695 40982 38771
rect 40610 38570 40703 38636
rect 40610 38554 40687 38570
tri 40687 38554 40703 38570 nw
rect 40739 38537 40853 38695
rect 40889 38570 40982 38636
tri 40889 38554 40905 38570 ne
rect 40905 38554 40982 38570
rect 40722 38455 40870 38537
rect 40610 38422 40687 38438
tri 40687 38422 40703 38438 sw
rect 40610 38356 40703 38422
rect 40610 38254 40703 38320
rect 40610 38238 40687 38254
tri 40687 38238 40703 38254 nw
rect 40739 38221 40853 38455
tri 40889 38422 40905 38438 se
rect 40905 38422 40982 38438
rect 40889 38356 40982 38422
rect 40889 38254 40982 38320
tri 40889 38238 40905 38254 ne
rect 40905 38238 40982 38254
rect 40722 38139 40870 38221
rect 40610 38106 40687 38122
tri 40687 38106 40703 38122 sw
rect 40610 38040 40703 38106
rect 40739 37981 40853 38139
tri 40889 38106 40905 38122 se
rect 40905 38106 40982 38122
rect 40889 38040 40982 38106
rect 40610 37905 40982 37981
rect 40610 37780 40703 37846
rect 40610 37764 40687 37780
tri 40687 37764 40703 37780 nw
rect 40739 37747 40853 37905
rect 40889 37780 40982 37846
tri 40889 37764 40905 37780 ne
rect 40905 37764 40982 37780
rect 40722 37665 40870 37747
rect 40610 37632 40687 37648
tri 40687 37632 40703 37648 sw
rect 40610 37566 40703 37632
rect 40610 37464 40703 37530
rect 40610 37448 40687 37464
tri 40687 37448 40703 37464 nw
rect 40739 37431 40853 37665
tri 40889 37632 40905 37648 se
rect 40905 37632 40982 37648
rect 40889 37566 40982 37632
rect 40889 37464 40982 37530
tri 40889 37448 40905 37464 ne
rect 40905 37448 40982 37464
rect 40722 37349 40870 37431
rect 40610 37316 40687 37332
tri 40687 37316 40703 37332 sw
rect 40610 37250 40703 37316
rect 40739 37191 40853 37349
tri 40889 37316 40905 37332 se
rect 40905 37316 40982 37332
rect 40889 37250 40982 37316
rect 40610 37115 40982 37191
rect 40610 36990 40703 37056
rect 40610 36974 40687 36990
tri 40687 36974 40703 36990 nw
rect 40739 36957 40853 37115
rect 40889 36990 40982 37056
tri 40889 36974 40905 36990 ne
rect 40905 36974 40982 36990
rect 40722 36875 40870 36957
rect 40610 36842 40687 36858
tri 40687 36842 40703 36858 sw
rect 40610 36776 40703 36842
rect 40610 36674 40703 36740
rect 40610 36658 40687 36674
tri 40687 36658 40703 36674 nw
rect 40739 36641 40853 36875
tri 40889 36842 40905 36858 se
rect 40905 36842 40982 36858
rect 40889 36776 40982 36842
rect 40889 36674 40982 36740
tri 40889 36658 40905 36674 ne
rect 40905 36658 40982 36674
rect 40722 36559 40870 36641
rect 40610 36526 40687 36542
tri 40687 36526 40703 36542 sw
rect 40610 36460 40703 36526
rect 40739 36401 40853 36559
tri 40889 36526 40905 36542 se
rect 40905 36526 40982 36542
rect 40889 36460 40982 36526
rect 40610 36325 40982 36401
rect 40610 36200 40703 36266
rect 40610 36184 40687 36200
tri 40687 36184 40703 36200 nw
rect 40739 36167 40853 36325
rect 40889 36200 40982 36266
tri 40889 36184 40905 36200 ne
rect 40905 36184 40982 36200
rect 40722 36085 40870 36167
rect 40610 36052 40687 36068
tri 40687 36052 40703 36068 sw
rect 40610 35986 40703 36052
rect 40610 35884 40703 35950
rect 40610 35868 40687 35884
tri 40687 35868 40703 35884 nw
rect 40739 35851 40853 36085
tri 40889 36052 40905 36068 se
rect 40905 36052 40982 36068
rect 40889 35986 40982 36052
rect 40889 35884 40982 35950
tri 40889 35868 40905 35884 ne
rect 40905 35868 40982 35884
rect 40722 35769 40870 35851
rect 40610 35736 40687 35752
tri 40687 35736 40703 35752 sw
rect 40610 35670 40703 35736
rect 40739 35611 40853 35769
tri 40889 35736 40905 35752 se
rect 40905 35736 40982 35752
rect 40889 35670 40982 35736
rect 40610 35535 40982 35611
rect 40610 35410 40703 35476
rect 40610 35394 40687 35410
tri 40687 35394 40703 35410 nw
rect 40739 35377 40853 35535
rect 40889 35410 40982 35476
tri 40889 35394 40905 35410 ne
rect 40905 35394 40982 35410
rect 40722 35295 40870 35377
rect 40610 35262 40687 35278
tri 40687 35262 40703 35278 sw
rect 40610 35196 40703 35262
rect 40610 35094 40703 35160
rect 40610 35078 40687 35094
tri 40687 35078 40703 35094 nw
rect 40739 35061 40853 35295
tri 40889 35262 40905 35278 se
rect 40905 35262 40982 35278
rect 40889 35196 40982 35262
rect 40889 35094 40982 35160
tri 40889 35078 40905 35094 ne
rect 40905 35078 40982 35094
rect 40722 34979 40870 35061
rect 40610 34946 40687 34962
tri 40687 34946 40703 34962 sw
rect 40610 34880 40703 34946
rect 40739 34821 40853 34979
tri 40889 34946 40905 34962 se
rect 40905 34946 40982 34962
rect 40889 34880 40982 34946
rect 40610 34745 40982 34821
rect 40610 34620 40703 34686
rect 40610 34604 40687 34620
tri 40687 34604 40703 34620 nw
rect 40739 34587 40853 34745
rect 40889 34620 40982 34686
tri 40889 34604 40905 34620 ne
rect 40905 34604 40982 34620
rect 40722 34505 40870 34587
rect 40610 34472 40687 34488
tri 40687 34472 40703 34488 sw
rect 40610 34406 40703 34472
rect 40610 34304 40703 34370
rect 40610 34288 40687 34304
tri 40687 34288 40703 34304 nw
rect 40739 34271 40853 34505
tri 40889 34472 40905 34488 se
rect 40905 34472 40982 34488
rect 40889 34406 40982 34472
rect 40889 34304 40982 34370
tri 40889 34288 40905 34304 ne
rect 40905 34288 40982 34304
rect 40722 34189 40870 34271
rect 40610 34156 40687 34172
tri 40687 34156 40703 34172 sw
rect 40610 34090 40703 34156
rect 40739 34031 40853 34189
tri 40889 34156 40905 34172 se
rect 40905 34156 40982 34172
rect 40889 34090 40982 34156
rect 40610 33955 40982 34031
rect 40610 33830 40703 33896
rect 40610 33814 40687 33830
tri 40687 33814 40703 33830 nw
rect 40739 33797 40853 33955
rect 40889 33830 40982 33896
tri 40889 33814 40905 33830 ne
rect 40905 33814 40982 33830
rect 40722 33715 40870 33797
rect 40610 33682 40687 33698
tri 40687 33682 40703 33698 sw
rect 40610 33616 40703 33682
rect 40610 33514 40703 33580
rect 40610 33498 40687 33514
tri 40687 33498 40703 33514 nw
rect 40739 33481 40853 33715
tri 40889 33682 40905 33698 se
rect 40905 33682 40982 33698
rect 40889 33616 40982 33682
rect 40889 33514 40982 33580
tri 40889 33498 40905 33514 ne
rect 40905 33498 40982 33514
rect 40722 33399 40870 33481
rect 40610 33366 40687 33382
tri 40687 33366 40703 33382 sw
rect 40610 33300 40703 33366
rect 40739 33241 40853 33399
tri 40889 33366 40905 33382 se
rect 40905 33366 40982 33382
rect 40889 33300 40982 33366
rect 40610 33165 40982 33241
rect 40610 33040 40703 33106
rect 40610 33024 40687 33040
tri 40687 33024 40703 33040 nw
rect 40739 33007 40853 33165
rect 40889 33040 40982 33106
tri 40889 33024 40905 33040 ne
rect 40905 33024 40982 33040
rect 40722 32925 40870 33007
rect 40610 32892 40687 32908
tri 40687 32892 40703 32908 sw
rect 40610 32826 40703 32892
rect 40610 32724 40703 32790
rect 40610 32708 40687 32724
tri 40687 32708 40703 32724 nw
rect 40739 32691 40853 32925
tri 40889 32892 40905 32908 se
rect 40905 32892 40982 32908
rect 40889 32826 40982 32892
rect 40889 32724 40982 32790
tri 40889 32708 40905 32724 ne
rect 40905 32708 40982 32724
rect 40722 32609 40870 32691
rect 40610 32576 40687 32592
tri 40687 32576 40703 32592 sw
rect 40610 32510 40703 32576
rect 40739 32451 40853 32609
tri 40889 32576 40905 32592 se
rect 40905 32576 40982 32592
rect 40889 32510 40982 32576
rect 40610 32375 40982 32451
rect 40610 32250 40703 32316
rect 40610 32234 40687 32250
tri 40687 32234 40703 32250 nw
rect 40739 32217 40853 32375
rect 40889 32250 40982 32316
tri 40889 32234 40905 32250 ne
rect 40905 32234 40982 32250
rect 40722 32135 40870 32217
rect 40610 32102 40687 32118
tri 40687 32102 40703 32118 sw
rect 40610 32036 40703 32102
rect 40610 31934 40703 32000
rect 40610 31918 40687 31934
tri 40687 31918 40703 31934 nw
rect 40739 31901 40853 32135
tri 40889 32102 40905 32118 se
rect 40905 32102 40982 32118
rect 40889 32036 40982 32102
rect 40889 31934 40982 32000
tri 40889 31918 40905 31934 ne
rect 40905 31918 40982 31934
rect 40722 31819 40870 31901
rect 40610 31786 40687 31802
tri 40687 31786 40703 31802 sw
rect 40610 31720 40703 31786
rect 40739 31661 40853 31819
tri 40889 31786 40905 31802 se
rect 40905 31786 40982 31802
rect 40889 31720 40982 31786
rect 40610 31585 40982 31661
rect 40610 31460 40703 31526
rect 40610 31444 40687 31460
tri 40687 31444 40703 31460 nw
rect 40739 31427 40853 31585
rect 40889 31460 40982 31526
tri 40889 31444 40905 31460 ne
rect 40905 31444 40982 31460
rect 40722 31345 40870 31427
rect 40610 31312 40687 31328
tri 40687 31312 40703 31328 sw
rect 40610 31246 40703 31312
rect 40610 31144 40703 31210
rect 40610 31128 40687 31144
tri 40687 31128 40703 31144 nw
rect 40739 31111 40853 31345
tri 40889 31312 40905 31328 se
rect 40905 31312 40982 31328
rect 40889 31246 40982 31312
rect 40889 31144 40982 31210
tri 40889 31128 40905 31144 ne
rect 40905 31128 40982 31144
rect 40722 31029 40870 31111
rect 40610 30996 40687 31012
tri 40687 30996 40703 31012 sw
rect 40610 30930 40703 30996
rect 40739 30871 40853 31029
tri 40889 30996 40905 31012 se
rect 40905 30996 40982 31012
rect 40889 30930 40982 30996
rect 40610 30795 40982 30871
rect 40610 30670 40703 30736
rect 40610 30654 40687 30670
tri 40687 30654 40703 30670 nw
rect 40739 30637 40853 30795
rect 40889 30670 40982 30736
tri 40889 30654 40905 30670 ne
rect 40905 30654 40982 30670
rect 40722 30555 40870 30637
rect 40610 30522 40687 30538
tri 40687 30522 40703 30538 sw
rect 40610 30456 40703 30522
rect 40610 30354 40703 30420
rect 40610 30338 40687 30354
tri 40687 30338 40703 30354 nw
rect 40739 30321 40853 30555
tri 40889 30522 40905 30538 se
rect 40905 30522 40982 30538
rect 40889 30456 40982 30522
rect 40889 30354 40982 30420
tri 40889 30338 40905 30354 ne
rect 40905 30338 40982 30354
rect 40722 30239 40870 30321
rect 40610 30206 40687 30222
tri 40687 30206 40703 30222 sw
rect 40610 30140 40703 30206
rect 40739 30081 40853 30239
tri 40889 30206 40905 30222 se
rect 40905 30206 40982 30222
rect 40889 30140 40982 30206
rect 40610 30005 40982 30081
rect 40610 29880 40703 29946
rect 40610 29864 40687 29880
tri 40687 29864 40703 29880 nw
rect 40739 29847 40853 30005
rect 40889 29880 40982 29946
tri 40889 29864 40905 29880 ne
rect 40905 29864 40982 29880
rect 40722 29765 40870 29847
rect 40610 29732 40687 29748
tri 40687 29732 40703 29748 sw
rect 40610 29666 40703 29732
rect 40610 29564 40703 29630
rect 40610 29548 40687 29564
tri 40687 29548 40703 29564 nw
rect 40739 29531 40853 29765
tri 40889 29732 40905 29748 se
rect 40905 29732 40982 29748
rect 40889 29666 40982 29732
rect 40889 29564 40982 29630
tri 40889 29548 40905 29564 ne
rect 40905 29548 40982 29564
rect 40722 29449 40870 29531
rect 40610 29416 40687 29432
tri 40687 29416 40703 29432 sw
rect 40610 29350 40703 29416
rect 40739 29291 40853 29449
tri 40889 29416 40905 29432 se
rect 40905 29416 40982 29432
rect 40889 29350 40982 29416
rect 40610 29215 40982 29291
rect 40610 29090 40703 29156
rect 40610 29074 40687 29090
tri 40687 29074 40703 29090 nw
rect 40739 29057 40853 29215
rect 40889 29090 40982 29156
tri 40889 29074 40905 29090 ne
rect 40905 29074 40982 29090
rect 40722 28975 40870 29057
rect 40610 28942 40687 28958
tri 40687 28942 40703 28958 sw
rect 40610 28876 40703 28942
rect 40739 28833 40853 28975
tri 40889 28942 40905 28958 se
rect 40905 28942 40982 28958
rect 40889 28876 40982 28942
rect 41018 28463 41054 80603
rect 41090 28463 41126 80603
rect 41162 80445 41198 80603
rect 41154 80303 41206 80445
rect 41162 28763 41198 80303
rect 41154 28621 41206 28763
rect 41162 28463 41198 28621
rect 41234 28463 41270 80603
rect 41306 28463 41342 80603
rect 41378 28833 41462 80233
rect 41498 28463 41534 80603
rect 41570 28463 41606 80603
rect 41642 80445 41678 80603
rect 41634 80303 41686 80445
rect 41642 28763 41678 80303
rect 41634 28621 41686 28763
rect 41642 28463 41678 28621
rect 41714 28463 41750 80603
rect 41786 28463 41822 80603
rect 41858 80124 41951 80190
rect 41858 80108 41935 80124
tri 41935 80108 41951 80124 nw
rect 41987 80091 42101 80233
rect 42137 80124 42230 80190
tri 42137 80108 42153 80124 ne
rect 42153 80108 42230 80124
rect 41970 80009 42118 80091
rect 41858 79976 41935 79992
tri 41935 79976 41951 79992 sw
rect 41858 79910 41951 79976
rect 41987 79851 42101 80009
tri 42137 79976 42153 79992 se
rect 42153 79976 42230 79992
rect 42137 79910 42230 79976
rect 41858 79775 42230 79851
rect 41858 79650 41951 79716
rect 41858 79634 41935 79650
tri 41935 79634 41951 79650 nw
rect 41987 79617 42101 79775
rect 42137 79650 42230 79716
tri 42137 79634 42153 79650 ne
rect 42153 79634 42230 79650
rect 41970 79535 42118 79617
rect 41858 79502 41935 79518
tri 41935 79502 41951 79518 sw
rect 41858 79436 41951 79502
rect 41858 79334 41951 79400
rect 41858 79318 41935 79334
tri 41935 79318 41951 79334 nw
rect 41987 79301 42101 79535
tri 42137 79502 42153 79518 se
rect 42153 79502 42230 79518
rect 42137 79436 42230 79502
rect 42137 79334 42230 79400
tri 42137 79318 42153 79334 ne
rect 42153 79318 42230 79334
rect 41970 79219 42118 79301
rect 41858 79186 41935 79202
tri 41935 79186 41951 79202 sw
rect 41858 79120 41951 79186
rect 41987 79061 42101 79219
tri 42137 79186 42153 79202 se
rect 42153 79186 42230 79202
rect 42137 79120 42230 79186
rect 41858 78985 42230 79061
rect 41858 78860 41951 78926
rect 41858 78844 41935 78860
tri 41935 78844 41951 78860 nw
rect 41987 78827 42101 78985
rect 42137 78860 42230 78926
tri 42137 78844 42153 78860 ne
rect 42153 78844 42230 78860
rect 41970 78745 42118 78827
rect 41858 78712 41935 78728
tri 41935 78712 41951 78728 sw
rect 41858 78646 41951 78712
rect 41858 78544 41951 78610
rect 41858 78528 41935 78544
tri 41935 78528 41951 78544 nw
rect 41987 78511 42101 78745
tri 42137 78712 42153 78728 se
rect 42153 78712 42230 78728
rect 42137 78646 42230 78712
rect 42137 78544 42230 78610
tri 42137 78528 42153 78544 ne
rect 42153 78528 42230 78544
rect 41970 78429 42118 78511
rect 41858 78396 41935 78412
tri 41935 78396 41951 78412 sw
rect 41858 78330 41951 78396
rect 41987 78271 42101 78429
tri 42137 78396 42153 78412 se
rect 42153 78396 42230 78412
rect 42137 78330 42230 78396
rect 41858 78195 42230 78271
rect 41858 78070 41951 78136
rect 41858 78054 41935 78070
tri 41935 78054 41951 78070 nw
rect 41987 78037 42101 78195
rect 42137 78070 42230 78136
tri 42137 78054 42153 78070 ne
rect 42153 78054 42230 78070
rect 41970 77955 42118 78037
rect 41858 77922 41935 77938
tri 41935 77922 41951 77938 sw
rect 41858 77856 41951 77922
rect 41858 77754 41951 77820
rect 41858 77738 41935 77754
tri 41935 77738 41951 77754 nw
rect 41987 77721 42101 77955
tri 42137 77922 42153 77938 se
rect 42153 77922 42230 77938
rect 42137 77856 42230 77922
rect 42137 77754 42230 77820
tri 42137 77738 42153 77754 ne
rect 42153 77738 42230 77754
rect 41970 77639 42118 77721
rect 41858 77606 41935 77622
tri 41935 77606 41951 77622 sw
rect 41858 77540 41951 77606
rect 41987 77481 42101 77639
tri 42137 77606 42153 77622 se
rect 42153 77606 42230 77622
rect 42137 77540 42230 77606
rect 41858 77405 42230 77481
rect 41858 77280 41951 77346
rect 41858 77264 41935 77280
tri 41935 77264 41951 77280 nw
rect 41987 77247 42101 77405
rect 42137 77280 42230 77346
tri 42137 77264 42153 77280 ne
rect 42153 77264 42230 77280
rect 41970 77165 42118 77247
rect 41858 77132 41935 77148
tri 41935 77132 41951 77148 sw
rect 41858 77066 41951 77132
rect 41858 76964 41951 77030
rect 41858 76948 41935 76964
tri 41935 76948 41951 76964 nw
rect 41987 76931 42101 77165
tri 42137 77132 42153 77148 se
rect 42153 77132 42230 77148
rect 42137 77066 42230 77132
rect 42137 76964 42230 77030
tri 42137 76948 42153 76964 ne
rect 42153 76948 42230 76964
rect 41970 76849 42118 76931
rect 41858 76816 41935 76832
tri 41935 76816 41951 76832 sw
rect 41858 76750 41951 76816
rect 41987 76691 42101 76849
tri 42137 76816 42153 76832 se
rect 42153 76816 42230 76832
rect 42137 76750 42230 76816
rect 41858 76615 42230 76691
rect 41858 76490 41951 76556
rect 41858 76474 41935 76490
tri 41935 76474 41951 76490 nw
rect 41987 76457 42101 76615
rect 42137 76490 42230 76556
tri 42137 76474 42153 76490 ne
rect 42153 76474 42230 76490
rect 41970 76375 42118 76457
rect 41858 76342 41935 76358
tri 41935 76342 41951 76358 sw
rect 41858 76276 41951 76342
rect 41858 76174 41951 76240
rect 41858 76158 41935 76174
tri 41935 76158 41951 76174 nw
rect 41987 76141 42101 76375
tri 42137 76342 42153 76358 se
rect 42153 76342 42230 76358
rect 42137 76276 42230 76342
rect 42137 76174 42230 76240
tri 42137 76158 42153 76174 ne
rect 42153 76158 42230 76174
rect 41970 76059 42118 76141
rect 41858 76026 41935 76042
tri 41935 76026 41951 76042 sw
rect 41858 75960 41951 76026
rect 41987 75901 42101 76059
tri 42137 76026 42153 76042 se
rect 42153 76026 42230 76042
rect 42137 75960 42230 76026
rect 41858 75825 42230 75901
rect 41858 75700 41951 75766
rect 41858 75684 41935 75700
tri 41935 75684 41951 75700 nw
rect 41987 75667 42101 75825
rect 42137 75700 42230 75766
tri 42137 75684 42153 75700 ne
rect 42153 75684 42230 75700
rect 41970 75585 42118 75667
rect 41858 75552 41935 75568
tri 41935 75552 41951 75568 sw
rect 41858 75486 41951 75552
rect 41858 75384 41951 75450
rect 41858 75368 41935 75384
tri 41935 75368 41951 75384 nw
rect 41987 75351 42101 75585
tri 42137 75552 42153 75568 se
rect 42153 75552 42230 75568
rect 42137 75486 42230 75552
rect 42137 75384 42230 75450
tri 42137 75368 42153 75384 ne
rect 42153 75368 42230 75384
rect 41970 75269 42118 75351
rect 41858 75236 41935 75252
tri 41935 75236 41951 75252 sw
rect 41858 75170 41951 75236
rect 41987 75111 42101 75269
tri 42137 75236 42153 75252 se
rect 42153 75236 42230 75252
rect 42137 75170 42230 75236
rect 41858 75035 42230 75111
rect 41858 74910 41951 74976
rect 41858 74894 41935 74910
tri 41935 74894 41951 74910 nw
rect 41987 74877 42101 75035
rect 42137 74910 42230 74976
tri 42137 74894 42153 74910 ne
rect 42153 74894 42230 74910
rect 41970 74795 42118 74877
rect 41858 74762 41935 74778
tri 41935 74762 41951 74778 sw
rect 41858 74696 41951 74762
rect 41858 74594 41951 74660
rect 41858 74578 41935 74594
tri 41935 74578 41951 74594 nw
rect 41987 74561 42101 74795
tri 42137 74762 42153 74778 se
rect 42153 74762 42230 74778
rect 42137 74696 42230 74762
rect 42137 74594 42230 74660
tri 42137 74578 42153 74594 ne
rect 42153 74578 42230 74594
rect 41970 74479 42118 74561
rect 41858 74446 41935 74462
tri 41935 74446 41951 74462 sw
rect 41858 74380 41951 74446
rect 41987 74321 42101 74479
tri 42137 74446 42153 74462 se
rect 42153 74446 42230 74462
rect 42137 74380 42230 74446
rect 41858 74245 42230 74321
rect 41858 74120 41951 74186
rect 41858 74104 41935 74120
tri 41935 74104 41951 74120 nw
rect 41987 74087 42101 74245
rect 42137 74120 42230 74186
tri 42137 74104 42153 74120 ne
rect 42153 74104 42230 74120
rect 41970 74005 42118 74087
rect 41858 73972 41935 73988
tri 41935 73972 41951 73988 sw
rect 41858 73906 41951 73972
rect 41858 73804 41951 73870
rect 41858 73788 41935 73804
tri 41935 73788 41951 73804 nw
rect 41987 73771 42101 74005
tri 42137 73972 42153 73988 se
rect 42153 73972 42230 73988
rect 42137 73906 42230 73972
rect 42137 73804 42230 73870
tri 42137 73788 42153 73804 ne
rect 42153 73788 42230 73804
rect 41970 73689 42118 73771
rect 41858 73656 41935 73672
tri 41935 73656 41951 73672 sw
rect 41858 73590 41951 73656
rect 41987 73531 42101 73689
tri 42137 73656 42153 73672 se
rect 42153 73656 42230 73672
rect 42137 73590 42230 73656
rect 41858 73455 42230 73531
rect 41858 73330 41951 73396
rect 41858 73314 41935 73330
tri 41935 73314 41951 73330 nw
rect 41987 73297 42101 73455
rect 42137 73330 42230 73396
tri 42137 73314 42153 73330 ne
rect 42153 73314 42230 73330
rect 41970 73215 42118 73297
rect 41858 73182 41935 73198
tri 41935 73182 41951 73198 sw
rect 41858 73116 41951 73182
rect 41858 73014 41951 73080
rect 41858 72998 41935 73014
tri 41935 72998 41951 73014 nw
rect 41987 72981 42101 73215
tri 42137 73182 42153 73198 se
rect 42153 73182 42230 73198
rect 42137 73116 42230 73182
rect 42137 73014 42230 73080
tri 42137 72998 42153 73014 ne
rect 42153 72998 42230 73014
rect 41970 72899 42118 72981
rect 41858 72866 41935 72882
tri 41935 72866 41951 72882 sw
rect 41858 72800 41951 72866
rect 41987 72741 42101 72899
tri 42137 72866 42153 72882 se
rect 42153 72866 42230 72882
rect 42137 72800 42230 72866
rect 41858 72665 42230 72741
rect 41858 72540 41951 72606
rect 41858 72524 41935 72540
tri 41935 72524 41951 72540 nw
rect 41987 72507 42101 72665
rect 42137 72540 42230 72606
tri 42137 72524 42153 72540 ne
rect 42153 72524 42230 72540
rect 41970 72425 42118 72507
rect 41858 72392 41935 72408
tri 41935 72392 41951 72408 sw
rect 41858 72326 41951 72392
rect 41858 72224 41951 72290
rect 41858 72208 41935 72224
tri 41935 72208 41951 72224 nw
rect 41987 72191 42101 72425
tri 42137 72392 42153 72408 se
rect 42153 72392 42230 72408
rect 42137 72326 42230 72392
rect 42137 72224 42230 72290
tri 42137 72208 42153 72224 ne
rect 42153 72208 42230 72224
rect 41970 72109 42118 72191
rect 41858 72076 41935 72092
tri 41935 72076 41951 72092 sw
rect 41858 72010 41951 72076
rect 41987 71951 42101 72109
tri 42137 72076 42153 72092 se
rect 42153 72076 42230 72092
rect 42137 72010 42230 72076
rect 41858 71875 42230 71951
rect 41858 71750 41951 71816
rect 41858 71734 41935 71750
tri 41935 71734 41951 71750 nw
rect 41987 71717 42101 71875
rect 42137 71750 42230 71816
tri 42137 71734 42153 71750 ne
rect 42153 71734 42230 71750
rect 41970 71635 42118 71717
rect 41858 71602 41935 71618
tri 41935 71602 41951 71618 sw
rect 41858 71536 41951 71602
rect 41858 71434 41951 71500
rect 41858 71418 41935 71434
tri 41935 71418 41951 71434 nw
rect 41987 71401 42101 71635
tri 42137 71602 42153 71618 se
rect 42153 71602 42230 71618
rect 42137 71536 42230 71602
rect 42137 71434 42230 71500
tri 42137 71418 42153 71434 ne
rect 42153 71418 42230 71434
rect 41970 71319 42118 71401
rect 41858 71286 41935 71302
tri 41935 71286 41951 71302 sw
rect 41858 71220 41951 71286
rect 41987 71161 42101 71319
tri 42137 71286 42153 71302 se
rect 42153 71286 42230 71302
rect 42137 71220 42230 71286
rect 41858 71085 42230 71161
rect 41858 70960 41951 71026
rect 41858 70944 41935 70960
tri 41935 70944 41951 70960 nw
rect 41987 70927 42101 71085
rect 42137 70960 42230 71026
tri 42137 70944 42153 70960 ne
rect 42153 70944 42230 70960
rect 41970 70845 42118 70927
rect 41858 70812 41935 70828
tri 41935 70812 41951 70828 sw
rect 41858 70746 41951 70812
rect 41858 70644 41951 70710
rect 41858 70628 41935 70644
tri 41935 70628 41951 70644 nw
rect 41987 70611 42101 70845
tri 42137 70812 42153 70828 se
rect 42153 70812 42230 70828
rect 42137 70746 42230 70812
rect 42137 70644 42230 70710
tri 42137 70628 42153 70644 ne
rect 42153 70628 42230 70644
rect 41970 70529 42118 70611
rect 41858 70496 41935 70512
tri 41935 70496 41951 70512 sw
rect 41858 70430 41951 70496
rect 41987 70371 42101 70529
tri 42137 70496 42153 70512 se
rect 42153 70496 42230 70512
rect 42137 70430 42230 70496
rect 41858 70295 42230 70371
rect 41858 70170 41951 70236
rect 41858 70154 41935 70170
tri 41935 70154 41951 70170 nw
rect 41987 70137 42101 70295
rect 42137 70170 42230 70236
tri 42137 70154 42153 70170 ne
rect 42153 70154 42230 70170
rect 41970 70055 42118 70137
rect 41858 70022 41935 70038
tri 41935 70022 41951 70038 sw
rect 41858 69956 41951 70022
rect 41858 69854 41951 69920
rect 41858 69838 41935 69854
tri 41935 69838 41951 69854 nw
rect 41987 69821 42101 70055
tri 42137 70022 42153 70038 se
rect 42153 70022 42230 70038
rect 42137 69956 42230 70022
rect 42137 69854 42230 69920
tri 42137 69838 42153 69854 ne
rect 42153 69838 42230 69854
rect 41970 69739 42118 69821
rect 41858 69706 41935 69722
tri 41935 69706 41951 69722 sw
rect 41858 69640 41951 69706
rect 41987 69581 42101 69739
tri 42137 69706 42153 69722 se
rect 42153 69706 42230 69722
rect 42137 69640 42230 69706
rect 41858 69505 42230 69581
rect 41858 69380 41951 69446
rect 41858 69364 41935 69380
tri 41935 69364 41951 69380 nw
rect 41987 69347 42101 69505
rect 42137 69380 42230 69446
tri 42137 69364 42153 69380 ne
rect 42153 69364 42230 69380
rect 41970 69265 42118 69347
rect 41858 69232 41935 69248
tri 41935 69232 41951 69248 sw
rect 41858 69166 41951 69232
rect 41858 69064 41951 69130
rect 41858 69048 41935 69064
tri 41935 69048 41951 69064 nw
rect 41987 69031 42101 69265
tri 42137 69232 42153 69248 se
rect 42153 69232 42230 69248
rect 42137 69166 42230 69232
rect 42137 69064 42230 69130
tri 42137 69048 42153 69064 ne
rect 42153 69048 42230 69064
rect 41970 68949 42118 69031
rect 41858 68916 41935 68932
tri 41935 68916 41951 68932 sw
rect 41858 68850 41951 68916
rect 41987 68791 42101 68949
tri 42137 68916 42153 68932 se
rect 42153 68916 42230 68932
rect 42137 68850 42230 68916
rect 41858 68715 42230 68791
rect 41858 68590 41951 68656
rect 41858 68574 41935 68590
tri 41935 68574 41951 68590 nw
rect 41987 68557 42101 68715
rect 42137 68590 42230 68656
tri 42137 68574 42153 68590 ne
rect 42153 68574 42230 68590
rect 41970 68475 42118 68557
rect 41858 68442 41935 68458
tri 41935 68442 41951 68458 sw
rect 41858 68376 41951 68442
rect 41858 68274 41951 68340
rect 41858 68258 41935 68274
tri 41935 68258 41951 68274 nw
rect 41987 68241 42101 68475
tri 42137 68442 42153 68458 se
rect 42153 68442 42230 68458
rect 42137 68376 42230 68442
rect 42137 68274 42230 68340
tri 42137 68258 42153 68274 ne
rect 42153 68258 42230 68274
rect 41970 68159 42118 68241
rect 41858 68126 41935 68142
tri 41935 68126 41951 68142 sw
rect 41858 68060 41951 68126
rect 41987 68001 42101 68159
tri 42137 68126 42153 68142 se
rect 42153 68126 42230 68142
rect 42137 68060 42230 68126
rect 41858 67925 42230 68001
rect 41858 67800 41951 67866
rect 41858 67784 41935 67800
tri 41935 67784 41951 67800 nw
rect 41987 67767 42101 67925
rect 42137 67800 42230 67866
tri 42137 67784 42153 67800 ne
rect 42153 67784 42230 67800
rect 41970 67685 42118 67767
rect 41858 67652 41935 67668
tri 41935 67652 41951 67668 sw
rect 41858 67586 41951 67652
rect 41858 67484 41951 67550
rect 41858 67468 41935 67484
tri 41935 67468 41951 67484 nw
rect 41987 67451 42101 67685
tri 42137 67652 42153 67668 se
rect 42153 67652 42230 67668
rect 42137 67586 42230 67652
rect 42137 67484 42230 67550
tri 42137 67468 42153 67484 ne
rect 42153 67468 42230 67484
rect 41970 67369 42118 67451
rect 41858 67336 41935 67352
tri 41935 67336 41951 67352 sw
rect 41858 67270 41951 67336
rect 41987 67211 42101 67369
tri 42137 67336 42153 67352 se
rect 42153 67336 42230 67352
rect 42137 67270 42230 67336
rect 41858 67135 42230 67211
rect 41858 67010 41951 67076
rect 41858 66994 41935 67010
tri 41935 66994 41951 67010 nw
rect 41987 66977 42101 67135
rect 42137 67010 42230 67076
tri 42137 66994 42153 67010 ne
rect 42153 66994 42230 67010
rect 41970 66895 42118 66977
rect 41858 66862 41935 66878
tri 41935 66862 41951 66878 sw
rect 41858 66796 41951 66862
rect 41858 66694 41951 66760
rect 41858 66678 41935 66694
tri 41935 66678 41951 66694 nw
rect 41987 66661 42101 66895
tri 42137 66862 42153 66878 se
rect 42153 66862 42230 66878
rect 42137 66796 42230 66862
rect 42137 66694 42230 66760
tri 42137 66678 42153 66694 ne
rect 42153 66678 42230 66694
rect 41970 66579 42118 66661
rect 41858 66546 41935 66562
tri 41935 66546 41951 66562 sw
rect 41858 66480 41951 66546
rect 41987 66421 42101 66579
tri 42137 66546 42153 66562 se
rect 42153 66546 42230 66562
rect 42137 66480 42230 66546
rect 41858 66345 42230 66421
rect 41858 66220 41951 66286
rect 41858 66204 41935 66220
tri 41935 66204 41951 66220 nw
rect 41987 66187 42101 66345
rect 42137 66220 42230 66286
tri 42137 66204 42153 66220 ne
rect 42153 66204 42230 66220
rect 41970 66105 42118 66187
rect 41858 66072 41935 66088
tri 41935 66072 41951 66088 sw
rect 41858 66006 41951 66072
rect 41858 65904 41951 65970
rect 41858 65888 41935 65904
tri 41935 65888 41951 65904 nw
rect 41987 65871 42101 66105
tri 42137 66072 42153 66088 se
rect 42153 66072 42230 66088
rect 42137 66006 42230 66072
rect 42137 65904 42230 65970
tri 42137 65888 42153 65904 ne
rect 42153 65888 42230 65904
rect 41970 65789 42118 65871
rect 41858 65756 41935 65772
tri 41935 65756 41951 65772 sw
rect 41858 65690 41951 65756
rect 41987 65631 42101 65789
tri 42137 65756 42153 65772 se
rect 42153 65756 42230 65772
rect 42137 65690 42230 65756
rect 41858 65555 42230 65631
rect 41858 65430 41951 65496
rect 41858 65414 41935 65430
tri 41935 65414 41951 65430 nw
rect 41987 65397 42101 65555
rect 42137 65430 42230 65496
tri 42137 65414 42153 65430 ne
rect 42153 65414 42230 65430
rect 41970 65315 42118 65397
rect 41858 65282 41935 65298
tri 41935 65282 41951 65298 sw
rect 41858 65216 41951 65282
rect 41858 65114 41951 65180
rect 41858 65098 41935 65114
tri 41935 65098 41951 65114 nw
rect 41987 65081 42101 65315
tri 42137 65282 42153 65298 se
rect 42153 65282 42230 65298
rect 42137 65216 42230 65282
rect 42137 65114 42230 65180
tri 42137 65098 42153 65114 ne
rect 42153 65098 42230 65114
rect 41970 64999 42118 65081
rect 41858 64966 41935 64982
tri 41935 64966 41951 64982 sw
rect 41858 64900 41951 64966
rect 41987 64841 42101 64999
tri 42137 64966 42153 64982 se
rect 42153 64966 42230 64982
rect 42137 64900 42230 64966
rect 41858 64765 42230 64841
rect 41858 64640 41951 64706
rect 41858 64624 41935 64640
tri 41935 64624 41951 64640 nw
rect 41987 64607 42101 64765
rect 42137 64640 42230 64706
tri 42137 64624 42153 64640 ne
rect 42153 64624 42230 64640
rect 41970 64525 42118 64607
rect 41858 64492 41935 64508
tri 41935 64492 41951 64508 sw
rect 41858 64426 41951 64492
rect 41858 64324 41951 64390
rect 41858 64308 41935 64324
tri 41935 64308 41951 64324 nw
rect 41987 64291 42101 64525
tri 42137 64492 42153 64508 se
rect 42153 64492 42230 64508
rect 42137 64426 42230 64492
rect 42137 64324 42230 64390
tri 42137 64308 42153 64324 ne
rect 42153 64308 42230 64324
rect 41970 64209 42118 64291
rect 41858 64176 41935 64192
tri 41935 64176 41951 64192 sw
rect 41858 64110 41951 64176
rect 41987 64051 42101 64209
tri 42137 64176 42153 64192 se
rect 42153 64176 42230 64192
rect 42137 64110 42230 64176
rect 41858 63975 42230 64051
rect 41858 63850 41951 63916
rect 41858 63834 41935 63850
tri 41935 63834 41951 63850 nw
rect 41987 63817 42101 63975
rect 42137 63850 42230 63916
tri 42137 63834 42153 63850 ne
rect 42153 63834 42230 63850
rect 41970 63735 42118 63817
rect 41858 63702 41935 63718
tri 41935 63702 41951 63718 sw
rect 41858 63636 41951 63702
rect 41858 63534 41951 63600
rect 41858 63518 41935 63534
tri 41935 63518 41951 63534 nw
rect 41987 63501 42101 63735
tri 42137 63702 42153 63718 se
rect 42153 63702 42230 63718
rect 42137 63636 42230 63702
rect 42137 63534 42230 63600
tri 42137 63518 42153 63534 ne
rect 42153 63518 42230 63534
rect 41970 63419 42118 63501
rect 41858 63386 41935 63402
tri 41935 63386 41951 63402 sw
rect 41858 63320 41951 63386
rect 41987 63261 42101 63419
tri 42137 63386 42153 63402 se
rect 42153 63386 42230 63402
rect 42137 63320 42230 63386
rect 41858 63185 42230 63261
rect 41858 63060 41951 63126
rect 41858 63044 41935 63060
tri 41935 63044 41951 63060 nw
rect 41987 63027 42101 63185
rect 42137 63060 42230 63126
tri 42137 63044 42153 63060 ne
rect 42153 63044 42230 63060
rect 41970 62945 42118 63027
rect 41858 62912 41935 62928
tri 41935 62912 41951 62928 sw
rect 41858 62846 41951 62912
rect 41858 62744 41951 62810
rect 41858 62728 41935 62744
tri 41935 62728 41951 62744 nw
rect 41987 62711 42101 62945
tri 42137 62912 42153 62928 se
rect 42153 62912 42230 62928
rect 42137 62846 42230 62912
rect 42137 62744 42230 62810
tri 42137 62728 42153 62744 ne
rect 42153 62728 42230 62744
rect 41970 62629 42118 62711
rect 41858 62596 41935 62612
tri 41935 62596 41951 62612 sw
rect 41858 62530 41951 62596
rect 41987 62471 42101 62629
tri 42137 62596 42153 62612 se
rect 42153 62596 42230 62612
rect 42137 62530 42230 62596
rect 41858 62395 42230 62471
rect 41858 62270 41951 62336
rect 41858 62254 41935 62270
tri 41935 62254 41951 62270 nw
rect 41987 62237 42101 62395
rect 42137 62270 42230 62336
tri 42137 62254 42153 62270 ne
rect 42153 62254 42230 62270
rect 41970 62155 42118 62237
rect 41858 62122 41935 62138
tri 41935 62122 41951 62138 sw
rect 41858 62056 41951 62122
rect 41858 61954 41951 62020
rect 41858 61938 41935 61954
tri 41935 61938 41951 61954 nw
rect 41987 61921 42101 62155
tri 42137 62122 42153 62138 se
rect 42153 62122 42230 62138
rect 42137 62056 42230 62122
rect 42137 61954 42230 62020
tri 42137 61938 42153 61954 ne
rect 42153 61938 42230 61954
rect 41970 61839 42118 61921
rect 41858 61806 41935 61822
tri 41935 61806 41951 61822 sw
rect 41858 61740 41951 61806
rect 41987 61681 42101 61839
tri 42137 61806 42153 61822 se
rect 42153 61806 42230 61822
rect 42137 61740 42230 61806
rect 41858 61605 42230 61681
rect 41858 61480 41951 61546
rect 41858 61464 41935 61480
tri 41935 61464 41951 61480 nw
rect 41987 61447 42101 61605
rect 42137 61480 42230 61546
tri 42137 61464 42153 61480 ne
rect 42153 61464 42230 61480
rect 41970 61365 42118 61447
rect 41858 61332 41935 61348
tri 41935 61332 41951 61348 sw
rect 41858 61266 41951 61332
rect 41858 61164 41951 61230
rect 41858 61148 41935 61164
tri 41935 61148 41951 61164 nw
rect 41987 61131 42101 61365
tri 42137 61332 42153 61348 se
rect 42153 61332 42230 61348
rect 42137 61266 42230 61332
rect 42137 61164 42230 61230
tri 42137 61148 42153 61164 ne
rect 42153 61148 42230 61164
rect 41970 61049 42118 61131
rect 41858 61016 41935 61032
tri 41935 61016 41951 61032 sw
rect 41858 60950 41951 61016
rect 41987 60891 42101 61049
tri 42137 61016 42153 61032 se
rect 42153 61016 42230 61032
rect 42137 60950 42230 61016
rect 41858 60815 42230 60891
rect 41858 60690 41951 60756
rect 41858 60674 41935 60690
tri 41935 60674 41951 60690 nw
rect 41987 60657 42101 60815
rect 42137 60690 42230 60756
tri 42137 60674 42153 60690 ne
rect 42153 60674 42230 60690
rect 41970 60575 42118 60657
rect 41858 60542 41935 60558
tri 41935 60542 41951 60558 sw
rect 41858 60476 41951 60542
rect 41858 60374 41951 60440
rect 41858 60358 41935 60374
tri 41935 60358 41951 60374 nw
rect 41987 60341 42101 60575
tri 42137 60542 42153 60558 se
rect 42153 60542 42230 60558
rect 42137 60476 42230 60542
rect 42137 60374 42230 60440
tri 42137 60358 42153 60374 ne
rect 42153 60358 42230 60374
rect 41970 60259 42118 60341
rect 41858 60226 41935 60242
tri 41935 60226 41951 60242 sw
rect 41858 60160 41951 60226
rect 41987 60101 42101 60259
tri 42137 60226 42153 60242 se
rect 42153 60226 42230 60242
rect 42137 60160 42230 60226
rect 41858 60025 42230 60101
rect 41858 59900 41951 59966
rect 41858 59884 41935 59900
tri 41935 59884 41951 59900 nw
rect 41987 59867 42101 60025
rect 42137 59900 42230 59966
tri 42137 59884 42153 59900 ne
rect 42153 59884 42230 59900
rect 41970 59785 42118 59867
rect 41858 59752 41935 59768
tri 41935 59752 41951 59768 sw
rect 41858 59686 41951 59752
rect 41858 59584 41951 59650
rect 41858 59568 41935 59584
tri 41935 59568 41951 59584 nw
rect 41987 59551 42101 59785
tri 42137 59752 42153 59768 se
rect 42153 59752 42230 59768
rect 42137 59686 42230 59752
rect 42137 59584 42230 59650
tri 42137 59568 42153 59584 ne
rect 42153 59568 42230 59584
rect 41970 59469 42118 59551
rect 41858 59436 41935 59452
tri 41935 59436 41951 59452 sw
rect 41858 59370 41951 59436
rect 41987 59311 42101 59469
tri 42137 59436 42153 59452 se
rect 42153 59436 42230 59452
rect 42137 59370 42230 59436
rect 41858 59235 42230 59311
rect 41858 59110 41951 59176
rect 41858 59094 41935 59110
tri 41935 59094 41951 59110 nw
rect 41987 59077 42101 59235
rect 42137 59110 42230 59176
tri 42137 59094 42153 59110 ne
rect 42153 59094 42230 59110
rect 41970 58995 42118 59077
rect 41858 58962 41935 58978
tri 41935 58962 41951 58978 sw
rect 41858 58896 41951 58962
rect 41858 58794 41951 58860
rect 41858 58778 41935 58794
tri 41935 58778 41951 58794 nw
rect 41987 58761 42101 58995
tri 42137 58962 42153 58978 se
rect 42153 58962 42230 58978
rect 42137 58896 42230 58962
rect 42137 58794 42230 58860
tri 42137 58778 42153 58794 ne
rect 42153 58778 42230 58794
rect 41970 58679 42118 58761
rect 41858 58646 41935 58662
tri 41935 58646 41951 58662 sw
rect 41858 58580 41951 58646
rect 41987 58521 42101 58679
tri 42137 58646 42153 58662 se
rect 42153 58646 42230 58662
rect 42137 58580 42230 58646
rect 41858 58445 42230 58521
rect 41858 58320 41951 58386
rect 41858 58304 41935 58320
tri 41935 58304 41951 58320 nw
rect 41987 58287 42101 58445
rect 42137 58320 42230 58386
tri 42137 58304 42153 58320 ne
rect 42153 58304 42230 58320
rect 41970 58205 42118 58287
rect 41858 58172 41935 58188
tri 41935 58172 41951 58188 sw
rect 41858 58106 41951 58172
rect 41858 58004 41951 58070
rect 41858 57988 41935 58004
tri 41935 57988 41951 58004 nw
rect 41987 57971 42101 58205
tri 42137 58172 42153 58188 se
rect 42153 58172 42230 58188
rect 42137 58106 42230 58172
rect 42137 58004 42230 58070
tri 42137 57988 42153 58004 ne
rect 42153 57988 42230 58004
rect 41970 57889 42118 57971
rect 41858 57856 41935 57872
tri 41935 57856 41951 57872 sw
rect 41858 57790 41951 57856
rect 41987 57731 42101 57889
tri 42137 57856 42153 57872 se
rect 42153 57856 42230 57872
rect 42137 57790 42230 57856
rect 41858 57655 42230 57731
rect 41858 57530 41951 57596
rect 41858 57514 41935 57530
tri 41935 57514 41951 57530 nw
rect 41987 57497 42101 57655
rect 42137 57530 42230 57596
tri 42137 57514 42153 57530 ne
rect 42153 57514 42230 57530
rect 41970 57415 42118 57497
rect 41858 57382 41935 57398
tri 41935 57382 41951 57398 sw
rect 41858 57316 41951 57382
rect 41858 57214 41951 57280
rect 41858 57198 41935 57214
tri 41935 57198 41951 57214 nw
rect 41987 57181 42101 57415
tri 42137 57382 42153 57398 se
rect 42153 57382 42230 57398
rect 42137 57316 42230 57382
rect 42137 57214 42230 57280
tri 42137 57198 42153 57214 ne
rect 42153 57198 42230 57214
rect 41970 57099 42118 57181
rect 41858 57066 41935 57082
tri 41935 57066 41951 57082 sw
rect 41858 57000 41951 57066
rect 41987 56941 42101 57099
tri 42137 57066 42153 57082 se
rect 42153 57066 42230 57082
rect 42137 57000 42230 57066
rect 41858 56865 42230 56941
rect 41858 56740 41951 56806
rect 41858 56724 41935 56740
tri 41935 56724 41951 56740 nw
rect 41987 56707 42101 56865
rect 42137 56740 42230 56806
tri 42137 56724 42153 56740 ne
rect 42153 56724 42230 56740
rect 41970 56625 42118 56707
rect 41858 56592 41935 56608
tri 41935 56592 41951 56608 sw
rect 41858 56526 41951 56592
rect 41858 56424 41951 56490
rect 41858 56408 41935 56424
tri 41935 56408 41951 56424 nw
rect 41987 56391 42101 56625
tri 42137 56592 42153 56608 se
rect 42153 56592 42230 56608
rect 42137 56526 42230 56592
rect 42137 56424 42230 56490
tri 42137 56408 42153 56424 ne
rect 42153 56408 42230 56424
rect 41970 56309 42118 56391
rect 41858 56276 41935 56292
tri 41935 56276 41951 56292 sw
rect 41858 56210 41951 56276
rect 41987 56151 42101 56309
tri 42137 56276 42153 56292 se
rect 42153 56276 42230 56292
rect 42137 56210 42230 56276
rect 41858 56075 42230 56151
rect 41858 55950 41951 56016
rect 41858 55934 41935 55950
tri 41935 55934 41951 55950 nw
rect 41987 55917 42101 56075
rect 42137 55950 42230 56016
tri 42137 55934 42153 55950 ne
rect 42153 55934 42230 55950
rect 41970 55835 42118 55917
rect 41858 55802 41935 55818
tri 41935 55802 41951 55818 sw
rect 41858 55736 41951 55802
rect 41858 55634 41951 55700
rect 41858 55618 41935 55634
tri 41935 55618 41951 55634 nw
rect 41987 55601 42101 55835
tri 42137 55802 42153 55818 se
rect 42153 55802 42230 55818
rect 42137 55736 42230 55802
rect 42137 55634 42230 55700
tri 42137 55618 42153 55634 ne
rect 42153 55618 42230 55634
rect 41970 55519 42118 55601
rect 41858 55486 41935 55502
tri 41935 55486 41951 55502 sw
rect 41858 55420 41951 55486
rect 41987 55361 42101 55519
tri 42137 55486 42153 55502 se
rect 42153 55486 42230 55502
rect 42137 55420 42230 55486
rect 41858 55285 42230 55361
rect 41858 55160 41951 55226
rect 41858 55144 41935 55160
tri 41935 55144 41951 55160 nw
rect 41987 55127 42101 55285
rect 42137 55160 42230 55226
tri 42137 55144 42153 55160 ne
rect 42153 55144 42230 55160
rect 41970 55045 42118 55127
rect 41858 55012 41935 55028
tri 41935 55012 41951 55028 sw
rect 41858 54946 41951 55012
rect 41858 54844 41951 54910
rect 41858 54828 41935 54844
tri 41935 54828 41951 54844 nw
rect 41987 54811 42101 55045
tri 42137 55012 42153 55028 se
rect 42153 55012 42230 55028
rect 42137 54946 42230 55012
rect 42137 54844 42230 54910
tri 42137 54828 42153 54844 ne
rect 42153 54828 42230 54844
rect 41970 54729 42118 54811
rect 41858 54696 41935 54712
tri 41935 54696 41951 54712 sw
rect 41858 54630 41951 54696
rect 41987 54571 42101 54729
tri 42137 54696 42153 54712 se
rect 42153 54696 42230 54712
rect 42137 54630 42230 54696
rect 41858 54495 42230 54571
rect 41858 54370 41951 54436
rect 41858 54354 41935 54370
tri 41935 54354 41951 54370 nw
rect 41987 54337 42101 54495
rect 42137 54370 42230 54436
tri 42137 54354 42153 54370 ne
rect 42153 54354 42230 54370
rect 41970 54255 42118 54337
rect 41858 54222 41935 54238
tri 41935 54222 41951 54238 sw
rect 41858 54156 41951 54222
rect 41858 54054 41951 54120
rect 41858 54038 41935 54054
tri 41935 54038 41951 54054 nw
rect 41987 54021 42101 54255
tri 42137 54222 42153 54238 se
rect 42153 54222 42230 54238
rect 42137 54156 42230 54222
rect 42137 54054 42230 54120
tri 42137 54038 42153 54054 ne
rect 42153 54038 42230 54054
rect 41970 53939 42118 54021
rect 41858 53906 41935 53922
tri 41935 53906 41951 53922 sw
rect 41858 53840 41951 53906
rect 41987 53781 42101 53939
tri 42137 53906 42153 53922 se
rect 42153 53906 42230 53922
rect 42137 53840 42230 53906
rect 41858 53705 42230 53781
rect 41858 53580 41951 53646
rect 41858 53564 41935 53580
tri 41935 53564 41951 53580 nw
rect 41987 53547 42101 53705
rect 42137 53580 42230 53646
tri 42137 53564 42153 53580 ne
rect 42153 53564 42230 53580
rect 41970 53465 42118 53547
rect 41858 53432 41935 53448
tri 41935 53432 41951 53448 sw
rect 41858 53366 41951 53432
rect 41858 53264 41951 53330
rect 41858 53248 41935 53264
tri 41935 53248 41951 53264 nw
rect 41987 53231 42101 53465
tri 42137 53432 42153 53448 se
rect 42153 53432 42230 53448
rect 42137 53366 42230 53432
rect 42137 53264 42230 53330
tri 42137 53248 42153 53264 ne
rect 42153 53248 42230 53264
rect 41970 53149 42118 53231
rect 41858 53116 41935 53132
tri 41935 53116 41951 53132 sw
rect 41858 53050 41951 53116
rect 41987 52991 42101 53149
tri 42137 53116 42153 53132 se
rect 42153 53116 42230 53132
rect 42137 53050 42230 53116
rect 41858 52915 42230 52991
rect 41858 52790 41951 52856
rect 41858 52774 41935 52790
tri 41935 52774 41951 52790 nw
rect 41987 52757 42101 52915
rect 42137 52790 42230 52856
tri 42137 52774 42153 52790 ne
rect 42153 52774 42230 52790
rect 41970 52675 42118 52757
rect 41858 52642 41935 52658
tri 41935 52642 41951 52658 sw
rect 41858 52576 41951 52642
rect 41858 52474 41951 52540
rect 41858 52458 41935 52474
tri 41935 52458 41951 52474 nw
rect 41987 52441 42101 52675
tri 42137 52642 42153 52658 se
rect 42153 52642 42230 52658
rect 42137 52576 42230 52642
rect 42137 52474 42230 52540
tri 42137 52458 42153 52474 ne
rect 42153 52458 42230 52474
rect 41970 52359 42118 52441
rect 41858 52326 41935 52342
tri 41935 52326 41951 52342 sw
rect 41858 52260 41951 52326
rect 41987 52201 42101 52359
tri 42137 52326 42153 52342 se
rect 42153 52326 42230 52342
rect 42137 52260 42230 52326
rect 41858 52125 42230 52201
rect 41858 52000 41951 52066
rect 41858 51984 41935 52000
tri 41935 51984 41951 52000 nw
rect 41987 51967 42101 52125
rect 42137 52000 42230 52066
tri 42137 51984 42153 52000 ne
rect 42153 51984 42230 52000
rect 41970 51885 42118 51967
rect 41858 51852 41935 51868
tri 41935 51852 41951 51868 sw
rect 41858 51786 41951 51852
rect 41858 51684 41951 51750
rect 41858 51668 41935 51684
tri 41935 51668 41951 51684 nw
rect 41987 51651 42101 51885
tri 42137 51852 42153 51868 se
rect 42153 51852 42230 51868
rect 42137 51786 42230 51852
rect 42137 51684 42230 51750
tri 42137 51668 42153 51684 ne
rect 42153 51668 42230 51684
rect 41970 51569 42118 51651
rect 41858 51536 41935 51552
tri 41935 51536 41951 51552 sw
rect 41858 51470 41951 51536
rect 41987 51411 42101 51569
tri 42137 51536 42153 51552 se
rect 42153 51536 42230 51552
rect 42137 51470 42230 51536
rect 41858 51335 42230 51411
rect 41858 51210 41951 51276
rect 41858 51194 41935 51210
tri 41935 51194 41951 51210 nw
rect 41987 51177 42101 51335
rect 42137 51210 42230 51276
tri 42137 51194 42153 51210 ne
rect 42153 51194 42230 51210
rect 41970 51095 42118 51177
rect 41858 51062 41935 51078
tri 41935 51062 41951 51078 sw
rect 41858 50996 41951 51062
rect 41858 50894 41951 50960
rect 41858 50878 41935 50894
tri 41935 50878 41951 50894 nw
rect 41987 50861 42101 51095
tri 42137 51062 42153 51078 se
rect 42153 51062 42230 51078
rect 42137 50996 42230 51062
rect 42137 50894 42230 50960
tri 42137 50878 42153 50894 ne
rect 42153 50878 42230 50894
rect 41970 50779 42118 50861
rect 41858 50746 41935 50762
tri 41935 50746 41951 50762 sw
rect 41858 50680 41951 50746
rect 41987 50621 42101 50779
tri 42137 50746 42153 50762 se
rect 42153 50746 42230 50762
rect 42137 50680 42230 50746
rect 41858 50545 42230 50621
rect 41858 50420 41951 50486
rect 41858 50404 41935 50420
tri 41935 50404 41951 50420 nw
rect 41987 50387 42101 50545
rect 42137 50420 42230 50486
tri 42137 50404 42153 50420 ne
rect 42153 50404 42230 50420
rect 41970 50305 42118 50387
rect 41858 50272 41935 50288
tri 41935 50272 41951 50288 sw
rect 41858 50206 41951 50272
rect 41858 50104 41951 50170
rect 41858 50088 41935 50104
tri 41935 50088 41951 50104 nw
rect 41987 50071 42101 50305
tri 42137 50272 42153 50288 se
rect 42153 50272 42230 50288
rect 42137 50206 42230 50272
rect 42137 50104 42230 50170
tri 42137 50088 42153 50104 ne
rect 42153 50088 42230 50104
rect 41970 49989 42118 50071
rect 41858 49956 41935 49972
tri 41935 49956 41951 49972 sw
rect 41858 49890 41951 49956
rect 41987 49831 42101 49989
tri 42137 49956 42153 49972 se
rect 42153 49956 42230 49972
rect 42137 49890 42230 49956
rect 41858 49755 42230 49831
rect 41858 49630 41951 49696
rect 41858 49614 41935 49630
tri 41935 49614 41951 49630 nw
rect 41987 49597 42101 49755
rect 42137 49630 42230 49696
tri 42137 49614 42153 49630 ne
rect 42153 49614 42230 49630
rect 41970 49515 42118 49597
rect 41858 49482 41935 49498
tri 41935 49482 41951 49498 sw
rect 41858 49416 41951 49482
rect 41858 49314 41951 49380
rect 41858 49298 41935 49314
tri 41935 49298 41951 49314 nw
rect 41987 49281 42101 49515
tri 42137 49482 42153 49498 se
rect 42153 49482 42230 49498
rect 42137 49416 42230 49482
rect 42137 49314 42230 49380
tri 42137 49298 42153 49314 ne
rect 42153 49298 42230 49314
rect 41970 49199 42118 49281
rect 41858 49166 41935 49182
tri 41935 49166 41951 49182 sw
rect 41858 49100 41951 49166
rect 41987 49041 42101 49199
tri 42137 49166 42153 49182 se
rect 42153 49166 42230 49182
rect 42137 49100 42230 49166
rect 41858 48965 42230 49041
rect 41858 48840 41951 48906
rect 41858 48824 41935 48840
tri 41935 48824 41951 48840 nw
rect 41987 48807 42101 48965
rect 42137 48840 42230 48906
tri 42137 48824 42153 48840 ne
rect 42153 48824 42230 48840
rect 41970 48725 42118 48807
rect 41858 48692 41935 48708
tri 41935 48692 41951 48708 sw
rect 41858 48626 41951 48692
rect 41858 48524 41951 48590
rect 41858 48508 41935 48524
tri 41935 48508 41951 48524 nw
rect 41987 48491 42101 48725
tri 42137 48692 42153 48708 se
rect 42153 48692 42230 48708
rect 42137 48626 42230 48692
rect 42137 48524 42230 48590
tri 42137 48508 42153 48524 ne
rect 42153 48508 42230 48524
rect 41970 48409 42118 48491
rect 41858 48376 41935 48392
tri 41935 48376 41951 48392 sw
rect 41858 48310 41951 48376
rect 41987 48251 42101 48409
tri 42137 48376 42153 48392 se
rect 42153 48376 42230 48392
rect 42137 48310 42230 48376
rect 41858 48175 42230 48251
rect 41858 48050 41951 48116
rect 41858 48034 41935 48050
tri 41935 48034 41951 48050 nw
rect 41987 48017 42101 48175
rect 42137 48050 42230 48116
tri 42137 48034 42153 48050 ne
rect 42153 48034 42230 48050
rect 41970 47935 42118 48017
rect 41858 47902 41935 47918
tri 41935 47902 41951 47918 sw
rect 41858 47836 41951 47902
rect 41858 47734 41951 47800
rect 41858 47718 41935 47734
tri 41935 47718 41951 47734 nw
rect 41987 47701 42101 47935
tri 42137 47902 42153 47918 se
rect 42153 47902 42230 47918
rect 42137 47836 42230 47902
rect 42137 47734 42230 47800
tri 42137 47718 42153 47734 ne
rect 42153 47718 42230 47734
rect 41970 47619 42118 47701
rect 41858 47586 41935 47602
tri 41935 47586 41951 47602 sw
rect 41858 47520 41951 47586
rect 41987 47461 42101 47619
tri 42137 47586 42153 47602 se
rect 42153 47586 42230 47602
rect 42137 47520 42230 47586
rect 41858 47385 42230 47461
rect 41858 47260 41951 47326
rect 41858 47244 41935 47260
tri 41935 47244 41951 47260 nw
rect 41987 47227 42101 47385
rect 42137 47260 42230 47326
tri 42137 47244 42153 47260 ne
rect 42153 47244 42230 47260
rect 41970 47145 42118 47227
rect 41858 47112 41935 47128
tri 41935 47112 41951 47128 sw
rect 41858 47046 41951 47112
rect 41858 46944 41951 47010
rect 41858 46928 41935 46944
tri 41935 46928 41951 46944 nw
rect 41987 46911 42101 47145
tri 42137 47112 42153 47128 se
rect 42153 47112 42230 47128
rect 42137 47046 42230 47112
rect 42137 46944 42230 47010
tri 42137 46928 42153 46944 ne
rect 42153 46928 42230 46944
rect 41970 46829 42118 46911
rect 41858 46796 41935 46812
tri 41935 46796 41951 46812 sw
rect 41858 46730 41951 46796
rect 41987 46671 42101 46829
tri 42137 46796 42153 46812 se
rect 42153 46796 42230 46812
rect 42137 46730 42230 46796
rect 41858 46595 42230 46671
rect 41858 46470 41951 46536
rect 41858 46454 41935 46470
tri 41935 46454 41951 46470 nw
rect 41987 46437 42101 46595
rect 42137 46470 42230 46536
tri 42137 46454 42153 46470 ne
rect 42153 46454 42230 46470
rect 41970 46355 42118 46437
rect 41858 46322 41935 46338
tri 41935 46322 41951 46338 sw
rect 41858 46256 41951 46322
rect 41858 46154 41951 46220
rect 41858 46138 41935 46154
tri 41935 46138 41951 46154 nw
rect 41987 46121 42101 46355
tri 42137 46322 42153 46338 se
rect 42153 46322 42230 46338
rect 42137 46256 42230 46322
rect 42137 46154 42230 46220
tri 42137 46138 42153 46154 ne
rect 42153 46138 42230 46154
rect 41970 46039 42118 46121
rect 41858 46006 41935 46022
tri 41935 46006 41951 46022 sw
rect 41858 45940 41951 46006
rect 41987 45881 42101 46039
tri 42137 46006 42153 46022 se
rect 42153 46006 42230 46022
rect 42137 45940 42230 46006
rect 41858 45805 42230 45881
rect 41858 45680 41951 45746
rect 41858 45664 41935 45680
tri 41935 45664 41951 45680 nw
rect 41987 45647 42101 45805
rect 42137 45680 42230 45746
tri 42137 45664 42153 45680 ne
rect 42153 45664 42230 45680
rect 41970 45565 42118 45647
rect 41858 45532 41935 45548
tri 41935 45532 41951 45548 sw
rect 41858 45466 41951 45532
rect 41858 45364 41951 45430
rect 41858 45348 41935 45364
tri 41935 45348 41951 45364 nw
rect 41987 45331 42101 45565
tri 42137 45532 42153 45548 se
rect 42153 45532 42230 45548
rect 42137 45466 42230 45532
rect 42137 45364 42230 45430
tri 42137 45348 42153 45364 ne
rect 42153 45348 42230 45364
rect 41970 45249 42118 45331
rect 41858 45216 41935 45232
tri 41935 45216 41951 45232 sw
rect 41858 45150 41951 45216
rect 41987 45091 42101 45249
tri 42137 45216 42153 45232 se
rect 42153 45216 42230 45232
rect 42137 45150 42230 45216
rect 41858 45015 42230 45091
rect 41858 44890 41951 44956
rect 41858 44874 41935 44890
tri 41935 44874 41951 44890 nw
rect 41987 44857 42101 45015
rect 42137 44890 42230 44956
tri 42137 44874 42153 44890 ne
rect 42153 44874 42230 44890
rect 41970 44775 42118 44857
rect 41858 44742 41935 44758
tri 41935 44742 41951 44758 sw
rect 41858 44676 41951 44742
rect 41858 44574 41951 44640
rect 41858 44558 41935 44574
tri 41935 44558 41951 44574 nw
rect 41987 44541 42101 44775
tri 42137 44742 42153 44758 se
rect 42153 44742 42230 44758
rect 42137 44676 42230 44742
rect 42137 44574 42230 44640
tri 42137 44558 42153 44574 ne
rect 42153 44558 42230 44574
rect 41970 44459 42118 44541
rect 41858 44426 41935 44442
tri 41935 44426 41951 44442 sw
rect 41858 44360 41951 44426
rect 41987 44301 42101 44459
tri 42137 44426 42153 44442 se
rect 42153 44426 42230 44442
rect 42137 44360 42230 44426
rect 41858 44225 42230 44301
rect 41858 44100 41951 44166
rect 41858 44084 41935 44100
tri 41935 44084 41951 44100 nw
rect 41987 44067 42101 44225
rect 42137 44100 42230 44166
tri 42137 44084 42153 44100 ne
rect 42153 44084 42230 44100
rect 41970 43985 42118 44067
rect 41858 43952 41935 43968
tri 41935 43952 41951 43968 sw
rect 41858 43886 41951 43952
rect 41858 43784 41951 43850
rect 41858 43768 41935 43784
tri 41935 43768 41951 43784 nw
rect 41987 43751 42101 43985
tri 42137 43952 42153 43968 se
rect 42153 43952 42230 43968
rect 42137 43886 42230 43952
rect 42137 43784 42230 43850
tri 42137 43768 42153 43784 ne
rect 42153 43768 42230 43784
rect 41970 43669 42118 43751
rect 41858 43636 41935 43652
tri 41935 43636 41951 43652 sw
rect 41858 43570 41951 43636
rect 41987 43511 42101 43669
tri 42137 43636 42153 43652 se
rect 42153 43636 42230 43652
rect 42137 43570 42230 43636
rect 41858 43435 42230 43511
rect 41858 43310 41951 43376
rect 41858 43294 41935 43310
tri 41935 43294 41951 43310 nw
rect 41987 43277 42101 43435
rect 42137 43310 42230 43376
tri 42137 43294 42153 43310 ne
rect 42153 43294 42230 43310
rect 41970 43195 42118 43277
rect 41858 43162 41935 43178
tri 41935 43162 41951 43178 sw
rect 41858 43096 41951 43162
rect 41858 42994 41951 43060
rect 41858 42978 41935 42994
tri 41935 42978 41951 42994 nw
rect 41987 42961 42101 43195
tri 42137 43162 42153 43178 se
rect 42153 43162 42230 43178
rect 42137 43096 42230 43162
rect 42137 42994 42230 43060
tri 42137 42978 42153 42994 ne
rect 42153 42978 42230 42994
rect 41970 42879 42118 42961
rect 41858 42846 41935 42862
tri 41935 42846 41951 42862 sw
rect 41858 42780 41951 42846
rect 41987 42721 42101 42879
tri 42137 42846 42153 42862 se
rect 42153 42846 42230 42862
rect 42137 42780 42230 42846
rect 41858 42645 42230 42721
rect 41858 42520 41951 42586
rect 41858 42504 41935 42520
tri 41935 42504 41951 42520 nw
rect 41987 42487 42101 42645
rect 42137 42520 42230 42586
tri 42137 42504 42153 42520 ne
rect 42153 42504 42230 42520
rect 41970 42405 42118 42487
rect 41858 42372 41935 42388
tri 41935 42372 41951 42388 sw
rect 41858 42306 41951 42372
rect 41858 42204 41951 42270
rect 41858 42188 41935 42204
tri 41935 42188 41951 42204 nw
rect 41987 42171 42101 42405
tri 42137 42372 42153 42388 se
rect 42153 42372 42230 42388
rect 42137 42306 42230 42372
rect 42137 42204 42230 42270
tri 42137 42188 42153 42204 ne
rect 42153 42188 42230 42204
rect 41970 42089 42118 42171
rect 41858 42056 41935 42072
tri 41935 42056 41951 42072 sw
rect 41858 41990 41951 42056
rect 41987 41931 42101 42089
tri 42137 42056 42153 42072 se
rect 42153 42056 42230 42072
rect 42137 41990 42230 42056
rect 41858 41855 42230 41931
rect 41858 41730 41951 41796
rect 41858 41714 41935 41730
tri 41935 41714 41951 41730 nw
rect 41987 41697 42101 41855
rect 42137 41730 42230 41796
tri 42137 41714 42153 41730 ne
rect 42153 41714 42230 41730
rect 41970 41615 42118 41697
rect 41858 41582 41935 41598
tri 41935 41582 41951 41598 sw
rect 41858 41516 41951 41582
rect 41858 41414 41951 41480
rect 41858 41398 41935 41414
tri 41935 41398 41951 41414 nw
rect 41987 41381 42101 41615
tri 42137 41582 42153 41598 se
rect 42153 41582 42230 41598
rect 42137 41516 42230 41582
rect 42137 41414 42230 41480
tri 42137 41398 42153 41414 ne
rect 42153 41398 42230 41414
rect 41970 41299 42118 41381
rect 41858 41266 41935 41282
tri 41935 41266 41951 41282 sw
rect 41858 41200 41951 41266
rect 41987 41141 42101 41299
tri 42137 41266 42153 41282 se
rect 42153 41266 42230 41282
rect 42137 41200 42230 41266
rect 41858 41065 42230 41141
rect 41858 40940 41951 41006
rect 41858 40924 41935 40940
tri 41935 40924 41951 40940 nw
rect 41987 40907 42101 41065
rect 42137 40940 42230 41006
tri 42137 40924 42153 40940 ne
rect 42153 40924 42230 40940
rect 41970 40825 42118 40907
rect 41858 40792 41935 40808
tri 41935 40792 41951 40808 sw
rect 41858 40726 41951 40792
rect 41858 40624 41951 40690
rect 41858 40608 41935 40624
tri 41935 40608 41951 40624 nw
rect 41987 40591 42101 40825
tri 42137 40792 42153 40808 se
rect 42153 40792 42230 40808
rect 42137 40726 42230 40792
rect 42137 40624 42230 40690
tri 42137 40608 42153 40624 ne
rect 42153 40608 42230 40624
rect 41970 40509 42118 40591
rect 41858 40476 41935 40492
tri 41935 40476 41951 40492 sw
rect 41858 40410 41951 40476
rect 41987 40351 42101 40509
tri 42137 40476 42153 40492 se
rect 42153 40476 42230 40492
rect 42137 40410 42230 40476
rect 41858 40275 42230 40351
rect 41858 40150 41951 40216
rect 41858 40134 41935 40150
tri 41935 40134 41951 40150 nw
rect 41987 40117 42101 40275
rect 42137 40150 42230 40216
tri 42137 40134 42153 40150 ne
rect 42153 40134 42230 40150
rect 41970 40035 42118 40117
rect 41858 40002 41935 40018
tri 41935 40002 41951 40018 sw
rect 41858 39936 41951 40002
rect 41858 39834 41951 39900
rect 41858 39818 41935 39834
tri 41935 39818 41951 39834 nw
rect 41987 39801 42101 40035
tri 42137 40002 42153 40018 se
rect 42153 40002 42230 40018
rect 42137 39936 42230 40002
rect 42137 39834 42230 39900
tri 42137 39818 42153 39834 ne
rect 42153 39818 42230 39834
rect 41970 39719 42118 39801
rect 41858 39686 41935 39702
tri 41935 39686 41951 39702 sw
rect 41858 39620 41951 39686
rect 41987 39561 42101 39719
tri 42137 39686 42153 39702 se
rect 42153 39686 42230 39702
rect 42137 39620 42230 39686
rect 41858 39485 42230 39561
rect 41858 39360 41951 39426
rect 41858 39344 41935 39360
tri 41935 39344 41951 39360 nw
rect 41987 39327 42101 39485
rect 42137 39360 42230 39426
tri 42137 39344 42153 39360 ne
rect 42153 39344 42230 39360
rect 41970 39245 42118 39327
rect 41858 39212 41935 39228
tri 41935 39212 41951 39228 sw
rect 41858 39146 41951 39212
rect 41858 39044 41951 39110
rect 41858 39028 41935 39044
tri 41935 39028 41951 39044 nw
rect 41987 39011 42101 39245
tri 42137 39212 42153 39228 se
rect 42153 39212 42230 39228
rect 42137 39146 42230 39212
rect 42137 39044 42230 39110
tri 42137 39028 42153 39044 ne
rect 42153 39028 42230 39044
rect 41970 38929 42118 39011
rect 41858 38896 41935 38912
tri 41935 38896 41951 38912 sw
rect 41858 38830 41951 38896
rect 41987 38771 42101 38929
tri 42137 38896 42153 38912 se
rect 42153 38896 42230 38912
rect 42137 38830 42230 38896
rect 41858 38695 42230 38771
rect 41858 38570 41951 38636
rect 41858 38554 41935 38570
tri 41935 38554 41951 38570 nw
rect 41987 38537 42101 38695
rect 42137 38570 42230 38636
tri 42137 38554 42153 38570 ne
rect 42153 38554 42230 38570
rect 41970 38455 42118 38537
rect 41858 38422 41935 38438
tri 41935 38422 41951 38438 sw
rect 41858 38356 41951 38422
rect 41858 38254 41951 38320
rect 41858 38238 41935 38254
tri 41935 38238 41951 38254 nw
rect 41987 38221 42101 38455
tri 42137 38422 42153 38438 se
rect 42153 38422 42230 38438
rect 42137 38356 42230 38422
rect 42137 38254 42230 38320
tri 42137 38238 42153 38254 ne
rect 42153 38238 42230 38254
rect 41970 38139 42118 38221
rect 41858 38106 41935 38122
tri 41935 38106 41951 38122 sw
rect 41858 38040 41951 38106
rect 41987 37981 42101 38139
tri 42137 38106 42153 38122 se
rect 42153 38106 42230 38122
rect 42137 38040 42230 38106
rect 41858 37905 42230 37981
rect 41858 37780 41951 37846
rect 41858 37764 41935 37780
tri 41935 37764 41951 37780 nw
rect 41987 37747 42101 37905
rect 42137 37780 42230 37846
tri 42137 37764 42153 37780 ne
rect 42153 37764 42230 37780
rect 41970 37665 42118 37747
rect 41858 37632 41935 37648
tri 41935 37632 41951 37648 sw
rect 41858 37566 41951 37632
rect 41858 37464 41951 37530
rect 41858 37448 41935 37464
tri 41935 37448 41951 37464 nw
rect 41987 37431 42101 37665
tri 42137 37632 42153 37648 se
rect 42153 37632 42230 37648
rect 42137 37566 42230 37632
rect 42137 37464 42230 37530
tri 42137 37448 42153 37464 ne
rect 42153 37448 42230 37464
rect 41970 37349 42118 37431
rect 41858 37316 41935 37332
tri 41935 37316 41951 37332 sw
rect 41858 37250 41951 37316
rect 41987 37191 42101 37349
tri 42137 37316 42153 37332 se
rect 42153 37316 42230 37332
rect 42137 37250 42230 37316
rect 41858 37115 42230 37191
rect 41858 36990 41951 37056
rect 41858 36974 41935 36990
tri 41935 36974 41951 36990 nw
rect 41987 36957 42101 37115
rect 42137 36990 42230 37056
tri 42137 36974 42153 36990 ne
rect 42153 36974 42230 36990
rect 41970 36875 42118 36957
rect 41858 36842 41935 36858
tri 41935 36842 41951 36858 sw
rect 41858 36776 41951 36842
rect 41858 36674 41951 36740
rect 41858 36658 41935 36674
tri 41935 36658 41951 36674 nw
rect 41987 36641 42101 36875
tri 42137 36842 42153 36858 se
rect 42153 36842 42230 36858
rect 42137 36776 42230 36842
rect 42137 36674 42230 36740
tri 42137 36658 42153 36674 ne
rect 42153 36658 42230 36674
rect 41970 36559 42118 36641
rect 41858 36526 41935 36542
tri 41935 36526 41951 36542 sw
rect 41858 36460 41951 36526
rect 41987 36401 42101 36559
tri 42137 36526 42153 36542 se
rect 42153 36526 42230 36542
rect 42137 36460 42230 36526
rect 41858 36325 42230 36401
rect 41858 36200 41951 36266
rect 41858 36184 41935 36200
tri 41935 36184 41951 36200 nw
rect 41987 36167 42101 36325
rect 42137 36200 42230 36266
tri 42137 36184 42153 36200 ne
rect 42153 36184 42230 36200
rect 41970 36085 42118 36167
rect 41858 36052 41935 36068
tri 41935 36052 41951 36068 sw
rect 41858 35986 41951 36052
rect 41858 35884 41951 35950
rect 41858 35868 41935 35884
tri 41935 35868 41951 35884 nw
rect 41987 35851 42101 36085
tri 42137 36052 42153 36068 se
rect 42153 36052 42230 36068
rect 42137 35986 42230 36052
rect 42137 35884 42230 35950
tri 42137 35868 42153 35884 ne
rect 42153 35868 42230 35884
rect 41970 35769 42118 35851
rect 41858 35736 41935 35752
tri 41935 35736 41951 35752 sw
rect 41858 35670 41951 35736
rect 41987 35611 42101 35769
tri 42137 35736 42153 35752 se
rect 42153 35736 42230 35752
rect 42137 35670 42230 35736
rect 41858 35535 42230 35611
rect 41858 35410 41951 35476
rect 41858 35394 41935 35410
tri 41935 35394 41951 35410 nw
rect 41987 35377 42101 35535
rect 42137 35410 42230 35476
tri 42137 35394 42153 35410 ne
rect 42153 35394 42230 35410
rect 41970 35295 42118 35377
rect 41858 35262 41935 35278
tri 41935 35262 41951 35278 sw
rect 41858 35196 41951 35262
rect 41858 35094 41951 35160
rect 41858 35078 41935 35094
tri 41935 35078 41951 35094 nw
rect 41987 35061 42101 35295
tri 42137 35262 42153 35278 se
rect 42153 35262 42230 35278
rect 42137 35196 42230 35262
rect 42137 35094 42230 35160
tri 42137 35078 42153 35094 ne
rect 42153 35078 42230 35094
rect 41970 34979 42118 35061
rect 41858 34946 41935 34962
tri 41935 34946 41951 34962 sw
rect 41858 34880 41951 34946
rect 41987 34821 42101 34979
tri 42137 34946 42153 34962 se
rect 42153 34946 42230 34962
rect 42137 34880 42230 34946
rect 41858 34745 42230 34821
rect 41858 34620 41951 34686
rect 41858 34604 41935 34620
tri 41935 34604 41951 34620 nw
rect 41987 34587 42101 34745
rect 42137 34620 42230 34686
tri 42137 34604 42153 34620 ne
rect 42153 34604 42230 34620
rect 41970 34505 42118 34587
rect 41858 34472 41935 34488
tri 41935 34472 41951 34488 sw
rect 41858 34406 41951 34472
rect 41858 34304 41951 34370
rect 41858 34288 41935 34304
tri 41935 34288 41951 34304 nw
rect 41987 34271 42101 34505
tri 42137 34472 42153 34488 se
rect 42153 34472 42230 34488
rect 42137 34406 42230 34472
rect 42137 34304 42230 34370
tri 42137 34288 42153 34304 ne
rect 42153 34288 42230 34304
rect 41970 34189 42118 34271
rect 41858 34156 41935 34172
tri 41935 34156 41951 34172 sw
rect 41858 34090 41951 34156
rect 41987 34031 42101 34189
tri 42137 34156 42153 34172 se
rect 42153 34156 42230 34172
rect 42137 34090 42230 34156
rect 41858 33955 42230 34031
rect 41858 33830 41951 33896
rect 41858 33814 41935 33830
tri 41935 33814 41951 33830 nw
rect 41987 33797 42101 33955
rect 42137 33830 42230 33896
tri 42137 33814 42153 33830 ne
rect 42153 33814 42230 33830
rect 41970 33715 42118 33797
rect 41858 33682 41935 33698
tri 41935 33682 41951 33698 sw
rect 41858 33616 41951 33682
rect 41858 33514 41951 33580
rect 41858 33498 41935 33514
tri 41935 33498 41951 33514 nw
rect 41987 33481 42101 33715
tri 42137 33682 42153 33698 se
rect 42153 33682 42230 33698
rect 42137 33616 42230 33682
rect 42137 33514 42230 33580
tri 42137 33498 42153 33514 ne
rect 42153 33498 42230 33514
rect 41970 33399 42118 33481
rect 41858 33366 41935 33382
tri 41935 33366 41951 33382 sw
rect 41858 33300 41951 33366
rect 41987 33241 42101 33399
tri 42137 33366 42153 33382 se
rect 42153 33366 42230 33382
rect 42137 33300 42230 33366
rect 41858 33165 42230 33241
rect 41858 33040 41951 33106
rect 41858 33024 41935 33040
tri 41935 33024 41951 33040 nw
rect 41987 33007 42101 33165
rect 42137 33040 42230 33106
tri 42137 33024 42153 33040 ne
rect 42153 33024 42230 33040
rect 41970 32925 42118 33007
rect 41858 32892 41935 32908
tri 41935 32892 41951 32908 sw
rect 41858 32826 41951 32892
rect 41858 32724 41951 32790
rect 41858 32708 41935 32724
tri 41935 32708 41951 32724 nw
rect 41987 32691 42101 32925
tri 42137 32892 42153 32908 se
rect 42153 32892 42230 32908
rect 42137 32826 42230 32892
rect 42137 32724 42230 32790
tri 42137 32708 42153 32724 ne
rect 42153 32708 42230 32724
rect 41970 32609 42118 32691
rect 41858 32576 41935 32592
tri 41935 32576 41951 32592 sw
rect 41858 32510 41951 32576
rect 41987 32451 42101 32609
tri 42137 32576 42153 32592 se
rect 42153 32576 42230 32592
rect 42137 32510 42230 32576
rect 41858 32375 42230 32451
rect 41858 32250 41951 32316
rect 41858 32234 41935 32250
tri 41935 32234 41951 32250 nw
rect 41987 32217 42101 32375
rect 42137 32250 42230 32316
tri 42137 32234 42153 32250 ne
rect 42153 32234 42230 32250
rect 41970 32135 42118 32217
rect 41858 32102 41935 32118
tri 41935 32102 41951 32118 sw
rect 41858 32036 41951 32102
rect 41858 31934 41951 32000
rect 41858 31918 41935 31934
tri 41935 31918 41951 31934 nw
rect 41987 31901 42101 32135
tri 42137 32102 42153 32118 se
rect 42153 32102 42230 32118
rect 42137 32036 42230 32102
rect 42137 31934 42230 32000
tri 42137 31918 42153 31934 ne
rect 42153 31918 42230 31934
rect 41970 31819 42118 31901
rect 41858 31786 41935 31802
tri 41935 31786 41951 31802 sw
rect 41858 31720 41951 31786
rect 41987 31661 42101 31819
tri 42137 31786 42153 31802 se
rect 42153 31786 42230 31802
rect 42137 31720 42230 31786
rect 41858 31585 42230 31661
rect 41858 31460 41951 31526
rect 41858 31444 41935 31460
tri 41935 31444 41951 31460 nw
rect 41987 31427 42101 31585
rect 42137 31460 42230 31526
tri 42137 31444 42153 31460 ne
rect 42153 31444 42230 31460
rect 41970 31345 42118 31427
rect 41858 31312 41935 31328
tri 41935 31312 41951 31328 sw
rect 41858 31246 41951 31312
rect 41858 31144 41951 31210
rect 41858 31128 41935 31144
tri 41935 31128 41951 31144 nw
rect 41987 31111 42101 31345
tri 42137 31312 42153 31328 se
rect 42153 31312 42230 31328
rect 42137 31246 42230 31312
rect 42137 31144 42230 31210
tri 42137 31128 42153 31144 ne
rect 42153 31128 42230 31144
rect 41970 31029 42118 31111
rect 41858 30996 41935 31012
tri 41935 30996 41951 31012 sw
rect 41858 30930 41951 30996
rect 41987 30871 42101 31029
tri 42137 30996 42153 31012 se
rect 42153 30996 42230 31012
rect 42137 30930 42230 30996
rect 41858 30795 42230 30871
rect 41858 30670 41951 30736
rect 41858 30654 41935 30670
tri 41935 30654 41951 30670 nw
rect 41987 30637 42101 30795
rect 42137 30670 42230 30736
tri 42137 30654 42153 30670 ne
rect 42153 30654 42230 30670
rect 41970 30555 42118 30637
rect 41858 30522 41935 30538
tri 41935 30522 41951 30538 sw
rect 41858 30456 41951 30522
rect 41858 30354 41951 30420
rect 41858 30338 41935 30354
tri 41935 30338 41951 30354 nw
rect 41987 30321 42101 30555
tri 42137 30522 42153 30538 se
rect 42153 30522 42230 30538
rect 42137 30456 42230 30522
rect 42137 30354 42230 30420
tri 42137 30338 42153 30354 ne
rect 42153 30338 42230 30354
rect 41970 30239 42118 30321
rect 41858 30206 41935 30222
tri 41935 30206 41951 30222 sw
rect 41858 30140 41951 30206
rect 41987 30081 42101 30239
tri 42137 30206 42153 30222 se
rect 42153 30206 42230 30222
rect 42137 30140 42230 30206
rect 41858 30005 42230 30081
rect 41858 29880 41951 29946
rect 41858 29864 41935 29880
tri 41935 29864 41951 29880 nw
rect 41987 29847 42101 30005
rect 42137 29880 42230 29946
tri 42137 29864 42153 29880 ne
rect 42153 29864 42230 29880
rect 41970 29765 42118 29847
rect 41858 29732 41935 29748
tri 41935 29732 41951 29748 sw
rect 41858 29666 41951 29732
rect 41858 29564 41951 29630
rect 41858 29548 41935 29564
tri 41935 29548 41951 29564 nw
rect 41987 29531 42101 29765
tri 42137 29732 42153 29748 se
rect 42153 29732 42230 29748
rect 42137 29666 42230 29732
rect 42137 29564 42230 29630
tri 42137 29548 42153 29564 ne
rect 42153 29548 42230 29564
rect 41970 29449 42118 29531
rect 41858 29416 41935 29432
tri 41935 29416 41951 29432 sw
rect 41858 29350 41951 29416
rect 41987 29291 42101 29449
tri 42137 29416 42153 29432 se
rect 42153 29416 42230 29432
rect 42137 29350 42230 29416
rect 41858 29215 42230 29291
rect 41858 29090 41951 29156
rect 41858 29074 41935 29090
tri 41935 29074 41951 29090 nw
rect 41987 29057 42101 29215
rect 42137 29090 42230 29156
tri 42137 29074 42153 29090 ne
rect 42153 29074 42230 29090
rect 41970 28975 42118 29057
rect 41858 28942 41935 28958
tri 41935 28942 41951 28958 sw
rect 41858 28876 41951 28942
rect 41987 28833 42101 28975
tri 42137 28942 42153 28958 se
rect 42153 28942 42230 28958
rect 42137 28876 42230 28942
rect 42266 28463 42302 80603
rect 42338 28463 42374 80603
rect 42410 80445 42446 80603
rect 42402 80303 42454 80445
rect 42410 28763 42446 80303
rect 42402 28621 42454 28763
rect 42410 28463 42446 28621
rect 42482 28463 42518 80603
rect 42554 28463 42590 80603
rect 42626 28833 42710 80233
rect 42746 28463 42782 80603
rect 42818 28463 42854 80603
rect 42890 80445 42926 80603
rect 42882 80303 42934 80445
rect 42890 28763 42926 80303
rect 42882 28621 42934 28763
rect 42890 28463 42926 28621
rect 42962 28463 42998 80603
rect 43034 28463 43070 80603
rect 43106 80124 43199 80190
rect 43106 80108 43183 80124
tri 43183 80108 43199 80124 nw
rect 43235 80091 43349 80233
rect 43385 80124 43478 80190
tri 43385 80108 43401 80124 ne
rect 43401 80108 43478 80124
rect 43218 80009 43366 80091
rect 43106 79976 43183 79992
tri 43183 79976 43199 79992 sw
rect 43106 79910 43199 79976
rect 43235 79851 43349 80009
tri 43385 79976 43401 79992 se
rect 43401 79976 43478 79992
rect 43385 79910 43478 79976
rect 43106 79775 43478 79851
rect 43106 79650 43199 79716
rect 43106 79634 43183 79650
tri 43183 79634 43199 79650 nw
rect 43235 79617 43349 79775
rect 43385 79650 43478 79716
tri 43385 79634 43401 79650 ne
rect 43401 79634 43478 79650
rect 43218 79535 43366 79617
rect 43106 79502 43183 79518
tri 43183 79502 43199 79518 sw
rect 43106 79436 43199 79502
rect 43106 79334 43199 79400
rect 43106 79318 43183 79334
tri 43183 79318 43199 79334 nw
rect 43235 79301 43349 79535
tri 43385 79502 43401 79518 se
rect 43401 79502 43478 79518
rect 43385 79436 43478 79502
rect 43385 79334 43478 79400
tri 43385 79318 43401 79334 ne
rect 43401 79318 43478 79334
rect 43218 79219 43366 79301
rect 43106 79186 43183 79202
tri 43183 79186 43199 79202 sw
rect 43106 79120 43199 79186
rect 43235 79061 43349 79219
tri 43385 79186 43401 79202 se
rect 43401 79186 43478 79202
rect 43385 79120 43478 79186
rect 43106 78985 43478 79061
rect 43106 78860 43199 78926
rect 43106 78844 43183 78860
tri 43183 78844 43199 78860 nw
rect 43235 78827 43349 78985
rect 43385 78860 43478 78926
tri 43385 78844 43401 78860 ne
rect 43401 78844 43478 78860
rect 43218 78745 43366 78827
rect 43106 78712 43183 78728
tri 43183 78712 43199 78728 sw
rect 43106 78646 43199 78712
rect 43106 78544 43199 78610
rect 43106 78528 43183 78544
tri 43183 78528 43199 78544 nw
rect 43235 78511 43349 78745
tri 43385 78712 43401 78728 se
rect 43401 78712 43478 78728
rect 43385 78646 43478 78712
rect 43385 78544 43478 78610
tri 43385 78528 43401 78544 ne
rect 43401 78528 43478 78544
rect 43218 78429 43366 78511
rect 43106 78396 43183 78412
tri 43183 78396 43199 78412 sw
rect 43106 78330 43199 78396
rect 43235 78271 43349 78429
tri 43385 78396 43401 78412 se
rect 43401 78396 43478 78412
rect 43385 78330 43478 78396
rect 43106 78195 43478 78271
rect 43106 78070 43199 78136
rect 43106 78054 43183 78070
tri 43183 78054 43199 78070 nw
rect 43235 78037 43349 78195
rect 43385 78070 43478 78136
tri 43385 78054 43401 78070 ne
rect 43401 78054 43478 78070
rect 43218 77955 43366 78037
rect 43106 77922 43183 77938
tri 43183 77922 43199 77938 sw
rect 43106 77856 43199 77922
rect 43106 77754 43199 77820
rect 43106 77738 43183 77754
tri 43183 77738 43199 77754 nw
rect 43235 77721 43349 77955
tri 43385 77922 43401 77938 se
rect 43401 77922 43478 77938
rect 43385 77856 43478 77922
rect 43385 77754 43478 77820
tri 43385 77738 43401 77754 ne
rect 43401 77738 43478 77754
rect 43218 77639 43366 77721
rect 43106 77606 43183 77622
tri 43183 77606 43199 77622 sw
rect 43106 77540 43199 77606
rect 43235 77481 43349 77639
tri 43385 77606 43401 77622 se
rect 43401 77606 43478 77622
rect 43385 77540 43478 77606
rect 43106 77405 43478 77481
rect 43106 77280 43199 77346
rect 43106 77264 43183 77280
tri 43183 77264 43199 77280 nw
rect 43235 77247 43349 77405
rect 43385 77280 43478 77346
tri 43385 77264 43401 77280 ne
rect 43401 77264 43478 77280
rect 43218 77165 43366 77247
rect 43106 77132 43183 77148
tri 43183 77132 43199 77148 sw
rect 43106 77066 43199 77132
rect 43106 76964 43199 77030
rect 43106 76948 43183 76964
tri 43183 76948 43199 76964 nw
rect 43235 76931 43349 77165
tri 43385 77132 43401 77148 se
rect 43401 77132 43478 77148
rect 43385 77066 43478 77132
rect 43385 76964 43478 77030
tri 43385 76948 43401 76964 ne
rect 43401 76948 43478 76964
rect 43218 76849 43366 76931
rect 43106 76816 43183 76832
tri 43183 76816 43199 76832 sw
rect 43106 76750 43199 76816
rect 43235 76691 43349 76849
tri 43385 76816 43401 76832 se
rect 43401 76816 43478 76832
rect 43385 76750 43478 76816
rect 43106 76615 43478 76691
rect 43106 76490 43199 76556
rect 43106 76474 43183 76490
tri 43183 76474 43199 76490 nw
rect 43235 76457 43349 76615
rect 43385 76490 43478 76556
tri 43385 76474 43401 76490 ne
rect 43401 76474 43478 76490
rect 43218 76375 43366 76457
rect 43106 76342 43183 76358
tri 43183 76342 43199 76358 sw
rect 43106 76276 43199 76342
rect 43106 76174 43199 76240
rect 43106 76158 43183 76174
tri 43183 76158 43199 76174 nw
rect 43235 76141 43349 76375
tri 43385 76342 43401 76358 se
rect 43401 76342 43478 76358
rect 43385 76276 43478 76342
rect 43385 76174 43478 76240
tri 43385 76158 43401 76174 ne
rect 43401 76158 43478 76174
rect 43218 76059 43366 76141
rect 43106 76026 43183 76042
tri 43183 76026 43199 76042 sw
rect 43106 75960 43199 76026
rect 43235 75901 43349 76059
tri 43385 76026 43401 76042 se
rect 43401 76026 43478 76042
rect 43385 75960 43478 76026
rect 43106 75825 43478 75901
rect 43106 75700 43199 75766
rect 43106 75684 43183 75700
tri 43183 75684 43199 75700 nw
rect 43235 75667 43349 75825
rect 43385 75700 43478 75766
tri 43385 75684 43401 75700 ne
rect 43401 75684 43478 75700
rect 43218 75585 43366 75667
rect 43106 75552 43183 75568
tri 43183 75552 43199 75568 sw
rect 43106 75486 43199 75552
rect 43106 75384 43199 75450
rect 43106 75368 43183 75384
tri 43183 75368 43199 75384 nw
rect 43235 75351 43349 75585
tri 43385 75552 43401 75568 se
rect 43401 75552 43478 75568
rect 43385 75486 43478 75552
rect 43385 75384 43478 75450
tri 43385 75368 43401 75384 ne
rect 43401 75368 43478 75384
rect 43218 75269 43366 75351
rect 43106 75236 43183 75252
tri 43183 75236 43199 75252 sw
rect 43106 75170 43199 75236
rect 43235 75111 43349 75269
tri 43385 75236 43401 75252 se
rect 43401 75236 43478 75252
rect 43385 75170 43478 75236
rect 43106 75035 43478 75111
rect 43106 74910 43199 74976
rect 43106 74894 43183 74910
tri 43183 74894 43199 74910 nw
rect 43235 74877 43349 75035
rect 43385 74910 43478 74976
tri 43385 74894 43401 74910 ne
rect 43401 74894 43478 74910
rect 43218 74795 43366 74877
rect 43106 74762 43183 74778
tri 43183 74762 43199 74778 sw
rect 43106 74696 43199 74762
rect 43106 74594 43199 74660
rect 43106 74578 43183 74594
tri 43183 74578 43199 74594 nw
rect 43235 74561 43349 74795
tri 43385 74762 43401 74778 se
rect 43401 74762 43478 74778
rect 43385 74696 43478 74762
rect 43385 74594 43478 74660
tri 43385 74578 43401 74594 ne
rect 43401 74578 43478 74594
rect 43218 74479 43366 74561
rect 43106 74446 43183 74462
tri 43183 74446 43199 74462 sw
rect 43106 74380 43199 74446
rect 43235 74321 43349 74479
tri 43385 74446 43401 74462 se
rect 43401 74446 43478 74462
rect 43385 74380 43478 74446
rect 43106 74245 43478 74321
rect 43106 74120 43199 74186
rect 43106 74104 43183 74120
tri 43183 74104 43199 74120 nw
rect 43235 74087 43349 74245
rect 43385 74120 43478 74186
tri 43385 74104 43401 74120 ne
rect 43401 74104 43478 74120
rect 43218 74005 43366 74087
rect 43106 73972 43183 73988
tri 43183 73972 43199 73988 sw
rect 43106 73906 43199 73972
rect 43106 73804 43199 73870
rect 43106 73788 43183 73804
tri 43183 73788 43199 73804 nw
rect 43235 73771 43349 74005
tri 43385 73972 43401 73988 se
rect 43401 73972 43478 73988
rect 43385 73906 43478 73972
rect 43385 73804 43478 73870
tri 43385 73788 43401 73804 ne
rect 43401 73788 43478 73804
rect 43218 73689 43366 73771
rect 43106 73656 43183 73672
tri 43183 73656 43199 73672 sw
rect 43106 73590 43199 73656
rect 43235 73531 43349 73689
tri 43385 73656 43401 73672 se
rect 43401 73656 43478 73672
rect 43385 73590 43478 73656
rect 43106 73455 43478 73531
rect 43106 73330 43199 73396
rect 43106 73314 43183 73330
tri 43183 73314 43199 73330 nw
rect 43235 73297 43349 73455
rect 43385 73330 43478 73396
tri 43385 73314 43401 73330 ne
rect 43401 73314 43478 73330
rect 43218 73215 43366 73297
rect 43106 73182 43183 73198
tri 43183 73182 43199 73198 sw
rect 43106 73116 43199 73182
rect 43106 73014 43199 73080
rect 43106 72998 43183 73014
tri 43183 72998 43199 73014 nw
rect 43235 72981 43349 73215
tri 43385 73182 43401 73198 se
rect 43401 73182 43478 73198
rect 43385 73116 43478 73182
rect 43385 73014 43478 73080
tri 43385 72998 43401 73014 ne
rect 43401 72998 43478 73014
rect 43218 72899 43366 72981
rect 43106 72866 43183 72882
tri 43183 72866 43199 72882 sw
rect 43106 72800 43199 72866
rect 43235 72741 43349 72899
tri 43385 72866 43401 72882 se
rect 43401 72866 43478 72882
rect 43385 72800 43478 72866
rect 43106 72665 43478 72741
rect 43106 72540 43199 72606
rect 43106 72524 43183 72540
tri 43183 72524 43199 72540 nw
rect 43235 72507 43349 72665
rect 43385 72540 43478 72606
tri 43385 72524 43401 72540 ne
rect 43401 72524 43478 72540
rect 43218 72425 43366 72507
rect 43106 72392 43183 72408
tri 43183 72392 43199 72408 sw
rect 43106 72326 43199 72392
rect 43106 72224 43199 72290
rect 43106 72208 43183 72224
tri 43183 72208 43199 72224 nw
rect 43235 72191 43349 72425
tri 43385 72392 43401 72408 se
rect 43401 72392 43478 72408
rect 43385 72326 43478 72392
rect 43385 72224 43478 72290
tri 43385 72208 43401 72224 ne
rect 43401 72208 43478 72224
rect 43218 72109 43366 72191
rect 43106 72076 43183 72092
tri 43183 72076 43199 72092 sw
rect 43106 72010 43199 72076
rect 43235 71951 43349 72109
tri 43385 72076 43401 72092 se
rect 43401 72076 43478 72092
rect 43385 72010 43478 72076
rect 43106 71875 43478 71951
rect 43106 71750 43199 71816
rect 43106 71734 43183 71750
tri 43183 71734 43199 71750 nw
rect 43235 71717 43349 71875
rect 43385 71750 43478 71816
tri 43385 71734 43401 71750 ne
rect 43401 71734 43478 71750
rect 43218 71635 43366 71717
rect 43106 71602 43183 71618
tri 43183 71602 43199 71618 sw
rect 43106 71536 43199 71602
rect 43106 71434 43199 71500
rect 43106 71418 43183 71434
tri 43183 71418 43199 71434 nw
rect 43235 71401 43349 71635
tri 43385 71602 43401 71618 se
rect 43401 71602 43478 71618
rect 43385 71536 43478 71602
rect 43385 71434 43478 71500
tri 43385 71418 43401 71434 ne
rect 43401 71418 43478 71434
rect 43218 71319 43366 71401
rect 43106 71286 43183 71302
tri 43183 71286 43199 71302 sw
rect 43106 71220 43199 71286
rect 43235 71161 43349 71319
tri 43385 71286 43401 71302 se
rect 43401 71286 43478 71302
rect 43385 71220 43478 71286
rect 43106 71085 43478 71161
rect 43106 70960 43199 71026
rect 43106 70944 43183 70960
tri 43183 70944 43199 70960 nw
rect 43235 70927 43349 71085
rect 43385 70960 43478 71026
tri 43385 70944 43401 70960 ne
rect 43401 70944 43478 70960
rect 43218 70845 43366 70927
rect 43106 70812 43183 70828
tri 43183 70812 43199 70828 sw
rect 43106 70746 43199 70812
rect 43106 70644 43199 70710
rect 43106 70628 43183 70644
tri 43183 70628 43199 70644 nw
rect 43235 70611 43349 70845
tri 43385 70812 43401 70828 se
rect 43401 70812 43478 70828
rect 43385 70746 43478 70812
rect 43385 70644 43478 70710
tri 43385 70628 43401 70644 ne
rect 43401 70628 43478 70644
rect 43218 70529 43366 70611
rect 43106 70496 43183 70512
tri 43183 70496 43199 70512 sw
rect 43106 70430 43199 70496
rect 43235 70371 43349 70529
tri 43385 70496 43401 70512 se
rect 43401 70496 43478 70512
rect 43385 70430 43478 70496
rect 43106 70295 43478 70371
rect 43106 70170 43199 70236
rect 43106 70154 43183 70170
tri 43183 70154 43199 70170 nw
rect 43235 70137 43349 70295
rect 43385 70170 43478 70236
tri 43385 70154 43401 70170 ne
rect 43401 70154 43478 70170
rect 43218 70055 43366 70137
rect 43106 70022 43183 70038
tri 43183 70022 43199 70038 sw
rect 43106 69956 43199 70022
rect 43106 69854 43199 69920
rect 43106 69838 43183 69854
tri 43183 69838 43199 69854 nw
rect 43235 69821 43349 70055
tri 43385 70022 43401 70038 se
rect 43401 70022 43478 70038
rect 43385 69956 43478 70022
rect 43385 69854 43478 69920
tri 43385 69838 43401 69854 ne
rect 43401 69838 43478 69854
rect 43218 69739 43366 69821
rect 43106 69706 43183 69722
tri 43183 69706 43199 69722 sw
rect 43106 69640 43199 69706
rect 43235 69581 43349 69739
tri 43385 69706 43401 69722 se
rect 43401 69706 43478 69722
rect 43385 69640 43478 69706
rect 43106 69505 43478 69581
rect 43106 69380 43199 69446
rect 43106 69364 43183 69380
tri 43183 69364 43199 69380 nw
rect 43235 69347 43349 69505
rect 43385 69380 43478 69446
tri 43385 69364 43401 69380 ne
rect 43401 69364 43478 69380
rect 43218 69265 43366 69347
rect 43106 69232 43183 69248
tri 43183 69232 43199 69248 sw
rect 43106 69166 43199 69232
rect 43106 69064 43199 69130
rect 43106 69048 43183 69064
tri 43183 69048 43199 69064 nw
rect 43235 69031 43349 69265
tri 43385 69232 43401 69248 se
rect 43401 69232 43478 69248
rect 43385 69166 43478 69232
rect 43385 69064 43478 69130
tri 43385 69048 43401 69064 ne
rect 43401 69048 43478 69064
rect 43218 68949 43366 69031
rect 43106 68916 43183 68932
tri 43183 68916 43199 68932 sw
rect 43106 68850 43199 68916
rect 43235 68791 43349 68949
tri 43385 68916 43401 68932 se
rect 43401 68916 43478 68932
rect 43385 68850 43478 68916
rect 43106 68715 43478 68791
rect 43106 68590 43199 68656
rect 43106 68574 43183 68590
tri 43183 68574 43199 68590 nw
rect 43235 68557 43349 68715
rect 43385 68590 43478 68656
tri 43385 68574 43401 68590 ne
rect 43401 68574 43478 68590
rect 43218 68475 43366 68557
rect 43106 68442 43183 68458
tri 43183 68442 43199 68458 sw
rect 43106 68376 43199 68442
rect 43106 68274 43199 68340
rect 43106 68258 43183 68274
tri 43183 68258 43199 68274 nw
rect 43235 68241 43349 68475
tri 43385 68442 43401 68458 se
rect 43401 68442 43478 68458
rect 43385 68376 43478 68442
rect 43385 68274 43478 68340
tri 43385 68258 43401 68274 ne
rect 43401 68258 43478 68274
rect 43218 68159 43366 68241
rect 43106 68126 43183 68142
tri 43183 68126 43199 68142 sw
rect 43106 68060 43199 68126
rect 43235 68001 43349 68159
tri 43385 68126 43401 68142 se
rect 43401 68126 43478 68142
rect 43385 68060 43478 68126
rect 43106 67925 43478 68001
rect 43106 67800 43199 67866
rect 43106 67784 43183 67800
tri 43183 67784 43199 67800 nw
rect 43235 67767 43349 67925
rect 43385 67800 43478 67866
tri 43385 67784 43401 67800 ne
rect 43401 67784 43478 67800
rect 43218 67685 43366 67767
rect 43106 67652 43183 67668
tri 43183 67652 43199 67668 sw
rect 43106 67586 43199 67652
rect 43106 67484 43199 67550
rect 43106 67468 43183 67484
tri 43183 67468 43199 67484 nw
rect 43235 67451 43349 67685
tri 43385 67652 43401 67668 se
rect 43401 67652 43478 67668
rect 43385 67586 43478 67652
rect 43385 67484 43478 67550
tri 43385 67468 43401 67484 ne
rect 43401 67468 43478 67484
rect 43218 67369 43366 67451
rect 43106 67336 43183 67352
tri 43183 67336 43199 67352 sw
rect 43106 67270 43199 67336
rect 43235 67211 43349 67369
tri 43385 67336 43401 67352 se
rect 43401 67336 43478 67352
rect 43385 67270 43478 67336
rect 43106 67135 43478 67211
rect 43106 67010 43199 67076
rect 43106 66994 43183 67010
tri 43183 66994 43199 67010 nw
rect 43235 66977 43349 67135
rect 43385 67010 43478 67076
tri 43385 66994 43401 67010 ne
rect 43401 66994 43478 67010
rect 43218 66895 43366 66977
rect 43106 66862 43183 66878
tri 43183 66862 43199 66878 sw
rect 43106 66796 43199 66862
rect 43106 66694 43199 66760
rect 43106 66678 43183 66694
tri 43183 66678 43199 66694 nw
rect 43235 66661 43349 66895
tri 43385 66862 43401 66878 se
rect 43401 66862 43478 66878
rect 43385 66796 43478 66862
rect 43385 66694 43478 66760
tri 43385 66678 43401 66694 ne
rect 43401 66678 43478 66694
rect 43218 66579 43366 66661
rect 43106 66546 43183 66562
tri 43183 66546 43199 66562 sw
rect 43106 66480 43199 66546
rect 43235 66421 43349 66579
tri 43385 66546 43401 66562 se
rect 43401 66546 43478 66562
rect 43385 66480 43478 66546
rect 43106 66345 43478 66421
rect 43106 66220 43199 66286
rect 43106 66204 43183 66220
tri 43183 66204 43199 66220 nw
rect 43235 66187 43349 66345
rect 43385 66220 43478 66286
tri 43385 66204 43401 66220 ne
rect 43401 66204 43478 66220
rect 43218 66105 43366 66187
rect 43106 66072 43183 66088
tri 43183 66072 43199 66088 sw
rect 43106 66006 43199 66072
rect 43106 65904 43199 65970
rect 43106 65888 43183 65904
tri 43183 65888 43199 65904 nw
rect 43235 65871 43349 66105
tri 43385 66072 43401 66088 se
rect 43401 66072 43478 66088
rect 43385 66006 43478 66072
rect 43385 65904 43478 65970
tri 43385 65888 43401 65904 ne
rect 43401 65888 43478 65904
rect 43218 65789 43366 65871
rect 43106 65756 43183 65772
tri 43183 65756 43199 65772 sw
rect 43106 65690 43199 65756
rect 43235 65631 43349 65789
tri 43385 65756 43401 65772 se
rect 43401 65756 43478 65772
rect 43385 65690 43478 65756
rect 43106 65555 43478 65631
rect 43106 65430 43199 65496
rect 43106 65414 43183 65430
tri 43183 65414 43199 65430 nw
rect 43235 65397 43349 65555
rect 43385 65430 43478 65496
tri 43385 65414 43401 65430 ne
rect 43401 65414 43478 65430
rect 43218 65315 43366 65397
rect 43106 65282 43183 65298
tri 43183 65282 43199 65298 sw
rect 43106 65216 43199 65282
rect 43106 65114 43199 65180
rect 43106 65098 43183 65114
tri 43183 65098 43199 65114 nw
rect 43235 65081 43349 65315
tri 43385 65282 43401 65298 se
rect 43401 65282 43478 65298
rect 43385 65216 43478 65282
rect 43385 65114 43478 65180
tri 43385 65098 43401 65114 ne
rect 43401 65098 43478 65114
rect 43218 64999 43366 65081
rect 43106 64966 43183 64982
tri 43183 64966 43199 64982 sw
rect 43106 64900 43199 64966
rect 43235 64841 43349 64999
tri 43385 64966 43401 64982 se
rect 43401 64966 43478 64982
rect 43385 64900 43478 64966
rect 43106 64765 43478 64841
rect 43106 64640 43199 64706
rect 43106 64624 43183 64640
tri 43183 64624 43199 64640 nw
rect 43235 64607 43349 64765
rect 43385 64640 43478 64706
tri 43385 64624 43401 64640 ne
rect 43401 64624 43478 64640
rect 43218 64525 43366 64607
rect 43106 64492 43183 64508
tri 43183 64492 43199 64508 sw
rect 43106 64426 43199 64492
rect 43106 64324 43199 64390
rect 43106 64308 43183 64324
tri 43183 64308 43199 64324 nw
rect 43235 64291 43349 64525
tri 43385 64492 43401 64508 se
rect 43401 64492 43478 64508
rect 43385 64426 43478 64492
rect 43385 64324 43478 64390
tri 43385 64308 43401 64324 ne
rect 43401 64308 43478 64324
rect 43218 64209 43366 64291
rect 43106 64176 43183 64192
tri 43183 64176 43199 64192 sw
rect 43106 64110 43199 64176
rect 43235 64051 43349 64209
tri 43385 64176 43401 64192 se
rect 43401 64176 43478 64192
rect 43385 64110 43478 64176
rect 43106 63975 43478 64051
rect 43106 63850 43199 63916
rect 43106 63834 43183 63850
tri 43183 63834 43199 63850 nw
rect 43235 63817 43349 63975
rect 43385 63850 43478 63916
tri 43385 63834 43401 63850 ne
rect 43401 63834 43478 63850
rect 43218 63735 43366 63817
rect 43106 63702 43183 63718
tri 43183 63702 43199 63718 sw
rect 43106 63636 43199 63702
rect 43106 63534 43199 63600
rect 43106 63518 43183 63534
tri 43183 63518 43199 63534 nw
rect 43235 63501 43349 63735
tri 43385 63702 43401 63718 se
rect 43401 63702 43478 63718
rect 43385 63636 43478 63702
rect 43385 63534 43478 63600
tri 43385 63518 43401 63534 ne
rect 43401 63518 43478 63534
rect 43218 63419 43366 63501
rect 43106 63386 43183 63402
tri 43183 63386 43199 63402 sw
rect 43106 63320 43199 63386
rect 43235 63261 43349 63419
tri 43385 63386 43401 63402 se
rect 43401 63386 43478 63402
rect 43385 63320 43478 63386
rect 43106 63185 43478 63261
rect 43106 63060 43199 63126
rect 43106 63044 43183 63060
tri 43183 63044 43199 63060 nw
rect 43235 63027 43349 63185
rect 43385 63060 43478 63126
tri 43385 63044 43401 63060 ne
rect 43401 63044 43478 63060
rect 43218 62945 43366 63027
rect 43106 62912 43183 62928
tri 43183 62912 43199 62928 sw
rect 43106 62846 43199 62912
rect 43106 62744 43199 62810
rect 43106 62728 43183 62744
tri 43183 62728 43199 62744 nw
rect 43235 62711 43349 62945
tri 43385 62912 43401 62928 se
rect 43401 62912 43478 62928
rect 43385 62846 43478 62912
rect 43385 62744 43478 62810
tri 43385 62728 43401 62744 ne
rect 43401 62728 43478 62744
rect 43218 62629 43366 62711
rect 43106 62596 43183 62612
tri 43183 62596 43199 62612 sw
rect 43106 62530 43199 62596
rect 43235 62471 43349 62629
tri 43385 62596 43401 62612 se
rect 43401 62596 43478 62612
rect 43385 62530 43478 62596
rect 43106 62395 43478 62471
rect 43106 62270 43199 62336
rect 43106 62254 43183 62270
tri 43183 62254 43199 62270 nw
rect 43235 62237 43349 62395
rect 43385 62270 43478 62336
tri 43385 62254 43401 62270 ne
rect 43401 62254 43478 62270
rect 43218 62155 43366 62237
rect 43106 62122 43183 62138
tri 43183 62122 43199 62138 sw
rect 43106 62056 43199 62122
rect 43106 61954 43199 62020
rect 43106 61938 43183 61954
tri 43183 61938 43199 61954 nw
rect 43235 61921 43349 62155
tri 43385 62122 43401 62138 se
rect 43401 62122 43478 62138
rect 43385 62056 43478 62122
rect 43385 61954 43478 62020
tri 43385 61938 43401 61954 ne
rect 43401 61938 43478 61954
rect 43218 61839 43366 61921
rect 43106 61806 43183 61822
tri 43183 61806 43199 61822 sw
rect 43106 61740 43199 61806
rect 43235 61681 43349 61839
tri 43385 61806 43401 61822 se
rect 43401 61806 43478 61822
rect 43385 61740 43478 61806
rect 43106 61605 43478 61681
rect 43106 61480 43199 61546
rect 43106 61464 43183 61480
tri 43183 61464 43199 61480 nw
rect 43235 61447 43349 61605
rect 43385 61480 43478 61546
tri 43385 61464 43401 61480 ne
rect 43401 61464 43478 61480
rect 43218 61365 43366 61447
rect 43106 61332 43183 61348
tri 43183 61332 43199 61348 sw
rect 43106 61266 43199 61332
rect 43106 61164 43199 61230
rect 43106 61148 43183 61164
tri 43183 61148 43199 61164 nw
rect 43235 61131 43349 61365
tri 43385 61332 43401 61348 se
rect 43401 61332 43478 61348
rect 43385 61266 43478 61332
rect 43385 61164 43478 61230
tri 43385 61148 43401 61164 ne
rect 43401 61148 43478 61164
rect 43218 61049 43366 61131
rect 43106 61016 43183 61032
tri 43183 61016 43199 61032 sw
rect 43106 60950 43199 61016
rect 43235 60891 43349 61049
tri 43385 61016 43401 61032 se
rect 43401 61016 43478 61032
rect 43385 60950 43478 61016
rect 43106 60815 43478 60891
rect 43106 60690 43199 60756
rect 43106 60674 43183 60690
tri 43183 60674 43199 60690 nw
rect 43235 60657 43349 60815
rect 43385 60690 43478 60756
tri 43385 60674 43401 60690 ne
rect 43401 60674 43478 60690
rect 43218 60575 43366 60657
rect 43106 60542 43183 60558
tri 43183 60542 43199 60558 sw
rect 43106 60476 43199 60542
rect 43106 60374 43199 60440
rect 43106 60358 43183 60374
tri 43183 60358 43199 60374 nw
rect 43235 60341 43349 60575
tri 43385 60542 43401 60558 se
rect 43401 60542 43478 60558
rect 43385 60476 43478 60542
rect 43385 60374 43478 60440
tri 43385 60358 43401 60374 ne
rect 43401 60358 43478 60374
rect 43218 60259 43366 60341
rect 43106 60226 43183 60242
tri 43183 60226 43199 60242 sw
rect 43106 60160 43199 60226
rect 43235 60101 43349 60259
tri 43385 60226 43401 60242 se
rect 43401 60226 43478 60242
rect 43385 60160 43478 60226
rect 43106 60025 43478 60101
rect 43106 59900 43199 59966
rect 43106 59884 43183 59900
tri 43183 59884 43199 59900 nw
rect 43235 59867 43349 60025
rect 43385 59900 43478 59966
tri 43385 59884 43401 59900 ne
rect 43401 59884 43478 59900
rect 43218 59785 43366 59867
rect 43106 59752 43183 59768
tri 43183 59752 43199 59768 sw
rect 43106 59686 43199 59752
rect 43106 59584 43199 59650
rect 43106 59568 43183 59584
tri 43183 59568 43199 59584 nw
rect 43235 59551 43349 59785
tri 43385 59752 43401 59768 se
rect 43401 59752 43478 59768
rect 43385 59686 43478 59752
rect 43385 59584 43478 59650
tri 43385 59568 43401 59584 ne
rect 43401 59568 43478 59584
rect 43218 59469 43366 59551
rect 43106 59436 43183 59452
tri 43183 59436 43199 59452 sw
rect 43106 59370 43199 59436
rect 43235 59311 43349 59469
tri 43385 59436 43401 59452 se
rect 43401 59436 43478 59452
rect 43385 59370 43478 59436
rect 43106 59235 43478 59311
rect 43106 59110 43199 59176
rect 43106 59094 43183 59110
tri 43183 59094 43199 59110 nw
rect 43235 59077 43349 59235
rect 43385 59110 43478 59176
tri 43385 59094 43401 59110 ne
rect 43401 59094 43478 59110
rect 43218 58995 43366 59077
rect 43106 58962 43183 58978
tri 43183 58962 43199 58978 sw
rect 43106 58896 43199 58962
rect 43106 58794 43199 58860
rect 43106 58778 43183 58794
tri 43183 58778 43199 58794 nw
rect 43235 58761 43349 58995
tri 43385 58962 43401 58978 se
rect 43401 58962 43478 58978
rect 43385 58896 43478 58962
rect 43385 58794 43478 58860
tri 43385 58778 43401 58794 ne
rect 43401 58778 43478 58794
rect 43218 58679 43366 58761
rect 43106 58646 43183 58662
tri 43183 58646 43199 58662 sw
rect 43106 58580 43199 58646
rect 43235 58521 43349 58679
tri 43385 58646 43401 58662 se
rect 43401 58646 43478 58662
rect 43385 58580 43478 58646
rect 43106 58445 43478 58521
rect 43106 58320 43199 58386
rect 43106 58304 43183 58320
tri 43183 58304 43199 58320 nw
rect 43235 58287 43349 58445
rect 43385 58320 43478 58386
tri 43385 58304 43401 58320 ne
rect 43401 58304 43478 58320
rect 43218 58205 43366 58287
rect 43106 58172 43183 58188
tri 43183 58172 43199 58188 sw
rect 43106 58106 43199 58172
rect 43106 58004 43199 58070
rect 43106 57988 43183 58004
tri 43183 57988 43199 58004 nw
rect 43235 57971 43349 58205
tri 43385 58172 43401 58188 se
rect 43401 58172 43478 58188
rect 43385 58106 43478 58172
rect 43385 58004 43478 58070
tri 43385 57988 43401 58004 ne
rect 43401 57988 43478 58004
rect 43218 57889 43366 57971
rect 43106 57856 43183 57872
tri 43183 57856 43199 57872 sw
rect 43106 57790 43199 57856
rect 43235 57731 43349 57889
tri 43385 57856 43401 57872 se
rect 43401 57856 43478 57872
rect 43385 57790 43478 57856
rect 43106 57655 43478 57731
rect 43106 57530 43199 57596
rect 43106 57514 43183 57530
tri 43183 57514 43199 57530 nw
rect 43235 57497 43349 57655
rect 43385 57530 43478 57596
tri 43385 57514 43401 57530 ne
rect 43401 57514 43478 57530
rect 43218 57415 43366 57497
rect 43106 57382 43183 57398
tri 43183 57382 43199 57398 sw
rect 43106 57316 43199 57382
rect 43106 57214 43199 57280
rect 43106 57198 43183 57214
tri 43183 57198 43199 57214 nw
rect 43235 57181 43349 57415
tri 43385 57382 43401 57398 se
rect 43401 57382 43478 57398
rect 43385 57316 43478 57382
rect 43385 57214 43478 57280
tri 43385 57198 43401 57214 ne
rect 43401 57198 43478 57214
rect 43218 57099 43366 57181
rect 43106 57066 43183 57082
tri 43183 57066 43199 57082 sw
rect 43106 57000 43199 57066
rect 43235 56941 43349 57099
tri 43385 57066 43401 57082 se
rect 43401 57066 43478 57082
rect 43385 57000 43478 57066
rect 43106 56865 43478 56941
rect 43106 56740 43199 56806
rect 43106 56724 43183 56740
tri 43183 56724 43199 56740 nw
rect 43235 56707 43349 56865
rect 43385 56740 43478 56806
tri 43385 56724 43401 56740 ne
rect 43401 56724 43478 56740
rect 43218 56625 43366 56707
rect 43106 56592 43183 56608
tri 43183 56592 43199 56608 sw
rect 43106 56526 43199 56592
rect 43106 56424 43199 56490
rect 43106 56408 43183 56424
tri 43183 56408 43199 56424 nw
rect 43235 56391 43349 56625
tri 43385 56592 43401 56608 se
rect 43401 56592 43478 56608
rect 43385 56526 43478 56592
rect 43385 56424 43478 56490
tri 43385 56408 43401 56424 ne
rect 43401 56408 43478 56424
rect 43218 56309 43366 56391
rect 43106 56276 43183 56292
tri 43183 56276 43199 56292 sw
rect 43106 56210 43199 56276
rect 43235 56151 43349 56309
tri 43385 56276 43401 56292 se
rect 43401 56276 43478 56292
rect 43385 56210 43478 56276
rect 43106 56075 43478 56151
rect 43106 55950 43199 56016
rect 43106 55934 43183 55950
tri 43183 55934 43199 55950 nw
rect 43235 55917 43349 56075
rect 43385 55950 43478 56016
tri 43385 55934 43401 55950 ne
rect 43401 55934 43478 55950
rect 43218 55835 43366 55917
rect 43106 55802 43183 55818
tri 43183 55802 43199 55818 sw
rect 43106 55736 43199 55802
rect 43106 55634 43199 55700
rect 43106 55618 43183 55634
tri 43183 55618 43199 55634 nw
rect 43235 55601 43349 55835
tri 43385 55802 43401 55818 se
rect 43401 55802 43478 55818
rect 43385 55736 43478 55802
rect 43385 55634 43478 55700
tri 43385 55618 43401 55634 ne
rect 43401 55618 43478 55634
rect 43218 55519 43366 55601
rect 43106 55486 43183 55502
tri 43183 55486 43199 55502 sw
rect 43106 55420 43199 55486
rect 43235 55361 43349 55519
tri 43385 55486 43401 55502 se
rect 43401 55486 43478 55502
rect 43385 55420 43478 55486
rect 43106 55285 43478 55361
rect 43106 55160 43199 55226
rect 43106 55144 43183 55160
tri 43183 55144 43199 55160 nw
rect 43235 55127 43349 55285
rect 43385 55160 43478 55226
tri 43385 55144 43401 55160 ne
rect 43401 55144 43478 55160
rect 43218 55045 43366 55127
rect 43106 55012 43183 55028
tri 43183 55012 43199 55028 sw
rect 43106 54946 43199 55012
rect 43106 54844 43199 54910
rect 43106 54828 43183 54844
tri 43183 54828 43199 54844 nw
rect 43235 54811 43349 55045
tri 43385 55012 43401 55028 se
rect 43401 55012 43478 55028
rect 43385 54946 43478 55012
rect 43385 54844 43478 54910
tri 43385 54828 43401 54844 ne
rect 43401 54828 43478 54844
rect 43218 54729 43366 54811
rect 43106 54696 43183 54712
tri 43183 54696 43199 54712 sw
rect 43106 54630 43199 54696
rect 43235 54571 43349 54729
tri 43385 54696 43401 54712 se
rect 43401 54696 43478 54712
rect 43385 54630 43478 54696
rect 43106 54495 43478 54571
rect 43106 54370 43199 54436
rect 43106 54354 43183 54370
tri 43183 54354 43199 54370 nw
rect 43235 54337 43349 54495
rect 43385 54370 43478 54436
tri 43385 54354 43401 54370 ne
rect 43401 54354 43478 54370
rect 43218 54255 43366 54337
rect 43106 54222 43183 54238
tri 43183 54222 43199 54238 sw
rect 43106 54156 43199 54222
rect 43106 54054 43199 54120
rect 43106 54038 43183 54054
tri 43183 54038 43199 54054 nw
rect 43235 54021 43349 54255
tri 43385 54222 43401 54238 se
rect 43401 54222 43478 54238
rect 43385 54156 43478 54222
rect 43385 54054 43478 54120
tri 43385 54038 43401 54054 ne
rect 43401 54038 43478 54054
rect 43218 53939 43366 54021
rect 43106 53906 43183 53922
tri 43183 53906 43199 53922 sw
rect 43106 53840 43199 53906
rect 43235 53781 43349 53939
tri 43385 53906 43401 53922 se
rect 43401 53906 43478 53922
rect 43385 53840 43478 53906
rect 43106 53705 43478 53781
rect 43106 53580 43199 53646
rect 43106 53564 43183 53580
tri 43183 53564 43199 53580 nw
rect 43235 53547 43349 53705
rect 43385 53580 43478 53646
tri 43385 53564 43401 53580 ne
rect 43401 53564 43478 53580
rect 43218 53465 43366 53547
rect 43106 53432 43183 53448
tri 43183 53432 43199 53448 sw
rect 43106 53366 43199 53432
rect 43106 53264 43199 53330
rect 43106 53248 43183 53264
tri 43183 53248 43199 53264 nw
rect 43235 53231 43349 53465
tri 43385 53432 43401 53448 se
rect 43401 53432 43478 53448
rect 43385 53366 43478 53432
rect 43385 53264 43478 53330
tri 43385 53248 43401 53264 ne
rect 43401 53248 43478 53264
rect 43218 53149 43366 53231
rect 43106 53116 43183 53132
tri 43183 53116 43199 53132 sw
rect 43106 53050 43199 53116
rect 43235 52991 43349 53149
tri 43385 53116 43401 53132 se
rect 43401 53116 43478 53132
rect 43385 53050 43478 53116
rect 43106 52915 43478 52991
rect 43106 52790 43199 52856
rect 43106 52774 43183 52790
tri 43183 52774 43199 52790 nw
rect 43235 52757 43349 52915
rect 43385 52790 43478 52856
tri 43385 52774 43401 52790 ne
rect 43401 52774 43478 52790
rect 43218 52675 43366 52757
rect 43106 52642 43183 52658
tri 43183 52642 43199 52658 sw
rect 43106 52576 43199 52642
rect 43106 52474 43199 52540
rect 43106 52458 43183 52474
tri 43183 52458 43199 52474 nw
rect 43235 52441 43349 52675
tri 43385 52642 43401 52658 se
rect 43401 52642 43478 52658
rect 43385 52576 43478 52642
rect 43385 52474 43478 52540
tri 43385 52458 43401 52474 ne
rect 43401 52458 43478 52474
rect 43218 52359 43366 52441
rect 43106 52326 43183 52342
tri 43183 52326 43199 52342 sw
rect 43106 52260 43199 52326
rect 43235 52201 43349 52359
tri 43385 52326 43401 52342 se
rect 43401 52326 43478 52342
rect 43385 52260 43478 52326
rect 43106 52125 43478 52201
rect 43106 52000 43199 52066
rect 43106 51984 43183 52000
tri 43183 51984 43199 52000 nw
rect 43235 51967 43349 52125
rect 43385 52000 43478 52066
tri 43385 51984 43401 52000 ne
rect 43401 51984 43478 52000
rect 43218 51885 43366 51967
rect 43106 51852 43183 51868
tri 43183 51852 43199 51868 sw
rect 43106 51786 43199 51852
rect 43106 51684 43199 51750
rect 43106 51668 43183 51684
tri 43183 51668 43199 51684 nw
rect 43235 51651 43349 51885
tri 43385 51852 43401 51868 se
rect 43401 51852 43478 51868
rect 43385 51786 43478 51852
rect 43385 51684 43478 51750
tri 43385 51668 43401 51684 ne
rect 43401 51668 43478 51684
rect 43218 51569 43366 51651
rect 43106 51536 43183 51552
tri 43183 51536 43199 51552 sw
rect 43106 51470 43199 51536
rect 43235 51411 43349 51569
tri 43385 51536 43401 51552 se
rect 43401 51536 43478 51552
rect 43385 51470 43478 51536
rect 43106 51335 43478 51411
rect 43106 51210 43199 51276
rect 43106 51194 43183 51210
tri 43183 51194 43199 51210 nw
rect 43235 51177 43349 51335
rect 43385 51210 43478 51276
tri 43385 51194 43401 51210 ne
rect 43401 51194 43478 51210
rect 43218 51095 43366 51177
rect 43106 51062 43183 51078
tri 43183 51062 43199 51078 sw
rect 43106 50996 43199 51062
rect 43106 50894 43199 50960
rect 43106 50878 43183 50894
tri 43183 50878 43199 50894 nw
rect 43235 50861 43349 51095
tri 43385 51062 43401 51078 se
rect 43401 51062 43478 51078
rect 43385 50996 43478 51062
rect 43385 50894 43478 50960
tri 43385 50878 43401 50894 ne
rect 43401 50878 43478 50894
rect 43218 50779 43366 50861
rect 43106 50746 43183 50762
tri 43183 50746 43199 50762 sw
rect 43106 50680 43199 50746
rect 43235 50621 43349 50779
tri 43385 50746 43401 50762 se
rect 43401 50746 43478 50762
rect 43385 50680 43478 50746
rect 43106 50545 43478 50621
rect 43106 50420 43199 50486
rect 43106 50404 43183 50420
tri 43183 50404 43199 50420 nw
rect 43235 50387 43349 50545
rect 43385 50420 43478 50486
tri 43385 50404 43401 50420 ne
rect 43401 50404 43478 50420
rect 43218 50305 43366 50387
rect 43106 50272 43183 50288
tri 43183 50272 43199 50288 sw
rect 43106 50206 43199 50272
rect 43106 50104 43199 50170
rect 43106 50088 43183 50104
tri 43183 50088 43199 50104 nw
rect 43235 50071 43349 50305
tri 43385 50272 43401 50288 se
rect 43401 50272 43478 50288
rect 43385 50206 43478 50272
rect 43385 50104 43478 50170
tri 43385 50088 43401 50104 ne
rect 43401 50088 43478 50104
rect 43218 49989 43366 50071
rect 43106 49956 43183 49972
tri 43183 49956 43199 49972 sw
rect 43106 49890 43199 49956
rect 43235 49831 43349 49989
tri 43385 49956 43401 49972 se
rect 43401 49956 43478 49972
rect 43385 49890 43478 49956
rect 43106 49755 43478 49831
rect 43106 49630 43199 49696
rect 43106 49614 43183 49630
tri 43183 49614 43199 49630 nw
rect 43235 49597 43349 49755
rect 43385 49630 43478 49696
tri 43385 49614 43401 49630 ne
rect 43401 49614 43478 49630
rect 43218 49515 43366 49597
rect 43106 49482 43183 49498
tri 43183 49482 43199 49498 sw
rect 43106 49416 43199 49482
rect 43106 49314 43199 49380
rect 43106 49298 43183 49314
tri 43183 49298 43199 49314 nw
rect 43235 49281 43349 49515
tri 43385 49482 43401 49498 se
rect 43401 49482 43478 49498
rect 43385 49416 43478 49482
rect 43385 49314 43478 49380
tri 43385 49298 43401 49314 ne
rect 43401 49298 43478 49314
rect 43218 49199 43366 49281
rect 43106 49166 43183 49182
tri 43183 49166 43199 49182 sw
rect 43106 49100 43199 49166
rect 43235 49041 43349 49199
tri 43385 49166 43401 49182 se
rect 43401 49166 43478 49182
rect 43385 49100 43478 49166
rect 43106 48965 43478 49041
rect 43106 48840 43199 48906
rect 43106 48824 43183 48840
tri 43183 48824 43199 48840 nw
rect 43235 48807 43349 48965
rect 43385 48840 43478 48906
tri 43385 48824 43401 48840 ne
rect 43401 48824 43478 48840
rect 43218 48725 43366 48807
rect 43106 48692 43183 48708
tri 43183 48692 43199 48708 sw
rect 43106 48626 43199 48692
rect 43106 48524 43199 48590
rect 43106 48508 43183 48524
tri 43183 48508 43199 48524 nw
rect 43235 48491 43349 48725
tri 43385 48692 43401 48708 se
rect 43401 48692 43478 48708
rect 43385 48626 43478 48692
rect 43385 48524 43478 48590
tri 43385 48508 43401 48524 ne
rect 43401 48508 43478 48524
rect 43218 48409 43366 48491
rect 43106 48376 43183 48392
tri 43183 48376 43199 48392 sw
rect 43106 48310 43199 48376
rect 43235 48251 43349 48409
tri 43385 48376 43401 48392 se
rect 43401 48376 43478 48392
rect 43385 48310 43478 48376
rect 43106 48175 43478 48251
rect 43106 48050 43199 48116
rect 43106 48034 43183 48050
tri 43183 48034 43199 48050 nw
rect 43235 48017 43349 48175
rect 43385 48050 43478 48116
tri 43385 48034 43401 48050 ne
rect 43401 48034 43478 48050
rect 43218 47935 43366 48017
rect 43106 47902 43183 47918
tri 43183 47902 43199 47918 sw
rect 43106 47836 43199 47902
rect 43106 47734 43199 47800
rect 43106 47718 43183 47734
tri 43183 47718 43199 47734 nw
rect 43235 47701 43349 47935
tri 43385 47902 43401 47918 se
rect 43401 47902 43478 47918
rect 43385 47836 43478 47902
rect 43385 47734 43478 47800
tri 43385 47718 43401 47734 ne
rect 43401 47718 43478 47734
rect 43218 47619 43366 47701
rect 43106 47586 43183 47602
tri 43183 47586 43199 47602 sw
rect 43106 47520 43199 47586
rect 43235 47461 43349 47619
tri 43385 47586 43401 47602 se
rect 43401 47586 43478 47602
rect 43385 47520 43478 47586
rect 43106 47385 43478 47461
rect 43106 47260 43199 47326
rect 43106 47244 43183 47260
tri 43183 47244 43199 47260 nw
rect 43235 47227 43349 47385
rect 43385 47260 43478 47326
tri 43385 47244 43401 47260 ne
rect 43401 47244 43478 47260
rect 43218 47145 43366 47227
rect 43106 47112 43183 47128
tri 43183 47112 43199 47128 sw
rect 43106 47046 43199 47112
rect 43106 46944 43199 47010
rect 43106 46928 43183 46944
tri 43183 46928 43199 46944 nw
rect 43235 46911 43349 47145
tri 43385 47112 43401 47128 se
rect 43401 47112 43478 47128
rect 43385 47046 43478 47112
rect 43385 46944 43478 47010
tri 43385 46928 43401 46944 ne
rect 43401 46928 43478 46944
rect 43218 46829 43366 46911
rect 43106 46796 43183 46812
tri 43183 46796 43199 46812 sw
rect 43106 46730 43199 46796
rect 43235 46671 43349 46829
tri 43385 46796 43401 46812 se
rect 43401 46796 43478 46812
rect 43385 46730 43478 46796
rect 43106 46595 43478 46671
rect 43106 46470 43199 46536
rect 43106 46454 43183 46470
tri 43183 46454 43199 46470 nw
rect 43235 46437 43349 46595
rect 43385 46470 43478 46536
tri 43385 46454 43401 46470 ne
rect 43401 46454 43478 46470
rect 43218 46355 43366 46437
rect 43106 46322 43183 46338
tri 43183 46322 43199 46338 sw
rect 43106 46256 43199 46322
rect 43106 46154 43199 46220
rect 43106 46138 43183 46154
tri 43183 46138 43199 46154 nw
rect 43235 46121 43349 46355
tri 43385 46322 43401 46338 se
rect 43401 46322 43478 46338
rect 43385 46256 43478 46322
rect 43385 46154 43478 46220
tri 43385 46138 43401 46154 ne
rect 43401 46138 43478 46154
rect 43218 46039 43366 46121
rect 43106 46006 43183 46022
tri 43183 46006 43199 46022 sw
rect 43106 45940 43199 46006
rect 43235 45881 43349 46039
tri 43385 46006 43401 46022 se
rect 43401 46006 43478 46022
rect 43385 45940 43478 46006
rect 43106 45805 43478 45881
rect 43106 45680 43199 45746
rect 43106 45664 43183 45680
tri 43183 45664 43199 45680 nw
rect 43235 45647 43349 45805
rect 43385 45680 43478 45746
tri 43385 45664 43401 45680 ne
rect 43401 45664 43478 45680
rect 43218 45565 43366 45647
rect 43106 45532 43183 45548
tri 43183 45532 43199 45548 sw
rect 43106 45466 43199 45532
rect 43106 45364 43199 45430
rect 43106 45348 43183 45364
tri 43183 45348 43199 45364 nw
rect 43235 45331 43349 45565
tri 43385 45532 43401 45548 se
rect 43401 45532 43478 45548
rect 43385 45466 43478 45532
rect 43385 45364 43478 45430
tri 43385 45348 43401 45364 ne
rect 43401 45348 43478 45364
rect 43218 45249 43366 45331
rect 43106 45216 43183 45232
tri 43183 45216 43199 45232 sw
rect 43106 45150 43199 45216
rect 43235 45091 43349 45249
tri 43385 45216 43401 45232 se
rect 43401 45216 43478 45232
rect 43385 45150 43478 45216
rect 43106 45015 43478 45091
rect 43106 44890 43199 44956
rect 43106 44874 43183 44890
tri 43183 44874 43199 44890 nw
rect 43235 44857 43349 45015
rect 43385 44890 43478 44956
tri 43385 44874 43401 44890 ne
rect 43401 44874 43478 44890
rect 43218 44775 43366 44857
rect 43106 44742 43183 44758
tri 43183 44742 43199 44758 sw
rect 43106 44676 43199 44742
rect 43106 44574 43199 44640
rect 43106 44558 43183 44574
tri 43183 44558 43199 44574 nw
rect 43235 44541 43349 44775
tri 43385 44742 43401 44758 se
rect 43401 44742 43478 44758
rect 43385 44676 43478 44742
rect 43385 44574 43478 44640
tri 43385 44558 43401 44574 ne
rect 43401 44558 43478 44574
rect 43218 44459 43366 44541
rect 43106 44426 43183 44442
tri 43183 44426 43199 44442 sw
rect 43106 44360 43199 44426
rect 43235 44301 43349 44459
tri 43385 44426 43401 44442 se
rect 43401 44426 43478 44442
rect 43385 44360 43478 44426
rect 43106 44225 43478 44301
rect 43106 44100 43199 44166
rect 43106 44084 43183 44100
tri 43183 44084 43199 44100 nw
rect 43235 44067 43349 44225
rect 43385 44100 43478 44166
tri 43385 44084 43401 44100 ne
rect 43401 44084 43478 44100
rect 43218 43985 43366 44067
rect 43106 43952 43183 43968
tri 43183 43952 43199 43968 sw
rect 43106 43886 43199 43952
rect 43106 43784 43199 43850
rect 43106 43768 43183 43784
tri 43183 43768 43199 43784 nw
rect 43235 43751 43349 43985
tri 43385 43952 43401 43968 se
rect 43401 43952 43478 43968
rect 43385 43886 43478 43952
rect 43385 43784 43478 43850
tri 43385 43768 43401 43784 ne
rect 43401 43768 43478 43784
rect 43218 43669 43366 43751
rect 43106 43636 43183 43652
tri 43183 43636 43199 43652 sw
rect 43106 43570 43199 43636
rect 43235 43511 43349 43669
tri 43385 43636 43401 43652 se
rect 43401 43636 43478 43652
rect 43385 43570 43478 43636
rect 43106 43435 43478 43511
rect 43106 43310 43199 43376
rect 43106 43294 43183 43310
tri 43183 43294 43199 43310 nw
rect 43235 43277 43349 43435
rect 43385 43310 43478 43376
tri 43385 43294 43401 43310 ne
rect 43401 43294 43478 43310
rect 43218 43195 43366 43277
rect 43106 43162 43183 43178
tri 43183 43162 43199 43178 sw
rect 43106 43096 43199 43162
rect 43106 42994 43199 43060
rect 43106 42978 43183 42994
tri 43183 42978 43199 42994 nw
rect 43235 42961 43349 43195
tri 43385 43162 43401 43178 se
rect 43401 43162 43478 43178
rect 43385 43096 43478 43162
rect 43385 42994 43478 43060
tri 43385 42978 43401 42994 ne
rect 43401 42978 43478 42994
rect 43218 42879 43366 42961
rect 43106 42846 43183 42862
tri 43183 42846 43199 42862 sw
rect 43106 42780 43199 42846
rect 43235 42721 43349 42879
tri 43385 42846 43401 42862 se
rect 43401 42846 43478 42862
rect 43385 42780 43478 42846
rect 43106 42645 43478 42721
rect 43106 42520 43199 42586
rect 43106 42504 43183 42520
tri 43183 42504 43199 42520 nw
rect 43235 42487 43349 42645
rect 43385 42520 43478 42586
tri 43385 42504 43401 42520 ne
rect 43401 42504 43478 42520
rect 43218 42405 43366 42487
rect 43106 42372 43183 42388
tri 43183 42372 43199 42388 sw
rect 43106 42306 43199 42372
rect 43106 42204 43199 42270
rect 43106 42188 43183 42204
tri 43183 42188 43199 42204 nw
rect 43235 42171 43349 42405
tri 43385 42372 43401 42388 se
rect 43401 42372 43478 42388
rect 43385 42306 43478 42372
rect 43385 42204 43478 42270
tri 43385 42188 43401 42204 ne
rect 43401 42188 43478 42204
rect 43218 42089 43366 42171
rect 43106 42056 43183 42072
tri 43183 42056 43199 42072 sw
rect 43106 41990 43199 42056
rect 43235 41931 43349 42089
tri 43385 42056 43401 42072 se
rect 43401 42056 43478 42072
rect 43385 41990 43478 42056
rect 43106 41855 43478 41931
rect 43106 41730 43199 41796
rect 43106 41714 43183 41730
tri 43183 41714 43199 41730 nw
rect 43235 41697 43349 41855
rect 43385 41730 43478 41796
tri 43385 41714 43401 41730 ne
rect 43401 41714 43478 41730
rect 43218 41615 43366 41697
rect 43106 41582 43183 41598
tri 43183 41582 43199 41598 sw
rect 43106 41516 43199 41582
rect 43106 41414 43199 41480
rect 43106 41398 43183 41414
tri 43183 41398 43199 41414 nw
rect 43235 41381 43349 41615
tri 43385 41582 43401 41598 se
rect 43401 41582 43478 41598
rect 43385 41516 43478 41582
rect 43385 41414 43478 41480
tri 43385 41398 43401 41414 ne
rect 43401 41398 43478 41414
rect 43218 41299 43366 41381
rect 43106 41266 43183 41282
tri 43183 41266 43199 41282 sw
rect 43106 41200 43199 41266
rect 43235 41141 43349 41299
tri 43385 41266 43401 41282 se
rect 43401 41266 43478 41282
rect 43385 41200 43478 41266
rect 43106 41065 43478 41141
rect 43106 40940 43199 41006
rect 43106 40924 43183 40940
tri 43183 40924 43199 40940 nw
rect 43235 40907 43349 41065
rect 43385 40940 43478 41006
tri 43385 40924 43401 40940 ne
rect 43401 40924 43478 40940
rect 43218 40825 43366 40907
rect 43106 40792 43183 40808
tri 43183 40792 43199 40808 sw
rect 43106 40726 43199 40792
rect 43106 40624 43199 40690
rect 43106 40608 43183 40624
tri 43183 40608 43199 40624 nw
rect 43235 40591 43349 40825
tri 43385 40792 43401 40808 se
rect 43401 40792 43478 40808
rect 43385 40726 43478 40792
rect 43385 40624 43478 40690
tri 43385 40608 43401 40624 ne
rect 43401 40608 43478 40624
rect 43218 40509 43366 40591
rect 43106 40476 43183 40492
tri 43183 40476 43199 40492 sw
rect 43106 40410 43199 40476
rect 43235 40351 43349 40509
tri 43385 40476 43401 40492 se
rect 43401 40476 43478 40492
rect 43385 40410 43478 40476
rect 43106 40275 43478 40351
rect 43106 40150 43199 40216
rect 43106 40134 43183 40150
tri 43183 40134 43199 40150 nw
rect 43235 40117 43349 40275
rect 43385 40150 43478 40216
tri 43385 40134 43401 40150 ne
rect 43401 40134 43478 40150
rect 43218 40035 43366 40117
rect 43106 40002 43183 40018
tri 43183 40002 43199 40018 sw
rect 43106 39936 43199 40002
rect 43106 39834 43199 39900
rect 43106 39818 43183 39834
tri 43183 39818 43199 39834 nw
rect 43235 39801 43349 40035
tri 43385 40002 43401 40018 se
rect 43401 40002 43478 40018
rect 43385 39936 43478 40002
rect 43385 39834 43478 39900
tri 43385 39818 43401 39834 ne
rect 43401 39818 43478 39834
rect 43218 39719 43366 39801
rect 43106 39686 43183 39702
tri 43183 39686 43199 39702 sw
rect 43106 39620 43199 39686
rect 43235 39561 43349 39719
tri 43385 39686 43401 39702 se
rect 43401 39686 43478 39702
rect 43385 39620 43478 39686
rect 43106 39485 43478 39561
rect 43106 39360 43199 39426
rect 43106 39344 43183 39360
tri 43183 39344 43199 39360 nw
rect 43235 39327 43349 39485
rect 43385 39360 43478 39426
tri 43385 39344 43401 39360 ne
rect 43401 39344 43478 39360
rect 43218 39245 43366 39327
rect 43106 39212 43183 39228
tri 43183 39212 43199 39228 sw
rect 43106 39146 43199 39212
rect 43106 39044 43199 39110
rect 43106 39028 43183 39044
tri 43183 39028 43199 39044 nw
rect 43235 39011 43349 39245
tri 43385 39212 43401 39228 se
rect 43401 39212 43478 39228
rect 43385 39146 43478 39212
rect 43385 39044 43478 39110
tri 43385 39028 43401 39044 ne
rect 43401 39028 43478 39044
rect 43218 38929 43366 39011
rect 43106 38896 43183 38912
tri 43183 38896 43199 38912 sw
rect 43106 38830 43199 38896
rect 43235 38771 43349 38929
tri 43385 38896 43401 38912 se
rect 43401 38896 43478 38912
rect 43385 38830 43478 38896
rect 43106 38695 43478 38771
rect 43106 38570 43199 38636
rect 43106 38554 43183 38570
tri 43183 38554 43199 38570 nw
rect 43235 38537 43349 38695
rect 43385 38570 43478 38636
tri 43385 38554 43401 38570 ne
rect 43401 38554 43478 38570
rect 43218 38455 43366 38537
rect 43106 38422 43183 38438
tri 43183 38422 43199 38438 sw
rect 43106 38356 43199 38422
rect 43106 38254 43199 38320
rect 43106 38238 43183 38254
tri 43183 38238 43199 38254 nw
rect 43235 38221 43349 38455
tri 43385 38422 43401 38438 se
rect 43401 38422 43478 38438
rect 43385 38356 43478 38422
rect 43385 38254 43478 38320
tri 43385 38238 43401 38254 ne
rect 43401 38238 43478 38254
rect 43218 38139 43366 38221
rect 43106 38106 43183 38122
tri 43183 38106 43199 38122 sw
rect 43106 38040 43199 38106
rect 43235 37981 43349 38139
tri 43385 38106 43401 38122 se
rect 43401 38106 43478 38122
rect 43385 38040 43478 38106
rect 43106 37905 43478 37981
rect 43106 37780 43199 37846
rect 43106 37764 43183 37780
tri 43183 37764 43199 37780 nw
rect 43235 37747 43349 37905
rect 43385 37780 43478 37846
tri 43385 37764 43401 37780 ne
rect 43401 37764 43478 37780
rect 43218 37665 43366 37747
rect 43106 37632 43183 37648
tri 43183 37632 43199 37648 sw
rect 43106 37566 43199 37632
rect 43106 37464 43199 37530
rect 43106 37448 43183 37464
tri 43183 37448 43199 37464 nw
rect 43235 37431 43349 37665
tri 43385 37632 43401 37648 se
rect 43401 37632 43478 37648
rect 43385 37566 43478 37632
rect 43385 37464 43478 37530
tri 43385 37448 43401 37464 ne
rect 43401 37448 43478 37464
rect 43218 37349 43366 37431
rect 43106 37316 43183 37332
tri 43183 37316 43199 37332 sw
rect 43106 37250 43199 37316
rect 43235 37191 43349 37349
tri 43385 37316 43401 37332 se
rect 43401 37316 43478 37332
rect 43385 37250 43478 37316
rect 43106 37115 43478 37191
rect 43106 36990 43199 37056
rect 43106 36974 43183 36990
tri 43183 36974 43199 36990 nw
rect 43235 36957 43349 37115
rect 43385 36990 43478 37056
tri 43385 36974 43401 36990 ne
rect 43401 36974 43478 36990
rect 43218 36875 43366 36957
rect 43106 36842 43183 36858
tri 43183 36842 43199 36858 sw
rect 43106 36776 43199 36842
rect 43106 36674 43199 36740
rect 43106 36658 43183 36674
tri 43183 36658 43199 36674 nw
rect 43235 36641 43349 36875
tri 43385 36842 43401 36858 se
rect 43401 36842 43478 36858
rect 43385 36776 43478 36842
rect 43385 36674 43478 36740
tri 43385 36658 43401 36674 ne
rect 43401 36658 43478 36674
rect 43218 36559 43366 36641
rect 43106 36526 43183 36542
tri 43183 36526 43199 36542 sw
rect 43106 36460 43199 36526
rect 43235 36401 43349 36559
tri 43385 36526 43401 36542 se
rect 43401 36526 43478 36542
rect 43385 36460 43478 36526
rect 43106 36325 43478 36401
rect 43106 36200 43199 36266
rect 43106 36184 43183 36200
tri 43183 36184 43199 36200 nw
rect 43235 36167 43349 36325
rect 43385 36200 43478 36266
tri 43385 36184 43401 36200 ne
rect 43401 36184 43478 36200
rect 43218 36085 43366 36167
rect 43106 36052 43183 36068
tri 43183 36052 43199 36068 sw
rect 43106 35986 43199 36052
rect 43106 35884 43199 35950
rect 43106 35868 43183 35884
tri 43183 35868 43199 35884 nw
rect 43235 35851 43349 36085
tri 43385 36052 43401 36068 se
rect 43401 36052 43478 36068
rect 43385 35986 43478 36052
rect 43385 35884 43478 35950
tri 43385 35868 43401 35884 ne
rect 43401 35868 43478 35884
rect 43218 35769 43366 35851
rect 43106 35736 43183 35752
tri 43183 35736 43199 35752 sw
rect 43106 35670 43199 35736
rect 43235 35611 43349 35769
tri 43385 35736 43401 35752 se
rect 43401 35736 43478 35752
rect 43385 35670 43478 35736
rect 43106 35535 43478 35611
rect 43106 35410 43199 35476
rect 43106 35394 43183 35410
tri 43183 35394 43199 35410 nw
rect 43235 35377 43349 35535
rect 43385 35410 43478 35476
tri 43385 35394 43401 35410 ne
rect 43401 35394 43478 35410
rect 43218 35295 43366 35377
rect 43106 35262 43183 35278
tri 43183 35262 43199 35278 sw
rect 43106 35196 43199 35262
rect 43106 35094 43199 35160
rect 43106 35078 43183 35094
tri 43183 35078 43199 35094 nw
rect 43235 35061 43349 35295
tri 43385 35262 43401 35278 se
rect 43401 35262 43478 35278
rect 43385 35196 43478 35262
rect 43385 35094 43478 35160
tri 43385 35078 43401 35094 ne
rect 43401 35078 43478 35094
rect 43218 34979 43366 35061
rect 43106 34946 43183 34962
tri 43183 34946 43199 34962 sw
rect 43106 34880 43199 34946
rect 43235 34821 43349 34979
tri 43385 34946 43401 34962 se
rect 43401 34946 43478 34962
rect 43385 34880 43478 34946
rect 43106 34745 43478 34821
rect 43106 34620 43199 34686
rect 43106 34604 43183 34620
tri 43183 34604 43199 34620 nw
rect 43235 34587 43349 34745
rect 43385 34620 43478 34686
tri 43385 34604 43401 34620 ne
rect 43401 34604 43478 34620
rect 43218 34505 43366 34587
rect 43106 34472 43183 34488
tri 43183 34472 43199 34488 sw
rect 43106 34406 43199 34472
rect 43106 34304 43199 34370
rect 43106 34288 43183 34304
tri 43183 34288 43199 34304 nw
rect 43235 34271 43349 34505
tri 43385 34472 43401 34488 se
rect 43401 34472 43478 34488
rect 43385 34406 43478 34472
rect 43385 34304 43478 34370
tri 43385 34288 43401 34304 ne
rect 43401 34288 43478 34304
rect 43218 34189 43366 34271
rect 43106 34156 43183 34172
tri 43183 34156 43199 34172 sw
rect 43106 34090 43199 34156
rect 43235 34031 43349 34189
tri 43385 34156 43401 34172 se
rect 43401 34156 43478 34172
rect 43385 34090 43478 34156
rect 43106 33955 43478 34031
rect 43106 33830 43199 33896
rect 43106 33814 43183 33830
tri 43183 33814 43199 33830 nw
rect 43235 33797 43349 33955
rect 43385 33830 43478 33896
tri 43385 33814 43401 33830 ne
rect 43401 33814 43478 33830
rect 43218 33715 43366 33797
rect 43106 33682 43183 33698
tri 43183 33682 43199 33698 sw
rect 43106 33616 43199 33682
rect 43106 33514 43199 33580
rect 43106 33498 43183 33514
tri 43183 33498 43199 33514 nw
rect 43235 33481 43349 33715
tri 43385 33682 43401 33698 se
rect 43401 33682 43478 33698
rect 43385 33616 43478 33682
rect 43385 33514 43478 33580
tri 43385 33498 43401 33514 ne
rect 43401 33498 43478 33514
rect 43218 33399 43366 33481
rect 43106 33366 43183 33382
tri 43183 33366 43199 33382 sw
rect 43106 33300 43199 33366
rect 43235 33241 43349 33399
tri 43385 33366 43401 33382 se
rect 43401 33366 43478 33382
rect 43385 33300 43478 33366
rect 43106 33165 43478 33241
rect 43106 33040 43199 33106
rect 43106 33024 43183 33040
tri 43183 33024 43199 33040 nw
rect 43235 33007 43349 33165
rect 43385 33040 43478 33106
tri 43385 33024 43401 33040 ne
rect 43401 33024 43478 33040
rect 43218 32925 43366 33007
rect 43106 32892 43183 32908
tri 43183 32892 43199 32908 sw
rect 43106 32826 43199 32892
rect 43106 32724 43199 32790
rect 43106 32708 43183 32724
tri 43183 32708 43199 32724 nw
rect 43235 32691 43349 32925
tri 43385 32892 43401 32908 se
rect 43401 32892 43478 32908
rect 43385 32826 43478 32892
rect 43385 32724 43478 32790
tri 43385 32708 43401 32724 ne
rect 43401 32708 43478 32724
rect 43218 32609 43366 32691
rect 43106 32576 43183 32592
tri 43183 32576 43199 32592 sw
rect 43106 32510 43199 32576
rect 43235 32451 43349 32609
tri 43385 32576 43401 32592 se
rect 43401 32576 43478 32592
rect 43385 32510 43478 32576
rect 43106 32375 43478 32451
rect 43106 32250 43199 32316
rect 43106 32234 43183 32250
tri 43183 32234 43199 32250 nw
rect 43235 32217 43349 32375
rect 43385 32250 43478 32316
tri 43385 32234 43401 32250 ne
rect 43401 32234 43478 32250
rect 43218 32135 43366 32217
rect 43106 32102 43183 32118
tri 43183 32102 43199 32118 sw
rect 43106 32036 43199 32102
rect 43106 31934 43199 32000
rect 43106 31918 43183 31934
tri 43183 31918 43199 31934 nw
rect 43235 31901 43349 32135
tri 43385 32102 43401 32118 se
rect 43401 32102 43478 32118
rect 43385 32036 43478 32102
rect 43385 31934 43478 32000
tri 43385 31918 43401 31934 ne
rect 43401 31918 43478 31934
rect 43218 31819 43366 31901
rect 43106 31786 43183 31802
tri 43183 31786 43199 31802 sw
rect 43106 31720 43199 31786
rect 43235 31661 43349 31819
tri 43385 31786 43401 31802 se
rect 43401 31786 43478 31802
rect 43385 31720 43478 31786
rect 43106 31585 43478 31661
rect 43106 31460 43199 31526
rect 43106 31444 43183 31460
tri 43183 31444 43199 31460 nw
rect 43235 31427 43349 31585
rect 43385 31460 43478 31526
tri 43385 31444 43401 31460 ne
rect 43401 31444 43478 31460
rect 43218 31345 43366 31427
rect 43106 31312 43183 31328
tri 43183 31312 43199 31328 sw
rect 43106 31246 43199 31312
rect 43106 31144 43199 31210
rect 43106 31128 43183 31144
tri 43183 31128 43199 31144 nw
rect 43235 31111 43349 31345
tri 43385 31312 43401 31328 se
rect 43401 31312 43478 31328
rect 43385 31246 43478 31312
rect 43385 31144 43478 31210
tri 43385 31128 43401 31144 ne
rect 43401 31128 43478 31144
rect 43218 31029 43366 31111
rect 43106 30996 43183 31012
tri 43183 30996 43199 31012 sw
rect 43106 30930 43199 30996
rect 43235 30871 43349 31029
tri 43385 30996 43401 31012 se
rect 43401 30996 43478 31012
rect 43385 30930 43478 30996
rect 43106 30795 43478 30871
rect 43106 30670 43199 30736
rect 43106 30654 43183 30670
tri 43183 30654 43199 30670 nw
rect 43235 30637 43349 30795
rect 43385 30670 43478 30736
tri 43385 30654 43401 30670 ne
rect 43401 30654 43478 30670
rect 43218 30555 43366 30637
rect 43106 30522 43183 30538
tri 43183 30522 43199 30538 sw
rect 43106 30456 43199 30522
rect 43106 30354 43199 30420
rect 43106 30338 43183 30354
tri 43183 30338 43199 30354 nw
rect 43235 30321 43349 30555
tri 43385 30522 43401 30538 se
rect 43401 30522 43478 30538
rect 43385 30456 43478 30522
rect 43385 30354 43478 30420
tri 43385 30338 43401 30354 ne
rect 43401 30338 43478 30354
rect 43218 30239 43366 30321
rect 43106 30206 43183 30222
tri 43183 30206 43199 30222 sw
rect 43106 30140 43199 30206
rect 43235 30081 43349 30239
tri 43385 30206 43401 30222 se
rect 43401 30206 43478 30222
rect 43385 30140 43478 30206
rect 43106 30005 43478 30081
rect 43106 29880 43199 29946
rect 43106 29864 43183 29880
tri 43183 29864 43199 29880 nw
rect 43235 29847 43349 30005
rect 43385 29880 43478 29946
tri 43385 29864 43401 29880 ne
rect 43401 29864 43478 29880
rect 43218 29765 43366 29847
rect 43106 29732 43183 29748
tri 43183 29732 43199 29748 sw
rect 43106 29666 43199 29732
rect 43106 29564 43199 29630
rect 43106 29548 43183 29564
tri 43183 29548 43199 29564 nw
rect 43235 29531 43349 29765
tri 43385 29732 43401 29748 se
rect 43401 29732 43478 29748
rect 43385 29666 43478 29732
rect 43385 29564 43478 29630
tri 43385 29548 43401 29564 ne
rect 43401 29548 43478 29564
rect 43218 29449 43366 29531
rect 43106 29416 43183 29432
tri 43183 29416 43199 29432 sw
rect 43106 29350 43199 29416
rect 43235 29291 43349 29449
tri 43385 29416 43401 29432 se
rect 43401 29416 43478 29432
rect 43385 29350 43478 29416
rect 43106 29215 43478 29291
rect 43106 29090 43199 29156
rect 43106 29074 43183 29090
tri 43183 29074 43199 29090 nw
rect 43235 29057 43349 29215
rect 43385 29090 43478 29156
tri 43385 29074 43401 29090 ne
rect 43401 29074 43478 29090
rect 43218 28975 43366 29057
rect 43106 28942 43183 28958
tri 43183 28942 43199 28958 sw
rect 43106 28876 43199 28942
rect 43235 28833 43349 28975
tri 43385 28942 43401 28958 se
rect 43401 28942 43478 28958
rect 43385 28876 43478 28942
rect 43514 28463 43550 80603
rect 43586 28463 43622 80603
rect 43658 80445 43694 80603
rect 43650 80303 43702 80445
rect 43658 28763 43694 80303
rect 43650 28621 43702 28763
rect 43658 28463 43694 28621
rect 43730 28463 43766 80603
rect 43802 28463 43838 80603
rect 43874 28833 43958 80233
rect 43994 28463 44030 80603
rect 44066 28463 44102 80603
rect 44138 80445 44174 80603
rect 44130 80303 44182 80445
rect 44138 28763 44174 80303
rect 44130 28621 44182 28763
rect 44138 28463 44174 28621
rect 44210 28463 44246 80603
rect 44282 28463 44318 80603
rect 44354 80124 44447 80190
rect 44354 80108 44431 80124
tri 44431 80108 44447 80124 nw
rect 44483 80091 44597 80233
rect 44633 80124 44726 80190
tri 44633 80108 44649 80124 ne
rect 44649 80108 44726 80124
rect 44466 80009 44614 80091
rect 44354 79976 44431 79992
tri 44431 79976 44447 79992 sw
rect 44354 79910 44447 79976
rect 44483 79851 44597 80009
tri 44633 79976 44649 79992 se
rect 44649 79976 44726 79992
rect 44633 79910 44726 79976
rect 44354 79775 44726 79851
rect 44354 79650 44447 79716
rect 44354 79634 44431 79650
tri 44431 79634 44447 79650 nw
rect 44483 79617 44597 79775
rect 44633 79650 44726 79716
tri 44633 79634 44649 79650 ne
rect 44649 79634 44726 79650
rect 44466 79535 44614 79617
rect 44354 79502 44431 79518
tri 44431 79502 44447 79518 sw
rect 44354 79436 44447 79502
rect 44354 79334 44447 79400
rect 44354 79318 44431 79334
tri 44431 79318 44447 79334 nw
rect 44483 79301 44597 79535
tri 44633 79502 44649 79518 se
rect 44649 79502 44726 79518
rect 44633 79436 44726 79502
rect 44633 79334 44726 79400
tri 44633 79318 44649 79334 ne
rect 44649 79318 44726 79334
rect 44466 79219 44614 79301
rect 44354 79186 44431 79202
tri 44431 79186 44447 79202 sw
rect 44354 79120 44447 79186
rect 44483 79061 44597 79219
tri 44633 79186 44649 79202 se
rect 44649 79186 44726 79202
rect 44633 79120 44726 79186
rect 44354 78985 44726 79061
rect 44354 78860 44447 78926
rect 44354 78844 44431 78860
tri 44431 78844 44447 78860 nw
rect 44483 78827 44597 78985
rect 44633 78860 44726 78926
tri 44633 78844 44649 78860 ne
rect 44649 78844 44726 78860
rect 44466 78745 44614 78827
rect 44354 78712 44431 78728
tri 44431 78712 44447 78728 sw
rect 44354 78646 44447 78712
rect 44354 78544 44447 78610
rect 44354 78528 44431 78544
tri 44431 78528 44447 78544 nw
rect 44483 78511 44597 78745
tri 44633 78712 44649 78728 se
rect 44649 78712 44726 78728
rect 44633 78646 44726 78712
rect 44633 78544 44726 78610
tri 44633 78528 44649 78544 ne
rect 44649 78528 44726 78544
rect 44466 78429 44614 78511
rect 44354 78396 44431 78412
tri 44431 78396 44447 78412 sw
rect 44354 78330 44447 78396
rect 44483 78271 44597 78429
tri 44633 78396 44649 78412 se
rect 44649 78396 44726 78412
rect 44633 78330 44726 78396
rect 44354 78195 44726 78271
rect 44354 78070 44447 78136
rect 44354 78054 44431 78070
tri 44431 78054 44447 78070 nw
rect 44483 78037 44597 78195
rect 44633 78070 44726 78136
tri 44633 78054 44649 78070 ne
rect 44649 78054 44726 78070
rect 44466 77955 44614 78037
rect 44354 77922 44431 77938
tri 44431 77922 44447 77938 sw
rect 44354 77856 44447 77922
rect 44354 77754 44447 77820
rect 44354 77738 44431 77754
tri 44431 77738 44447 77754 nw
rect 44483 77721 44597 77955
tri 44633 77922 44649 77938 se
rect 44649 77922 44726 77938
rect 44633 77856 44726 77922
rect 44633 77754 44726 77820
tri 44633 77738 44649 77754 ne
rect 44649 77738 44726 77754
rect 44466 77639 44614 77721
rect 44354 77606 44431 77622
tri 44431 77606 44447 77622 sw
rect 44354 77540 44447 77606
rect 44483 77481 44597 77639
tri 44633 77606 44649 77622 se
rect 44649 77606 44726 77622
rect 44633 77540 44726 77606
rect 44354 77405 44726 77481
rect 44354 77280 44447 77346
rect 44354 77264 44431 77280
tri 44431 77264 44447 77280 nw
rect 44483 77247 44597 77405
rect 44633 77280 44726 77346
tri 44633 77264 44649 77280 ne
rect 44649 77264 44726 77280
rect 44466 77165 44614 77247
rect 44354 77132 44431 77148
tri 44431 77132 44447 77148 sw
rect 44354 77066 44447 77132
rect 44354 76964 44447 77030
rect 44354 76948 44431 76964
tri 44431 76948 44447 76964 nw
rect 44483 76931 44597 77165
tri 44633 77132 44649 77148 se
rect 44649 77132 44726 77148
rect 44633 77066 44726 77132
rect 44633 76964 44726 77030
tri 44633 76948 44649 76964 ne
rect 44649 76948 44726 76964
rect 44466 76849 44614 76931
rect 44354 76816 44431 76832
tri 44431 76816 44447 76832 sw
rect 44354 76750 44447 76816
rect 44483 76691 44597 76849
tri 44633 76816 44649 76832 se
rect 44649 76816 44726 76832
rect 44633 76750 44726 76816
rect 44354 76615 44726 76691
rect 44354 76490 44447 76556
rect 44354 76474 44431 76490
tri 44431 76474 44447 76490 nw
rect 44483 76457 44597 76615
rect 44633 76490 44726 76556
tri 44633 76474 44649 76490 ne
rect 44649 76474 44726 76490
rect 44466 76375 44614 76457
rect 44354 76342 44431 76358
tri 44431 76342 44447 76358 sw
rect 44354 76276 44447 76342
rect 44354 76174 44447 76240
rect 44354 76158 44431 76174
tri 44431 76158 44447 76174 nw
rect 44483 76141 44597 76375
tri 44633 76342 44649 76358 se
rect 44649 76342 44726 76358
rect 44633 76276 44726 76342
rect 44633 76174 44726 76240
tri 44633 76158 44649 76174 ne
rect 44649 76158 44726 76174
rect 44466 76059 44614 76141
rect 44354 76026 44431 76042
tri 44431 76026 44447 76042 sw
rect 44354 75960 44447 76026
rect 44483 75901 44597 76059
tri 44633 76026 44649 76042 se
rect 44649 76026 44726 76042
rect 44633 75960 44726 76026
rect 44354 75825 44726 75901
rect 44354 75700 44447 75766
rect 44354 75684 44431 75700
tri 44431 75684 44447 75700 nw
rect 44483 75667 44597 75825
rect 44633 75700 44726 75766
tri 44633 75684 44649 75700 ne
rect 44649 75684 44726 75700
rect 44466 75585 44614 75667
rect 44354 75552 44431 75568
tri 44431 75552 44447 75568 sw
rect 44354 75486 44447 75552
rect 44354 75384 44447 75450
rect 44354 75368 44431 75384
tri 44431 75368 44447 75384 nw
rect 44483 75351 44597 75585
tri 44633 75552 44649 75568 se
rect 44649 75552 44726 75568
rect 44633 75486 44726 75552
rect 44633 75384 44726 75450
tri 44633 75368 44649 75384 ne
rect 44649 75368 44726 75384
rect 44466 75269 44614 75351
rect 44354 75236 44431 75252
tri 44431 75236 44447 75252 sw
rect 44354 75170 44447 75236
rect 44483 75111 44597 75269
tri 44633 75236 44649 75252 se
rect 44649 75236 44726 75252
rect 44633 75170 44726 75236
rect 44354 75035 44726 75111
rect 44354 74910 44447 74976
rect 44354 74894 44431 74910
tri 44431 74894 44447 74910 nw
rect 44483 74877 44597 75035
rect 44633 74910 44726 74976
tri 44633 74894 44649 74910 ne
rect 44649 74894 44726 74910
rect 44466 74795 44614 74877
rect 44354 74762 44431 74778
tri 44431 74762 44447 74778 sw
rect 44354 74696 44447 74762
rect 44354 74594 44447 74660
rect 44354 74578 44431 74594
tri 44431 74578 44447 74594 nw
rect 44483 74561 44597 74795
tri 44633 74762 44649 74778 se
rect 44649 74762 44726 74778
rect 44633 74696 44726 74762
rect 44633 74594 44726 74660
tri 44633 74578 44649 74594 ne
rect 44649 74578 44726 74594
rect 44466 74479 44614 74561
rect 44354 74446 44431 74462
tri 44431 74446 44447 74462 sw
rect 44354 74380 44447 74446
rect 44483 74321 44597 74479
tri 44633 74446 44649 74462 se
rect 44649 74446 44726 74462
rect 44633 74380 44726 74446
rect 44354 74245 44726 74321
rect 44354 74120 44447 74186
rect 44354 74104 44431 74120
tri 44431 74104 44447 74120 nw
rect 44483 74087 44597 74245
rect 44633 74120 44726 74186
tri 44633 74104 44649 74120 ne
rect 44649 74104 44726 74120
rect 44466 74005 44614 74087
rect 44354 73972 44431 73988
tri 44431 73972 44447 73988 sw
rect 44354 73906 44447 73972
rect 44354 73804 44447 73870
rect 44354 73788 44431 73804
tri 44431 73788 44447 73804 nw
rect 44483 73771 44597 74005
tri 44633 73972 44649 73988 se
rect 44649 73972 44726 73988
rect 44633 73906 44726 73972
rect 44633 73804 44726 73870
tri 44633 73788 44649 73804 ne
rect 44649 73788 44726 73804
rect 44466 73689 44614 73771
rect 44354 73656 44431 73672
tri 44431 73656 44447 73672 sw
rect 44354 73590 44447 73656
rect 44483 73531 44597 73689
tri 44633 73656 44649 73672 se
rect 44649 73656 44726 73672
rect 44633 73590 44726 73656
rect 44354 73455 44726 73531
rect 44354 73330 44447 73396
rect 44354 73314 44431 73330
tri 44431 73314 44447 73330 nw
rect 44483 73297 44597 73455
rect 44633 73330 44726 73396
tri 44633 73314 44649 73330 ne
rect 44649 73314 44726 73330
rect 44466 73215 44614 73297
rect 44354 73182 44431 73198
tri 44431 73182 44447 73198 sw
rect 44354 73116 44447 73182
rect 44354 73014 44447 73080
rect 44354 72998 44431 73014
tri 44431 72998 44447 73014 nw
rect 44483 72981 44597 73215
tri 44633 73182 44649 73198 se
rect 44649 73182 44726 73198
rect 44633 73116 44726 73182
rect 44633 73014 44726 73080
tri 44633 72998 44649 73014 ne
rect 44649 72998 44726 73014
rect 44466 72899 44614 72981
rect 44354 72866 44431 72882
tri 44431 72866 44447 72882 sw
rect 44354 72800 44447 72866
rect 44483 72741 44597 72899
tri 44633 72866 44649 72882 se
rect 44649 72866 44726 72882
rect 44633 72800 44726 72866
rect 44354 72665 44726 72741
rect 44354 72540 44447 72606
rect 44354 72524 44431 72540
tri 44431 72524 44447 72540 nw
rect 44483 72507 44597 72665
rect 44633 72540 44726 72606
tri 44633 72524 44649 72540 ne
rect 44649 72524 44726 72540
rect 44466 72425 44614 72507
rect 44354 72392 44431 72408
tri 44431 72392 44447 72408 sw
rect 44354 72326 44447 72392
rect 44354 72224 44447 72290
rect 44354 72208 44431 72224
tri 44431 72208 44447 72224 nw
rect 44483 72191 44597 72425
tri 44633 72392 44649 72408 se
rect 44649 72392 44726 72408
rect 44633 72326 44726 72392
rect 44633 72224 44726 72290
tri 44633 72208 44649 72224 ne
rect 44649 72208 44726 72224
rect 44466 72109 44614 72191
rect 44354 72076 44431 72092
tri 44431 72076 44447 72092 sw
rect 44354 72010 44447 72076
rect 44483 71951 44597 72109
tri 44633 72076 44649 72092 se
rect 44649 72076 44726 72092
rect 44633 72010 44726 72076
rect 44354 71875 44726 71951
rect 44354 71750 44447 71816
rect 44354 71734 44431 71750
tri 44431 71734 44447 71750 nw
rect 44483 71717 44597 71875
rect 44633 71750 44726 71816
tri 44633 71734 44649 71750 ne
rect 44649 71734 44726 71750
rect 44466 71635 44614 71717
rect 44354 71602 44431 71618
tri 44431 71602 44447 71618 sw
rect 44354 71536 44447 71602
rect 44354 71434 44447 71500
rect 44354 71418 44431 71434
tri 44431 71418 44447 71434 nw
rect 44483 71401 44597 71635
tri 44633 71602 44649 71618 se
rect 44649 71602 44726 71618
rect 44633 71536 44726 71602
rect 44633 71434 44726 71500
tri 44633 71418 44649 71434 ne
rect 44649 71418 44726 71434
rect 44466 71319 44614 71401
rect 44354 71286 44431 71302
tri 44431 71286 44447 71302 sw
rect 44354 71220 44447 71286
rect 44483 71161 44597 71319
tri 44633 71286 44649 71302 se
rect 44649 71286 44726 71302
rect 44633 71220 44726 71286
rect 44354 71085 44726 71161
rect 44354 70960 44447 71026
rect 44354 70944 44431 70960
tri 44431 70944 44447 70960 nw
rect 44483 70927 44597 71085
rect 44633 70960 44726 71026
tri 44633 70944 44649 70960 ne
rect 44649 70944 44726 70960
rect 44466 70845 44614 70927
rect 44354 70812 44431 70828
tri 44431 70812 44447 70828 sw
rect 44354 70746 44447 70812
rect 44354 70644 44447 70710
rect 44354 70628 44431 70644
tri 44431 70628 44447 70644 nw
rect 44483 70611 44597 70845
tri 44633 70812 44649 70828 se
rect 44649 70812 44726 70828
rect 44633 70746 44726 70812
rect 44633 70644 44726 70710
tri 44633 70628 44649 70644 ne
rect 44649 70628 44726 70644
rect 44466 70529 44614 70611
rect 44354 70496 44431 70512
tri 44431 70496 44447 70512 sw
rect 44354 70430 44447 70496
rect 44483 70371 44597 70529
tri 44633 70496 44649 70512 se
rect 44649 70496 44726 70512
rect 44633 70430 44726 70496
rect 44354 70295 44726 70371
rect 44354 70170 44447 70236
rect 44354 70154 44431 70170
tri 44431 70154 44447 70170 nw
rect 44483 70137 44597 70295
rect 44633 70170 44726 70236
tri 44633 70154 44649 70170 ne
rect 44649 70154 44726 70170
rect 44466 70055 44614 70137
rect 44354 70022 44431 70038
tri 44431 70022 44447 70038 sw
rect 44354 69956 44447 70022
rect 44354 69854 44447 69920
rect 44354 69838 44431 69854
tri 44431 69838 44447 69854 nw
rect 44483 69821 44597 70055
tri 44633 70022 44649 70038 se
rect 44649 70022 44726 70038
rect 44633 69956 44726 70022
rect 44633 69854 44726 69920
tri 44633 69838 44649 69854 ne
rect 44649 69838 44726 69854
rect 44466 69739 44614 69821
rect 44354 69706 44431 69722
tri 44431 69706 44447 69722 sw
rect 44354 69640 44447 69706
rect 44483 69581 44597 69739
tri 44633 69706 44649 69722 se
rect 44649 69706 44726 69722
rect 44633 69640 44726 69706
rect 44354 69505 44726 69581
rect 44354 69380 44447 69446
rect 44354 69364 44431 69380
tri 44431 69364 44447 69380 nw
rect 44483 69347 44597 69505
rect 44633 69380 44726 69446
tri 44633 69364 44649 69380 ne
rect 44649 69364 44726 69380
rect 44466 69265 44614 69347
rect 44354 69232 44431 69248
tri 44431 69232 44447 69248 sw
rect 44354 69166 44447 69232
rect 44354 69064 44447 69130
rect 44354 69048 44431 69064
tri 44431 69048 44447 69064 nw
rect 44483 69031 44597 69265
tri 44633 69232 44649 69248 se
rect 44649 69232 44726 69248
rect 44633 69166 44726 69232
rect 44633 69064 44726 69130
tri 44633 69048 44649 69064 ne
rect 44649 69048 44726 69064
rect 44466 68949 44614 69031
rect 44354 68916 44431 68932
tri 44431 68916 44447 68932 sw
rect 44354 68850 44447 68916
rect 44483 68791 44597 68949
tri 44633 68916 44649 68932 se
rect 44649 68916 44726 68932
rect 44633 68850 44726 68916
rect 44354 68715 44726 68791
rect 44354 68590 44447 68656
rect 44354 68574 44431 68590
tri 44431 68574 44447 68590 nw
rect 44483 68557 44597 68715
rect 44633 68590 44726 68656
tri 44633 68574 44649 68590 ne
rect 44649 68574 44726 68590
rect 44466 68475 44614 68557
rect 44354 68442 44431 68458
tri 44431 68442 44447 68458 sw
rect 44354 68376 44447 68442
rect 44354 68274 44447 68340
rect 44354 68258 44431 68274
tri 44431 68258 44447 68274 nw
rect 44483 68241 44597 68475
tri 44633 68442 44649 68458 se
rect 44649 68442 44726 68458
rect 44633 68376 44726 68442
rect 44633 68274 44726 68340
tri 44633 68258 44649 68274 ne
rect 44649 68258 44726 68274
rect 44466 68159 44614 68241
rect 44354 68126 44431 68142
tri 44431 68126 44447 68142 sw
rect 44354 68060 44447 68126
rect 44483 68001 44597 68159
tri 44633 68126 44649 68142 se
rect 44649 68126 44726 68142
rect 44633 68060 44726 68126
rect 44354 67925 44726 68001
rect 44354 67800 44447 67866
rect 44354 67784 44431 67800
tri 44431 67784 44447 67800 nw
rect 44483 67767 44597 67925
rect 44633 67800 44726 67866
tri 44633 67784 44649 67800 ne
rect 44649 67784 44726 67800
rect 44466 67685 44614 67767
rect 44354 67652 44431 67668
tri 44431 67652 44447 67668 sw
rect 44354 67586 44447 67652
rect 44354 67484 44447 67550
rect 44354 67468 44431 67484
tri 44431 67468 44447 67484 nw
rect 44483 67451 44597 67685
tri 44633 67652 44649 67668 se
rect 44649 67652 44726 67668
rect 44633 67586 44726 67652
rect 44633 67484 44726 67550
tri 44633 67468 44649 67484 ne
rect 44649 67468 44726 67484
rect 44466 67369 44614 67451
rect 44354 67336 44431 67352
tri 44431 67336 44447 67352 sw
rect 44354 67270 44447 67336
rect 44483 67211 44597 67369
tri 44633 67336 44649 67352 se
rect 44649 67336 44726 67352
rect 44633 67270 44726 67336
rect 44354 67135 44726 67211
rect 44354 67010 44447 67076
rect 44354 66994 44431 67010
tri 44431 66994 44447 67010 nw
rect 44483 66977 44597 67135
rect 44633 67010 44726 67076
tri 44633 66994 44649 67010 ne
rect 44649 66994 44726 67010
rect 44466 66895 44614 66977
rect 44354 66862 44431 66878
tri 44431 66862 44447 66878 sw
rect 44354 66796 44447 66862
rect 44354 66694 44447 66760
rect 44354 66678 44431 66694
tri 44431 66678 44447 66694 nw
rect 44483 66661 44597 66895
tri 44633 66862 44649 66878 se
rect 44649 66862 44726 66878
rect 44633 66796 44726 66862
rect 44633 66694 44726 66760
tri 44633 66678 44649 66694 ne
rect 44649 66678 44726 66694
rect 44466 66579 44614 66661
rect 44354 66546 44431 66562
tri 44431 66546 44447 66562 sw
rect 44354 66480 44447 66546
rect 44483 66421 44597 66579
tri 44633 66546 44649 66562 se
rect 44649 66546 44726 66562
rect 44633 66480 44726 66546
rect 44354 66345 44726 66421
rect 44354 66220 44447 66286
rect 44354 66204 44431 66220
tri 44431 66204 44447 66220 nw
rect 44483 66187 44597 66345
rect 44633 66220 44726 66286
tri 44633 66204 44649 66220 ne
rect 44649 66204 44726 66220
rect 44466 66105 44614 66187
rect 44354 66072 44431 66088
tri 44431 66072 44447 66088 sw
rect 44354 66006 44447 66072
rect 44354 65904 44447 65970
rect 44354 65888 44431 65904
tri 44431 65888 44447 65904 nw
rect 44483 65871 44597 66105
tri 44633 66072 44649 66088 se
rect 44649 66072 44726 66088
rect 44633 66006 44726 66072
rect 44633 65904 44726 65970
tri 44633 65888 44649 65904 ne
rect 44649 65888 44726 65904
rect 44466 65789 44614 65871
rect 44354 65756 44431 65772
tri 44431 65756 44447 65772 sw
rect 44354 65690 44447 65756
rect 44483 65631 44597 65789
tri 44633 65756 44649 65772 se
rect 44649 65756 44726 65772
rect 44633 65690 44726 65756
rect 44354 65555 44726 65631
rect 44354 65430 44447 65496
rect 44354 65414 44431 65430
tri 44431 65414 44447 65430 nw
rect 44483 65397 44597 65555
rect 44633 65430 44726 65496
tri 44633 65414 44649 65430 ne
rect 44649 65414 44726 65430
rect 44466 65315 44614 65397
rect 44354 65282 44431 65298
tri 44431 65282 44447 65298 sw
rect 44354 65216 44447 65282
rect 44354 65114 44447 65180
rect 44354 65098 44431 65114
tri 44431 65098 44447 65114 nw
rect 44483 65081 44597 65315
tri 44633 65282 44649 65298 se
rect 44649 65282 44726 65298
rect 44633 65216 44726 65282
rect 44633 65114 44726 65180
tri 44633 65098 44649 65114 ne
rect 44649 65098 44726 65114
rect 44466 64999 44614 65081
rect 44354 64966 44431 64982
tri 44431 64966 44447 64982 sw
rect 44354 64900 44447 64966
rect 44483 64841 44597 64999
tri 44633 64966 44649 64982 se
rect 44649 64966 44726 64982
rect 44633 64900 44726 64966
rect 44354 64765 44726 64841
rect 44354 64640 44447 64706
rect 44354 64624 44431 64640
tri 44431 64624 44447 64640 nw
rect 44483 64607 44597 64765
rect 44633 64640 44726 64706
tri 44633 64624 44649 64640 ne
rect 44649 64624 44726 64640
rect 44466 64525 44614 64607
rect 44354 64492 44431 64508
tri 44431 64492 44447 64508 sw
rect 44354 64426 44447 64492
rect 44354 64324 44447 64390
rect 44354 64308 44431 64324
tri 44431 64308 44447 64324 nw
rect 44483 64291 44597 64525
tri 44633 64492 44649 64508 se
rect 44649 64492 44726 64508
rect 44633 64426 44726 64492
rect 44633 64324 44726 64390
tri 44633 64308 44649 64324 ne
rect 44649 64308 44726 64324
rect 44466 64209 44614 64291
rect 44354 64176 44431 64192
tri 44431 64176 44447 64192 sw
rect 44354 64110 44447 64176
rect 44483 64051 44597 64209
tri 44633 64176 44649 64192 se
rect 44649 64176 44726 64192
rect 44633 64110 44726 64176
rect 44354 63975 44726 64051
rect 44354 63850 44447 63916
rect 44354 63834 44431 63850
tri 44431 63834 44447 63850 nw
rect 44483 63817 44597 63975
rect 44633 63850 44726 63916
tri 44633 63834 44649 63850 ne
rect 44649 63834 44726 63850
rect 44466 63735 44614 63817
rect 44354 63702 44431 63718
tri 44431 63702 44447 63718 sw
rect 44354 63636 44447 63702
rect 44354 63534 44447 63600
rect 44354 63518 44431 63534
tri 44431 63518 44447 63534 nw
rect 44483 63501 44597 63735
tri 44633 63702 44649 63718 se
rect 44649 63702 44726 63718
rect 44633 63636 44726 63702
rect 44633 63534 44726 63600
tri 44633 63518 44649 63534 ne
rect 44649 63518 44726 63534
rect 44466 63419 44614 63501
rect 44354 63386 44431 63402
tri 44431 63386 44447 63402 sw
rect 44354 63320 44447 63386
rect 44483 63261 44597 63419
tri 44633 63386 44649 63402 se
rect 44649 63386 44726 63402
rect 44633 63320 44726 63386
rect 44354 63185 44726 63261
rect 44354 63060 44447 63126
rect 44354 63044 44431 63060
tri 44431 63044 44447 63060 nw
rect 44483 63027 44597 63185
rect 44633 63060 44726 63126
tri 44633 63044 44649 63060 ne
rect 44649 63044 44726 63060
rect 44466 62945 44614 63027
rect 44354 62912 44431 62928
tri 44431 62912 44447 62928 sw
rect 44354 62846 44447 62912
rect 44354 62744 44447 62810
rect 44354 62728 44431 62744
tri 44431 62728 44447 62744 nw
rect 44483 62711 44597 62945
tri 44633 62912 44649 62928 se
rect 44649 62912 44726 62928
rect 44633 62846 44726 62912
rect 44633 62744 44726 62810
tri 44633 62728 44649 62744 ne
rect 44649 62728 44726 62744
rect 44466 62629 44614 62711
rect 44354 62596 44431 62612
tri 44431 62596 44447 62612 sw
rect 44354 62530 44447 62596
rect 44483 62471 44597 62629
tri 44633 62596 44649 62612 se
rect 44649 62596 44726 62612
rect 44633 62530 44726 62596
rect 44354 62395 44726 62471
rect 44354 62270 44447 62336
rect 44354 62254 44431 62270
tri 44431 62254 44447 62270 nw
rect 44483 62237 44597 62395
rect 44633 62270 44726 62336
tri 44633 62254 44649 62270 ne
rect 44649 62254 44726 62270
rect 44466 62155 44614 62237
rect 44354 62122 44431 62138
tri 44431 62122 44447 62138 sw
rect 44354 62056 44447 62122
rect 44354 61954 44447 62020
rect 44354 61938 44431 61954
tri 44431 61938 44447 61954 nw
rect 44483 61921 44597 62155
tri 44633 62122 44649 62138 se
rect 44649 62122 44726 62138
rect 44633 62056 44726 62122
rect 44633 61954 44726 62020
tri 44633 61938 44649 61954 ne
rect 44649 61938 44726 61954
rect 44466 61839 44614 61921
rect 44354 61806 44431 61822
tri 44431 61806 44447 61822 sw
rect 44354 61740 44447 61806
rect 44483 61681 44597 61839
tri 44633 61806 44649 61822 se
rect 44649 61806 44726 61822
rect 44633 61740 44726 61806
rect 44354 61605 44726 61681
rect 44354 61480 44447 61546
rect 44354 61464 44431 61480
tri 44431 61464 44447 61480 nw
rect 44483 61447 44597 61605
rect 44633 61480 44726 61546
tri 44633 61464 44649 61480 ne
rect 44649 61464 44726 61480
rect 44466 61365 44614 61447
rect 44354 61332 44431 61348
tri 44431 61332 44447 61348 sw
rect 44354 61266 44447 61332
rect 44354 61164 44447 61230
rect 44354 61148 44431 61164
tri 44431 61148 44447 61164 nw
rect 44483 61131 44597 61365
tri 44633 61332 44649 61348 se
rect 44649 61332 44726 61348
rect 44633 61266 44726 61332
rect 44633 61164 44726 61230
tri 44633 61148 44649 61164 ne
rect 44649 61148 44726 61164
rect 44466 61049 44614 61131
rect 44354 61016 44431 61032
tri 44431 61016 44447 61032 sw
rect 44354 60950 44447 61016
rect 44483 60891 44597 61049
tri 44633 61016 44649 61032 se
rect 44649 61016 44726 61032
rect 44633 60950 44726 61016
rect 44354 60815 44726 60891
rect 44354 60690 44447 60756
rect 44354 60674 44431 60690
tri 44431 60674 44447 60690 nw
rect 44483 60657 44597 60815
rect 44633 60690 44726 60756
tri 44633 60674 44649 60690 ne
rect 44649 60674 44726 60690
rect 44466 60575 44614 60657
rect 44354 60542 44431 60558
tri 44431 60542 44447 60558 sw
rect 44354 60476 44447 60542
rect 44354 60374 44447 60440
rect 44354 60358 44431 60374
tri 44431 60358 44447 60374 nw
rect 44483 60341 44597 60575
tri 44633 60542 44649 60558 se
rect 44649 60542 44726 60558
rect 44633 60476 44726 60542
rect 44633 60374 44726 60440
tri 44633 60358 44649 60374 ne
rect 44649 60358 44726 60374
rect 44466 60259 44614 60341
rect 44354 60226 44431 60242
tri 44431 60226 44447 60242 sw
rect 44354 60160 44447 60226
rect 44483 60101 44597 60259
tri 44633 60226 44649 60242 se
rect 44649 60226 44726 60242
rect 44633 60160 44726 60226
rect 44354 60025 44726 60101
rect 44354 59900 44447 59966
rect 44354 59884 44431 59900
tri 44431 59884 44447 59900 nw
rect 44483 59867 44597 60025
rect 44633 59900 44726 59966
tri 44633 59884 44649 59900 ne
rect 44649 59884 44726 59900
rect 44466 59785 44614 59867
rect 44354 59752 44431 59768
tri 44431 59752 44447 59768 sw
rect 44354 59686 44447 59752
rect 44354 59584 44447 59650
rect 44354 59568 44431 59584
tri 44431 59568 44447 59584 nw
rect 44483 59551 44597 59785
tri 44633 59752 44649 59768 se
rect 44649 59752 44726 59768
rect 44633 59686 44726 59752
rect 44633 59584 44726 59650
tri 44633 59568 44649 59584 ne
rect 44649 59568 44726 59584
rect 44466 59469 44614 59551
rect 44354 59436 44431 59452
tri 44431 59436 44447 59452 sw
rect 44354 59370 44447 59436
rect 44483 59311 44597 59469
tri 44633 59436 44649 59452 se
rect 44649 59436 44726 59452
rect 44633 59370 44726 59436
rect 44354 59235 44726 59311
rect 44354 59110 44447 59176
rect 44354 59094 44431 59110
tri 44431 59094 44447 59110 nw
rect 44483 59077 44597 59235
rect 44633 59110 44726 59176
tri 44633 59094 44649 59110 ne
rect 44649 59094 44726 59110
rect 44466 58995 44614 59077
rect 44354 58962 44431 58978
tri 44431 58962 44447 58978 sw
rect 44354 58896 44447 58962
rect 44354 58794 44447 58860
rect 44354 58778 44431 58794
tri 44431 58778 44447 58794 nw
rect 44483 58761 44597 58995
tri 44633 58962 44649 58978 se
rect 44649 58962 44726 58978
rect 44633 58896 44726 58962
rect 44633 58794 44726 58860
tri 44633 58778 44649 58794 ne
rect 44649 58778 44726 58794
rect 44466 58679 44614 58761
rect 44354 58646 44431 58662
tri 44431 58646 44447 58662 sw
rect 44354 58580 44447 58646
rect 44483 58521 44597 58679
tri 44633 58646 44649 58662 se
rect 44649 58646 44726 58662
rect 44633 58580 44726 58646
rect 44354 58445 44726 58521
rect 44354 58320 44447 58386
rect 44354 58304 44431 58320
tri 44431 58304 44447 58320 nw
rect 44483 58287 44597 58445
rect 44633 58320 44726 58386
tri 44633 58304 44649 58320 ne
rect 44649 58304 44726 58320
rect 44466 58205 44614 58287
rect 44354 58172 44431 58188
tri 44431 58172 44447 58188 sw
rect 44354 58106 44447 58172
rect 44354 58004 44447 58070
rect 44354 57988 44431 58004
tri 44431 57988 44447 58004 nw
rect 44483 57971 44597 58205
tri 44633 58172 44649 58188 se
rect 44649 58172 44726 58188
rect 44633 58106 44726 58172
rect 44633 58004 44726 58070
tri 44633 57988 44649 58004 ne
rect 44649 57988 44726 58004
rect 44466 57889 44614 57971
rect 44354 57856 44431 57872
tri 44431 57856 44447 57872 sw
rect 44354 57790 44447 57856
rect 44483 57731 44597 57889
tri 44633 57856 44649 57872 se
rect 44649 57856 44726 57872
rect 44633 57790 44726 57856
rect 44354 57655 44726 57731
rect 44354 57530 44447 57596
rect 44354 57514 44431 57530
tri 44431 57514 44447 57530 nw
rect 44483 57497 44597 57655
rect 44633 57530 44726 57596
tri 44633 57514 44649 57530 ne
rect 44649 57514 44726 57530
rect 44466 57415 44614 57497
rect 44354 57382 44431 57398
tri 44431 57382 44447 57398 sw
rect 44354 57316 44447 57382
rect 44354 57214 44447 57280
rect 44354 57198 44431 57214
tri 44431 57198 44447 57214 nw
rect 44483 57181 44597 57415
tri 44633 57382 44649 57398 se
rect 44649 57382 44726 57398
rect 44633 57316 44726 57382
rect 44633 57214 44726 57280
tri 44633 57198 44649 57214 ne
rect 44649 57198 44726 57214
rect 44466 57099 44614 57181
rect 44354 57066 44431 57082
tri 44431 57066 44447 57082 sw
rect 44354 57000 44447 57066
rect 44483 56941 44597 57099
tri 44633 57066 44649 57082 se
rect 44649 57066 44726 57082
rect 44633 57000 44726 57066
rect 44354 56865 44726 56941
rect 44354 56740 44447 56806
rect 44354 56724 44431 56740
tri 44431 56724 44447 56740 nw
rect 44483 56707 44597 56865
rect 44633 56740 44726 56806
tri 44633 56724 44649 56740 ne
rect 44649 56724 44726 56740
rect 44466 56625 44614 56707
rect 44354 56592 44431 56608
tri 44431 56592 44447 56608 sw
rect 44354 56526 44447 56592
rect 44354 56424 44447 56490
rect 44354 56408 44431 56424
tri 44431 56408 44447 56424 nw
rect 44483 56391 44597 56625
tri 44633 56592 44649 56608 se
rect 44649 56592 44726 56608
rect 44633 56526 44726 56592
rect 44633 56424 44726 56490
tri 44633 56408 44649 56424 ne
rect 44649 56408 44726 56424
rect 44466 56309 44614 56391
rect 44354 56276 44431 56292
tri 44431 56276 44447 56292 sw
rect 44354 56210 44447 56276
rect 44483 56151 44597 56309
tri 44633 56276 44649 56292 se
rect 44649 56276 44726 56292
rect 44633 56210 44726 56276
rect 44354 56075 44726 56151
rect 44354 55950 44447 56016
rect 44354 55934 44431 55950
tri 44431 55934 44447 55950 nw
rect 44483 55917 44597 56075
rect 44633 55950 44726 56016
tri 44633 55934 44649 55950 ne
rect 44649 55934 44726 55950
rect 44466 55835 44614 55917
rect 44354 55802 44431 55818
tri 44431 55802 44447 55818 sw
rect 44354 55736 44447 55802
rect 44354 55634 44447 55700
rect 44354 55618 44431 55634
tri 44431 55618 44447 55634 nw
rect 44483 55601 44597 55835
tri 44633 55802 44649 55818 se
rect 44649 55802 44726 55818
rect 44633 55736 44726 55802
rect 44633 55634 44726 55700
tri 44633 55618 44649 55634 ne
rect 44649 55618 44726 55634
rect 44466 55519 44614 55601
rect 44354 55486 44431 55502
tri 44431 55486 44447 55502 sw
rect 44354 55420 44447 55486
rect 44483 55361 44597 55519
tri 44633 55486 44649 55502 se
rect 44649 55486 44726 55502
rect 44633 55420 44726 55486
rect 44354 55285 44726 55361
rect 44354 55160 44447 55226
rect 44354 55144 44431 55160
tri 44431 55144 44447 55160 nw
rect 44483 55127 44597 55285
rect 44633 55160 44726 55226
tri 44633 55144 44649 55160 ne
rect 44649 55144 44726 55160
rect 44466 55045 44614 55127
rect 44354 55012 44431 55028
tri 44431 55012 44447 55028 sw
rect 44354 54946 44447 55012
rect 44354 54844 44447 54910
rect 44354 54828 44431 54844
tri 44431 54828 44447 54844 nw
rect 44483 54811 44597 55045
tri 44633 55012 44649 55028 se
rect 44649 55012 44726 55028
rect 44633 54946 44726 55012
rect 44633 54844 44726 54910
tri 44633 54828 44649 54844 ne
rect 44649 54828 44726 54844
rect 44466 54729 44614 54811
rect 44354 54696 44431 54712
tri 44431 54696 44447 54712 sw
rect 44354 54630 44447 54696
rect 44483 54571 44597 54729
tri 44633 54696 44649 54712 se
rect 44649 54696 44726 54712
rect 44633 54630 44726 54696
rect 44354 54495 44726 54571
rect 44354 54370 44447 54436
rect 44354 54354 44431 54370
tri 44431 54354 44447 54370 nw
rect 44483 54337 44597 54495
rect 44633 54370 44726 54436
tri 44633 54354 44649 54370 ne
rect 44649 54354 44726 54370
rect 44466 54255 44614 54337
rect 44354 54222 44431 54238
tri 44431 54222 44447 54238 sw
rect 44354 54156 44447 54222
rect 44354 54054 44447 54120
rect 44354 54038 44431 54054
tri 44431 54038 44447 54054 nw
rect 44483 54021 44597 54255
tri 44633 54222 44649 54238 se
rect 44649 54222 44726 54238
rect 44633 54156 44726 54222
rect 44633 54054 44726 54120
tri 44633 54038 44649 54054 ne
rect 44649 54038 44726 54054
rect 44466 53939 44614 54021
rect 44354 53906 44431 53922
tri 44431 53906 44447 53922 sw
rect 44354 53840 44447 53906
rect 44483 53781 44597 53939
tri 44633 53906 44649 53922 se
rect 44649 53906 44726 53922
rect 44633 53840 44726 53906
rect 44354 53705 44726 53781
rect 44354 53580 44447 53646
rect 44354 53564 44431 53580
tri 44431 53564 44447 53580 nw
rect 44483 53547 44597 53705
rect 44633 53580 44726 53646
tri 44633 53564 44649 53580 ne
rect 44649 53564 44726 53580
rect 44466 53465 44614 53547
rect 44354 53432 44431 53448
tri 44431 53432 44447 53448 sw
rect 44354 53366 44447 53432
rect 44354 53264 44447 53330
rect 44354 53248 44431 53264
tri 44431 53248 44447 53264 nw
rect 44483 53231 44597 53465
tri 44633 53432 44649 53448 se
rect 44649 53432 44726 53448
rect 44633 53366 44726 53432
rect 44633 53264 44726 53330
tri 44633 53248 44649 53264 ne
rect 44649 53248 44726 53264
rect 44466 53149 44614 53231
rect 44354 53116 44431 53132
tri 44431 53116 44447 53132 sw
rect 44354 53050 44447 53116
rect 44483 52991 44597 53149
tri 44633 53116 44649 53132 se
rect 44649 53116 44726 53132
rect 44633 53050 44726 53116
rect 44354 52915 44726 52991
rect 44354 52790 44447 52856
rect 44354 52774 44431 52790
tri 44431 52774 44447 52790 nw
rect 44483 52757 44597 52915
rect 44633 52790 44726 52856
tri 44633 52774 44649 52790 ne
rect 44649 52774 44726 52790
rect 44466 52675 44614 52757
rect 44354 52642 44431 52658
tri 44431 52642 44447 52658 sw
rect 44354 52576 44447 52642
rect 44354 52474 44447 52540
rect 44354 52458 44431 52474
tri 44431 52458 44447 52474 nw
rect 44483 52441 44597 52675
tri 44633 52642 44649 52658 se
rect 44649 52642 44726 52658
rect 44633 52576 44726 52642
rect 44633 52474 44726 52540
tri 44633 52458 44649 52474 ne
rect 44649 52458 44726 52474
rect 44466 52359 44614 52441
rect 44354 52326 44431 52342
tri 44431 52326 44447 52342 sw
rect 44354 52260 44447 52326
rect 44483 52201 44597 52359
tri 44633 52326 44649 52342 se
rect 44649 52326 44726 52342
rect 44633 52260 44726 52326
rect 44354 52125 44726 52201
rect 44354 52000 44447 52066
rect 44354 51984 44431 52000
tri 44431 51984 44447 52000 nw
rect 44483 51967 44597 52125
rect 44633 52000 44726 52066
tri 44633 51984 44649 52000 ne
rect 44649 51984 44726 52000
rect 44466 51885 44614 51967
rect 44354 51852 44431 51868
tri 44431 51852 44447 51868 sw
rect 44354 51786 44447 51852
rect 44354 51684 44447 51750
rect 44354 51668 44431 51684
tri 44431 51668 44447 51684 nw
rect 44483 51651 44597 51885
tri 44633 51852 44649 51868 se
rect 44649 51852 44726 51868
rect 44633 51786 44726 51852
rect 44633 51684 44726 51750
tri 44633 51668 44649 51684 ne
rect 44649 51668 44726 51684
rect 44466 51569 44614 51651
rect 44354 51536 44431 51552
tri 44431 51536 44447 51552 sw
rect 44354 51470 44447 51536
rect 44483 51411 44597 51569
tri 44633 51536 44649 51552 se
rect 44649 51536 44726 51552
rect 44633 51470 44726 51536
rect 44354 51335 44726 51411
rect 44354 51210 44447 51276
rect 44354 51194 44431 51210
tri 44431 51194 44447 51210 nw
rect 44483 51177 44597 51335
rect 44633 51210 44726 51276
tri 44633 51194 44649 51210 ne
rect 44649 51194 44726 51210
rect 44466 51095 44614 51177
rect 44354 51062 44431 51078
tri 44431 51062 44447 51078 sw
rect 44354 50996 44447 51062
rect 44354 50894 44447 50960
rect 44354 50878 44431 50894
tri 44431 50878 44447 50894 nw
rect 44483 50861 44597 51095
tri 44633 51062 44649 51078 se
rect 44649 51062 44726 51078
rect 44633 50996 44726 51062
rect 44633 50894 44726 50960
tri 44633 50878 44649 50894 ne
rect 44649 50878 44726 50894
rect 44466 50779 44614 50861
rect 44354 50746 44431 50762
tri 44431 50746 44447 50762 sw
rect 44354 50680 44447 50746
rect 44483 50621 44597 50779
tri 44633 50746 44649 50762 se
rect 44649 50746 44726 50762
rect 44633 50680 44726 50746
rect 44354 50545 44726 50621
rect 44354 50420 44447 50486
rect 44354 50404 44431 50420
tri 44431 50404 44447 50420 nw
rect 44483 50387 44597 50545
rect 44633 50420 44726 50486
tri 44633 50404 44649 50420 ne
rect 44649 50404 44726 50420
rect 44466 50305 44614 50387
rect 44354 50272 44431 50288
tri 44431 50272 44447 50288 sw
rect 44354 50206 44447 50272
rect 44354 50104 44447 50170
rect 44354 50088 44431 50104
tri 44431 50088 44447 50104 nw
rect 44483 50071 44597 50305
tri 44633 50272 44649 50288 se
rect 44649 50272 44726 50288
rect 44633 50206 44726 50272
rect 44633 50104 44726 50170
tri 44633 50088 44649 50104 ne
rect 44649 50088 44726 50104
rect 44466 49989 44614 50071
rect 44354 49956 44431 49972
tri 44431 49956 44447 49972 sw
rect 44354 49890 44447 49956
rect 44483 49831 44597 49989
tri 44633 49956 44649 49972 se
rect 44649 49956 44726 49972
rect 44633 49890 44726 49956
rect 44354 49755 44726 49831
rect 44354 49630 44447 49696
rect 44354 49614 44431 49630
tri 44431 49614 44447 49630 nw
rect 44483 49597 44597 49755
rect 44633 49630 44726 49696
tri 44633 49614 44649 49630 ne
rect 44649 49614 44726 49630
rect 44466 49515 44614 49597
rect 44354 49482 44431 49498
tri 44431 49482 44447 49498 sw
rect 44354 49416 44447 49482
rect 44354 49314 44447 49380
rect 44354 49298 44431 49314
tri 44431 49298 44447 49314 nw
rect 44483 49281 44597 49515
tri 44633 49482 44649 49498 se
rect 44649 49482 44726 49498
rect 44633 49416 44726 49482
rect 44633 49314 44726 49380
tri 44633 49298 44649 49314 ne
rect 44649 49298 44726 49314
rect 44466 49199 44614 49281
rect 44354 49166 44431 49182
tri 44431 49166 44447 49182 sw
rect 44354 49100 44447 49166
rect 44483 49041 44597 49199
tri 44633 49166 44649 49182 se
rect 44649 49166 44726 49182
rect 44633 49100 44726 49166
rect 44354 48965 44726 49041
rect 44354 48840 44447 48906
rect 44354 48824 44431 48840
tri 44431 48824 44447 48840 nw
rect 44483 48807 44597 48965
rect 44633 48840 44726 48906
tri 44633 48824 44649 48840 ne
rect 44649 48824 44726 48840
rect 44466 48725 44614 48807
rect 44354 48692 44431 48708
tri 44431 48692 44447 48708 sw
rect 44354 48626 44447 48692
rect 44354 48524 44447 48590
rect 44354 48508 44431 48524
tri 44431 48508 44447 48524 nw
rect 44483 48491 44597 48725
tri 44633 48692 44649 48708 se
rect 44649 48692 44726 48708
rect 44633 48626 44726 48692
rect 44633 48524 44726 48590
tri 44633 48508 44649 48524 ne
rect 44649 48508 44726 48524
rect 44466 48409 44614 48491
rect 44354 48376 44431 48392
tri 44431 48376 44447 48392 sw
rect 44354 48310 44447 48376
rect 44483 48251 44597 48409
tri 44633 48376 44649 48392 se
rect 44649 48376 44726 48392
rect 44633 48310 44726 48376
rect 44354 48175 44726 48251
rect 44354 48050 44447 48116
rect 44354 48034 44431 48050
tri 44431 48034 44447 48050 nw
rect 44483 48017 44597 48175
rect 44633 48050 44726 48116
tri 44633 48034 44649 48050 ne
rect 44649 48034 44726 48050
rect 44466 47935 44614 48017
rect 44354 47902 44431 47918
tri 44431 47902 44447 47918 sw
rect 44354 47836 44447 47902
rect 44354 47734 44447 47800
rect 44354 47718 44431 47734
tri 44431 47718 44447 47734 nw
rect 44483 47701 44597 47935
tri 44633 47902 44649 47918 se
rect 44649 47902 44726 47918
rect 44633 47836 44726 47902
rect 44633 47734 44726 47800
tri 44633 47718 44649 47734 ne
rect 44649 47718 44726 47734
rect 44466 47619 44614 47701
rect 44354 47586 44431 47602
tri 44431 47586 44447 47602 sw
rect 44354 47520 44447 47586
rect 44483 47461 44597 47619
tri 44633 47586 44649 47602 se
rect 44649 47586 44726 47602
rect 44633 47520 44726 47586
rect 44354 47385 44726 47461
rect 44354 47260 44447 47326
rect 44354 47244 44431 47260
tri 44431 47244 44447 47260 nw
rect 44483 47227 44597 47385
rect 44633 47260 44726 47326
tri 44633 47244 44649 47260 ne
rect 44649 47244 44726 47260
rect 44466 47145 44614 47227
rect 44354 47112 44431 47128
tri 44431 47112 44447 47128 sw
rect 44354 47046 44447 47112
rect 44354 46944 44447 47010
rect 44354 46928 44431 46944
tri 44431 46928 44447 46944 nw
rect 44483 46911 44597 47145
tri 44633 47112 44649 47128 se
rect 44649 47112 44726 47128
rect 44633 47046 44726 47112
rect 44633 46944 44726 47010
tri 44633 46928 44649 46944 ne
rect 44649 46928 44726 46944
rect 44466 46829 44614 46911
rect 44354 46796 44431 46812
tri 44431 46796 44447 46812 sw
rect 44354 46730 44447 46796
rect 44483 46671 44597 46829
tri 44633 46796 44649 46812 se
rect 44649 46796 44726 46812
rect 44633 46730 44726 46796
rect 44354 46595 44726 46671
rect 44354 46470 44447 46536
rect 44354 46454 44431 46470
tri 44431 46454 44447 46470 nw
rect 44483 46437 44597 46595
rect 44633 46470 44726 46536
tri 44633 46454 44649 46470 ne
rect 44649 46454 44726 46470
rect 44466 46355 44614 46437
rect 44354 46322 44431 46338
tri 44431 46322 44447 46338 sw
rect 44354 46256 44447 46322
rect 44354 46154 44447 46220
rect 44354 46138 44431 46154
tri 44431 46138 44447 46154 nw
rect 44483 46121 44597 46355
tri 44633 46322 44649 46338 se
rect 44649 46322 44726 46338
rect 44633 46256 44726 46322
rect 44633 46154 44726 46220
tri 44633 46138 44649 46154 ne
rect 44649 46138 44726 46154
rect 44466 46039 44614 46121
rect 44354 46006 44431 46022
tri 44431 46006 44447 46022 sw
rect 44354 45940 44447 46006
rect 44483 45881 44597 46039
tri 44633 46006 44649 46022 se
rect 44649 46006 44726 46022
rect 44633 45940 44726 46006
rect 44354 45805 44726 45881
rect 44354 45680 44447 45746
rect 44354 45664 44431 45680
tri 44431 45664 44447 45680 nw
rect 44483 45647 44597 45805
rect 44633 45680 44726 45746
tri 44633 45664 44649 45680 ne
rect 44649 45664 44726 45680
rect 44466 45565 44614 45647
rect 44354 45532 44431 45548
tri 44431 45532 44447 45548 sw
rect 44354 45466 44447 45532
rect 44354 45364 44447 45430
rect 44354 45348 44431 45364
tri 44431 45348 44447 45364 nw
rect 44483 45331 44597 45565
tri 44633 45532 44649 45548 se
rect 44649 45532 44726 45548
rect 44633 45466 44726 45532
rect 44633 45364 44726 45430
tri 44633 45348 44649 45364 ne
rect 44649 45348 44726 45364
rect 44466 45249 44614 45331
rect 44354 45216 44431 45232
tri 44431 45216 44447 45232 sw
rect 44354 45150 44447 45216
rect 44483 45091 44597 45249
tri 44633 45216 44649 45232 se
rect 44649 45216 44726 45232
rect 44633 45150 44726 45216
rect 44354 45015 44726 45091
rect 44354 44890 44447 44956
rect 44354 44874 44431 44890
tri 44431 44874 44447 44890 nw
rect 44483 44857 44597 45015
rect 44633 44890 44726 44956
tri 44633 44874 44649 44890 ne
rect 44649 44874 44726 44890
rect 44466 44775 44614 44857
rect 44354 44742 44431 44758
tri 44431 44742 44447 44758 sw
rect 44354 44676 44447 44742
rect 44354 44574 44447 44640
rect 44354 44558 44431 44574
tri 44431 44558 44447 44574 nw
rect 44483 44541 44597 44775
tri 44633 44742 44649 44758 se
rect 44649 44742 44726 44758
rect 44633 44676 44726 44742
rect 44633 44574 44726 44640
tri 44633 44558 44649 44574 ne
rect 44649 44558 44726 44574
rect 44466 44459 44614 44541
rect 44354 44426 44431 44442
tri 44431 44426 44447 44442 sw
rect 44354 44360 44447 44426
rect 44483 44301 44597 44459
tri 44633 44426 44649 44442 se
rect 44649 44426 44726 44442
rect 44633 44360 44726 44426
rect 44354 44225 44726 44301
rect 44354 44100 44447 44166
rect 44354 44084 44431 44100
tri 44431 44084 44447 44100 nw
rect 44483 44067 44597 44225
rect 44633 44100 44726 44166
tri 44633 44084 44649 44100 ne
rect 44649 44084 44726 44100
rect 44466 43985 44614 44067
rect 44354 43952 44431 43968
tri 44431 43952 44447 43968 sw
rect 44354 43886 44447 43952
rect 44354 43784 44447 43850
rect 44354 43768 44431 43784
tri 44431 43768 44447 43784 nw
rect 44483 43751 44597 43985
tri 44633 43952 44649 43968 se
rect 44649 43952 44726 43968
rect 44633 43886 44726 43952
rect 44633 43784 44726 43850
tri 44633 43768 44649 43784 ne
rect 44649 43768 44726 43784
rect 44466 43669 44614 43751
rect 44354 43636 44431 43652
tri 44431 43636 44447 43652 sw
rect 44354 43570 44447 43636
rect 44483 43511 44597 43669
tri 44633 43636 44649 43652 se
rect 44649 43636 44726 43652
rect 44633 43570 44726 43636
rect 44354 43435 44726 43511
rect 44354 43310 44447 43376
rect 44354 43294 44431 43310
tri 44431 43294 44447 43310 nw
rect 44483 43277 44597 43435
rect 44633 43310 44726 43376
tri 44633 43294 44649 43310 ne
rect 44649 43294 44726 43310
rect 44466 43195 44614 43277
rect 44354 43162 44431 43178
tri 44431 43162 44447 43178 sw
rect 44354 43096 44447 43162
rect 44354 42994 44447 43060
rect 44354 42978 44431 42994
tri 44431 42978 44447 42994 nw
rect 44483 42961 44597 43195
tri 44633 43162 44649 43178 se
rect 44649 43162 44726 43178
rect 44633 43096 44726 43162
rect 44633 42994 44726 43060
tri 44633 42978 44649 42994 ne
rect 44649 42978 44726 42994
rect 44466 42879 44614 42961
rect 44354 42846 44431 42862
tri 44431 42846 44447 42862 sw
rect 44354 42780 44447 42846
rect 44483 42721 44597 42879
tri 44633 42846 44649 42862 se
rect 44649 42846 44726 42862
rect 44633 42780 44726 42846
rect 44354 42645 44726 42721
rect 44354 42520 44447 42586
rect 44354 42504 44431 42520
tri 44431 42504 44447 42520 nw
rect 44483 42487 44597 42645
rect 44633 42520 44726 42586
tri 44633 42504 44649 42520 ne
rect 44649 42504 44726 42520
rect 44466 42405 44614 42487
rect 44354 42372 44431 42388
tri 44431 42372 44447 42388 sw
rect 44354 42306 44447 42372
rect 44354 42204 44447 42270
rect 44354 42188 44431 42204
tri 44431 42188 44447 42204 nw
rect 44483 42171 44597 42405
tri 44633 42372 44649 42388 se
rect 44649 42372 44726 42388
rect 44633 42306 44726 42372
rect 44633 42204 44726 42270
tri 44633 42188 44649 42204 ne
rect 44649 42188 44726 42204
rect 44466 42089 44614 42171
rect 44354 42056 44431 42072
tri 44431 42056 44447 42072 sw
rect 44354 41990 44447 42056
rect 44483 41931 44597 42089
tri 44633 42056 44649 42072 se
rect 44649 42056 44726 42072
rect 44633 41990 44726 42056
rect 44354 41855 44726 41931
rect 44354 41730 44447 41796
rect 44354 41714 44431 41730
tri 44431 41714 44447 41730 nw
rect 44483 41697 44597 41855
rect 44633 41730 44726 41796
tri 44633 41714 44649 41730 ne
rect 44649 41714 44726 41730
rect 44466 41615 44614 41697
rect 44354 41582 44431 41598
tri 44431 41582 44447 41598 sw
rect 44354 41516 44447 41582
rect 44354 41414 44447 41480
rect 44354 41398 44431 41414
tri 44431 41398 44447 41414 nw
rect 44483 41381 44597 41615
tri 44633 41582 44649 41598 se
rect 44649 41582 44726 41598
rect 44633 41516 44726 41582
rect 44633 41414 44726 41480
tri 44633 41398 44649 41414 ne
rect 44649 41398 44726 41414
rect 44466 41299 44614 41381
rect 44354 41266 44431 41282
tri 44431 41266 44447 41282 sw
rect 44354 41200 44447 41266
rect 44483 41141 44597 41299
tri 44633 41266 44649 41282 se
rect 44649 41266 44726 41282
rect 44633 41200 44726 41266
rect 44354 41065 44726 41141
rect 44354 40940 44447 41006
rect 44354 40924 44431 40940
tri 44431 40924 44447 40940 nw
rect 44483 40907 44597 41065
rect 44633 40940 44726 41006
tri 44633 40924 44649 40940 ne
rect 44649 40924 44726 40940
rect 44466 40825 44614 40907
rect 44354 40792 44431 40808
tri 44431 40792 44447 40808 sw
rect 44354 40726 44447 40792
rect 44354 40624 44447 40690
rect 44354 40608 44431 40624
tri 44431 40608 44447 40624 nw
rect 44483 40591 44597 40825
tri 44633 40792 44649 40808 se
rect 44649 40792 44726 40808
rect 44633 40726 44726 40792
rect 44633 40624 44726 40690
tri 44633 40608 44649 40624 ne
rect 44649 40608 44726 40624
rect 44466 40509 44614 40591
rect 44354 40476 44431 40492
tri 44431 40476 44447 40492 sw
rect 44354 40410 44447 40476
rect 44483 40351 44597 40509
tri 44633 40476 44649 40492 se
rect 44649 40476 44726 40492
rect 44633 40410 44726 40476
rect 44354 40275 44726 40351
rect 44354 40150 44447 40216
rect 44354 40134 44431 40150
tri 44431 40134 44447 40150 nw
rect 44483 40117 44597 40275
rect 44633 40150 44726 40216
tri 44633 40134 44649 40150 ne
rect 44649 40134 44726 40150
rect 44466 40035 44614 40117
rect 44354 40002 44431 40018
tri 44431 40002 44447 40018 sw
rect 44354 39936 44447 40002
rect 44354 39834 44447 39900
rect 44354 39818 44431 39834
tri 44431 39818 44447 39834 nw
rect 44483 39801 44597 40035
tri 44633 40002 44649 40018 se
rect 44649 40002 44726 40018
rect 44633 39936 44726 40002
rect 44633 39834 44726 39900
tri 44633 39818 44649 39834 ne
rect 44649 39818 44726 39834
rect 44466 39719 44614 39801
rect 44354 39686 44431 39702
tri 44431 39686 44447 39702 sw
rect 44354 39620 44447 39686
rect 44483 39561 44597 39719
tri 44633 39686 44649 39702 se
rect 44649 39686 44726 39702
rect 44633 39620 44726 39686
rect 44354 39485 44726 39561
rect 44354 39360 44447 39426
rect 44354 39344 44431 39360
tri 44431 39344 44447 39360 nw
rect 44483 39327 44597 39485
rect 44633 39360 44726 39426
tri 44633 39344 44649 39360 ne
rect 44649 39344 44726 39360
rect 44466 39245 44614 39327
rect 44354 39212 44431 39228
tri 44431 39212 44447 39228 sw
rect 44354 39146 44447 39212
rect 44354 39044 44447 39110
rect 44354 39028 44431 39044
tri 44431 39028 44447 39044 nw
rect 44483 39011 44597 39245
tri 44633 39212 44649 39228 se
rect 44649 39212 44726 39228
rect 44633 39146 44726 39212
rect 44633 39044 44726 39110
tri 44633 39028 44649 39044 ne
rect 44649 39028 44726 39044
rect 44466 38929 44614 39011
rect 44354 38896 44431 38912
tri 44431 38896 44447 38912 sw
rect 44354 38830 44447 38896
rect 44483 38771 44597 38929
tri 44633 38896 44649 38912 se
rect 44649 38896 44726 38912
rect 44633 38830 44726 38896
rect 44354 38695 44726 38771
rect 44354 38570 44447 38636
rect 44354 38554 44431 38570
tri 44431 38554 44447 38570 nw
rect 44483 38537 44597 38695
rect 44633 38570 44726 38636
tri 44633 38554 44649 38570 ne
rect 44649 38554 44726 38570
rect 44466 38455 44614 38537
rect 44354 38422 44431 38438
tri 44431 38422 44447 38438 sw
rect 44354 38356 44447 38422
rect 44354 38254 44447 38320
rect 44354 38238 44431 38254
tri 44431 38238 44447 38254 nw
rect 44483 38221 44597 38455
tri 44633 38422 44649 38438 se
rect 44649 38422 44726 38438
rect 44633 38356 44726 38422
rect 44633 38254 44726 38320
tri 44633 38238 44649 38254 ne
rect 44649 38238 44726 38254
rect 44466 38139 44614 38221
rect 44354 38106 44431 38122
tri 44431 38106 44447 38122 sw
rect 44354 38040 44447 38106
rect 44483 37981 44597 38139
tri 44633 38106 44649 38122 se
rect 44649 38106 44726 38122
rect 44633 38040 44726 38106
rect 44354 37905 44726 37981
rect 44354 37780 44447 37846
rect 44354 37764 44431 37780
tri 44431 37764 44447 37780 nw
rect 44483 37747 44597 37905
rect 44633 37780 44726 37846
tri 44633 37764 44649 37780 ne
rect 44649 37764 44726 37780
rect 44466 37665 44614 37747
rect 44354 37632 44431 37648
tri 44431 37632 44447 37648 sw
rect 44354 37566 44447 37632
rect 44354 37464 44447 37530
rect 44354 37448 44431 37464
tri 44431 37448 44447 37464 nw
rect 44483 37431 44597 37665
tri 44633 37632 44649 37648 se
rect 44649 37632 44726 37648
rect 44633 37566 44726 37632
rect 44633 37464 44726 37530
tri 44633 37448 44649 37464 ne
rect 44649 37448 44726 37464
rect 44466 37349 44614 37431
rect 44354 37316 44431 37332
tri 44431 37316 44447 37332 sw
rect 44354 37250 44447 37316
rect 44483 37191 44597 37349
tri 44633 37316 44649 37332 se
rect 44649 37316 44726 37332
rect 44633 37250 44726 37316
rect 44354 37115 44726 37191
rect 44354 36990 44447 37056
rect 44354 36974 44431 36990
tri 44431 36974 44447 36990 nw
rect 44483 36957 44597 37115
rect 44633 36990 44726 37056
tri 44633 36974 44649 36990 ne
rect 44649 36974 44726 36990
rect 44466 36875 44614 36957
rect 44354 36842 44431 36858
tri 44431 36842 44447 36858 sw
rect 44354 36776 44447 36842
rect 44354 36674 44447 36740
rect 44354 36658 44431 36674
tri 44431 36658 44447 36674 nw
rect 44483 36641 44597 36875
tri 44633 36842 44649 36858 se
rect 44649 36842 44726 36858
rect 44633 36776 44726 36842
rect 44633 36674 44726 36740
tri 44633 36658 44649 36674 ne
rect 44649 36658 44726 36674
rect 44466 36559 44614 36641
rect 44354 36526 44431 36542
tri 44431 36526 44447 36542 sw
rect 44354 36460 44447 36526
rect 44483 36401 44597 36559
tri 44633 36526 44649 36542 se
rect 44649 36526 44726 36542
rect 44633 36460 44726 36526
rect 44354 36325 44726 36401
rect 44354 36200 44447 36266
rect 44354 36184 44431 36200
tri 44431 36184 44447 36200 nw
rect 44483 36167 44597 36325
rect 44633 36200 44726 36266
tri 44633 36184 44649 36200 ne
rect 44649 36184 44726 36200
rect 44466 36085 44614 36167
rect 44354 36052 44431 36068
tri 44431 36052 44447 36068 sw
rect 44354 35986 44447 36052
rect 44354 35884 44447 35950
rect 44354 35868 44431 35884
tri 44431 35868 44447 35884 nw
rect 44483 35851 44597 36085
tri 44633 36052 44649 36068 se
rect 44649 36052 44726 36068
rect 44633 35986 44726 36052
rect 44633 35884 44726 35950
tri 44633 35868 44649 35884 ne
rect 44649 35868 44726 35884
rect 44466 35769 44614 35851
rect 44354 35736 44431 35752
tri 44431 35736 44447 35752 sw
rect 44354 35670 44447 35736
rect 44483 35611 44597 35769
tri 44633 35736 44649 35752 se
rect 44649 35736 44726 35752
rect 44633 35670 44726 35736
rect 44354 35535 44726 35611
rect 44354 35410 44447 35476
rect 44354 35394 44431 35410
tri 44431 35394 44447 35410 nw
rect 44483 35377 44597 35535
rect 44633 35410 44726 35476
tri 44633 35394 44649 35410 ne
rect 44649 35394 44726 35410
rect 44466 35295 44614 35377
rect 44354 35262 44431 35278
tri 44431 35262 44447 35278 sw
rect 44354 35196 44447 35262
rect 44354 35094 44447 35160
rect 44354 35078 44431 35094
tri 44431 35078 44447 35094 nw
rect 44483 35061 44597 35295
tri 44633 35262 44649 35278 se
rect 44649 35262 44726 35278
rect 44633 35196 44726 35262
rect 44633 35094 44726 35160
tri 44633 35078 44649 35094 ne
rect 44649 35078 44726 35094
rect 44466 34979 44614 35061
rect 44354 34946 44431 34962
tri 44431 34946 44447 34962 sw
rect 44354 34880 44447 34946
rect 44483 34821 44597 34979
tri 44633 34946 44649 34962 se
rect 44649 34946 44726 34962
rect 44633 34880 44726 34946
rect 44354 34745 44726 34821
rect 44354 34620 44447 34686
rect 44354 34604 44431 34620
tri 44431 34604 44447 34620 nw
rect 44483 34587 44597 34745
rect 44633 34620 44726 34686
tri 44633 34604 44649 34620 ne
rect 44649 34604 44726 34620
rect 44466 34505 44614 34587
rect 44354 34472 44431 34488
tri 44431 34472 44447 34488 sw
rect 44354 34406 44447 34472
rect 44354 34304 44447 34370
rect 44354 34288 44431 34304
tri 44431 34288 44447 34304 nw
rect 44483 34271 44597 34505
tri 44633 34472 44649 34488 se
rect 44649 34472 44726 34488
rect 44633 34406 44726 34472
rect 44633 34304 44726 34370
tri 44633 34288 44649 34304 ne
rect 44649 34288 44726 34304
rect 44466 34189 44614 34271
rect 44354 34156 44431 34172
tri 44431 34156 44447 34172 sw
rect 44354 34090 44447 34156
rect 44483 34031 44597 34189
tri 44633 34156 44649 34172 se
rect 44649 34156 44726 34172
rect 44633 34090 44726 34156
rect 44354 33955 44726 34031
rect 44354 33830 44447 33896
rect 44354 33814 44431 33830
tri 44431 33814 44447 33830 nw
rect 44483 33797 44597 33955
rect 44633 33830 44726 33896
tri 44633 33814 44649 33830 ne
rect 44649 33814 44726 33830
rect 44466 33715 44614 33797
rect 44354 33682 44431 33698
tri 44431 33682 44447 33698 sw
rect 44354 33616 44447 33682
rect 44354 33514 44447 33580
rect 44354 33498 44431 33514
tri 44431 33498 44447 33514 nw
rect 44483 33481 44597 33715
tri 44633 33682 44649 33698 se
rect 44649 33682 44726 33698
rect 44633 33616 44726 33682
rect 44633 33514 44726 33580
tri 44633 33498 44649 33514 ne
rect 44649 33498 44726 33514
rect 44466 33399 44614 33481
rect 44354 33366 44431 33382
tri 44431 33366 44447 33382 sw
rect 44354 33300 44447 33366
rect 44483 33241 44597 33399
tri 44633 33366 44649 33382 se
rect 44649 33366 44726 33382
rect 44633 33300 44726 33366
rect 44354 33165 44726 33241
rect 44354 33040 44447 33106
rect 44354 33024 44431 33040
tri 44431 33024 44447 33040 nw
rect 44483 33007 44597 33165
rect 44633 33040 44726 33106
tri 44633 33024 44649 33040 ne
rect 44649 33024 44726 33040
rect 44466 32925 44614 33007
rect 44354 32892 44431 32908
tri 44431 32892 44447 32908 sw
rect 44354 32826 44447 32892
rect 44354 32724 44447 32790
rect 44354 32708 44431 32724
tri 44431 32708 44447 32724 nw
rect 44483 32691 44597 32925
tri 44633 32892 44649 32908 se
rect 44649 32892 44726 32908
rect 44633 32826 44726 32892
rect 44633 32724 44726 32790
tri 44633 32708 44649 32724 ne
rect 44649 32708 44726 32724
rect 44466 32609 44614 32691
rect 44354 32576 44431 32592
tri 44431 32576 44447 32592 sw
rect 44354 32510 44447 32576
rect 44483 32451 44597 32609
tri 44633 32576 44649 32592 se
rect 44649 32576 44726 32592
rect 44633 32510 44726 32576
rect 44354 32375 44726 32451
rect 44354 32250 44447 32316
rect 44354 32234 44431 32250
tri 44431 32234 44447 32250 nw
rect 44483 32217 44597 32375
rect 44633 32250 44726 32316
tri 44633 32234 44649 32250 ne
rect 44649 32234 44726 32250
rect 44466 32135 44614 32217
rect 44354 32102 44431 32118
tri 44431 32102 44447 32118 sw
rect 44354 32036 44447 32102
rect 44354 31934 44447 32000
rect 44354 31918 44431 31934
tri 44431 31918 44447 31934 nw
rect 44483 31901 44597 32135
tri 44633 32102 44649 32118 se
rect 44649 32102 44726 32118
rect 44633 32036 44726 32102
rect 44633 31934 44726 32000
tri 44633 31918 44649 31934 ne
rect 44649 31918 44726 31934
rect 44466 31819 44614 31901
rect 44354 31786 44431 31802
tri 44431 31786 44447 31802 sw
rect 44354 31720 44447 31786
rect 44483 31661 44597 31819
tri 44633 31786 44649 31802 se
rect 44649 31786 44726 31802
rect 44633 31720 44726 31786
rect 44354 31585 44726 31661
rect 44354 31460 44447 31526
rect 44354 31444 44431 31460
tri 44431 31444 44447 31460 nw
rect 44483 31427 44597 31585
rect 44633 31460 44726 31526
tri 44633 31444 44649 31460 ne
rect 44649 31444 44726 31460
rect 44466 31345 44614 31427
rect 44354 31312 44431 31328
tri 44431 31312 44447 31328 sw
rect 44354 31246 44447 31312
rect 44354 31144 44447 31210
rect 44354 31128 44431 31144
tri 44431 31128 44447 31144 nw
rect 44483 31111 44597 31345
tri 44633 31312 44649 31328 se
rect 44649 31312 44726 31328
rect 44633 31246 44726 31312
rect 44633 31144 44726 31210
tri 44633 31128 44649 31144 ne
rect 44649 31128 44726 31144
rect 44466 31029 44614 31111
rect 44354 30996 44431 31012
tri 44431 30996 44447 31012 sw
rect 44354 30930 44447 30996
rect 44483 30871 44597 31029
tri 44633 30996 44649 31012 se
rect 44649 30996 44726 31012
rect 44633 30930 44726 30996
rect 44354 30795 44726 30871
rect 44354 30670 44447 30736
rect 44354 30654 44431 30670
tri 44431 30654 44447 30670 nw
rect 44483 30637 44597 30795
rect 44633 30670 44726 30736
tri 44633 30654 44649 30670 ne
rect 44649 30654 44726 30670
rect 44466 30555 44614 30637
rect 44354 30522 44431 30538
tri 44431 30522 44447 30538 sw
rect 44354 30456 44447 30522
rect 44354 30354 44447 30420
rect 44354 30338 44431 30354
tri 44431 30338 44447 30354 nw
rect 44483 30321 44597 30555
tri 44633 30522 44649 30538 se
rect 44649 30522 44726 30538
rect 44633 30456 44726 30522
rect 44633 30354 44726 30420
tri 44633 30338 44649 30354 ne
rect 44649 30338 44726 30354
rect 44466 30239 44614 30321
rect 44354 30206 44431 30222
tri 44431 30206 44447 30222 sw
rect 44354 30140 44447 30206
rect 44483 30081 44597 30239
tri 44633 30206 44649 30222 se
rect 44649 30206 44726 30222
rect 44633 30140 44726 30206
rect 44354 30005 44726 30081
rect 44354 29880 44447 29946
rect 44354 29864 44431 29880
tri 44431 29864 44447 29880 nw
rect 44483 29847 44597 30005
rect 44633 29880 44726 29946
tri 44633 29864 44649 29880 ne
rect 44649 29864 44726 29880
rect 44466 29765 44614 29847
rect 44354 29732 44431 29748
tri 44431 29732 44447 29748 sw
rect 44354 29666 44447 29732
rect 44354 29564 44447 29630
rect 44354 29548 44431 29564
tri 44431 29548 44447 29564 nw
rect 44483 29531 44597 29765
tri 44633 29732 44649 29748 se
rect 44649 29732 44726 29748
rect 44633 29666 44726 29732
rect 44633 29564 44726 29630
tri 44633 29548 44649 29564 ne
rect 44649 29548 44726 29564
rect 44466 29449 44614 29531
rect 44354 29416 44431 29432
tri 44431 29416 44447 29432 sw
rect 44354 29350 44447 29416
rect 44483 29291 44597 29449
tri 44633 29416 44649 29432 se
rect 44649 29416 44726 29432
rect 44633 29350 44726 29416
rect 44354 29215 44726 29291
rect 44354 29090 44447 29156
rect 44354 29074 44431 29090
tri 44431 29074 44447 29090 nw
rect 44483 29057 44597 29215
rect 44633 29090 44726 29156
tri 44633 29074 44649 29090 ne
rect 44649 29074 44726 29090
rect 44466 28975 44614 29057
rect 44354 28942 44431 28958
tri 44431 28942 44447 28958 sw
rect 44354 28876 44447 28942
rect 44483 28833 44597 28975
tri 44633 28942 44649 28958 se
rect 44649 28942 44726 28958
rect 44633 28876 44726 28942
rect 44762 28463 44798 80603
rect 44834 28463 44870 80603
rect 44906 80445 44942 80603
rect 44898 80303 44950 80445
rect 44906 28763 44942 80303
rect 44898 28621 44950 28763
rect 44906 28463 44942 28621
rect 44978 28463 45014 80603
rect 45050 28463 45086 80603
rect 45122 28833 45206 80233
rect 45242 28463 45278 80603
rect 45314 28463 45350 80603
rect 45386 80445 45422 80603
rect 45378 80303 45430 80445
rect 45386 28763 45422 80303
rect 45378 28621 45430 28763
rect 45386 28463 45422 28621
rect 45458 28463 45494 80603
rect 45530 28463 45566 80603
rect 45602 80124 45695 80190
rect 45602 80108 45679 80124
tri 45679 80108 45695 80124 nw
rect 45731 80091 45845 80233
rect 45881 80124 45974 80190
tri 45881 80108 45897 80124 ne
rect 45897 80108 45974 80124
rect 45714 80009 45862 80091
rect 45602 79976 45679 79992
tri 45679 79976 45695 79992 sw
rect 45602 79910 45695 79976
rect 45731 79851 45845 80009
tri 45881 79976 45897 79992 se
rect 45897 79976 45974 79992
rect 45881 79910 45974 79976
rect 45602 79775 45974 79851
rect 45602 79650 45695 79716
rect 45602 79634 45679 79650
tri 45679 79634 45695 79650 nw
rect 45731 79617 45845 79775
rect 45881 79650 45974 79716
tri 45881 79634 45897 79650 ne
rect 45897 79634 45974 79650
rect 45714 79535 45862 79617
rect 45602 79502 45679 79518
tri 45679 79502 45695 79518 sw
rect 45602 79436 45695 79502
rect 45602 79334 45695 79400
rect 45602 79318 45679 79334
tri 45679 79318 45695 79334 nw
rect 45731 79301 45845 79535
tri 45881 79502 45897 79518 se
rect 45897 79502 45974 79518
rect 45881 79436 45974 79502
rect 45881 79334 45974 79400
tri 45881 79318 45897 79334 ne
rect 45897 79318 45974 79334
rect 45714 79219 45862 79301
rect 45602 79186 45679 79202
tri 45679 79186 45695 79202 sw
rect 45602 79120 45695 79186
rect 45731 79061 45845 79219
tri 45881 79186 45897 79202 se
rect 45897 79186 45974 79202
rect 45881 79120 45974 79186
rect 45602 78985 45974 79061
rect 45602 78860 45695 78926
rect 45602 78844 45679 78860
tri 45679 78844 45695 78860 nw
rect 45731 78827 45845 78985
rect 45881 78860 45974 78926
tri 45881 78844 45897 78860 ne
rect 45897 78844 45974 78860
rect 45714 78745 45862 78827
rect 45602 78712 45679 78728
tri 45679 78712 45695 78728 sw
rect 45602 78646 45695 78712
rect 45602 78544 45695 78610
rect 45602 78528 45679 78544
tri 45679 78528 45695 78544 nw
rect 45731 78511 45845 78745
tri 45881 78712 45897 78728 se
rect 45897 78712 45974 78728
rect 45881 78646 45974 78712
rect 45881 78544 45974 78610
tri 45881 78528 45897 78544 ne
rect 45897 78528 45974 78544
rect 45714 78429 45862 78511
rect 45602 78396 45679 78412
tri 45679 78396 45695 78412 sw
rect 45602 78330 45695 78396
rect 45731 78271 45845 78429
tri 45881 78396 45897 78412 se
rect 45897 78396 45974 78412
rect 45881 78330 45974 78396
rect 45602 78195 45974 78271
rect 45602 78070 45695 78136
rect 45602 78054 45679 78070
tri 45679 78054 45695 78070 nw
rect 45731 78037 45845 78195
rect 45881 78070 45974 78136
tri 45881 78054 45897 78070 ne
rect 45897 78054 45974 78070
rect 45714 77955 45862 78037
rect 45602 77922 45679 77938
tri 45679 77922 45695 77938 sw
rect 45602 77856 45695 77922
rect 45602 77754 45695 77820
rect 45602 77738 45679 77754
tri 45679 77738 45695 77754 nw
rect 45731 77721 45845 77955
tri 45881 77922 45897 77938 se
rect 45897 77922 45974 77938
rect 45881 77856 45974 77922
rect 45881 77754 45974 77820
tri 45881 77738 45897 77754 ne
rect 45897 77738 45974 77754
rect 45714 77639 45862 77721
rect 45602 77606 45679 77622
tri 45679 77606 45695 77622 sw
rect 45602 77540 45695 77606
rect 45731 77481 45845 77639
tri 45881 77606 45897 77622 se
rect 45897 77606 45974 77622
rect 45881 77540 45974 77606
rect 45602 77405 45974 77481
rect 45602 77280 45695 77346
rect 45602 77264 45679 77280
tri 45679 77264 45695 77280 nw
rect 45731 77247 45845 77405
rect 45881 77280 45974 77346
tri 45881 77264 45897 77280 ne
rect 45897 77264 45974 77280
rect 45714 77165 45862 77247
rect 45602 77132 45679 77148
tri 45679 77132 45695 77148 sw
rect 45602 77066 45695 77132
rect 45602 76964 45695 77030
rect 45602 76948 45679 76964
tri 45679 76948 45695 76964 nw
rect 45731 76931 45845 77165
tri 45881 77132 45897 77148 se
rect 45897 77132 45974 77148
rect 45881 77066 45974 77132
rect 45881 76964 45974 77030
tri 45881 76948 45897 76964 ne
rect 45897 76948 45974 76964
rect 45714 76849 45862 76931
rect 45602 76816 45679 76832
tri 45679 76816 45695 76832 sw
rect 45602 76750 45695 76816
rect 45731 76691 45845 76849
tri 45881 76816 45897 76832 se
rect 45897 76816 45974 76832
rect 45881 76750 45974 76816
rect 45602 76615 45974 76691
rect 45602 76490 45695 76556
rect 45602 76474 45679 76490
tri 45679 76474 45695 76490 nw
rect 45731 76457 45845 76615
rect 45881 76490 45974 76556
tri 45881 76474 45897 76490 ne
rect 45897 76474 45974 76490
rect 45714 76375 45862 76457
rect 45602 76342 45679 76358
tri 45679 76342 45695 76358 sw
rect 45602 76276 45695 76342
rect 45602 76174 45695 76240
rect 45602 76158 45679 76174
tri 45679 76158 45695 76174 nw
rect 45731 76141 45845 76375
tri 45881 76342 45897 76358 se
rect 45897 76342 45974 76358
rect 45881 76276 45974 76342
rect 45881 76174 45974 76240
tri 45881 76158 45897 76174 ne
rect 45897 76158 45974 76174
rect 45714 76059 45862 76141
rect 45602 76026 45679 76042
tri 45679 76026 45695 76042 sw
rect 45602 75960 45695 76026
rect 45731 75901 45845 76059
tri 45881 76026 45897 76042 se
rect 45897 76026 45974 76042
rect 45881 75960 45974 76026
rect 45602 75825 45974 75901
rect 45602 75700 45695 75766
rect 45602 75684 45679 75700
tri 45679 75684 45695 75700 nw
rect 45731 75667 45845 75825
rect 45881 75700 45974 75766
tri 45881 75684 45897 75700 ne
rect 45897 75684 45974 75700
rect 45714 75585 45862 75667
rect 45602 75552 45679 75568
tri 45679 75552 45695 75568 sw
rect 45602 75486 45695 75552
rect 45602 75384 45695 75450
rect 45602 75368 45679 75384
tri 45679 75368 45695 75384 nw
rect 45731 75351 45845 75585
tri 45881 75552 45897 75568 se
rect 45897 75552 45974 75568
rect 45881 75486 45974 75552
rect 45881 75384 45974 75450
tri 45881 75368 45897 75384 ne
rect 45897 75368 45974 75384
rect 45714 75269 45862 75351
rect 45602 75236 45679 75252
tri 45679 75236 45695 75252 sw
rect 45602 75170 45695 75236
rect 45731 75111 45845 75269
tri 45881 75236 45897 75252 se
rect 45897 75236 45974 75252
rect 45881 75170 45974 75236
rect 45602 75035 45974 75111
rect 45602 74910 45695 74976
rect 45602 74894 45679 74910
tri 45679 74894 45695 74910 nw
rect 45731 74877 45845 75035
rect 45881 74910 45974 74976
tri 45881 74894 45897 74910 ne
rect 45897 74894 45974 74910
rect 45714 74795 45862 74877
rect 45602 74762 45679 74778
tri 45679 74762 45695 74778 sw
rect 45602 74696 45695 74762
rect 45602 74594 45695 74660
rect 45602 74578 45679 74594
tri 45679 74578 45695 74594 nw
rect 45731 74561 45845 74795
tri 45881 74762 45897 74778 se
rect 45897 74762 45974 74778
rect 45881 74696 45974 74762
rect 45881 74594 45974 74660
tri 45881 74578 45897 74594 ne
rect 45897 74578 45974 74594
rect 45714 74479 45862 74561
rect 45602 74446 45679 74462
tri 45679 74446 45695 74462 sw
rect 45602 74380 45695 74446
rect 45731 74321 45845 74479
tri 45881 74446 45897 74462 se
rect 45897 74446 45974 74462
rect 45881 74380 45974 74446
rect 45602 74245 45974 74321
rect 45602 74120 45695 74186
rect 45602 74104 45679 74120
tri 45679 74104 45695 74120 nw
rect 45731 74087 45845 74245
rect 45881 74120 45974 74186
tri 45881 74104 45897 74120 ne
rect 45897 74104 45974 74120
rect 45714 74005 45862 74087
rect 45602 73972 45679 73988
tri 45679 73972 45695 73988 sw
rect 45602 73906 45695 73972
rect 45602 73804 45695 73870
rect 45602 73788 45679 73804
tri 45679 73788 45695 73804 nw
rect 45731 73771 45845 74005
tri 45881 73972 45897 73988 se
rect 45897 73972 45974 73988
rect 45881 73906 45974 73972
rect 45881 73804 45974 73870
tri 45881 73788 45897 73804 ne
rect 45897 73788 45974 73804
rect 45714 73689 45862 73771
rect 45602 73656 45679 73672
tri 45679 73656 45695 73672 sw
rect 45602 73590 45695 73656
rect 45731 73531 45845 73689
tri 45881 73656 45897 73672 se
rect 45897 73656 45974 73672
rect 45881 73590 45974 73656
rect 45602 73455 45974 73531
rect 45602 73330 45695 73396
rect 45602 73314 45679 73330
tri 45679 73314 45695 73330 nw
rect 45731 73297 45845 73455
rect 45881 73330 45974 73396
tri 45881 73314 45897 73330 ne
rect 45897 73314 45974 73330
rect 45714 73215 45862 73297
rect 45602 73182 45679 73198
tri 45679 73182 45695 73198 sw
rect 45602 73116 45695 73182
rect 45602 73014 45695 73080
rect 45602 72998 45679 73014
tri 45679 72998 45695 73014 nw
rect 45731 72981 45845 73215
tri 45881 73182 45897 73198 se
rect 45897 73182 45974 73198
rect 45881 73116 45974 73182
rect 45881 73014 45974 73080
tri 45881 72998 45897 73014 ne
rect 45897 72998 45974 73014
rect 45714 72899 45862 72981
rect 45602 72866 45679 72882
tri 45679 72866 45695 72882 sw
rect 45602 72800 45695 72866
rect 45731 72741 45845 72899
tri 45881 72866 45897 72882 se
rect 45897 72866 45974 72882
rect 45881 72800 45974 72866
rect 45602 72665 45974 72741
rect 45602 72540 45695 72606
rect 45602 72524 45679 72540
tri 45679 72524 45695 72540 nw
rect 45731 72507 45845 72665
rect 45881 72540 45974 72606
tri 45881 72524 45897 72540 ne
rect 45897 72524 45974 72540
rect 45714 72425 45862 72507
rect 45602 72392 45679 72408
tri 45679 72392 45695 72408 sw
rect 45602 72326 45695 72392
rect 45602 72224 45695 72290
rect 45602 72208 45679 72224
tri 45679 72208 45695 72224 nw
rect 45731 72191 45845 72425
tri 45881 72392 45897 72408 se
rect 45897 72392 45974 72408
rect 45881 72326 45974 72392
rect 45881 72224 45974 72290
tri 45881 72208 45897 72224 ne
rect 45897 72208 45974 72224
rect 45714 72109 45862 72191
rect 45602 72076 45679 72092
tri 45679 72076 45695 72092 sw
rect 45602 72010 45695 72076
rect 45731 71951 45845 72109
tri 45881 72076 45897 72092 se
rect 45897 72076 45974 72092
rect 45881 72010 45974 72076
rect 45602 71875 45974 71951
rect 45602 71750 45695 71816
rect 45602 71734 45679 71750
tri 45679 71734 45695 71750 nw
rect 45731 71717 45845 71875
rect 45881 71750 45974 71816
tri 45881 71734 45897 71750 ne
rect 45897 71734 45974 71750
rect 45714 71635 45862 71717
rect 45602 71602 45679 71618
tri 45679 71602 45695 71618 sw
rect 45602 71536 45695 71602
rect 45602 71434 45695 71500
rect 45602 71418 45679 71434
tri 45679 71418 45695 71434 nw
rect 45731 71401 45845 71635
tri 45881 71602 45897 71618 se
rect 45897 71602 45974 71618
rect 45881 71536 45974 71602
rect 45881 71434 45974 71500
tri 45881 71418 45897 71434 ne
rect 45897 71418 45974 71434
rect 45714 71319 45862 71401
rect 45602 71286 45679 71302
tri 45679 71286 45695 71302 sw
rect 45602 71220 45695 71286
rect 45731 71161 45845 71319
tri 45881 71286 45897 71302 se
rect 45897 71286 45974 71302
rect 45881 71220 45974 71286
rect 45602 71085 45974 71161
rect 45602 70960 45695 71026
rect 45602 70944 45679 70960
tri 45679 70944 45695 70960 nw
rect 45731 70927 45845 71085
rect 45881 70960 45974 71026
tri 45881 70944 45897 70960 ne
rect 45897 70944 45974 70960
rect 45714 70845 45862 70927
rect 45602 70812 45679 70828
tri 45679 70812 45695 70828 sw
rect 45602 70746 45695 70812
rect 45602 70644 45695 70710
rect 45602 70628 45679 70644
tri 45679 70628 45695 70644 nw
rect 45731 70611 45845 70845
tri 45881 70812 45897 70828 se
rect 45897 70812 45974 70828
rect 45881 70746 45974 70812
rect 45881 70644 45974 70710
tri 45881 70628 45897 70644 ne
rect 45897 70628 45974 70644
rect 45714 70529 45862 70611
rect 45602 70496 45679 70512
tri 45679 70496 45695 70512 sw
rect 45602 70430 45695 70496
rect 45731 70371 45845 70529
tri 45881 70496 45897 70512 se
rect 45897 70496 45974 70512
rect 45881 70430 45974 70496
rect 45602 70295 45974 70371
rect 45602 70170 45695 70236
rect 45602 70154 45679 70170
tri 45679 70154 45695 70170 nw
rect 45731 70137 45845 70295
rect 45881 70170 45974 70236
tri 45881 70154 45897 70170 ne
rect 45897 70154 45974 70170
rect 45714 70055 45862 70137
rect 45602 70022 45679 70038
tri 45679 70022 45695 70038 sw
rect 45602 69956 45695 70022
rect 45602 69854 45695 69920
rect 45602 69838 45679 69854
tri 45679 69838 45695 69854 nw
rect 45731 69821 45845 70055
tri 45881 70022 45897 70038 se
rect 45897 70022 45974 70038
rect 45881 69956 45974 70022
rect 45881 69854 45974 69920
tri 45881 69838 45897 69854 ne
rect 45897 69838 45974 69854
rect 45714 69739 45862 69821
rect 45602 69706 45679 69722
tri 45679 69706 45695 69722 sw
rect 45602 69640 45695 69706
rect 45731 69581 45845 69739
tri 45881 69706 45897 69722 se
rect 45897 69706 45974 69722
rect 45881 69640 45974 69706
rect 45602 69505 45974 69581
rect 45602 69380 45695 69446
rect 45602 69364 45679 69380
tri 45679 69364 45695 69380 nw
rect 45731 69347 45845 69505
rect 45881 69380 45974 69446
tri 45881 69364 45897 69380 ne
rect 45897 69364 45974 69380
rect 45714 69265 45862 69347
rect 45602 69232 45679 69248
tri 45679 69232 45695 69248 sw
rect 45602 69166 45695 69232
rect 45602 69064 45695 69130
rect 45602 69048 45679 69064
tri 45679 69048 45695 69064 nw
rect 45731 69031 45845 69265
tri 45881 69232 45897 69248 se
rect 45897 69232 45974 69248
rect 45881 69166 45974 69232
rect 45881 69064 45974 69130
tri 45881 69048 45897 69064 ne
rect 45897 69048 45974 69064
rect 45714 68949 45862 69031
rect 45602 68916 45679 68932
tri 45679 68916 45695 68932 sw
rect 45602 68850 45695 68916
rect 45731 68791 45845 68949
tri 45881 68916 45897 68932 se
rect 45897 68916 45974 68932
rect 45881 68850 45974 68916
rect 45602 68715 45974 68791
rect 45602 68590 45695 68656
rect 45602 68574 45679 68590
tri 45679 68574 45695 68590 nw
rect 45731 68557 45845 68715
rect 45881 68590 45974 68656
tri 45881 68574 45897 68590 ne
rect 45897 68574 45974 68590
rect 45714 68475 45862 68557
rect 45602 68442 45679 68458
tri 45679 68442 45695 68458 sw
rect 45602 68376 45695 68442
rect 45602 68274 45695 68340
rect 45602 68258 45679 68274
tri 45679 68258 45695 68274 nw
rect 45731 68241 45845 68475
tri 45881 68442 45897 68458 se
rect 45897 68442 45974 68458
rect 45881 68376 45974 68442
rect 45881 68274 45974 68340
tri 45881 68258 45897 68274 ne
rect 45897 68258 45974 68274
rect 45714 68159 45862 68241
rect 45602 68126 45679 68142
tri 45679 68126 45695 68142 sw
rect 45602 68060 45695 68126
rect 45731 68001 45845 68159
tri 45881 68126 45897 68142 se
rect 45897 68126 45974 68142
rect 45881 68060 45974 68126
rect 45602 67925 45974 68001
rect 45602 67800 45695 67866
rect 45602 67784 45679 67800
tri 45679 67784 45695 67800 nw
rect 45731 67767 45845 67925
rect 45881 67800 45974 67866
tri 45881 67784 45897 67800 ne
rect 45897 67784 45974 67800
rect 45714 67685 45862 67767
rect 45602 67652 45679 67668
tri 45679 67652 45695 67668 sw
rect 45602 67586 45695 67652
rect 45602 67484 45695 67550
rect 45602 67468 45679 67484
tri 45679 67468 45695 67484 nw
rect 45731 67451 45845 67685
tri 45881 67652 45897 67668 se
rect 45897 67652 45974 67668
rect 45881 67586 45974 67652
rect 45881 67484 45974 67550
tri 45881 67468 45897 67484 ne
rect 45897 67468 45974 67484
rect 45714 67369 45862 67451
rect 45602 67336 45679 67352
tri 45679 67336 45695 67352 sw
rect 45602 67270 45695 67336
rect 45731 67211 45845 67369
tri 45881 67336 45897 67352 se
rect 45897 67336 45974 67352
rect 45881 67270 45974 67336
rect 45602 67135 45974 67211
rect 45602 67010 45695 67076
rect 45602 66994 45679 67010
tri 45679 66994 45695 67010 nw
rect 45731 66977 45845 67135
rect 45881 67010 45974 67076
tri 45881 66994 45897 67010 ne
rect 45897 66994 45974 67010
rect 45714 66895 45862 66977
rect 45602 66862 45679 66878
tri 45679 66862 45695 66878 sw
rect 45602 66796 45695 66862
rect 45602 66694 45695 66760
rect 45602 66678 45679 66694
tri 45679 66678 45695 66694 nw
rect 45731 66661 45845 66895
tri 45881 66862 45897 66878 se
rect 45897 66862 45974 66878
rect 45881 66796 45974 66862
rect 45881 66694 45974 66760
tri 45881 66678 45897 66694 ne
rect 45897 66678 45974 66694
rect 45714 66579 45862 66661
rect 45602 66546 45679 66562
tri 45679 66546 45695 66562 sw
rect 45602 66480 45695 66546
rect 45731 66421 45845 66579
tri 45881 66546 45897 66562 se
rect 45897 66546 45974 66562
rect 45881 66480 45974 66546
rect 45602 66345 45974 66421
rect 45602 66220 45695 66286
rect 45602 66204 45679 66220
tri 45679 66204 45695 66220 nw
rect 45731 66187 45845 66345
rect 45881 66220 45974 66286
tri 45881 66204 45897 66220 ne
rect 45897 66204 45974 66220
rect 45714 66105 45862 66187
rect 45602 66072 45679 66088
tri 45679 66072 45695 66088 sw
rect 45602 66006 45695 66072
rect 45602 65904 45695 65970
rect 45602 65888 45679 65904
tri 45679 65888 45695 65904 nw
rect 45731 65871 45845 66105
tri 45881 66072 45897 66088 se
rect 45897 66072 45974 66088
rect 45881 66006 45974 66072
rect 45881 65904 45974 65970
tri 45881 65888 45897 65904 ne
rect 45897 65888 45974 65904
rect 45714 65789 45862 65871
rect 45602 65756 45679 65772
tri 45679 65756 45695 65772 sw
rect 45602 65690 45695 65756
rect 45731 65631 45845 65789
tri 45881 65756 45897 65772 se
rect 45897 65756 45974 65772
rect 45881 65690 45974 65756
rect 45602 65555 45974 65631
rect 45602 65430 45695 65496
rect 45602 65414 45679 65430
tri 45679 65414 45695 65430 nw
rect 45731 65397 45845 65555
rect 45881 65430 45974 65496
tri 45881 65414 45897 65430 ne
rect 45897 65414 45974 65430
rect 45714 65315 45862 65397
rect 45602 65282 45679 65298
tri 45679 65282 45695 65298 sw
rect 45602 65216 45695 65282
rect 45602 65114 45695 65180
rect 45602 65098 45679 65114
tri 45679 65098 45695 65114 nw
rect 45731 65081 45845 65315
tri 45881 65282 45897 65298 se
rect 45897 65282 45974 65298
rect 45881 65216 45974 65282
rect 45881 65114 45974 65180
tri 45881 65098 45897 65114 ne
rect 45897 65098 45974 65114
rect 45714 64999 45862 65081
rect 45602 64966 45679 64982
tri 45679 64966 45695 64982 sw
rect 45602 64900 45695 64966
rect 45731 64841 45845 64999
tri 45881 64966 45897 64982 se
rect 45897 64966 45974 64982
rect 45881 64900 45974 64966
rect 45602 64765 45974 64841
rect 45602 64640 45695 64706
rect 45602 64624 45679 64640
tri 45679 64624 45695 64640 nw
rect 45731 64607 45845 64765
rect 45881 64640 45974 64706
tri 45881 64624 45897 64640 ne
rect 45897 64624 45974 64640
rect 45714 64525 45862 64607
rect 45602 64492 45679 64508
tri 45679 64492 45695 64508 sw
rect 45602 64426 45695 64492
rect 45602 64324 45695 64390
rect 45602 64308 45679 64324
tri 45679 64308 45695 64324 nw
rect 45731 64291 45845 64525
tri 45881 64492 45897 64508 se
rect 45897 64492 45974 64508
rect 45881 64426 45974 64492
rect 45881 64324 45974 64390
tri 45881 64308 45897 64324 ne
rect 45897 64308 45974 64324
rect 45714 64209 45862 64291
rect 45602 64176 45679 64192
tri 45679 64176 45695 64192 sw
rect 45602 64110 45695 64176
rect 45731 64051 45845 64209
tri 45881 64176 45897 64192 se
rect 45897 64176 45974 64192
rect 45881 64110 45974 64176
rect 45602 63975 45974 64051
rect 45602 63850 45695 63916
rect 45602 63834 45679 63850
tri 45679 63834 45695 63850 nw
rect 45731 63817 45845 63975
rect 45881 63850 45974 63916
tri 45881 63834 45897 63850 ne
rect 45897 63834 45974 63850
rect 45714 63735 45862 63817
rect 45602 63702 45679 63718
tri 45679 63702 45695 63718 sw
rect 45602 63636 45695 63702
rect 45602 63534 45695 63600
rect 45602 63518 45679 63534
tri 45679 63518 45695 63534 nw
rect 45731 63501 45845 63735
tri 45881 63702 45897 63718 se
rect 45897 63702 45974 63718
rect 45881 63636 45974 63702
rect 45881 63534 45974 63600
tri 45881 63518 45897 63534 ne
rect 45897 63518 45974 63534
rect 45714 63419 45862 63501
rect 45602 63386 45679 63402
tri 45679 63386 45695 63402 sw
rect 45602 63320 45695 63386
rect 45731 63261 45845 63419
tri 45881 63386 45897 63402 se
rect 45897 63386 45974 63402
rect 45881 63320 45974 63386
rect 45602 63185 45974 63261
rect 45602 63060 45695 63126
rect 45602 63044 45679 63060
tri 45679 63044 45695 63060 nw
rect 45731 63027 45845 63185
rect 45881 63060 45974 63126
tri 45881 63044 45897 63060 ne
rect 45897 63044 45974 63060
rect 45714 62945 45862 63027
rect 45602 62912 45679 62928
tri 45679 62912 45695 62928 sw
rect 45602 62846 45695 62912
rect 45602 62744 45695 62810
rect 45602 62728 45679 62744
tri 45679 62728 45695 62744 nw
rect 45731 62711 45845 62945
tri 45881 62912 45897 62928 se
rect 45897 62912 45974 62928
rect 45881 62846 45974 62912
rect 45881 62744 45974 62810
tri 45881 62728 45897 62744 ne
rect 45897 62728 45974 62744
rect 45714 62629 45862 62711
rect 45602 62596 45679 62612
tri 45679 62596 45695 62612 sw
rect 45602 62530 45695 62596
rect 45731 62471 45845 62629
tri 45881 62596 45897 62612 se
rect 45897 62596 45974 62612
rect 45881 62530 45974 62596
rect 45602 62395 45974 62471
rect 45602 62270 45695 62336
rect 45602 62254 45679 62270
tri 45679 62254 45695 62270 nw
rect 45731 62237 45845 62395
rect 45881 62270 45974 62336
tri 45881 62254 45897 62270 ne
rect 45897 62254 45974 62270
rect 45714 62155 45862 62237
rect 45602 62122 45679 62138
tri 45679 62122 45695 62138 sw
rect 45602 62056 45695 62122
rect 45602 61954 45695 62020
rect 45602 61938 45679 61954
tri 45679 61938 45695 61954 nw
rect 45731 61921 45845 62155
tri 45881 62122 45897 62138 se
rect 45897 62122 45974 62138
rect 45881 62056 45974 62122
rect 45881 61954 45974 62020
tri 45881 61938 45897 61954 ne
rect 45897 61938 45974 61954
rect 45714 61839 45862 61921
rect 45602 61806 45679 61822
tri 45679 61806 45695 61822 sw
rect 45602 61740 45695 61806
rect 45731 61681 45845 61839
tri 45881 61806 45897 61822 se
rect 45897 61806 45974 61822
rect 45881 61740 45974 61806
rect 45602 61605 45974 61681
rect 45602 61480 45695 61546
rect 45602 61464 45679 61480
tri 45679 61464 45695 61480 nw
rect 45731 61447 45845 61605
rect 45881 61480 45974 61546
tri 45881 61464 45897 61480 ne
rect 45897 61464 45974 61480
rect 45714 61365 45862 61447
rect 45602 61332 45679 61348
tri 45679 61332 45695 61348 sw
rect 45602 61266 45695 61332
rect 45602 61164 45695 61230
rect 45602 61148 45679 61164
tri 45679 61148 45695 61164 nw
rect 45731 61131 45845 61365
tri 45881 61332 45897 61348 se
rect 45897 61332 45974 61348
rect 45881 61266 45974 61332
rect 45881 61164 45974 61230
tri 45881 61148 45897 61164 ne
rect 45897 61148 45974 61164
rect 45714 61049 45862 61131
rect 45602 61016 45679 61032
tri 45679 61016 45695 61032 sw
rect 45602 60950 45695 61016
rect 45731 60891 45845 61049
tri 45881 61016 45897 61032 se
rect 45897 61016 45974 61032
rect 45881 60950 45974 61016
rect 45602 60815 45974 60891
rect 45602 60690 45695 60756
rect 45602 60674 45679 60690
tri 45679 60674 45695 60690 nw
rect 45731 60657 45845 60815
rect 45881 60690 45974 60756
tri 45881 60674 45897 60690 ne
rect 45897 60674 45974 60690
rect 45714 60575 45862 60657
rect 45602 60542 45679 60558
tri 45679 60542 45695 60558 sw
rect 45602 60476 45695 60542
rect 45602 60374 45695 60440
rect 45602 60358 45679 60374
tri 45679 60358 45695 60374 nw
rect 45731 60341 45845 60575
tri 45881 60542 45897 60558 se
rect 45897 60542 45974 60558
rect 45881 60476 45974 60542
rect 45881 60374 45974 60440
tri 45881 60358 45897 60374 ne
rect 45897 60358 45974 60374
rect 45714 60259 45862 60341
rect 45602 60226 45679 60242
tri 45679 60226 45695 60242 sw
rect 45602 60160 45695 60226
rect 45731 60101 45845 60259
tri 45881 60226 45897 60242 se
rect 45897 60226 45974 60242
rect 45881 60160 45974 60226
rect 45602 60025 45974 60101
rect 45602 59900 45695 59966
rect 45602 59884 45679 59900
tri 45679 59884 45695 59900 nw
rect 45731 59867 45845 60025
rect 45881 59900 45974 59966
tri 45881 59884 45897 59900 ne
rect 45897 59884 45974 59900
rect 45714 59785 45862 59867
rect 45602 59752 45679 59768
tri 45679 59752 45695 59768 sw
rect 45602 59686 45695 59752
rect 45602 59584 45695 59650
rect 45602 59568 45679 59584
tri 45679 59568 45695 59584 nw
rect 45731 59551 45845 59785
tri 45881 59752 45897 59768 se
rect 45897 59752 45974 59768
rect 45881 59686 45974 59752
rect 45881 59584 45974 59650
tri 45881 59568 45897 59584 ne
rect 45897 59568 45974 59584
rect 45714 59469 45862 59551
rect 45602 59436 45679 59452
tri 45679 59436 45695 59452 sw
rect 45602 59370 45695 59436
rect 45731 59311 45845 59469
tri 45881 59436 45897 59452 se
rect 45897 59436 45974 59452
rect 45881 59370 45974 59436
rect 45602 59235 45974 59311
rect 45602 59110 45695 59176
rect 45602 59094 45679 59110
tri 45679 59094 45695 59110 nw
rect 45731 59077 45845 59235
rect 45881 59110 45974 59176
tri 45881 59094 45897 59110 ne
rect 45897 59094 45974 59110
rect 45714 58995 45862 59077
rect 45602 58962 45679 58978
tri 45679 58962 45695 58978 sw
rect 45602 58896 45695 58962
rect 45602 58794 45695 58860
rect 45602 58778 45679 58794
tri 45679 58778 45695 58794 nw
rect 45731 58761 45845 58995
tri 45881 58962 45897 58978 se
rect 45897 58962 45974 58978
rect 45881 58896 45974 58962
rect 45881 58794 45974 58860
tri 45881 58778 45897 58794 ne
rect 45897 58778 45974 58794
rect 45714 58679 45862 58761
rect 45602 58646 45679 58662
tri 45679 58646 45695 58662 sw
rect 45602 58580 45695 58646
rect 45731 58521 45845 58679
tri 45881 58646 45897 58662 se
rect 45897 58646 45974 58662
rect 45881 58580 45974 58646
rect 45602 58445 45974 58521
rect 45602 58320 45695 58386
rect 45602 58304 45679 58320
tri 45679 58304 45695 58320 nw
rect 45731 58287 45845 58445
rect 45881 58320 45974 58386
tri 45881 58304 45897 58320 ne
rect 45897 58304 45974 58320
rect 45714 58205 45862 58287
rect 45602 58172 45679 58188
tri 45679 58172 45695 58188 sw
rect 45602 58106 45695 58172
rect 45602 58004 45695 58070
rect 45602 57988 45679 58004
tri 45679 57988 45695 58004 nw
rect 45731 57971 45845 58205
tri 45881 58172 45897 58188 se
rect 45897 58172 45974 58188
rect 45881 58106 45974 58172
rect 45881 58004 45974 58070
tri 45881 57988 45897 58004 ne
rect 45897 57988 45974 58004
rect 45714 57889 45862 57971
rect 45602 57856 45679 57872
tri 45679 57856 45695 57872 sw
rect 45602 57790 45695 57856
rect 45731 57731 45845 57889
tri 45881 57856 45897 57872 se
rect 45897 57856 45974 57872
rect 45881 57790 45974 57856
rect 45602 57655 45974 57731
rect 45602 57530 45695 57596
rect 45602 57514 45679 57530
tri 45679 57514 45695 57530 nw
rect 45731 57497 45845 57655
rect 45881 57530 45974 57596
tri 45881 57514 45897 57530 ne
rect 45897 57514 45974 57530
rect 45714 57415 45862 57497
rect 45602 57382 45679 57398
tri 45679 57382 45695 57398 sw
rect 45602 57316 45695 57382
rect 45602 57214 45695 57280
rect 45602 57198 45679 57214
tri 45679 57198 45695 57214 nw
rect 45731 57181 45845 57415
tri 45881 57382 45897 57398 se
rect 45897 57382 45974 57398
rect 45881 57316 45974 57382
rect 45881 57214 45974 57280
tri 45881 57198 45897 57214 ne
rect 45897 57198 45974 57214
rect 45714 57099 45862 57181
rect 45602 57066 45679 57082
tri 45679 57066 45695 57082 sw
rect 45602 57000 45695 57066
rect 45731 56941 45845 57099
tri 45881 57066 45897 57082 se
rect 45897 57066 45974 57082
rect 45881 57000 45974 57066
rect 45602 56865 45974 56941
rect 45602 56740 45695 56806
rect 45602 56724 45679 56740
tri 45679 56724 45695 56740 nw
rect 45731 56707 45845 56865
rect 45881 56740 45974 56806
tri 45881 56724 45897 56740 ne
rect 45897 56724 45974 56740
rect 45714 56625 45862 56707
rect 45602 56592 45679 56608
tri 45679 56592 45695 56608 sw
rect 45602 56526 45695 56592
rect 45602 56424 45695 56490
rect 45602 56408 45679 56424
tri 45679 56408 45695 56424 nw
rect 45731 56391 45845 56625
tri 45881 56592 45897 56608 se
rect 45897 56592 45974 56608
rect 45881 56526 45974 56592
rect 45881 56424 45974 56490
tri 45881 56408 45897 56424 ne
rect 45897 56408 45974 56424
rect 45714 56309 45862 56391
rect 45602 56276 45679 56292
tri 45679 56276 45695 56292 sw
rect 45602 56210 45695 56276
rect 45731 56151 45845 56309
tri 45881 56276 45897 56292 se
rect 45897 56276 45974 56292
rect 45881 56210 45974 56276
rect 45602 56075 45974 56151
rect 45602 55950 45695 56016
rect 45602 55934 45679 55950
tri 45679 55934 45695 55950 nw
rect 45731 55917 45845 56075
rect 45881 55950 45974 56016
tri 45881 55934 45897 55950 ne
rect 45897 55934 45974 55950
rect 45714 55835 45862 55917
rect 45602 55802 45679 55818
tri 45679 55802 45695 55818 sw
rect 45602 55736 45695 55802
rect 45602 55634 45695 55700
rect 45602 55618 45679 55634
tri 45679 55618 45695 55634 nw
rect 45731 55601 45845 55835
tri 45881 55802 45897 55818 se
rect 45897 55802 45974 55818
rect 45881 55736 45974 55802
rect 45881 55634 45974 55700
tri 45881 55618 45897 55634 ne
rect 45897 55618 45974 55634
rect 45714 55519 45862 55601
rect 45602 55486 45679 55502
tri 45679 55486 45695 55502 sw
rect 45602 55420 45695 55486
rect 45731 55361 45845 55519
tri 45881 55486 45897 55502 se
rect 45897 55486 45974 55502
rect 45881 55420 45974 55486
rect 45602 55285 45974 55361
rect 45602 55160 45695 55226
rect 45602 55144 45679 55160
tri 45679 55144 45695 55160 nw
rect 45731 55127 45845 55285
rect 45881 55160 45974 55226
tri 45881 55144 45897 55160 ne
rect 45897 55144 45974 55160
rect 45714 55045 45862 55127
rect 45602 55012 45679 55028
tri 45679 55012 45695 55028 sw
rect 45602 54946 45695 55012
rect 45602 54844 45695 54910
rect 45602 54828 45679 54844
tri 45679 54828 45695 54844 nw
rect 45731 54811 45845 55045
tri 45881 55012 45897 55028 se
rect 45897 55012 45974 55028
rect 45881 54946 45974 55012
rect 45881 54844 45974 54910
tri 45881 54828 45897 54844 ne
rect 45897 54828 45974 54844
rect 45714 54729 45862 54811
rect 45602 54696 45679 54712
tri 45679 54696 45695 54712 sw
rect 45602 54630 45695 54696
rect 45731 54571 45845 54729
tri 45881 54696 45897 54712 se
rect 45897 54696 45974 54712
rect 45881 54630 45974 54696
rect 45602 54495 45974 54571
rect 45602 54370 45695 54436
rect 45602 54354 45679 54370
tri 45679 54354 45695 54370 nw
rect 45731 54337 45845 54495
rect 45881 54370 45974 54436
tri 45881 54354 45897 54370 ne
rect 45897 54354 45974 54370
rect 45714 54255 45862 54337
rect 45602 54222 45679 54238
tri 45679 54222 45695 54238 sw
rect 45602 54156 45695 54222
rect 45602 54054 45695 54120
rect 45602 54038 45679 54054
tri 45679 54038 45695 54054 nw
rect 45731 54021 45845 54255
tri 45881 54222 45897 54238 se
rect 45897 54222 45974 54238
rect 45881 54156 45974 54222
rect 45881 54054 45974 54120
tri 45881 54038 45897 54054 ne
rect 45897 54038 45974 54054
rect 45714 53939 45862 54021
rect 45602 53906 45679 53922
tri 45679 53906 45695 53922 sw
rect 45602 53840 45695 53906
rect 45731 53781 45845 53939
tri 45881 53906 45897 53922 se
rect 45897 53906 45974 53922
rect 45881 53840 45974 53906
rect 45602 53705 45974 53781
rect 45602 53580 45695 53646
rect 45602 53564 45679 53580
tri 45679 53564 45695 53580 nw
rect 45731 53547 45845 53705
rect 45881 53580 45974 53646
tri 45881 53564 45897 53580 ne
rect 45897 53564 45974 53580
rect 45714 53465 45862 53547
rect 45602 53432 45679 53448
tri 45679 53432 45695 53448 sw
rect 45602 53366 45695 53432
rect 45602 53264 45695 53330
rect 45602 53248 45679 53264
tri 45679 53248 45695 53264 nw
rect 45731 53231 45845 53465
tri 45881 53432 45897 53448 se
rect 45897 53432 45974 53448
rect 45881 53366 45974 53432
rect 45881 53264 45974 53330
tri 45881 53248 45897 53264 ne
rect 45897 53248 45974 53264
rect 45714 53149 45862 53231
rect 45602 53116 45679 53132
tri 45679 53116 45695 53132 sw
rect 45602 53050 45695 53116
rect 45731 52991 45845 53149
tri 45881 53116 45897 53132 se
rect 45897 53116 45974 53132
rect 45881 53050 45974 53116
rect 45602 52915 45974 52991
rect 45602 52790 45695 52856
rect 45602 52774 45679 52790
tri 45679 52774 45695 52790 nw
rect 45731 52757 45845 52915
rect 45881 52790 45974 52856
tri 45881 52774 45897 52790 ne
rect 45897 52774 45974 52790
rect 45714 52675 45862 52757
rect 45602 52642 45679 52658
tri 45679 52642 45695 52658 sw
rect 45602 52576 45695 52642
rect 45602 52474 45695 52540
rect 45602 52458 45679 52474
tri 45679 52458 45695 52474 nw
rect 45731 52441 45845 52675
tri 45881 52642 45897 52658 se
rect 45897 52642 45974 52658
rect 45881 52576 45974 52642
rect 45881 52474 45974 52540
tri 45881 52458 45897 52474 ne
rect 45897 52458 45974 52474
rect 45714 52359 45862 52441
rect 45602 52326 45679 52342
tri 45679 52326 45695 52342 sw
rect 45602 52260 45695 52326
rect 45731 52201 45845 52359
tri 45881 52326 45897 52342 se
rect 45897 52326 45974 52342
rect 45881 52260 45974 52326
rect 45602 52125 45974 52201
rect 45602 52000 45695 52066
rect 45602 51984 45679 52000
tri 45679 51984 45695 52000 nw
rect 45731 51967 45845 52125
rect 45881 52000 45974 52066
tri 45881 51984 45897 52000 ne
rect 45897 51984 45974 52000
rect 45714 51885 45862 51967
rect 45602 51852 45679 51868
tri 45679 51852 45695 51868 sw
rect 45602 51786 45695 51852
rect 45602 51684 45695 51750
rect 45602 51668 45679 51684
tri 45679 51668 45695 51684 nw
rect 45731 51651 45845 51885
tri 45881 51852 45897 51868 se
rect 45897 51852 45974 51868
rect 45881 51786 45974 51852
rect 45881 51684 45974 51750
tri 45881 51668 45897 51684 ne
rect 45897 51668 45974 51684
rect 45714 51569 45862 51651
rect 45602 51536 45679 51552
tri 45679 51536 45695 51552 sw
rect 45602 51470 45695 51536
rect 45731 51411 45845 51569
tri 45881 51536 45897 51552 se
rect 45897 51536 45974 51552
rect 45881 51470 45974 51536
rect 45602 51335 45974 51411
rect 45602 51210 45695 51276
rect 45602 51194 45679 51210
tri 45679 51194 45695 51210 nw
rect 45731 51177 45845 51335
rect 45881 51210 45974 51276
tri 45881 51194 45897 51210 ne
rect 45897 51194 45974 51210
rect 45714 51095 45862 51177
rect 45602 51062 45679 51078
tri 45679 51062 45695 51078 sw
rect 45602 50996 45695 51062
rect 45602 50894 45695 50960
rect 45602 50878 45679 50894
tri 45679 50878 45695 50894 nw
rect 45731 50861 45845 51095
tri 45881 51062 45897 51078 se
rect 45897 51062 45974 51078
rect 45881 50996 45974 51062
rect 45881 50894 45974 50960
tri 45881 50878 45897 50894 ne
rect 45897 50878 45974 50894
rect 45714 50779 45862 50861
rect 45602 50746 45679 50762
tri 45679 50746 45695 50762 sw
rect 45602 50680 45695 50746
rect 45731 50621 45845 50779
tri 45881 50746 45897 50762 se
rect 45897 50746 45974 50762
rect 45881 50680 45974 50746
rect 45602 50545 45974 50621
rect 45602 50420 45695 50486
rect 45602 50404 45679 50420
tri 45679 50404 45695 50420 nw
rect 45731 50387 45845 50545
rect 45881 50420 45974 50486
tri 45881 50404 45897 50420 ne
rect 45897 50404 45974 50420
rect 45714 50305 45862 50387
rect 45602 50272 45679 50288
tri 45679 50272 45695 50288 sw
rect 45602 50206 45695 50272
rect 45602 50104 45695 50170
rect 45602 50088 45679 50104
tri 45679 50088 45695 50104 nw
rect 45731 50071 45845 50305
tri 45881 50272 45897 50288 se
rect 45897 50272 45974 50288
rect 45881 50206 45974 50272
rect 45881 50104 45974 50170
tri 45881 50088 45897 50104 ne
rect 45897 50088 45974 50104
rect 45714 49989 45862 50071
rect 45602 49956 45679 49972
tri 45679 49956 45695 49972 sw
rect 45602 49890 45695 49956
rect 45731 49831 45845 49989
tri 45881 49956 45897 49972 se
rect 45897 49956 45974 49972
rect 45881 49890 45974 49956
rect 45602 49755 45974 49831
rect 45602 49630 45695 49696
rect 45602 49614 45679 49630
tri 45679 49614 45695 49630 nw
rect 45731 49597 45845 49755
rect 45881 49630 45974 49696
tri 45881 49614 45897 49630 ne
rect 45897 49614 45974 49630
rect 45714 49515 45862 49597
rect 45602 49482 45679 49498
tri 45679 49482 45695 49498 sw
rect 45602 49416 45695 49482
rect 45602 49314 45695 49380
rect 45602 49298 45679 49314
tri 45679 49298 45695 49314 nw
rect 45731 49281 45845 49515
tri 45881 49482 45897 49498 se
rect 45897 49482 45974 49498
rect 45881 49416 45974 49482
rect 45881 49314 45974 49380
tri 45881 49298 45897 49314 ne
rect 45897 49298 45974 49314
rect 45714 49199 45862 49281
rect 45602 49166 45679 49182
tri 45679 49166 45695 49182 sw
rect 45602 49100 45695 49166
rect 45731 49041 45845 49199
tri 45881 49166 45897 49182 se
rect 45897 49166 45974 49182
rect 45881 49100 45974 49166
rect 45602 48965 45974 49041
rect 45602 48840 45695 48906
rect 45602 48824 45679 48840
tri 45679 48824 45695 48840 nw
rect 45731 48807 45845 48965
rect 45881 48840 45974 48906
tri 45881 48824 45897 48840 ne
rect 45897 48824 45974 48840
rect 45714 48725 45862 48807
rect 45602 48692 45679 48708
tri 45679 48692 45695 48708 sw
rect 45602 48626 45695 48692
rect 45602 48524 45695 48590
rect 45602 48508 45679 48524
tri 45679 48508 45695 48524 nw
rect 45731 48491 45845 48725
tri 45881 48692 45897 48708 se
rect 45897 48692 45974 48708
rect 45881 48626 45974 48692
rect 45881 48524 45974 48590
tri 45881 48508 45897 48524 ne
rect 45897 48508 45974 48524
rect 45714 48409 45862 48491
rect 45602 48376 45679 48392
tri 45679 48376 45695 48392 sw
rect 45602 48310 45695 48376
rect 45731 48251 45845 48409
tri 45881 48376 45897 48392 se
rect 45897 48376 45974 48392
rect 45881 48310 45974 48376
rect 45602 48175 45974 48251
rect 45602 48050 45695 48116
rect 45602 48034 45679 48050
tri 45679 48034 45695 48050 nw
rect 45731 48017 45845 48175
rect 45881 48050 45974 48116
tri 45881 48034 45897 48050 ne
rect 45897 48034 45974 48050
rect 45714 47935 45862 48017
rect 45602 47902 45679 47918
tri 45679 47902 45695 47918 sw
rect 45602 47836 45695 47902
rect 45602 47734 45695 47800
rect 45602 47718 45679 47734
tri 45679 47718 45695 47734 nw
rect 45731 47701 45845 47935
tri 45881 47902 45897 47918 se
rect 45897 47902 45974 47918
rect 45881 47836 45974 47902
rect 45881 47734 45974 47800
tri 45881 47718 45897 47734 ne
rect 45897 47718 45974 47734
rect 45714 47619 45862 47701
rect 45602 47586 45679 47602
tri 45679 47586 45695 47602 sw
rect 45602 47520 45695 47586
rect 45731 47461 45845 47619
tri 45881 47586 45897 47602 se
rect 45897 47586 45974 47602
rect 45881 47520 45974 47586
rect 45602 47385 45974 47461
rect 45602 47260 45695 47326
rect 45602 47244 45679 47260
tri 45679 47244 45695 47260 nw
rect 45731 47227 45845 47385
rect 45881 47260 45974 47326
tri 45881 47244 45897 47260 ne
rect 45897 47244 45974 47260
rect 45714 47145 45862 47227
rect 45602 47112 45679 47128
tri 45679 47112 45695 47128 sw
rect 45602 47046 45695 47112
rect 45602 46944 45695 47010
rect 45602 46928 45679 46944
tri 45679 46928 45695 46944 nw
rect 45731 46911 45845 47145
tri 45881 47112 45897 47128 se
rect 45897 47112 45974 47128
rect 45881 47046 45974 47112
rect 45881 46944 45974 47010
tri 45881 46928 45897 46944 ne
rect 45897 46928 45974 46944
rect 45714 46829 45862 46911
rect 45602 46796 45679 46812
tri 45679 46796 45695 46812 sw
rect 45602 46730 45695 46796
rect 45731 46671 45845 46829
tri 45881 46796 45897 46812 se
rect 45897 46796 45974 46812
rect 45881 46730 45974 46796
rect 45602 46595 45974 46671
rect 45602 46470 45695 46536
rect 45602 46454 45679 46470
tri 45679 46454 45695 46470 nw
rect 45731 46437 45845 46595
rect 45881 46470 45974 46536
tri 45881 46454 45897 46470 ne
rect 45897 46454 45974 46470
rect 45714 46355 45862 46437
rect 45602 46322 45679 46338
tri 45679 46322 45695 46338 sw
rect 45602 46256 45695 46322
rect 45602 46154 45695 46220
rect 45602 46138 45679 46154
tri 45679 46138 45695 46154 nw
rect 45731 46121 45845 46355
tri 45881 46322 45897 46338 se
rect 45897 46322 45974 46338
rect 45881 46256 45974 46322
rect 45881 46154 45974 46220
tri 45881 46138 45897 46154 ne
rect 45897 46138 45974 46154
rect 45714 46039 45862 46121
rect 45602 46006 45679 46022
tri 45679 46006 45695 46022 sw
rect 45602 45940 45695 46006
rect 45731 45881 45845 46039
tri 45881 46006 45897 46022 se
rect 45897 46006 45974 46022
rect 45881 45940 45974 46006
rect 45602 45805 45974 45881
rect 45602 45680 45695 45746
rect 45602 45664 45679 45680
tri 45679 45664 45695 45680 nw
rect 45731 45647 45845 45805
rect 45881 45680 45974 45746
tri 45881 45664 45897 45680 ne
rect 45897 45664 45974 45680
rect 45714 45565 45862 45647
rect 45602 45532 45679 45548
tri 45679 45532 45695 45548 sw
rect 45602 45466 45695 45532
rect 45602 45364 45695 45430
rect 45602 45348 45679 45364
tri 45679 45348 45695 45364 nw
rect 45731 45331 45845 45565
tri 45881 45532 45897 45548 se
rect 45897 45532 45974 45548
rect 45881 45466 45974 45532
rect 45881 45364 45974 45430
tri 45881 45348 45897 45364 ne
rect 45897 45348 45974 45364
rect 45714 45249 45862 45331
rect 45602 45216 45679 45232
tri 45679 45216 45695 45232 sw
rect 45602 45150 45695 45216
rect 45731 45091 45845 45249
tri 45881 45216 45897 45232 se
rect 45897 45216 45974 45232
rect 45881 45150 45974 45216
rect 45602 45015 45974 45091
rect 45602 44890 45695 44956
rect 45602 44874 45679 44890
tri 45679 44874 45695 44890 nw
rect 45731 44857 45845 45015
rect 45881 44890 45974 44956
tri 45881 44874 45897 44890 ne
rect 45897 44874 45974 44890
rect 45714 44775 45862 44857
rect 45602 44742 45679 44758
tri 45679 44742 45695 44758 sw
rect 45602 44676 45695 44742
rect 45602 44574 45695 44640
rect 45602 44558 45679 44574
tri 45679 44558 45695 44574 nw
rect 45731 44541 45845 44775
tri 45881 44742 45897 44758 se
rect 45897 44742 45974 44758
rect 45881 44676 45974 44742
rect 45881 44574 45974 44640
tri 45881 44558 45897 44574 ne
rect 45897 44558 45974 44574
rect 45714 44459 45862 44541
rect 45602 44426 45679 44442
tri 45679 44426 45695 44442 sw
rect 45602 44360 45695 44426
rect 45731 44301 45845 44459
tri 45881 44426 45897 44442 se
rect 45897 44426 45974 44442
rect 45881 44360 45974 44426
rect 45602 44225 45974 44301
rect 45602 44100 45695 44166
rect 45602 44084 45679 44100
tri 45679 44084 45695 44100 nw
rect 45731 44067 45845 44225
rect 45881 44100 45974 44166
tri 45881 44084 45897 44100 ne
rect 45897 44084 45974 44100
rect 45714 43985 45862 44067
rect 45602 43952 45679 43968
tri 45679 43952 45695 43968 sw
rect 45602 43886 45695 43952
rect 45602 43784 45695 43850
rect 45602 43768 45679 43784
tri 45679 43768 45695 43784 nw
rect 45731 43751 45845 43985
tri 45881 43952 45897 43968 se
rect 45897 43952 45974 43968
rect 45881 43886 45974 43952
rect 45881 43784 45974 43850
tri 45881 43768 45897 43784 ne
rect 45897 43768 45974 43784
rect 45714 43669 45862 43751
rect 45602 43636 45679 43652
tri 45679 43636 45695 43652 sw
rect 45602 43570 45695 43636
rect 45731 43511 45845 43669
tri 45881 43636 45897 43652 se
rect 45897 43636 45974 43652
rect 45881 43570 45974 43636
rect 45602 43435 45974 43511
rect 45602 43310 45695 43376
rect 45602 43294 45679 43310
tri 45679 43294 45695 43310 nw
rect 45731 43277 45845 43435
rect 45881 43310 45974 43376
tri 45881 43294 45897 43310 ne
rect 45897 43294 45974 43310
rect 45714 43195 45862 43277
rect 45602 43162 45679 43178
tri 45679 43162 45695 43178 sw
rect 45602 43096 45695 43162
rect 45602 42994 45695 43060
rect 45602 42978 45679 42994
tri 45679 42978 45695 42994 nw
rect 45731 42961 45845 43195
tri 45881 43162 45897 43178 se
rect 45897 43162 45974 43178
rect 45881 43096 45974 43162
rect 45881 42994 45974 43060
tri 45881 42978 45897 42994 ne
rect 45897 42978 45974 42994
rect 45714 42879 45862 42961
rect 45602 42846 45679 42862
tri 45679 42846 45695 42862 sw
rect 45602 42780 45695 42846
rect 45731 42721 45845 42879
tri 45881 42846 45897 42862 se
rect 45897 42846 45974 42862
rect 45881 42780 45974 42846
rect 45602 42645 45974 42721
rect 45602 42520 45695 42586
rect 45602 42504 45679 42520
tri 45679 42504 45695 42520 nw
rect 45731 42487 45845 42645
rect 45881 42520 45974 42586
tri 45881 42504 45897 42520 ne
rect 45897 42504 45974 42520
rect 45714 42405 45862 42487
rect 45602 42372 45679 42388
tri 45679 42372 45695 42388 sw
rect 45602 42306 45695 42372
rect 45602 42204 45695 42270
rect 45602 42188 45679 42204
tri 45679 42188 45695 42204 nw
rect 45731 42171 45845 42405
tri 45881 42372 45897 42388 se
rect 45897 42372 45974 42388
rect 45881 42306 45974 42372
rect 45881 42204 45974 42270
tri 45881 42188 45897 42204 ne
rect 45897 42188 45974 42204
rect 45714 42089 45862 42171
rect 45602 42056 45679 42072
tri 45679 42056 45695 42072 sw
rect 45602 41990 45695 42056
rect 45731 41931 45845 42089
tri 45881 42056 45897 42072 se
rect 45897 42056 45974 42072
rect 45881 41990 45974 42056
rect 45602 41855 45974 41931
rect 45602 41730 45695 41796
rect 45602 41714 45679 41730
tri 45679 41714 45695 41730 nw
rect 45731 41697 45845 41855
rect 45881 41730 45974 41796
tri 45881 41714 45897 41730 ne
rect 45897 41714 45974 41730
rect 45714 41615 45862 41697
rect 45602 41582 45679 41598
tri 45679 41582 45695 41598 sw
rect 45602 41516 45695 41582
rect 45602 41414 45695 41480
rect 45602 41398 45679 41414
tri 45679 41398 45695 41414 nw
rect 45731 41381 45845 41615
tri 45881 41582 45897 41598 se
rect 45897 41582 45974 41598
rect 45881 41516 45974 41582
rect 45881 41414 45974 41480
tri 45881 41398 45897 41414 ne
rect 45897 41398 45974 41414
rect 45714 41299 45862 41381
rect 45602 41266 45679 41282
tri 45679 41266 45695 41282 sw
rect 45602 41200 45695 41266
rect 45731 41141 45845 41299
tri 45881 41266 45897 41282 se
rect 45897 41266 45974 41282
rect 45881 41200 45974 41266
rect 45602 41065 45974 41141
rect 45602 40940 45695 41006
rect 45602 40924 45679 40940
tri 45679 40924 45695 40940 nw
rect 45731 40907 45845 41065
rect 45881 40940 45974 41006
tri 45881 40924 45897 40940 ne
rect 45897 40924 45974 40940
rect 45714 40825 45862 40907
rect 45602 40792 45679 40808
tri 45679 40792 45695 40808 sw
rect 45602 40726 45695 40792
rect 45602 40624 45695 40690
rect 45602 40608 45679 40624
tri 45679 40608 45695 40624 nw
rect 45731 40591 45845 40825
tri 45881 40792 45897 40808 se
rect 45897 40792 45974 40808
rect 45881 40726 45974 40792
rect 45881 40624 45974 40690
tri 45881 40608 45897 40624 ne
rect 45897 40608 45974 40624
rect 45714 40509 45862 40591
rect 45602 40476 45679 40492
tri 45679 40476 45695 40492 sw
rect 45602 40410 45695 40476
rect 45731 40351 45845 40509
tri 45881 40476 45897 40492 se
rect 45897 40476 45974 40492
rect 45881 40410 45974 40476
rect 45602 40275 45974 40351
rect 45602 40150 45695 40216
rect 45602 40134 45679 40150
tri 45679 40134 45695 40150 nw
rect 45731 40117 45845 40275
rect 45881 40150 45974 40216
tri 45881 40134 45897 40150 ne
rect 45897 40134 45974 40150
rect 45714 40035 45862 40117
rect 45602 40002 45679 40018
tri 45679 40002 45695 40018 sw
rect 45602 39936 45695 40002
rect 45602 39834 45695 39900
rect 45602 39818 45679 39834
tri 45679 39818 45695 39834 nw
rect 45731 39801 45845 40035
tri 45881 40002 45897 40018 se
rect 45897 40002 45974 40018
rect 45881 39936 45974 40002
rect 45881 39834 45974 39900
tri 45881 39818 45897 39834 ne
rect 45897 39818 45974 39834
rect 45714 39719 45862 39801
rect 45602 39686 45679 39702
tri 45679 39686 45695 39702 sw
rect 45602 39620 45695 39686
rect 45731 39561 45845 39719
tri 45881 39686 45897 39702 se
rect 45897 39686 45974 39702
rect 45881 39620 45974 39686
rect 45602 39485 45974 39561
rect 45602 39360 45695 39426
rect 45602 39344 45679 39360
tri 45679 39344 45695 39360 nw
rect 45731 39327 45845 39485
rect 45881 39360 45974 39426
tri 45881 39344 45897 39360 ne
rect 45897 39344 45974 39360
rect 45714 39245 45862 39327
rect 45602 39212 45679 39228
tri 45679 39212 45695 39228 sw
rect 45602 39146 45695 39212
rect 45602 39044 45695 39110
rect 45602 39028 45679 39044
tri 45679 39028 45695 39044 nw
rect 45731 39011 45845 39245
tri 45881 39212 45897 39228 se
rect 45897 39212 45974 39228
rect 45881 39146 45974 39212
rect 45881 39044 45974 39110
tri 45881 39028 45897 39044 ne
rect 45897 39028 45974 39044
rect 45714 38929 45862 39011
rect 45602 38896 45679 38912
tri 45679 38896 45695 38912 sw
rect 45602 38830 45695 38896
rect 45731 38771 45845 38929
tri 45881 38896 45897 38912 se
rect 45897 38896 45974 38912
rect 45881 38830 45974 38896
rect 45602 38695 45974 38771
rect 45602 38570 45695 38636
rect 45602 38554 45679 38570
tri 45679 38554 45695 38570 nw
rect 45731 38537 45845 38695
rect 45881 38570 45974 38636
tri 45881 38554 45897 38570 ne
rect 45897 38554 45974 38570
rect 45714 38455 45862 38537
rect 45602 38422 45679 38438
tri 45679 38422 45695 38438 sw
rect 45602 38356 45695 38422
rect 45602 38254 45695 38320
rect 45602 38238 45679 38254
tri 45679 38238 45695 38254 nw
rect 45731 38221 45845 38455
tri 45881 38422 45897 38438 se
rect 45897 38422 45974 38438
rect 45881 38356 45974 38422
rect 45881 38254 45974 38320
tri 45881 38238 45897 38254 ne
rect 45897 38238 45974 38254
rect 45714 38139 45862 38221
rect 45602 38106 45679 38122
tri 45679 38106 45695 38122 sw
rect 45602 38040 45695 38106
rect 45731 37981 45845 38139
tri 45881 38106 45897 38122 se
rect 45897 38106 45974 38122
rect 45881 38040 45974 38106
rect 45602 37905 45974 37981
rect 45602 37780 45695 37846
rect 45602 37764 45679 37780
tri 45679 37764 45695 37780 nw
rect 45731 37747 45845 37905
rect 45881 37780 45974 37846
tri 45881 37764 45897 37780 ne
rect 45897 37764 45974 37780
rect 45714 37665 45862 37747
rect 45602 37632 45679 37648
tri 45679 37632 45695 37648 sw
rect 45602 37566 45695 37632
rect 45602 37464 45695 37530
rect 45602 37448 45679 37464
tri 45679 37448 45695 37464 nw
rect 45731 37431 45845 37665
tri 45881 37632 45897 37648 se
rect 45897 37632 45974 37648
rect 45881 37566 45974 37632
rect 45881 37464 45974 37530
tri 45881 37448 45897 37464 ne
rect 45897 37448 45974 37464
rect 45714 37349 45862 37431
rect 45602 37316 45679 37332
tri 45679 37316 45695 37332 sw
rect 45602 37250 45695 37316
rect 45731 37191 45845 37349
tri 45881 37316 45897 37332 se
rect 45897 37316 45974 37332
rect 45881 37250 45974 37316
rect 45602 37115 45974 37191
rect 45602 36990 45695 37056
rect 45602 36974 45679 36990
tri 45679 36974 45695 36990 nw
rect 45731 36957 45845 37115
rect 45881 36990 45974 37056
tri 45881 36974 45897 36990 ne
rect 45897 36974 45974 36990
rect 45714 36875 45862 36957
rect 45602 36842 45679 36858
tri 45679 36842 45695 36858 sw
rect 45602 36776 45695 36842
rect 45602 36674 45695 36740
rect 45602 36658 45679 36674
tri 45679 36658 45695 36674 nw
rect 45731 36641 45845 36875
tri 45881 36842 45897 36858 se
rect 45897 36842 45974 36858
rect 45881 36776 45974 36842
rect 45881 36674 45974 36740
tri 45881 36658 45897 36674 ne
rect 45897 36658 45974 36674
rect 45714 36559 45862 36641
rect 45602 36526 45679 36542
tri 45679 36526 45695 36542 sw
rect 45602 36460 45695 36526
rect 45731 36401 45845 36559
tri 45881 36526 45897 36542 se
rect 45897 36526 45974 36542
rect 45881 36460 45974 36526
rect 45602 36325 45974 36401
rect 45602 36200 45695 36266
rect 45602 36184 45679 36200
tri 45679 36184 45695 36200 nw
rect 45731 36167 45845 36325
rect 45881 36200 45974 36266
tri 45881 36184 45897 36200 ne
rect 45897 36184 45974 36200
rect 45714 36085 45862 36167
rect 45602 36052 45679 36068
tri 45679 36052 45695 36068 sw
rect 45602 35986 45695 36052
rect 45602 35884 45695 35950
rect 45602 35868 45679 35884
tri 45679 35868 45695 35884 nw
rect 45731 35851 45845 36085
tri 45881 36052 45897 36068 se
rect 45897 36052 45974 36068
rect 45881 35986 45974 36052
rect 45881 35884 45974 35950
tri 45881 35868 45897 35884 ne
rect 45897 35868 45974 35884
rect 45714 35769 45862 35851
rect 45602 35736 45679 35752
tri 45679 35736 45695 35752 sw
rect 45602 35670 45695 35736
rect 45731 35611 45845 35769
tri 45881 35736 45897 35752 se
rect 45897 35736 45974 35752
rect 45881 35670 45974 35736
rect 45602 35535 45974 35611
rect 45602 35410 45695 35476
rect 45602 35394 45679 35410
tri 45679 35394 45695 35410 nw
rect 45731 35377 45845 35535
rect 45881 35410 45974 35476
tri 45881 35394 45897 35410 ne
rect 45897 35394 45974 35410
rect 45714 35295 45862 35377
rect 45602 35262 45679 35278
tri 45679 35262 45695 35278 sw
rect 45602 35196 45695 35262
rect 45602 35094 45695 35160
rect 45602 35078 45679 35094
tri 45679 35078 45695 35094 nw
rect 45731 35061 45845 35295
tri 45881 35262 45897 35278 se
rect 45897 35262 45974 35278
rect 45881 35196 45974 35262
rect 45881 35094 45974 35160
tri 45881 35078 45897 35094 ne
rect 45897 35078 45974 35094
rect 45714 34979 45862 35061
rect 45602 34946 45679 34962
tri 45679 34946 45695 34962 sw
rect 45602 34880 45695 34946
rect 45731 34821 45845 34979
tri 45881 34946 45897 34962 se
rect 45897 34946 45974 34962
rect 45881 34880 45974 34946
rect 45602 34745 45974 34821
rect 45602 34620 45695 34686
rect 45602 34604 45679 34620
tri 45679 34604 45695 34620 nw
rect 45731 34587 45845 34745
rect 45881 34620 45974 34686
tri 45881 34604 45897 34620 ne
rect 45897 34604 45974 34620
rect 45714 34505 45862 34587
rect 45602 34472 45679 34488
tri 45679 34472 45695 34488 sw
rect 45602 34406 45695 34472
rect 45602 34304 45695 34370
rect 45602 34288 45679 34304
tri 45679 34288 45695 34304 nw
rect 45731 34271 45845 34505
tri 45881 34472 45897 34488 se
rect 45897 34472 45974 34488
rect 45881 34406 45974 34472
rect 45881 34304 45974 34370
tri 45881 34288 45897 34304 ne
rect 45897 34288 45974 34304
rect 45714 34189 45862 34271
rect 45602 34156 45679 34172
tri 45679 34156 45695 34172 sw
rect 45602 34090 45695 34156
rect 45731 34031 45845 34189
tri 45881 34156 45897 34172 se
rect 45897 34156 45974 34172
rect 45881 34090 45974 34156
rect 45602 33955 45974 34031
rect 45602 33830 45695 33896
rect 45602 33814 45679 33830
tri 45679 33814 45695 33830 nw
rect 45731 33797 45845 33955
rect 45881 33830 45974 33896
tri 45881 33814 45897 33830 ne
rect 45897 33814 45974 33830
rect 45714 33715 45862 33797
rect 45602 33682 45679 33698
tri 45679 33682 45695 33698 sw
rect 45602 33616 45695 33682
rect 45602 33514 45695 33580
rect 45602 33498 45679 33514
tri 45679 33498 45695 33514 nw
rect 45731 33481 45845 33715
tri 45881 33682 45897 33698 se
rect 45897 33682 45974 33698
rect 45881 33616 45974 33682
rect 45881 33514 45974 33580
tri 45881 33498 45897 33514 ne
rect 45897 33498 45974 33514
rect 45714 33399 45862 33481
rect 45602 33366 45679 33382
tri 45679 33366 45695 33382 sw
rect 45602 33300 45695 33366
rect 45731 33241 45845 33399
tri 45881 33366 45897 33382 se
rect 45897 33366 45974 33382
rect 45881 33300 45974 33366
rect 45602 33165 45974 33241
rect 45602 33040 45695 33106
rect 45602 33024 45679 33040
tri 45679 33024 45695 33040 nw
rect 45731 33007 45845 33165
rect 45881 33040 45974 33106
tri 45881 33024 45897 33040 ne
rect 45897 33024 45974 33040
rect 45714 32925 45862 33007
rect 45602 32892 45679 32908
tri 45679 32892 45695 32908 sw
rect 45602 32826 45695 32892
rect 45602 32724 45695 32790
rect 45602 32708 45679 32724
tri 45679 32708 45695 32724 nw
rect 45731 32691 45845 32925
tri 45881 32892 45897 32908 se
rect 45897 32892 45974 32908
rect 45881 32826 45974 32892
rect 45881 32724 45974 32790
tri 45881 32708 45897 32724 ne
rect 45897 32708 45974 32724
rect 45714 32609 45862 32691
rect 45602 32576 45679 32592
tri 45679 32576 45695 32592 sw
rect 45602 32510 45695 32576
rect 45731 32451 45845 32609
tri 45881 32576 45897 32592 se
rect 45897 32576 45974 32592
rect 45881 32510 45974 32576
rect 45602 32375 45974 32451
rect 45602 32250 45695 32316
rect 45602 32234 45679 32250
tri 45679 32234 45695 32250 nw
rect 45731 32217 45845 32375
rect 45881 32250 45974 32316
tri 45881 32234 45897 32250 ne
rect 45897 32234 45974 32250
rect 45714 32135 45862 32217
rect 45602 32102 45679 32118
tri 45679 32102 45695 32118 sw
rect 45602 32036 45695 32102
rect 45602 31934 45695 32000
rect 45602 31918 45679 31934
tri 45679 31918 45695 31934 nw
rect 45731 31901 45845 32135
tri 45881 32102 45897 32118 se
rect 45897 32102 45974 32118
rect 45881 32036 45974 32102
rect 45881 31934 45974 32000
tri 45881 31918 45897 31934 ne
rect 45897 31918 45974 31934
rect 45714 31819 45862 31901
rect 45602 31786 45679 31802
tri 45679 31786 45695 31802 sw
rect 45602 31720 45695 31786
rect 45731 31661 45845 31819
tri 45881 31786 45897 31802 se
rect 45897 31786 45974 31802
rect 45881 31720 45974 31786
rect 45602 31585 45974 31661
rect 45602 31460 45695 31526
rect 45602 31444 45679 31460
tri 45679 31444 45695 31460 nw
rect 45731 31427 45845 31585
rect 45881 31460 45974 31526
tri 45881 31444 45897 31460 ne
rect 45897 31444 45974 31460
rect 45714 31345 45862 31427
rect 45602 31312 45679 31328
tri 45679 31312 45695 31328 sw
rect 45602 31246 45695 31312
rect 45602 31144 45695 31210
rect 45602 31128 45679 31144
tri 45679 31128 45695 31144 nw
rect 45731 31111 45845 31345
tri 45881 31312 45897 31328 se
rect 45897 31312 45974 31328
rect 45881 31246 45974 31312
rect 45881 31144 45974 31210
tri 45881 31128 45897 31144 ne
rect 45897 31128 45974 31144
rect 45714 31029 45862 31111
rect 45602 30996 45679 31012
tri 45679 30996 45695 31012 sw
rect 45602 30930 45695 30996
rect 45731 30871 45845 31029
tri 45881 30996 45897 31012 se
rect 45897 30996 45974 31012
rect 45881 30930 45974 30996
rect 45602 30795 45974 30871
rect 45602 30670 45695 30736
rect 45602 30654 45679 30670
tri 45679 30654 45695 30670 nw
rect 45731 30637 45845 30795
rect 45881 30670 45974 30736
tri 45881 30654 45897 30670 ne
rect 45897 30654 45974 30670
rect 45714 30555 45862 30637
rect 45602 30522 45679 30538
tri 45679 30522 45695 30538 sw
rect 45602 30456 45695 30522
rect 45602 30354 45695 30420
rect 45602 30338 45679 30354
tri 45679 30338 45695 30354 nw
rect 45731 30321 45845 30555
tri 45881 30522 45897 30538 se
rect 45897 30522 45974 30538
rect 45881 30456 45974 30522
rect 45881 30354 45974 30420
tri 45881 30338 45897 30354 ne
rect 45897 30338 45974 30354
rect 45714 30239 45862 30321
rect 45602 30206 45679 30222
tri 45679 30206 45695 30222 sw
rect 45602 30140 45695 30206
rect 45731 30081 45845 30239
tri 45881 30206 45897 30222 se
rect 45897 30206 45974 30222
rect 45881 30140 45974 30206
rect 45602 30005 45974 30081
rect 45602 29880 45695 29946
rect 45602 29864 45679 29880
tri 45679 29864 45695 29880 nw
rect 45731 29847 45845 30005
rect 45881 29880 45974 29946
tri 45881 29864 45897 29880 ne
rect 45897 29864 45974 29880
rect 45714 29765 45862 29847
rect 45602 29732 45679 29748
tri 45679 29732 45695 29748 sw
rect 45602 29666 45695 29732
rect 45602 29564 45695 29630
rect 45602 29548 45679 29564
tri 45679 29548 45695 29564 nw
rect 45731 29531 45845 29765
tri 45881 29732 45897 29748 se
rect 45897 29732 45974 29748
rect 45881 29666 45974 29732
rect 45881 29564 45974 29630
tri 45881 29548 45897 29564 ne
rect 45897 29548 45974 29564
rect 45714 29449 45862 29531
rect 45602 29416 45679 29432
tri 45679 29416 45695 29432 sw
rect 45602 29350 45695 29416
rect 45731 29291 45845 29449
tri 45881 29416 45897 29432 se
rect 45897 29416 45974 29432
rect 45881 29350 45974 29416
rect 45602 29215 45974 29291
rect 45602 29090 45695 29156
rect 45602 29074 45679 29090
tri 45679 29074 45695 29090 nw
rect 45731 29057 45845 29215
rect 45881 29090 45974 29156
tri 45881 29074 45897 29090 ne
rect 45897 29074 45974 29090
rect 45714 28975 45862 29057
rect 45602 28942 45679 28958
tri 45679 28942 45695 28958 sw
rect 45602 28876 45695 28942
rect 45731 28833 45845 28975
tri 45881 28942 45897 28958 se
rect 45897 28942 45974 28958
rect 45881 28876 45974 28942
rect 46010 28463 46046 80603
rect 46082 28463 46118 80603
rect 46154 80445 46190 80603
rect 46146 80303 46198 80445
rect 46154 28763 46190 80303
rect 46146 28621 46198 28763
rect 46154 28463 46190 28621
rect 46226 28463 46262 80603
rect 46298 28463 46334 80603
rect 46370 28833 46454 80233
rect 46490 28463 46526 80603
rect 46562 28463 46598 80603
rect 46634 80445 46670 80603
rect 46626 80303 46678 80445
rect 46634 28763 46670 80303
rect 46626 28621 46678 28763
rect 46634 28463 46670 28621
rect 46706 28463 46742 80603
rect 46778 28463 46814 80603
rect 46850 80124 46943 80190
rect 46850 80108 46927 80124
tri 46927 80108 46943 80124 nw
rect 46979 80091 47093 80233
rect 47129 80124 47222 80190
tri 47129 80108 47145 80124 ne
rect 47145 80108 47222 80124
rect 46962 80009 47110 80091
rect 46850 79976 46927 79992
tri 46927 79976 46943 79992 sw
rect 46850 79910 46943 79976
rect 46979 79851 47093 80009
tri 47129 79976 47145 79992 se
rect 47145 79976 47222 79992
rect 47129 79910 47222 79976
rect 46850 79775 47222 79851
rect 46850 79650 46943 79716
rect 46850 79634 46927 79650
tri 46927 79634 46943 79650 nw
rect 46979 79617 47093 79775
rect 47129 79650 47222 79716
tri 47129 79634 47145 79650 ne
rect 47145 79634 47222 79650
rect 46962 79535 47110 79617
rect 46850 79502 46927 79518
tri 46927 79502 46943 79518 sw
rect 46850 79436 46943 79502
rect 46850 79334 46943 79400
rect 46850 79318 46927 79334
tri 46927 79318 46943 79334 nw
rect 46979 79301 47093 79535
tri 47129 79502 47145 79518 se
rect 47145 79502 47222 79518
rect 47129 79436 47222 79502
rect 47129 79334 47222 79400
tri 47129 79318 47145 79334 ne
rect 47145 79318 47222 79334
rect 46962 79219 47110 79301
rect 46850 79186 46927 79202
tri 46927 79186 46943 79202 sw
rect 46850 79120 46943 79186
rect 46979 79061 47093 79219
tri 47129 79186 47145 79202 se
rect 47145 79186 47222 79202
rect 47129 79120 47222 79186
rect 46850 78985 47222 79061
rect 46850 78860 46943 78926
rect 46850 78844 46927 78860
tri 46927 78844 46943 78860 nw
rect 46979 78827 47093 78985
rect 47129 78860 47222 78926
tri 47129 78844 47145 78860 ne
rect 47145 78844 47222 78860
rect 46962 78745 47110 78827
rect 46850 78712 46927 78728
tri 46927 78712 46943 78728 sw
rect 46850 78646 46943 78712
rect 46850 78544 46943 78610
rect 46850 78528 46927 78544
tri 46927 78528 46943 78544 nw
rect 46979 78511 47093 78745
tri 47129 78712 47145 78728 se
rect 47145 78712 47222 78728
rect 47129 78646 47222 78712
rect 47129 78544 47222 78610
tri 47129 78528 47145 78544 ne
rect 47145 78528 47222 78544
rect 46962 78429 47110 78511
rect 46850 78396 46927 78412
tri 46927 78396 46943 78412 sw
rect 46850 78330 46943 78396
rect 46979 78271 47093 78429
tri 47129 78396 47145 78412 se
rect 47145 78396 47222 78412
rect 47129 78330 47222 78396
rect 46850 78195 47222 78271
rect 46850 78070 46943 78136
rect 46850 78054 46927 78070
tri 46927 78054 46943 78070 nw
rect 46979 78037 47093 78195
rect 47129 78070 47222 78136
tri 47129 78054 47145 78070 ne
rect 47145 78054 47222 78070
rect 46962 77955 47110 78037
rect 46850 77922 46927 77938
tri 46927 77922 46943 77938 sw
rect 46850 77856 46943 77922
rect 46850 77754 46943 77820
rect 46850 77738 46927 77754
tri 46927 77738 46943 77754 nw
rect 46979 77721 47093 77955
tri 47129 77922 47145 77938 se
rect 47145 77922 47222 77938
rect 47129 77856 47222 77922
rect 47129 77754 47222 77820
tri 47129 77738 47145 77754 ne
rect 47145 77738 47222 77754
rect 46962 77639 47110 77721
rect 46850 77606 46927 77622
tri 46927 77606 46943 77622 sw
rect 46850 77540 46943 77606
rect 46979 77481 47093 77639
tri 47129 77606 47145 77622 se
rect 47145 77606 47222 77622
rect 47129 77540 47222 77606
rect 46850 77405 47222 77481
rect 46850 77280 46943 77346
rect 46850 77264 46927 77280
tri 46927 77264 46943 77280 nw
rect 46979 77247 47093 77405
rect 47129 77280 47222 77346
tri 47129 77264 47145 77280 ne
rect 47145 77264 47222 77280
rect 46962 77165 47110 77247
rect 46850 77132 46927 77148
tri 46927 77132 46943 77148 sw
rect 46850 77066 46943 77132
rect 46850 76964 46943 77030
rect 46850 76948 46927 76964
tri 46927 76948 46943 76964 nw
rect 46979 76931 47093 77165
tri 47129 77132 47145 77148 se
rect 47145 77132 47222 77148
rect 47129 77066 47222 77132
rect 47129 76964 47222 77030
tri 47129 76948 47145 76964 ne
rect 47145 76948 47222 76964
rect 46962 76849 47110 76931
rect 46850 76816 46927 76832
tri 46927 76816 46943 76832 sw
rect 46850 76750 46943 76816
rect 46979 76691 47093 76849
tri 47129 76816 47145 76832 se
rect 47145 76816 47222 76832
rect 47129 76750 47222 76816
rect 46850 76615 47222 76691
rect 46850 76490 46943 76556
rect 46850 76474 46927 76490
tri 46927 76474 46943 76490 nw
rect 46979 76457 47093 76615
rect 47129 76490 47222 76556
tri 47129 76474 47145 76490 ne
rect 47145 76474 47222 76490
rect 46962 76375 47110 76457
rect 46850 76342 46927 76358
tri 46927 76342 46943 76358 sw
rect 46850 76276 46943 76342
rect 46850 76174 46943 76240
rect 46850 76158 46927 76174
tri 46927 76158 46943 76174 nw
rect 46979 76141 47093 76375
tri 47129 76342 47145 76358 se
rect 47145 76342 47222 76358
rect 47129 76276 47222 76342
rect 47129 76174 47222 76240
tri 47129 76158 47145 76174 ne
rect 47145 76158 47222 76174
rect 46962 76059 47110 76141
rect 46850 76026 46927 76042
tri 46927 76026 46943 76042 sw
rect 46850 75960 46943 76026
rect 46979 75901 47093 76059
tri 47129 76026 47145 76042 se
rect 47145 76026 47222 76042
rect 47129 75960 47222 76026
rect 46850 75825 47222 75901
rect 46850 75700 46943 75766
rect 46850 75684 46927 75700
tri 46927 75684 46943 75700 nw
rect 46979 75667 47093 75825
rect 47129 75700 47222 75766
tri 47129 75684 47145 75700 ne
rect 47145 75684 47222 75700
rect 46962 75585 47110 75667
rect 46850 75552 46927 75568
tri 46927 75552 46943 75568 sw
rect 46850 75486 46943 75552
rect 46850 75384 46943 75450
rect 46850 75368 46927 75384
tri 46927 75368 46943 75384 nw
rect 46979 75351 47093 75585
tri 47129 75552 47145 75568 se
rect 47145 75552 47222 75568
rect 47129 75486 47222 75552
rect 47129 75384 47222 75450
tri 47129 75368 47145 75384 ne
rect 47145 75368 47222 75384
rect 46962 75269 47110 75351
rect 46850 75236 46927 75252
tri 46927 75236 46943 75252 sw
rect 46850 75170 46943 75236
rect 46979 75111 47093 75269
tri 47129 75236 47145 75252 se
rect 47145 75236 47222 75252
rect 47129 75170 47222 75236
rect 46850 75035 47222 75111
rect 46850 74910 46943 74976
rect 46850 74894 46927 74910
tri 46927 74894 46943 74910 nw
rect 46979 74877 47093 75035
rect 47129 74910 47222 74976
tri 47129 74894 47145 74910 ne
rect 47145 74894 47222 74910
rect 46962 74795 47110 74877
rect 46850 74762 46927 74778
tri 46927 74762 46943 74778 sw
rect 46850 74696 46943 74762
rect 46850 74594 46943 74660
rect 46850 74578 46927 74594
tri 46927 74578 46943 74594 nw
rect 46979 74561 47093 74795
tri 47129 74762 47145 74778 se
rect 47145 74762 47222 74778
rect 47129 74696 47222 74762
rect 47129 74594 47222 74660
tri 47129 74578 47145 74594 ne
rect 47145 74578 47222 74594
rect 46962 74479 47110 74561
rect 46850 74446 46927 74462
tri 46927 74446 46943 74462 sw
rect 46850 74380 46943 74446
rect 46979 74321 47093 74479
tri 47129 74446 47145 74462 se
rect 47145 74446 47222 74462
rect 47129 74380 47222 74446
rect 46850 74245 47222 74321
rect 46850 74120 46943 74186
rect 46850 74104 46927 74120
tri 46927 74104 46943 74120 nw
rect 46979 74087 47093 74245
rect 47129 74120 47222 74186
tri 47129 74104 47145 74120 ne
rect 47145 74104 47222 74120
rect 46962 74005 47110 74087
rect 46850 73972 46927 73988
tri 46927 73972 46943 73988 sw
rect 46850 73906 46943 73972
rect 46850 73804 46943 73870
rect 46850 73788 46927 73804
tri 46927 73788 46943 73804 nw
rect 46979 73771 47093 74005
tri 47129 73972 47145 73988 se
rect 47145 73972 47222 73988
rect 47129 73906 47222 73972
rect 47129 73804 47222 73870
tri 47129 73788 47145 73804 ne
rect 47145 73788 47222 73804
rect 46962 73689 47110 73771
rect 46850 73656 46927 73672
tri 46927 73656 46943 73672 sw
rect 46850 73590 46943 73656
rect 46979 73531 47093 73689
tri 47129 73656 47145 73672 se
rect 47145 73656 47222 73672
rect 47129 73590 47222 73656
rect 46850 73455 47222 73531
rect 46850 73330 46943 73396
rect 46850 73314 46927 73330
tri 46927 73314 46943 73330 nw
rect 46979 73297 47093 73455
rect 47129 73330 47222 73396
tri 47129 73314 47145 73330 ne
rect 47145 73314 47222 73330
rect 46962 73215 47110 73297
rect 46850 73182 46927 73198
tri 46927 73182 46943 73198 sw
rect 46850 73116 46943 73182
rect 46850 73014 46943 73080
rect 46850 72998 46927 73014
tri 46927 72998 46943 73014 nw
rect 46979 72981 47093 73215
tri 47129 73182 47145 73198 se
rect 47145 73182 47222 73198
rect 47129 73116 47222 73182
rect 47129 73014 47222 73080
tri 47129 72998 47145 73014 ne
rect 47145 72998 47222 73014
rect 46962 72899 47110 72981
rect 46850 72866 46927 72882
tri 46927 72866 46943 72882 sw
rect 46850 72800 46943 72866
rect 46979 72741 47093 72899
tri 47129 72866 47145 72882 se
rect 47145 72866 47222 72882
rect 47129 72800 47222 72866
rect 46850 72665 47222 72741
rect 46850 72540 46943 72606
rect 46850 72524 46927 72540
tri 46927 72524 46943 72540 nw
rect 46979 72507 47093 72665
rect 47129 72540 47222 72606
tri 47129 72524 47145 72540 ne
rect 47145 72524 47222 72540
rect 46962 72425 47110 72507
rect 46850 72392 46927 72408
tri 46927 72392 46943 72408 sw
rect 46850 72326 46943 72392
rect 46850 72224 46943 72290
rect 46850 72208 46927 72224
tri 46927 72208 46943 72224 nw
rect 46979 72191 47093 72425
tri 47129 72392 47145 72408 se
rect 47145 72392 47222 72408
rect 47129 72326 47222 72392
rect 47129 72224 47222 72290
tri 47129 72208 47145 72224 ne
rect 47145 72208 47222 72224
rect 46962 72109 47110 72191
rect 46850 72076 46927 72092
tri 46927 72076 46943 72092 sw
rect 46850 72010 46943 72076
rect 46979 71951 47093 72109
tri 47129 72076 47145 72092 se
rect 47145 72076 47222 72092
rect 47129 72010 47222 72076
rect 46850 71875 47222 71951
rect 46850 71750 46943 71816
rect 46850 71734 46927 71750
tri 46927 71734 46943 71750 nw
rect 46979 71717 47093 71875
rect 47129 71750 47222 71816
tri 47129 71734 47145 71750 ne
rect 47145 71734 47222 71750
rect 46962 71635 47110 71717
rect 46850 71602 46927 71618
tri 46927 71602 46943 71618 sw
rect 46850 71536 46943 71602
rect 46850 71434 46943 71500
rect 46850 71418 46927 71434
tri 46927 71418 46943 71434 nw
rect 46979 71401 47093 71635
tri 47129 71602 47145 71618 se
rect 47145 71602 47222 71618
rect 47129 71536 47222 71602
rect 47129 71434 47222 71500
tri 47129 71418 47145 71434 ne
rect 47145 71418 47222 71434
rect 46962 71319 47110 71401
rect 46850 71286 46927 71302
tri 46927 71286 46943 71302 sw
rect 46850 71220 46943 71286
rect 46979 71161 47093 71319
tri 47129 71286 47145 71302 se
rect 47145 71286 47222 71302
rect 47129 71220 47222 71286
rect 46850 71085 47222 71161
rect 46850 70960 46943 71026
rect 46850 70944 46927 70960
tri 46927 70944 46943 70960 nw
rect 46979 70927 47093 71085
rect 47129 70960 47222 71026
tri 47129 70944 47145 70960 ne
rect 47145 70944 47222 70960
rect 46962 70845 47110 70927
rect 46850 70812 46927 70828
tri 46927 70812 46943 70828 sw
rect 46850 70746 46943 70812
rect 46850 70644 46943 70710
rect 46850 70628 46927 70644
tri 46927 70628 46943 70644 nw
rect 46979 70611 47093 70845
tri 47129 70812 47145 70828 se
rect 47145 70812 47222 70828
rect 47129 70746 47222 70812
rect 47129 70644 47222 70710
tri 47129 70628 47145 70644 ne
rect 47145 70628 47222 70644
rect 46962 70529 47110 70611
rect 46850 70496 46927 70512
tri 46927 70496 46943 70512 sw
rect 46850 70430 46943 70496
rect 46979 70371 47093 70529
tri 47129 70496 47145 70512 se
rect 47145 70496 47222 70512
rect 47129 70430 47222 70496
rect 46850 70295 47222 70371
rect 46850 70170 46943 70236
rect 46850 70154 46927 70170
tri 46927 70154 46943 70170 nw
rect 46979 70137 47093 70295
rect 47129 70170 47222 70236
tri 47129 70154 47145 70170 ne
rect 47145 70154 47222 70170
rect 46962 70055 47110 70137
rect 46850 70022 46927 70038
tri 46927 70022 46943 70038 sw
rect 46850 69956 46943 70022
rect 46850 69854 46943 69920
rect 46850 69838 46927 69854
tri 46927 69838 46943 69854 nw
rect 46979 69821 47093 70055
tri 47129 70022 47145 70038 se
rect 47145 70022 47222 70038
rect 47129 69956 47222 70022
rect 47129 69854 47222 69920
tri 47129 69838 47145 69854 ne
rect 47145 69838 47222 69854
rect 46962 69739 47110 69821
rect 46850 69706 46927 69722
tri 46927 69706 46943 69722 sw
rect 46850 69640 46943 69706
rect 46979 69581 47093 69739
tri 47129 69706 47145 69722 se
rect 47145 69706 47222 69722
rect 47129 69640 47222 69706
rect 46850 69505 47222 69581
rect 46850 69380 46943 69446
rect 46850 69364 46927 69380
tri 46927 69364 46943 69380 nw
rect 46979 69347 47093 69505
rect 47129 69380 47222 69446
tri 47129 69364 47145 69380 ne
rect 47145 69364 47222 69380
rect 46962 69265 47110 69347
rect 46850 69232 46927 69248
tri 46927 69232 46943 69248 sw
rect 46850 69166 46943 69232
rect 46850 69064 46943 69130
rect 46850 69048 46927 69064
tri 46927 69048 46943 69064 nw
rect 46979 69031 47093 69265
tri 47129 69232 47145 69248 se
rect 47145 69232 47222 69248
rect 47129 69166 47222 69232
rect 47129 69064 47222 69130
tri 47129 69048 47145 69064 ne
rect 47145 69048 47222 69064
rect 46962 68949 47110 69031
rect 46850 68916 46927 68932
tri 46927 68916 46943 68932 sw
rect 46850 68850 46943 68916
rect 46979 68791 47093 68949
tri 47129 68916 47145 68932 se
rect 47145 68916 47222 68932
rect 47129 68850 47222 68916
rect 46850 68715 47222 68791
rect 46850 68590 46943 68656
rect 46850 68574 46927 68590
tri 46927 68574 46943 68590 nw
rect 46979 68557 47093 68715
rect 47129 68590 47222 68656
tri 47129 68574 47145 68590 ne
rect 47145 68574 47222 68590
rect 46962 68475 47110 68557
rect 46850 68442 46927 68458
tri 46927 68442 46943 68458 sw
rect 46850 68376 46943 68442
rect 46850 68274 46943 68340
rect 46850 68258 46927 68274
tri 46927 68258 46943 68274 nw
rect 46979 68241 47093 68475
tri 47129 68442 47145 68458 se
rect 47145 68442 47222 68458
rect 47129 68376 47222 68442
rect 47129 68274 47222 68340
tri 47129 68258 47145 68274 ne
rect 47145 68258 47222 68274
rect 46962 68159 47110 68241
rect 46850 68126 46927 68142
tri 46927 68126 46943 68142 sw
rect 46850 68060 46943 68126
rect 46979 68001 47093 68159
tri 47129 68126 47145 68142 se
rect 47145 68126 47222 68142
rect 47129 68060 47222 68126
rect 46850 67925 47222 68001
rect 46850 67800 46943 67866
rect 46850 67784 46927 67800
tri 46927 67784 46943 67800 nw
rect 46979 67767 47093 67925
rect 47129 67800 47222 67866
tri 47129 67784 47145 67800 ne
rect 47145 67784 47222 67800
rect 46962 67685 47110 67767
rect 46850 67652 46927 67668
tri 46927 67652 46943 67668 sw
rect 46850 67586 46943 67652
rect 46850 67484 46943 67550
rect 46850 67468 46927 67484
tri 46927 67468 46943 67484 nw
rect 46979 67451 47093 67685
tri 47129 67652 47145 67668 se
rect 47145 67652 47222 67668
rect 47129 67586 47222 67652
rect 47129 67484 47222 67550
tri 47129 67468 47145 67484 ne
rect 47145 67468 47222 67484
rect 46962 67369 47110 67451
rect 46850 67336 46927 67352
tri 46927 67336 46943 67352 sw
rect 46850 67270 46943 67336
rect 46979 67211 47093 67369
tri 47129 67336 47145 67352 se
rect 47145 67336 47222 67352
rect 47129 67270 47222 67336
rect 46850 67135 47222 67211
rect 46850 67010 46943 67076
rect 46850 66994 46927 67010
tri 46927 66994 46943 67010 nw
rect 46979 66977 47093 67135
rect 47129 67010 47222 67076
tri 47129 66994 47145 67010 ne
rect 47145 66994 47222 67010
rect 46962 66895 47110 66977
rect 46850 66862 46927 66878
tri 46927 66862 46943 66878 sw
rect 46850 66796 46943 66862
rect 46850 66694 46943 66760
rect 46850 66678 46927 66694
tri 46927 66678 46943 66694 nw
rect 46979 66661 47093 66895
tri 47129 66862 47145 66878 se
rect 47145 66862 47222 66878
rect 47129 66796 47222 66862
rect 47129 66694 47222 66760
tri 47129 66678 47145 66694 ne
rect 47145 66678 47222 66694
rect 46962 66579 47110 66661
rect 46850 66546 46927 66562
tri 46927 66546 46943 66562 sw
rect 46850 66480 46943 66546
rect 46979 66421 47093 66579
tri 47129 66546 47145 66562 se
rect 47145 66546 47222 66562
rect 47129 66480 47222 66546
rect 46850 66345 47222 66421
rect 46850 66220 46943 66286
rect 46850 66204 46927 66220
tri 46927 66204 46943 66220 nw
rect 46979 66187 47093 66345
rect 47129 66220 47222 66286
tri 47129 66204 47145 66220 ne
rect 47145 66204 47222 66220
rect 46962 66105 47110 66187
rect 46850 66072 46927 66088
tri 46927 66072 46943 66088 sw
rect 46850 66006 46943 66072
rect 46850 65904 46943 65970
rect 46850 65888 46927 65904
tri 46927 65888 46943 65904 nw
rect 46979 65871 47093 66105
tri 47129 66072 47145 66088 se
rect 47145 66072 47222 66088
rect 47129 66006 47222 66072
rect 47129 65904 47222 65970
tri 47129 65888 47145 65904 ne
rect 47145 65888 47222 65904
rect 46962 65789 47110 65871
rect 46850 65756 46927 65772
tri 46927 65756 46943 65772 sw
rect 46850 65690 46943 65756
rect 46979 65631 47093 65789
tri 47129 65756 47145 65772 se
rect 47145 65756 47222 65772
rect 47129 65690 47222 65756
rect 46850 65555 47222 65631
rect 46850 65430 46943 65496
rect 46850 65414 46927 65430
tri 46927 65414 46943 65430 nw
rect 46979 65397 47093 65555
rect 47129 65430 47222 65496
tri 47129 65414 47145 65430 ne
rect 47145 65414 47222 65430
rect 46962 65315 47110 65397
rect 46850 65282 46927 65298
tri 46927 65282 46943 65298 sw
rect 46850 65216 46943 65282
rect 46850 65114 46943 65180
rect 46850 65098 46927 65114
tri 46927 65098 46943 65114 nw
rect 46979 65081 47093 65315
tri 47129 65282 47145 65298 se
rect 47145 65282 47222 65298
rect 47129 65216 47222 65282
rect 47129 65114 47222 65180
tri 47129 65098 47145 65114 ne
rect 47145 65098 47222 65114
rect 46962 64999 47110 65081
rect 46850 64966 46927 64982
tri 46927 64966 46943 64982 sw
rect 46850 64900 46943 64966
rect 46979 64841 47093 64999
tri 47129 64966 47145 64982 se
rect 47145 64966 47222 64982
rect 47129 64900 47222 64966
rect 46850 64765 47222 64841
rect 46850 64640 46943 64706
rect 46850 64624 46927 64640
tri 46927 64624 46943 64640 nw
rect 46979 64607 47093 64765
rect 47129 64640 47222 64706
tri 47129 64624 47145 64640 ne
rect 47145 64624 47222 64640
rect 46962 64525 47110 64607
rect 46850 64492 46927 64508
tri 46927 64492 46943 64508 sw
rect 46850 64426 46943 64492
rect 46850 64324 46943 64390
rect 46850 64308 46927 64324
tri 46927 64308 46943 64324 nw
rect 46979 64291 47093 64525
tri 47129 64492 47145 64508 se
rect 47145 64492 47222 64508
rect 47129 64426 47222 64492
rect 47129 64324 47222 64390
tri 47129 64308 47145 64324 ne
rect 47145 64308 47222 64324
rect 46962 64209 47110 64291
rect 46850 64176 46927 64192
tri 46927 64176 46943 64192 sw
rect 46850 64110 46943 64176
rect 46979 64051 47093 64209
tri 47129 64176 47145 64192 se
rect 47145 64176 47222 64192
rect 47129 64110 47222 64176
rect 46850 63975 47222 64051
rect 46850 63850 46943 63916
rect 46850 63834 46927 63850
tri 46927 63834 46943 63850 nw
rect 46979 63817 47093 63975
rect 47129 63850 47222 63916
tri 47129 63834 47145 63850 ne
rect 47145 63834 47222 63850
rect 46962 63735 47110 63817
rect 46850 63702 46927 63718
tri 46927 63702 46943 63718 sw
rect 46850 63636 46943 63702
rect 46850 63534 46943 63600
rect 46850 63518 46927 63534
tri 46927 63518 46943 63534 nw
rect 46979 63501 47093 63735
tri 47129 63702 47145 63718 se
rect 47145 63702 47222 63718
rect 47129 63636 47222 63702
rect 47129 63534 47222 63600
tri 47129 63518 47145 63534 ne
rect 47145 63518 47222 63534
rect 46962 63419 47110 63501
rect 46850 63386 46927 63402
tri 46927 63386 46943 63402 sw
rect 46850 63320 46943 63386
rect 46979 63261 47093 63419
tri 47129 63386 47145 63402 se
rect 47145 63386 47222 63402
rect 47129 63320 47222 63386
rect 46850 63185 47222 63261
rect 46850 63060 46943 63126
rect 46850 63044 46927 63060
tri 46927 63044 46943 63060 nw
rect 46979 63027 47093 63185
rect 47129 63060 47222 63126
tri 47129 63044 47145 63060 ne
rect 47145 63044 47222 63060
rect 46962 62945 47110 63027
rect 46850 62912 46927 62928
tri 46927 62912 46943 62928 sw
rect 46850 62846 46943 62912
rect 46850 62744 46943 62810
rect 46850 62728 46927 62744
tri 46927 62728 46943 62744 nw
rect 46979 62711 47093 62945
tri 47129 62912 47145 62928 se
rect 47145 62912 47222 62928
rect 47129 62846 47222 62912
rect 47129 62744 47222 62810
tri 47129 62728 47145 62744 ne
rect 47145 62728 47222 62744
rect 46962 62629 47110 62711
rect 46850 62596 46927 62612
tri 46927 62596 46943 62612 sw
rect 46850 62530 46943 62596
rect 46979 62471 47093 62629
tri 47129 62596 47145 62612 se
rect 47145 62596 47222 62612
rect 47129 62530 47222 62596
rect 46850 62395 47222 62471
rect 46850 62270 46943 62336
rect 46850 62254 46927 62270
tri 46927 62254 46943 62270 nw
rect 46979 62237 47093 62395
rect 47129 62270 47222 62336
tri 47129 62254 47145 62270 ne
rect 47145 62254 47222 62270
rect 46962 62155 47110 62237
rect 46850 62122 46927 62138
tri 46927 62122 46943 62138 sw
rect 46850 62056 46943 62122
rect 46850 61954 46943 62020
rect 46850 61938 46927 61954
tri 46927 61938 46943 61954 nw
rect 46979 61921 47093 62155
tri 47129 62122 47145 62138 se
rect 47145 62122 47222 62138
rect 47129 62056 47222 62122
rect 47129 61954 47222 62020
tri 47129 61938 47145 61954 ne
rect 47145 61938 47222 61954
rect 46962 61839 47110 61921
rect 46850 61806 46927 61822
tri 46927 61806 46943 61822 sw
rect 46850 61740 46943 61806
rect 46979 61681 47093 61839
tri 47129 61806 47145 61822 se
rect 47145 61806 47222 61822
rect 47129 61740 47222 61806
rect 46850 61605 47222 61681
rect 46850 61480 46943 61546
rect 46850 61464 46927 61480
tri 46927 61464 46943 61480 nw
rect 46979 61447 47093 61605
rect 47129 61480 47222 61546
tri 47129 61464 47145 61480 ne
rect 47145 61464 47222 61480
rect 46962 61365 47110 61447
rect 46850 61332 46927 61348
tri 46927 61332 46943 61348 sw
rect 46850 61266 46943 61332
rect 46850 61164 46943 61230
rect 46850 61148 46927 61164
tri 46927 61148 46943 61164 nw
rect 46979 61131 47093 61365
tri 47129 61332 47145 61348 se
rect 47145 61332 47222 61348
rect 47129 61266 47222 61332
rect 47129 61164 47222 61230
tri 47129 61148 47145 61164 ne
rect 47145 61148 47222 61164
rect 46962 61049 47110 61131
rect 46850 61016 46927 61032
tri 46927 61016 46943 61032 sw
rect 46850 60950 46943 61016
rect 46979 60891 47093 61049
tri 47129 61016 47145 61032 se
rect 47145 61016 47222 61032
rect 47129 60950 47222 61016
rect 46850 60815 47222 60891
rect 46850 60690 46943 60756
rect 46850 60674 46927 60690
tri 46927 60674 46943 60690 nw
rect 46979 60657 47093 60815
rect 47129 60690 47222 60756
tri 47129 60674 47145 60690 ne
rect 47145 60674 47222 60690
rect 46962 60575 47110 60657
rect 46850 60542 46927 60558
tri 46927 60542 46943 60558 sw
rect 46850 60476 46943 60542
rect 46850 60374 46943 60440
rect 46850 60358 46927 60374
tri 46927 60358 46943 60374 nw
rect 46979 60341 47093 60575
tri 47129 60542 47145 60558 se
rect 47145 60542 47222 60558
rect 47129 60476 47222 60542
rect 47129 60374 47222 60440
tri 47129 60358 47145 60374 ne
rect 47145 60358 47222 60374
rect 46962 60259 47110 60341
rect 46850 60226 46927 60242
tri 46927 60226 46943 60242 sw
rect 46850 60160 46943 60226
rect 46979 60101 47093 60259
tri 47129 60226 47145 60242 se
rect 47145 60226 47222 60242
rect 47129 60160 47222 60226
rect 46850 60025 47222 60101
rect 46850 59900 46943 59966
rect 46850 59884 46927 59900
tri 46927 59884 46943 59900 nw
rect 46979 59867 47093 60025
rect 47129 59900 47222 59966
tri 47129 59884 47145 59900 ne
rect 47145 59884 47222 59900
rect 46962 59785 47110 59867
rect 46850 59752 46927 59768
tri 46927 59752 46943 59768 sw
rect 46850 59686 46943 59752
rect 46850 59584 46943 59650
rect 46850 59568 46927 59584
tri 46927 59568 46943 59584 nw
rect 46979 59551 47093 59785
tri 47129 59752 47145 59768 se
rect 47145 59752 47222 59768
rect 47129 59686 47222 59752
rect 47129 59584 47222 59650
tri 47129 59568 47145 59584 ne
rect 47145 59568 47222 59584
rect 46962 59469 47110 59551
rect 46850 59436 46927 59452
tri 46927 59436 46943 59452 sw
rect 46850 59370 46943 59436
rect 46979 59311 47093 59469
tri 47129 59436 47145 59452 se
rect 47145 59436 47222 59452
rect 47129 59370 47222 59436
rect 46850 59235 47222 59311
rect 46850 59110 46943 59176
rect 46850 59094 46927 59110
tri 46927 59094 46943 59110 nw
rect 46979 59077 47093 59235
rect 47129 59110 47222 59176
tri 47129 59094 47145 59110 ne
rect 47145 59094 47222 59110
rect 46962 58995 47110 59077
rect 46850 58962 46927 58978
tri 46927 58962 46943 58978 sw
rect 46850 58896 46943 58962
rect 46850 58794 46943 58860
rect 46850 58778 46927 58794
tri 46927 58778 46943 58794 nw
rect 46979 58761 47093 58995
tri 47129 58962 47145 58978 se
rect 47145 58962 47222 58978
rect 47129 58896 47222 58962
rect 47129 58794 47222 58860
tri 47129 58778 47145 58794 ne
rect 47145 58778 47222 58794
rect 46962 58679 47110 58761
rect 46850 58646 46927 58662
tri 46927 58646 46943 58662 sw
rect 46850 58580 46943 58646
rect 46979 58521 47093 58679
tri 47129 58646 47145 58662 se
rect 47145 58646 47222 58662
rect 47129 58580 47222 58646
rect 46850 58445 47222 58521
rect 46850 58320 46943 58386
rect 46850 58304 46927 58320
tri 46927 58304 46943 58320 nw
rect 46979 58287 47093 58445
rect 47129 58320 47222 58386
tri 47129 58304 47145 58320 ne
rect 47145 58304 47222 58320
rect 46962 58205 47110 58287
rect 46850 58172 46927 58188
tri 46927 58172 46943 58188 sw
rect 46850 58106 46943 58172
rect 46850 58004 46943 58070
rect 46850 57988 46927 58004
tri 46927 57988 46943 58004 nw
rect 46979 57971 47093 58205
tri 47129 58172 47145 58188 se
rect 47145 58172 47222 58188
rect 47129 58106 47222 58172
rect 47129 58004 47222 58070
tri 47129 57988 47145 58004 ne
rect 47145 57988 47222 58004
rect 46962 57889 47110 57971
rect 46850 57856 46927 57872
tri 46927 57856 46943 57872 sw
rect 46850 57790 46943 57856
rect 46979 57731 47093 57889
tri 47129 57856 47145 57872 se
rect 47145 57856 47222 57872
rect 47129 57790 47222 57856
rect 46850 57655 47222 57731
rect 46850 57530 46943 57596
rect 46850 57514 46927 57530
tri 46927 57514 46943 57530 nw
rect 46979 57497 47093 57655
rect 47129 57530 47222 57596
tri 47129 57514 47145 57530 ne
rect 47145 57514 47222 57530
rect 46962 57415 47110 57497
rect 46850 57382 46927 57398
tri 46927 57382 46943 57398 sw
rect 46850 57316 46943 57382
rect 46850 57214 46943 57280
rect 46850 57198 46927 57214
tri 46927 57198 46943 57214 nw
rect 46979 57181 47093 57415
tri 47129 57382 47145 57398 se
rect 47145 57382 47222 57398
rect 47129 57316 47222 57382
rect 47129 57214 47222 57280
tri 47129 57198 47145 57214 ne
rect 47145 57198 47222 57214
rect 46962 57099 47110 57181
rect 46850 57066 46927 57082
tri 46927 57066 46943 57082 sw
rect 46850 57000 46943 57066
rect 46979 56941 47093 57099
tri 47129 57066 47145 57082 se
rect 47145 57066 47222 57082
rect 47129 57000 47222 57066
rect 46850 56865 47222 56941
rect 46850 56740 46943 56806
rect 46850 56724 46927 56740
tri 46927 56724 46943 56740 nw
rect 46979 56707 47093 56865
rect 47129 56740 47222 56806
tri 47129 56724 47145 56740 ne
rect 47145 56724 47222 56740
rect 46962 56625 47110 56707
rect 46850 56592 46927 56608
tri 46927 56592 46943 56608 sw
rect 46850 56526 46943 56592
rect 46850 56424 46943 56490
rect 46850 56408 46927 56424
tri 46927 56408 46943 56424 nw
rect 46979 56391 47093 56625
tri 47129 56592 47145 56608 se
rect 47145 56592 47222 56608
rect 47129 56526 47222 56592
rect 47129 56424 47222 56490
tri 47129 56408 47145 56424 ne
rect 47145 56408 47222 56424
rect 46962 56309 47110 56391
rect 46850 56276 46927 56292
tri 46927 56276 46943 56292 sw
rect 46850 56210 46943 56276
rect 46979 56151 47093 56309
tri 47129 56276 47145 56292 se
rect 47145 56276 47222 56292
rect 47129 56210 47222 56276
rect 46850 56075 47222 56151
rect 46850 55950 46943 56016
rect 46850 55934 46927 55950
tri 46927 55934 46943 55950 nw
rect 46979 55917 47093 56075
rect 47129 55950 47222 56016
tri 47129 55934 47145 55950 ne
rect 47145 55934 47222 55950
rect 46962 55835 47110 55917
rect 46850 55802 46927 55818
tri 46927 55802 46943 55818 sw
rect 46850 55736 46943 55802
rect 46850 55634 46943 55700
rect 46850 55618 46927 55634
tri 46927 55618 46943 55634 nw
rect 46979 55601 47093 55835
tri 47129 55802 47145 55818 se
rect 47145 55802 47222 55818
rect 47129 55736 47222 55802
rect 47129 55634 47222 55700
tri 47129 55618 47145 55634 ne
rect 47145 55618 47222 55634
rect 46962 55519 47110 55601
rect 46850 55486 46927 55502
tri 46927 55486 46943 55502 sw
rect 46850 55420 46943 55486
rect 46979 55361 47093 55519
tri 47129 55486 47145 55502 se
rect 47145 55486 47222 55502
rect 47129 55420 47222 55486
rect 46850 55285 47222 55361
rect 46850 55160 46943 55226
rect 46850 55144 46927 55160
tri 46927 55144 46943 55160 nw
rect 46979 55127 47093 55285
rect 47129 55160 47222 55226
tri 47129 55144 47145 55160 ne
rect 47145 55144 47222 55160
rect 46962 55045 47110 55127
rect 46850 55012 46927 55028
tri 46927 55012 46943 55028 sw
rect 46850 54946 46943 55012
rect 46850 54844 46943 54910
rect 46850 54828 46927 54844
tri 46927 54828 46943 54844 nw
rect 46979 54811 47093 55045
tri 47129 55012 47145 55028 se
rect 47145 55012 47222 55028
rect 47129 54946 47222 55012
rect 47129 54844 47222 54910
tri 47129 54828 47145 54844 ne
rect 47145 54828 47222 54844
rect 46962 54729 47110 54811
rect 46850 54696 46927 54712
tri 46927 54696 46943 54712 sw
rect 46850 54630 46943 54696
rect 46979 54571 47093 54729
tri 47129 54696 47145 54712 se
rect 47145 54696 47222 54712
rect 47129 54630 47222 54696
rect 46850 54495 47222 54571
rect 46850 54370 46943 54436
rect 46850 54354 46927 54370
tri 46927 54354 46943 54370 nw
rect 46979 54337 47093 54495
rect 47129 54370 47222 54436
tri 47129 54354 47145 54370 ne
rect 47145 54354 47222 54370
rect 46962 54255 47110 54337
rect 46850 54222 46927 54238
tri 46927 54222 46943 54238 sw
rect 46850 54156 46943 54222
rect 46850 54054 46943 54120
rect 46850 54038 46927 54054
tri 46927 54038 46943 54054 nw
rect 46979 54021 47093 54255
tri 47129 54222 47145 54238 se
rect 47145 54222 47222 54238
rect 47129 54156 47222 54222
rect 47129 54054 47222 54120
tri 47129 54038 47145 54054 ne
rect 47145 54038 47222 54054
rect 46962 53939 47110 54021
rect 46850 53906 46927 53922
tri 46927 53906 46943 53922 sw
rect 46850 53840 46943 53906
rect 46979 53781 47093 53939
tri 47129 53906 47145 53922 se
rect 47145 53906 47222 53922
rect 47129 53840 47222 53906
rect 46850 53705 47222 53781
rect 46850 53580 46943 53646
rect 46850 53564 46927 53580
tri 46927 53564 46943 53580 nw
rect 46979 53547 47093 53705
rect 47129 53580 47222 53646
tri 47129 53564 47145 53580 ne
rect 47145 53564 47222 53580
rect 46962 53465 47110 53547
rect 46850 53432 46927 53448
tri 46927 53432 46943 53448 sw
rect 46850 53366 46943 53432
rect 46850 53264 46943 53330
rect 46850 53248 46927 53264
tri 46927 53248 46943 53264 nw
rect 46979 53231 47093 53465
tri 47129 53432 47145 53448 se
rect 47145 53432 47222 53448
rect 47129 53366 47222 53432
rect 47129 53264 47222 53330
tri 47129 53248 47145 53264 ne
rect 47145 53248 47222 53264
rect 46962 53149 47110 53231
rect 46850 53116 46927 53132
tri 46927 53116 46943 53132 sw
rect 46850 53050 46943 53116
rect 46979 52991 47093 53149
tri 47129 53116 47145 53132 se
rect 47145 53116 47222 53132
rect 47129 53050 47222 53116
rect 46850 52915 47222 52991
rect 46850 52790 46943 52856
rect 46850 52774 46927 52790
tri 46927 52774 46943 52790 nw
rect 46979 52757 47093 52915
rect 47129 52790 47222 52856
tri 47129 52774 47145 52790 ne
rect 47145 52774 47222 52790
rect 46962 52675 47110 52757
rect 46850 52642 46927 52658
tri 46927 52642 46943 52658 sw
rect 46850 52576 46943 52642
rect 46850 52474 46943 52540
rect 46850 52458 46927 52474
tri 46927 52458 46943 52474 nw
rect 46979 52441 47093 52675
tri 47129 52642 47145 52658 se
rect 47145 52642 47222 52658
rect 47129 52576 47222 52642
rect 47129 52474 47222 52540
tri 47129 52458 47145 52474 ne
rect 47145 52458 47222 52474
rect 46962 52359 47110 52441
rect 46850 52326 46927 52342
tri 46927 52326 46943 52342 sw
rect 46850 52260 46943 52326
rect 46979 52201 47093 52359
tri 47129 52326 47145 52342 se
rect 47145 52326 47222 52342
rect 47129 52260 47222 52326
rect 46850 52125 47222 52201
rect 46850 52000 46943 52066
rect 46850 51984 46927 52000
tri 46927 51984 46943 52000 nw
rect 46979 51967 47093 52125
rect 47129 52000 47222 52066
tri 47129 51984 47145 52000 ne
rect 47145 51984 47222 52000
rect 46962 51885 47110 51967
rect 46850 51852 46927 51868
tri 46927 51852 46943 51868 sw
rect 46850 51786 46943 51852
rect 46850 51684 46943 51750
rect 46850 51668 46927 51684
tri 46927 51668 46943 51684 nw
rect 46979 51651 47093 51885
tri 47129 51852 47145 51868 se
rect 47145 51852 47222 51868
rect 47129 51786 47222 51852
rect 47129 51684 47222 51750
tri 47129 51668 47145 51684 ne
rect 47145 51668 47222 51684
rect 46962 51569 47110 51651
rect 46850 51536 46927 51552
tri 46927 51536 46943 51552 sw
rect 46850 51470 46943 51536
rect 46979 51411 47093 51569
tri 47129 51536 47145 51552 se
rect 47145 51536 47222 51552
rect 47129 51470 47222 51536
rect 46850 51335 47222 51411
rect 46850 51210 46943 51276
rect 46850 51194 46927 51210
tri 46927 51194 46943 51210 nw
rect 46979 51177 47093 51335
rect 47129 51210 47222 51276
tri 47129 51194 47145 51210 ne
rect 47145 51194 47222 51210
rect 46962 51095 47110 51177
rect 46850 51062 46927 51078
tri 46927 51062 46943 51078 sw
rect 46850 50996 46943 51062
rect 46850 50894 46943 50960
rect 46850 50878 46927 50894
tri 46927 50878 46943 50894 nw
rect 46979 50861 47093 51095
tri 47129 51062 47145 51078 se
rect 47145 51062 47222 51078
rect 47129 50996 47222 51062
rect 47129 50894 47222 50960
tri 47129 50878 47145 50894 ne
rect 47145 50878 47222 50894
rect 46962 50779 47110 50861
rect 46850 50746 46927 50762
tri 46927 50746 46943 50762 sw
rect 46850 50680 46943 50746
rect 46979 50621 47093 50779
tri 47129 50746 47145 50762 se
rect 47145 50746 47222 50762
rect 47129 50680 47222 50746
rect 46850 50545 47222 50621
rect 46850 50420 46943 50486
rect 46850 50404 46927 50420
tri 46927 50404 46943 50420 nw
rect 46979 50387 47093 50545
rect 47129 50420 47222 50486
tri 47129 50404 47145 50420 ne
rect 47145 50404 47222 50420
rect 46962 50305 47110 50387
rect 46850 50272 46927 50288
tri 46927 50272 46943 50288 sw
rect 46850 50206 46943 50272
rect 46850 50104 46943 50170
rect 46850 50088 46927 50104
tri 46927 50088 46943 50104 nw
rect 46979 50071 47093 50305
tri 47129 50272 47145 50288 se
rect 47145 50272 47222 50288
rect 47129 50206 47222 50272
rect 47129 50104 47222 50170
tri 47129 50088 47145 50104 ne
rect 47145 50088 47222 50104
rect 46962 49989 47110 50071
rect 46850 49956 46927 49972
tri 46927 49956 46943 49972 sw
rect 46850 49890 46943 49956
rect 46979 49831 47093 49989
tri 47129 49956 47145 49972 se
rect 47145 49956 47222 49972
rect 47129 49890 47222 49956
rect 46850 49755 47222 49831
rect 46850 49630 46943 49696
rect 46850 49614 46927 49630
tri 46927 49614 46943 49630 nw
rect 46979 49597 47093 49755
rect 47129 49630 47222 49696
tri 47129 49614 47145 49630 ne
rect 47145 49614 47222 49630
rect 46962 49515 47110 49597
rect 46850 49482 46927 49498
tri 46927 49482 46943 49498 sw
rect 46850 49416 46943 49482
rect 46850 49314 46943 49380
rect 46850 49298 46927 49314
tri 46927 49298 46943 49314 nw
rect 46979 49281 47093 49515
tri 47129 49482 47145 49498 se
rect 47145 49482 47222 49498
rect 47129 49416 47222 49482
rect 47129 49314 47222 49380
tri 47129 49298 47145 49314 ne
rect 47145 49298 47222 49314
rect 46962 49199 47110 49281
rect 46850 49166 46927 49182
tri 46927 49166 46943 49182 sw
rect 46850 49100 46943 49166
rect 46979 49041 47093 49199
tri 47129 49166 47145 49182 se
rect 47145 49166 47222 49182
rect 47129 49100 47222 49166
rect 46850 48965 47222 49041
rect 46850 48840 46943 48906
rect 46850 48824 46927 48840
tri 46927 48824 46943 48840 nw
rect 46979 48807 47093 48965
rect 47129 48840 47222 48906
tri 47129 48824 47145 48840 ne
rect 47145 48824 47222 48840
rect 46962 48725 47110 48807
rect 46850 48692 46927 48708
tri 46927 48692 46943 48708 sw
rect 46850 48626 46943 48692
rect 46850 48524 46943 48590
rect 46850 48508 46927 48524
tri 46927 48508 46943 48524 nw
rect 46979 48491 47093 48725
tri 47129 48692 47145 48708 se
rect 47145 48692 47222 48708
rect 47129 48626 47222 48692
rect 47129 48524 47222 48590
tri 47129 48508 47145 48524 ne
rect 47145 48508 47222 48524
rect 46962 48409 47110 48491
rect 46850 48376 46927 48392
tri 46927 48376 46943 48392 sw
rect 46850 48310 46943 48376
rect 46979 48251 47093 48409
tri 47129 48376 47145 48392 se
rect 47145 48376 47222 48392
rect 47129 48310 47222 48376
rect 46850 48175 47222 48251
rect 46850 48050 46943 48116
rect 46850 48034 46927 48050
tri 46927 48034 46943 48050 nw
rect 46979 48017 47093 48175
rect 47129 48050 47222 48116
tri 47129 48034 47145 48050 ne
rect 47145 48034 47222 48050
rect 46962 47935 47110 48017
rect 46850 47902 46927 47918
tri 46927 47902 46943 47918 sw
rect 46850 47836 46943 47902
rect 46850 47734 46943 47800
rect 46850 47718 46927 47734
tri 46927 47718 46943 47734 nw
rect 46979 47701 47093 47935
tri 47129 47902 47145 47918 se
rect 47145 47902 47222 47918
rect 47129 47836 47222 47902
rect 47129 47734 47222 47800
tri 47129 47718 47145 47734 ne
rect 47145 47718 47222 47734
rect 46962 47619 47110 47701
rect 46850 47586 46927 47602
tri 46927 47586 46943 47602 sw
rect 46850 47520 46943 47586
rect 46979 47461 47093 47619
tri 47129 47586 47145 47602 se
rect 47145 47586 47222 47602
rect 47129 47520 47222 47586
rect 46850 47385 47222 47461
rect 46850 47260 46943 47326
rect 46850 47244 46927 47260
tri 46927 47244 46943 47260 nw
rect 46979 47227 47093 47385
rect 47129 47260 47222 47326
tri 47129 47244 47145 47260 ne
rect 47145 47244 47222 47260
rect 46962 47145 47110 47227
rect 46850 47112 46927 47128
tri 46927 47112 46943 47128 sw
rect 46850 47046 46943 47112
rect 46850 46944 46943 47010
rect 46850 46928 46927 46944
tri 46927 46928 46943 46944 nw
rect 46979 46911 47093 47145
tri 47129 47112 47145 47128 se
rect 47145 47112 47222 47128
rect 47129 47046 47222 47112
rect 47129 46944 47222 47010
tri 47129 46928 47145 46944 ne
rect 47145 46928 47222 46944
rect 46962 46829 47110 46911
rect 46850 46796 46927 46812
tri 46927 46796 46943 46812 sw
rect 46850 46730 46943 46796
rect 46979 46671 47093 46829
tri 47129 46796 47145 46812 se
rect 47145 46796 47222 46812
rect 47129 46730 47222 46796
rect 46850 46595 47222 46671
rect 46850 46470 46943 46536
rect 46850 46454 46927 46470
tri 46927 46454 46943 46470 nw
rect 46979 46437 47093 46595
rect 47129 46470 47222 46536
tri 47129 46454 47145 46470 ne
rect 47145 46454 47222 46470
rect 46962 46355 47110 46437
rect 46850 46322 46927 46338
tri 46927 46322 46943 46338 sw
rect 46850 46256 46943 46322
rect 46850 46154 46943 46220
rect 46850 46138 46927 46154
tri 46927 46138 46943 46154 nw
rect 46979 46121 47093 46355
tri 47129 46322 47145 46338 se
rect 47145 46322 47222 46338
rect 47129 46256 47222 46322
rect 47129 46154 47222 46220
tri 47129 46138 47145 46154 ne
rect 47145 46138 47222 46154
rect 46962 46039 47110 46121
rect 46850 46006 46927 46022
tri 46927 46006 46943 46022 sw
rect 46850 45940 46943 46006
rect 46979 45881 47093 46039
tri 47129 46006 47145 46022 se
rect 47145 46006 47222 46022
rect 47129 45940 47222 46006
rect 46850 45805 47222 45881
rect 46850 45680 46943 45746
rect 46850 45664 46927 45680
tri 46927 45664 46943 45680 nw
rect 46979 45647 47093 45805
rect 47129 45680 47222 45746
tri 47129 45664 47145 45680 ne
rect 47145 45664 47222 45680
rect 46962 45565 47110 45647
rect 46850 45532 46927 45548
tri 46927 45532 46943 45548 sw
rect 46850 45466 46943 45532
rect 46850 45364 46943 45430
rect 46850 45348 46927 45364
tri 46927 45348 46943 45364 nw
rect 46979 45331 47093 45565
tri 47129 45532 47145 45548 se
rect 47145 45532 47222 45548
rect 47129 45466 47222 45532
rect 47129 45364 47222 45430
tri 47129 45348 47145 45364 ne
rect 47145 45348 47222 45364
rect 46962 45249 47110 45331
rect 46850 45216 46927 45232
tri 46927 45216 46943 45232 sw
rect 46850 45150 46943 45216
rect 46979 45091 47093 45249
tri 47129 45216 47145 45232 se
rect 47145 45216 47222 45232
rect 47129 45150 47222 45216
rect 46850 45015 47222 45091
rect 46850 44890 46943 44956
rect 46850 44874 46927 44890
tri 46927 44874 46943 44890 nw
rect 46979 44857 47093 45015
rect 47129 44890 47222 44956
tri 47129 44874 47145 44890 ne
rect 47145 44874 47222 44890
rect 46962 44775 47110 44857
rect 46850 44742 46927 44758
tri 46927 44742 46943 44758 sw
rect 46850 44676 46943 44742
rect 46850 44574 46943 44640
rect 46850 44558 46927 44574
tri 46927 44558 46943 44574 nw
rect 46979 44541 47093 44775
tri 47129 44742 47145 44758 se
rect 47145 44742 47222 44758
rect 47129 44676 47222 44742
rect 47129 44574 47222 44640
tri 47129 44558 47145 44574 ne
rect 47145 44558 47222 44574
rect 46962 44459 47110 44541
rect 46850 44426 46927 44442
tri 46927 44426 46943 44442 sw
rect 46850 44360 46943 44426
rect 46979 44301 47093 44459
tri 47129 44426 47145 44442 se
rect 47145 44426 47222 44442
rect 47129 44360 47222 44426
rect 46850 44225 47222 44301
rect 46850 44100 46943 44166
rect 46850 44084 46927 44100
tri 46927 44084 46943 44100 nw
rect 46979 44067 47093 44225
rect 47129 44100 47222 44166
tri 47129 44084 47145 44100 ne
rect 47145 44084 47222 44100
rect 46962 43985 47110 44067
rect 46850 43952 46927 43968
tri 46927 43952 46943 43968 sw
rect 46850 43886 46943 43952
rect 46850 43784 46943 43850
rect 46850 43768 46927 43784
tri 46927 43768 46943 43784 nw
rect 46979 43751 47093 43985
tri 47129 43952 47145 43968 se
rect 47145 43952 47222 43968
rect 47129 43886 47222 43952
rect 47129 43784 47222 43850
tri 47129 43768 47145 43784 ne
rect 47145 43768 47222 43784
rect 46962 43669 47110 43751
rect 46850 43636 46927 43652
tri 46927 43636 46943 43652 sw
rect 46850 43570 46943 43636
rect 46979 43511 47093 43669
tri 47129 43636 47145 43652 se
rect 47145 43636 47222 43652
rect 47129 43570 47222 43636
rect 46850 43435 47222 43511
rect 46850 43310 46943 43376
rect 46850 43294 46927 43310
tri 46927 43294 46943 43310 nw
rect 46979 43277 47093 43435
rect 47129 43310 47222 43376
tri 47129 43294 47145 43310 ne
rect 47145 43294 47222 43310
rect 46962 43195 47110 43277
rect 46850 43162 46927 43178
tri 46927 43162 46943 43178 sw
rect 46850 43096 46943 43162
rect 46850 42994 46943 43060
rect 46850 42978 46927 42994
tri 46927 42978 46943 42994 nw
rect 46979 42961 47093 43195
tri 47129 43162 47145 43178 se
rect 47145 43162 47222 43178
rect 47129 43096 47222 43162
rect 47129 42994 47222 43060
tri 47129 42978 47145 42994 ne
rect 47145 42978 47222 42994
rect 46962 42879 47110 42961
rect 46850 42846 46927 42862
tri 46927 42846 46943 42862 sw
rect 46850 42780 46943 42846
rect 46979 42721 47093 42879
tri 47129 42846 47145 42862 se
rect 47145 42846 47222 42862
rect 47129 42780 47222 42846
rect 46850 42645 47222 42721
rect 46850 42520 46943 42586
rect 46850 42504 46927 42520
tri 46927 42504 46943 42520 nw
rect 46979 42487 47093 42645
rect 47129 42520 47222 42586
tri 47129 42504 47145 42520 ne
rect 47145 42504 47222 42520
rect 46962 42405 47110 42487
rect 46850 42372 46927 42388
tri 46927 42372 46943 42388 sw
rect 46850 42306 46943 42372
rect 46850 42204 46943 42270
rect 46850 42188 46927 42204
tri 46927 42188 46943 42204 nw
rect 46979 42171 47093 42405
tri 47129 42372 47145 42388 se
rect 47145 42372 47222 42388
rect 47129 42306 47222 42372
rect 47129 42204 47222 42270
tri 47129 42188 47145 42204 ne
rect 47145 42188 47222 42204
rect 46962 42089 47110 42171
rect 46850 42056 46927 42072
tri 46927 42056 46943 42072 sw
rect 46850 41990 46943 42056
rect 46979 41931 47093 42089
tri 47129 42056 47145 42072 se
rect 47145 42056 47222 42072
rect 47129 41990 47222 42056
rect 46850 41855 47222 41931
rect 46850 41730 46943 41796
rect 46850 41714 46927 41730
tri 46927 41714 46943 41730 nw
rect 46979 41697 47093 41855
rect 47129 41730 47222 41796
tri 47129 41714 47145 41730 ne
rect 47145 41714 47222 41730
rect 46962 41615 47110 41697
rect 46850 41582 46927 41598
tri 46927 41582 46943 41598 sw
rect 46850 41516 46943 41582
rect 46850 41414 46943 41480
rect 46850 41398 46927 41414
tri 46927 41398 46943 41414 nw
rect 46979 41381 47093 41615
tri 47129 41582 47145 41598 se
rect 47145 41582 47222 41598
rect 47129 41516 47222 41582
rect 47129 41414 47222 41480
tri 47129 41398 47145 41414 ne
rect 47145 41398 47222 41414
rect 46962 41299 47110 41381
rect 46850 41266 46927 41282
tri 46927 41266 46943 41282 sw
rect 46850 41200 46943 41266
rect 46979 41141 47093 41299
tri 47129 41266 47145 41282 se
rect 47145 41266 47222 41282
rect 47129 41200 47222 41266
rect 46850 41065 47222 41141
rect 46850 40940 46943 41006
rect 46850 40924 46927 40940
tri 46927 40924 46943 40940 nw
rect 46979 40907 47093 41065
rect 47129 40940 47222 41006
tri 47129 40924 47145 40940 ne
rect 47145 40924 47222 40940
rect 46962 40825 47110 40907
rect 46850 40792 46927 40808
tri 46927 40792 46943 40808 sw
rect 46850 40726 46943 40792
rect 46850 40624 46943 40690
rect 46850 40608 46927 40624
tri 46927 40608 46943 40624 nw
rect 46979 40591 47093 40825
tri 47129 40792 47145 40808 se
rect 47145 40792 47222 40808
rect 47129 40726 47222 40792
rect 47129 40624 47222 40690
tri 47129 40608 47145 40624 ne
rect 47145 40608 47222 40624
rect 46962 40509 47110 40591
rect 46850 40476 46927 40492
tri 46927 40476 46943 40492 sw
rect 46850 40410 46943 40476
rect 46979 40351 47093 40509
tri 47129 40476 47145 40492 se
rect 47145 40476 47222 40492
rect 47129 40410 47222 40476
rect 46850 40275 47222 40351
rect 46850 40150 46943 40216
rect 46850 40134 46927 40150
tri 46927 40134 46943 40150 nw
rect 46979 40117 47093 40275
rect 47129 40150 47222 40216
tri 47129 40134 47145 40150 ne
rect 47145 40134 47222 40150
rect 46962 40035 47110 40117
rect 46850 40002 46927 40018
tri 46927 40002 46943 40018 sw
rect 46850 39936 46943 40002
rect 46850 39834 46943 39900
rect 46850 39818 46927 39834
tri 46927 39818 46943 39834 nw
rect 46979 39801 47093 40035
tri 47129 40002 47145 40018 se
rect 47145 40002 47222 40018
rect 47129 39936 47222 40002
rect 47129 39834 47222 39900
tri 47129 39818 47145 39834 ne
rect 47145 39818 47222 39834
rect 46962 39719 47110 39801
rect 46850 39686 46927 39702
tri 46927 39686 46943 39702 sw
rect 46850 39620 46943 39686
rect 46979 39561 47093 39719
tri 47129 39686 47145 39702 se
rect 47145 39686 47222 39702
rect 47129 39620 47222 39686
rect 46850 39485 47222 39561
rect 46850 39360 46943 39426
rect 46850 39344 46927 39360
tri 46927 39344 46943 39360 nw
rect 46979 39327 47093 39485
rect 47129 39360 47222 39426
tri 47129 39344 47145 39360 ne
rect 47145 39344 47222 39360
rect 46962 39245 47110 39327
rect 46850 39212 46927 39228
tri 46927 39212 46943 39228 sw
rect 46850 39146 46943 39212
rect 46850 39044 46943 39110
rect 46850 39028 46927 39044
tri 46927 39028 46943 39044 nw
rect 46979 39011 47093 39245
tri 47129 39212 47145 39228 se
rect 47145 39212 47222 39228
rect 47129 39146 47222 39212
rect 47129 39044 47222 39110
tri 47129 39028 47145 39044 ne
rect 47145 39028 47222 39044
rect 46962 38929 47110 39011
rect 46850 38896 46927 38912
tri 46927 38896 46943 38912 sw
rect 46850 38830 46943 38896
rect 46979 38771 47093 38929
tri 47129 38896 47145 38912 se
rect 47145 38896 47222 38912
rect 47129 38830 47222 38896
rect 46850 38695 47222 38771
rect 46850 38570 46943 38636
rect 46850 38554 46927 38570
tri 46927 38554 46943 38570 nw
rect 46979 38537 47093 38695
rect 47129 38570 47222 38636
tri 47129 38554 47145 38570 ne
rect 47145 38554 47222 38570
rect 46962 38455 47110 38537
rect 46850 38422 46927 38438
tri 46927 38422 46943 38438 sw
rect 46850 38356 46943 38422
rect 46850 38254 46943 38320
rect 46850 38238 46927 38254
tri 46927 38238 46943 38254 nw
rect 46979 38221 47093 38455
tri 47129 38422 47145 38438 se
rect 47145 38422 47222 38438
rect 47129 38356 47222 38422
rect 47129 38254 47222 38320
tri 47129 38238 47145 38254 ne
rect 47145 38238 47222 38254
rect 46962 38139 47110 38221
rect 46850 38106 46927 38122
tri 46927 38106 46943 38122 sw
rect 46850 38040 46943 38106
rect 46979 37981 47093 38139
tri 47129 38106 47145 38122 se
rect 47145 38106 47222 38122
rect 47129 38040 47222 38106
rect 46850 37905 47222 37981
rect 46850 37780 46943 37846
rect 46850 37764 46927 37780
tri 46927 37764 46943 37780 nw
rect 46979 37747 47093 37905
rect 47129 37780 47222 37846
tri 47129 37764 47145 37780 ne
rect 47145 37764 47222 37780
rect 46962 37665 47110 37747
rect 46850 37632 46927 37648
tri 46927 37632 46943 37648 sw
rect 46850 37566 46943 37632
rect 46850 37464 46943 37530
rect 46850 37448 46927 37464
tri 46927 37448 46943 37464 nw
rect 46979 37431 47093 37665
tri 47129 37632 47145 37648 se
rect 47145 37632 47222 37648
rect 47129 37566 47222 37632
rect 47129 37464 47222 37530
tri 47129 37448 47145 37464 ne
rect 47145 37448 47222 37464
rect 46962 37349 47110 37431
rect 46850 37316 46927 37332
tri 46927 37316 46943 37332 sw
rect 46850 37250 46943 37316
rect 46979 37191 47093 37349
tri 47129 37316 47145 37332 se
rect 47145 37316 47222 37332
rect 47129 37250 47222 37316
rect 46850 37115 47222 37191
rect 46850 36990 46943 37056
rect 46850 36974 46927 36990
tri 46927 36974 46943 36990 nw
rect 46979 36957 47093 37115
rect 47129 36990 47222 37056
tri 47129 36974 47145 36990 ne
rect 47145 36974 47222 36990
rect 46962 36875 47110 36957
rect 46850 36842 46927 36858
tri 46927 36842 46943 36858 sw
rect 46850 36776 46943 36842
rect 46850 36674 46943 36740
rect 46850 36658 46927 36674
tri 46927 36658 46943 36674 nw
rect 46979 36641 47093 36875
tri 47129 36842 47145 36858 se
rect 47145 36842 47222 36858
rect 47129 36776 47222 36842
rect 47129 36674 47222 36740
tri 47129 36658 47145 36674 ne
rect 47145 36658 47222 36674
rect 46962 36559 47110 36641
rect 46850 36526 46927 36542
tri 46927 36526 46943 36542 sw
rect 46850 36460 46943 36526
rect 46979 36401 47093 36559
tri 47129 36526 47145 36542 se
rect 47145 36526 47222 36542
rect 47129 36460 47222 36526
rect 46850 36325 47222 36401
rect 46850 36200 46943 36266
rect 46850 36184 46927 36200
tri 46927 36184 46943 36200 nw
rect 46979 36167 47093 36325
rect 47129 36200 47222 36266
tri 47129 36184 47145 36200 ne
rect 47145 36184 47222 36200
rect 46962 36085 47110 36167
rect 46850 36052 46927 36068
tri 46927 36052 46943 36068 sw
rect 46850 35986 46943 36052
rect 46850 35884 46943 35950
rect 46850 35868 46927 35884
tri 46927 35868 46943 35884 nw
rect 46979 35851 47093 36085
tri 47129 36052 47145 36068 se
rect 47145 36052 47222 36068
rect 47129 35986 47222 36052
rect 47129 35884 47222 35950
tri 47129 35868 47145 35884 ne
rect 47145 35868 47222 35884
rect 46962 35769 47110 35851
rect 46850 35736 46927 35752
tri 46927 35736 46943 35752 sw
rect 46850 35670 46943 35736
rect 46979 35611 47093 35769
tri 47129 35736 47145 35752 se
rect 47145 35736 47222 35752
rect 47129 35670 47222 35736
rect 46850 35535 47222 35611
rect 46850 35410 46943 35476
rect 46850 35394 46927 35410
tri 46927 35394 46943 35410 nw
rect 46979 35377 47093 35535
rect 47129 35410 47222 35476
tri 47129 35394 47145 35410 ne
rect 47145 35394 47222 35410
rect 46962 35295 47110 35377
rect 46850 35262 46927 35278
tri 46927 35262 46943 35278 sw
rect 46850 35196 46943 35262
rect 46850 35094 46943 35160
rect 46850 35078 46927 35094
tri 46927 35078 46943 35094 nw
rect 46979 35061 47093 35295
tri 47129 35262 47145 35278 se
rect 47145 35262 47222 35278
rect 47129 35196 47222 35262
rect 47129 35094 47222 35160
tri 47129 35078 47145 35094 ne
rect 47145 35078 47222 35094
rect 46962 34979 47110 35061
rect 46850 34946 46927 34962
tri 46927 34946 46943 34962 sw
rect 46850 34880 46943 34946
rect 46979 34821 47093 34979
tri 47129 34946 47145 34962 se
rect 47145 34946 47222 34962
rect 47129 34880 47222 34946
rect 46850 34745 47222 34821
rect 46850 34620 46943 34686
rect 46850 34604 46927 34620
tri 46927 34604 46943 34620 nw
rect 46979 34587 47093 34745
rect 47129 34620 47222 34686
tri 47129 34604 47145 34620 ne
rect 47145 34604 47222 34620
rect 46962 34505 47110 34587
rect 46850 34472 46927 34488
tri 46927 34472 46943 34488 sw
rect 46850 34406 46943 34472
rect 46850 34304 46943 34370
rect 46850 34288 46927 34304
tri 46927 34288 46943 34304 nw
rect 46979 34271 47093 34505
tri 47129 34472 47145 34488 se
rect 47145 34472 47222 34488
rect 47129 34406 47222 34472
rect 47129 34304 47222 34370
tri 47129 34288 47145 34304 ne
rect 47145 34288 47222 34304
rect 46962 34189 47110 34271
rect 46850 34156 46927 34172
tri 46927 34156 46943 34172 sw
rect 46850 34090 46943 34156
rect 46979 34031 47093 34189
tri 47129 34156 47145 34172 se
rect 47145 34156 47222 34172
rect 47129 34090 47222 34156
rect 46850 33955 47222 34031
rect 46850 33830 46943 33896
rect 46850 33814 46927 33830
tri 46927 33814 46943 33830 nw
rect 46979 33797 47093 33955
rect 47129 33830 47222 33896
tri 47129 33814 47145 33830 ne
rect 47145 33814 47222 33830
rect 46962 33715 47110 33797
rect 46850 33682 46927 33698
tri 46927 33682 46943 33698 sw
rect 46850 33616 46943 33682
rect 46850 33514 46943 33580
rect 46850 33498 46927 33514
tri 46927 33498 46943 33514 nw
rect 46979 33481 47093 33715
tri 47129 33682 47145 33698 se
rect 47145 33682 47222 33698
rect 47129 33616 47222 33682
rect 47129 33514 47222 33580
tri 47129 33498 47145 33514 ne
rect 47145 33498 47222 33514
rect 46962 33399 47110 33481
rect 46850 33366 46927 33382
tri 46927 33366 46943 33382 sw
rect 46850 33300 46943 33366
rect 46979 33241 47093 33399
tri 47129 33366 47145 33382 se
rect 47145 33366 47222 33382
rect 47129 33300 47222 33366
rect 46850 33165 47222 33241
rect 46850 33040 46943 33106
rect 46850 33024 46927 33040
tri 46927 33024 46943 33040 nw
rect 46979 33007 47093 33165
rect 47129 33040 47222 33106
tri 47129 33024 47145 33040 ne
rect 47145 33024 47222 33040
rect 46962 32925 47110 33007
rect 46850 32892 46927 32908
tri 46927 32892 46943 32908 sw
rect 46850 32826 46943 32892
rect 46850 32724 46943 32790
rect 46850 32708 46927 32724
tri 46927 32708 46943 32724 nw
rect 46979 32691 47093 32925
tri 47129 32892 47145 32908 se
rect 47145 32892 47222 32908
rect 47129 32826 47222 32892
rect 47129 32724 47222 32790
tri 47129 32708 47145 32724 ne
rect 47145 32708 47222 32724
rect 46962 32609 47110 32691
rect 46850 32576 46927 32592
tri 46927 32576 46943 32592 sw
rect 46850 32510 46943 32576
rect 46979 32451 47093 32609
tri 47129 32576 47145 32592 se
rect 47145 32576 47222 32592
rect 47129 32510 47222 32576
rect 46850 32375 47222 32451
rect 46850 32250 46943 32316
rect 46850 32234 46927 32250
tri 46927 32234 46943 32250 nw
rect 46979 32217 47093 32375
rect 47129 32250 47222 32316
tri 47129 32234 47145 32250 ne
rect 47145 32234 47222 32250
rect 46962 32135 47110 32217
rect 46850 32102 46927 32118
tri 46927 32102 46943 32118 sw
rect 46850 32036 46943 32102
rect 46850 31934 46943 32000
rect 46850 31918 46927 31934
tri 46927 31918 46943 31934 nw
rect 46979 31901 47093 32135
tri 47129 32102 47145 32118 se
rect 47145 32102 47222 32118
rect 47129 32036 47222 32102
rect 47129 31934 47222 32000
tri 47129 31918 47145 31934 ne
rect 47145 31918 47222 31934
rect 46962 31819 47110 31901
rect 46850 31786 46927 31802
tri 46927 31786 46943 31802 sw
rect 46850 31720 46943 31786
rect 46979 31661 47093 31819
tri 47129 31786 47145 31802 se
rect 47145 31786 47222 31802
rect 47129 31720 47222 31786
rect 46850 31585 47222 31661
rect 46850 31460 46943 31526
rect 46850 31444 46927 31460
tri 46927 31444 46943 31460 nw
rect 46979 31427 47093 31585
rect 47129 31460 47222 31526
tri 47129 31444 47145 31460 ne
rect 47145 31444 47222 31460
rect 46962 31345 47110 31427
rect 46850 31312 46927 31328
tri 46927 31312 46943 31328 sw
rect 46850 31246 46943 31312
rect 46850 31144 46943 31210
rect 46850 31128 46927 31144
tri 46927 31128 46943 31144 nw
rect 46979 31111 47093 31345
tri 47129 31312 47145 31328 se
rect 47145 31312 47222 31328
rect 47129 31246 47222 31312
rect 47129 31144 47222 31210
tri 47129 31128 47145 31144 ne
rect 47145 31128 47222 31144
rect 46962 31029 47110 31111
rect 46850 30996 46927 31012
tri 46927 30996 46943 31012 sw
rect 46850 30930 46943 30996
rect 46979 30871 47093 31029
tri 47129 30996 47145 31012 se
rect 47145 30996 47222 31012
rect 47129 30930 47222 30996
rect 46850 30795 47222 30871
rect 46850 30670 46943 30736
rect 46850 30654 46927 30670
tri 46927 30654 46943 30670 nw
rect 46979 30637 47093 30795
rect 47129 30670 47222 30736
tri 47129 30654 47145 30670 ne
rect 47145 30654 47222 30670
rect 46962 30555 47110 30637
rect 46850 30522 46927 30538
tri 46927 30522 46943 30538 sw
rect 46850 30456 46943 30522
rect 46850 30354 46943 30420
rect 46850 30338 46927 30354
tri 46927 30338 46943 30354 nw
rect 46979 30321 47093 30555
tri 47129 30522 47145 30538 se
rect 47145 30522 47222 30538
rect 47129 30456 47222 30522
rect 47129 30354 47222 30420
tri 47129 30338 47145 30354 ne
rect 47145 30338 47222 30354
rect 46962 30239 47110 30321
rect 46850 30206 46927 30222
tri 46927 30206 46943 30222 sw
rect 46850 30140 46943 30206
rect 46979 30081 47093 30239
tri 47129 30206 47145 30222 se
rect 47145 30206 47222 30222
rect 47129 30140 47222 30206
rect 46850 30005 47222 30081
rect 46850 29880 46943 29946
rect 46850 29864 46927 29880
tri 46927 29864 46943 29880 nw
rect 46979 29847 47093 30005
rect 47129 29880 47222 29946
tri 47129 29864 47145 29880 ne
rect 47145 29864 47222 29880
rect 46962 29765 47110 29847
rect 46850 29732 46927 29748
tri 46927 29732 46943 29748 sw
rect 46850 29666 46943 29732
rect 46850 29564 46943 29630
rect 46850 29548 46927 29564
tri 46927 29548 46943 29564 nw
rect 46979 29531 47093 29765
tri 47129 29732 47145 29748 se
rect 47145 29732 47222 29748
rect 47129 29666 47222 29732
rect 47129 29564 47222 29630
tri 47129 29548 47145 29564 ne
rect 47145 29548 47222 29564
rect 46962 29449 47110 29531
rect 46850 29416 46927 29432
tri 46927 29416 46943 29432 sw
rect 46850 29350 46943 29416
rect 46979 29291 47093 29449
tri 47129 29416 47145 29432 se
rect 47145 29416 47222 29432
rect 47129 29350 47222 29416
rect 46850 29215 47222 29291
rect 46850 29090 46943 29156
rect 46850 29074 46927 29090
tri 46927 29074 46943 29090 nw
rect 46979 29057 47093 29215
rect 47129 29090 47222 29156
tri 47129 29074 47145 29090 ne
rect 47145 29074 47222 29090
rect 46962 28975 47110 29057
rect 46850 28942 46927 28958
tri 46927 28942 46943 28958 sw
rect 46850 28876 46943 28942
rect 46979 28833 47093 28975
tri 47129 28942 47145 28958 se
rect 47145 28942 47222 28958
rect 47129 28876 47222 28942
rect 47258 28463 47294 80603
rect 47330 28463 47366 80603
rect 47402 80445 47438 80603
rect 47394 80303 47446 80445
rect 47402 28763 47438 80303
rect 47394 28621 47446 28763
rect 47402 28463 47438 28621
rect 47474 28463 47510 80603
rect 47546 28463 47582 80603
rect 47618 28833 47702 80233
rect 47738 28463 47774 80603
rect 47810 28463 47846 80603
rect 47882 80445 47918 80603
rect 47874 80303 47926 80445
rect 47882 28763 47918 80303
rect 47874 28621 47926 28763
rect 47882 28463 47918 28621
rect 47954 28463 47990 80603
rect 48026 28463 48062 80603
rect 48098 80124 48191 80190
rect 48098 80108 48175 80124
tri 48175 80108 48191 80124 nw
rect 48227 80091 48341 80233
rect 48377 80124 48470 80190
tri 48377 80108 48393 80124 ne
rect 48393 80108 48470 80124
rect 48210 80009 48358 80091
rect 48098 79976 48175 79992
tri 48175 79976 48191 79992 sw
rect 48098 79910 48191 79976
rect 48227 79851 48341 80009
tri 48377 79976 48393 79992 se
rect 48393 79976 48470 79992
rect 48377 79910 48470 79976
rect 48098 79775 48470 79851
rect 48098 79650 48191 79716
rect 48098 79634 48175 79650
tri 48175 79634 48191 79650 nw
rect 48227 79617 48341 79775
rect 48377 79650 48470 79716
tri 48377 79634 48393 79650 ne
rect 48393 79634 48470 79650
rect 48210 79535 48358 79617
rect 48098 79502 48175 79518
tri 48175 79502 48191 79518 sw
rect 48098 79436 48191 79502
rect 48098 79334 48191 79400
rect 48098 79318 48175 79334
tri 48175 79318 48191 79334 nw
rect 48227 79301 48341 79535
tri 48377 79502 48393 79518 se
rect 48393 79502 48470 79518
rect 48377 79436 48470 79502
rect 48377 79334 48470 79400
tri 48377 79318 48393 79334 ne
rect 48393 79318 48470 79334
rect 48210 79219 48358 79301
rect 48098 79186 48175 79202
tri 48175 79186 48191 79202 sw
rect 48098 79120 48191 79186
rect 48227 79061 48341 79219
tri 48377 79186 48393 79202 se
rect 48393 79186 48470 79202
rect 48377 79120 48470 79186
rect 48098 78985 48470 79061
rect 48098 78860 48191 78926
rect 48098 78844 48175 78860
tri 48175 78844 48191 78860 nw
rect 48227 78827 48341 78985
rect 48377 78860 48470 78926
tri 48377 78844 48393 78860 ne
rect 48393 78844 48470 78860
rect 48210 78745 48358 78827
rect 48098 78712 48175 78728
tri 48175 78712 48191 78728 sw
rect 48098 78646 48191 78712
rect 48098 78544 48191 78610
rect 48098 78528 48175 78544
tri 48175 78528 48191 78544 nw
rect 48227 78511 48341 78745
tri 48377 78712 48393 78728 se
rect 48393 78712 48470 78728
rect 48377 78646 48470 78712
rect 48377 78544 48470 78610
tri 48377 78528 48393 78544 ne
rect 48393 78528 48470 78544
rect 48210 78429 48358 78511
rect 48098 78396 48175 78412
tri 48175 78396 48191 78412 sw
rect 48098 78330 48191 78396
rect 48227 78271 48341 78429
tri 48377 78396 48393 78412 se
rect 48393 78396 48470 78412
rect 48377 78330 48470 78396
rect 48098 78195 48470 78271
rect 48098 78070 48191 78136
rect 48098 78054 48175 78070
tri 48175 78054 48191 78070 nw
rect 48227 78037 48341 78195
rect 48377 78070 48470 78136
tri 48377 78054 48393 78070 ne
rect 48393 78054 48470 78070
rect 48210 77955 48358 78037
rect 48098 77922 48175 77938
tri 48175 77922 48191 77938 sw
rect 48098 77856 48191 77922
rect 48098 77754 48191 77820
rect 48098 77738 48175 77754
tri 48175 77738 48191 77754 nw
rect 48227 77721 48341 77955
tri 48377 77922 48393 77938 se
rect 48393 77922 48470 77938
rect 48377 77856 48470 77922
rect 48377 77754 48470 77820
tri 48377 77738 48393 77754 ne
rect 48393 77738 48470 77754
rect 48210 77639 48358 77721
rect 48098 77606 48175 77622
tri 48175 77606 48191 77622 sw
rect 48098 77540 48191 77606
rect 48227 77481 48341 77639
tri 48377 77606 48393 77622 se
rect 48393 77606 48470 77622
rect 48377 77540 48470 77606
rect 48098 77405 48470 77481
rect 48098 77280 48191 77346
rect 48098 77264 48175 77280
tri 48175 77264 48191 77280 nw
rect 48227 77247 48341 77405
rect 48377 77280 48470 77346
tri 48377 77264 48393 77280 ne
rect 48393 77264 48470 77280
rect 48210 77165 48358 77247
rect 48098 77132 48175 77148
tri 48175 77132 48191 77148 sw
rect 48098 77066 48191 77132
rect 48098 76964 48191 77030
rect 48098 76948 48175 76964
tri 48175 76948 48191 76964 nw
rect 48227 76931 48341 77165
tri 48377 77132 48393 77148 se
rect 48393 77132 48470 77148
rect 48377 77066 48470 77132
rect 48377 76964 48470 77030
tri 48377 76948 48393 76964 ne
rect 48393 76948 48470 76964
rect 48210 76849 48358 76931
rect 48098 76816 48175 76832
tri 48175 76816 48191 76832 sw
rect 48098 76750 48191 76816
rect 48227 76691 48341 76849
tri 48377 76816 48393 76832 se
rect 48393 76816 48470 76832
rect 48377 76750 48470 76816
rect 48098 76615 48470 76691
rect 48098 76490 48191 76556
rect 48098 76474 48175 76490
tri 48175 76474 48191 76490 nw
rect 48227 76457 48341 76615
rect 48377 76490 48470 76556
tri 48377 76474 48393 76490 ne
rect 48393 76474 48470 76490
rect 48210 76375 48358 76457
rect 48098 76342 48175 76358
tri 48175 76342 48191 76358 sw
rect 48098 76276 48191 76342
rect 48098 76174 48191 76240
rect 48098 76158 48175 76174
tri 48175 76158 48191 76174 nw
rect 48227 76141 48341 76375
tri 48377 76342 48393 76358 se
rect 48393 76342 48470 76358
rect 48377 76276 48470 76342
rect 48377 76174 48470 76240
tri 48377 76158 48393 76174 ne
rect 48393 76158 48470 76174
rect 48210 76059 48358 76141
rect 48098 76026 48175 76042
tri 48175 76026 48191 76042 sw
rect 48098 75960 48191 76026
rect 48227 75901 48341 76059
tri 48377 76026 48393 76042 se
rect 48393 76026 48470 76042
rect 48377 75960 48470 76026
rect 48098 75825 48470 75901
rect 48098 75700 48191 75766
rect 48098 75684 48175 75700
tri 48175 75684 48191 75700 nw
rect 48227 75667 48341 75825
rect 48377 75700 48470 75766
tri 48377 75684 48393 75700 ne
rect 48393 75684 48470 75700
rect 48210 75585 48358 75667
rect 48098 75552 48175 75568
tri 48175 75552 48191 75568 sw
rect 48098 75486 48191 75552
rect 48098 75384 48191 75450
rect 48098 75368 48175 75384
tri 48175 75368 48191 75384 nw
rect 48227 75351 48341 75585
tri 48377 75552 48393 75568 se
rect 48393 75552 48470 75568
rect 48377 75486 48470 75552
rect 48377 75384 48470 75450
tri 48377 75368 48393 75384 ne
rect 48393 75368 48470 75384
rect 48210 75269 48358 75351
rect 48098 75236 48175 75252
tri 48175 75236 48191 75252 sw
rect 48098 75170 48191 75236
rect 48227 75111 48341 75269
tri 48377 75236 48393 75252 se
rect 48393 75236 48470 75252
rect 48377 75170 48470 75236
rect 48098 75035 48470 75111
rect 48098 74910 48191 74976
rect 48098 74894 48175 74910
tri 48175 74894 48191 74910 nw
rect 48227 74877 48341 75035
rect 48377 74910 48470 74976
tri 48377 74894 48393 74910 ne
rect 48393 74894 48470 74910
rect 48210 74795 48358 74877
rect 48098 74762 48175 74778
tri 48175 74762 48191 74778 sw
rect 48098 74696 48191 74762
rect 48098 74594 48191 74660
rect 48098 74578 48175 74594
tri 48175 74578 48191 74594 nw
rect 48227 74561 48341 74795
tri 48377 74762 48393 74778 se
rect 48393 74762 48470 74778
rect 48377 74696 48470 74762
rect 48377 74594 48470 74660
tri 48377 74578 48393 74594 ne
rect 48393 74578 48470 74594
rect 48210 74479 48358 74561
rect 48098 74446 48175 74462
tri 48175 74446 48191 74462 sw
rect 48098 74380 48191 74446
rect 48227 74321 48341 74479
tri 48377 74446 48393 74462 se
rect 48393 74446 48470 74462
rect 48377 74380 48470 74446
rect 48098 74245 48470 74321
rect 48098 74120 48191 74186
rect 48098 74104 48175 74120
tri 48175 74104 48191 74120 nw
rect 48227 74087 48341 74245
rect 48377 74120 48470 74186
tri 48377 74104 48393 74120 ne
rect 48393 74104 48470 74120
rect 48210 74005 48358 74087
rect 48098 73972 48175 73988
tri 48175 73972 48191 73988 sw
rect 48098 73906 48191 73972
rect 48098 73804 48191 73870
rect 48098 73788 48175 73804
tri 48175 73788 48191 73804 nw
rect 48227 73771 48341 74005
tri 48377 73972 48393 73988 se
rect 48393 73972 48470 73988
rect 48377 73906 48470 73972
rect 48377 73804 48470 73870
tri 48377 73788 48393 73804 ne
rect 48393 73788 48470 73804
rect 48210 73689 48358 73771
rect 48098 73656 48175 73672
tri 48175 73656 48191 73672 sw
rect 48098 73590 48191 73656
rect 48227 73531 48341 73689
tri 48377 73656 48393 73672 se
rect 48393 73656 48470 73672
rect 48377 73590 48470 73656
rect 48098 73455 48470 73531
rect 48098 73330 48191 73396
rect 48098 73314 48175 73330
tri 48175 73314 48191 73330 nw
rect 48227 73297 48341 73455
rect 48377 73330 48470 73396
tri 48377 73314 48393 73330 ne
rect 48393 73314 48470 73330
rect 48210 73215 48358 73297
rect 48098 73182 48175 73198
tri 48175 73182 48191 73198 sw
rect 48098 73116 48191 73182
rect 48098 73014 48191 73080
rect 48098 72998 48175 73014
tri 48175 72998 48191 73014 nw
rect 48227 72981 48341 73215
tri 48377 73182 48393 73198 se
rect 48393 73182 48470 73198
rect 48377 73116 48470 73182
rect 48377 73014 48470 73080
tri 48377 72998 48393 73014 ne
rect 48393 72998 48470 73014
rect 48210 72899 48358 72981
rect 48098 72866 48175 72882
tri 48175 72866 48191 72882 sw
rect 48098 72800 48191 72866
rect 48227 72741 48341 72899
tri 48377 72866 48393 72882 se
rect 48393 72866 48470 72882
rect 48377 72800 48470 72866
rect 48098 72665 48470 72741
rect 48098 72540 48191 72606
rect 48098 72524 48175 72540
tri 48175 72524 48191 72540 nw
rect 48227 72507 48341 72665
rect 48377 72540 48470 72606
tri 48377 72524 48393 72540 ne
rect 48393 72524 48470 72540
rect 48210 72425 48358 72507
rect 48098 72392 48175 72408
tri 48175 72392 48191 72408 sw
rect 48098 72326 48191 72392
rect 48098 72224 48191 72290
rect 48098 72208 48175 72224
tri 48175 72208 48191 72224 nw
rect 48227 72191 48341 72425
tri 48377 72392 48393 72408 se
rect 48393 72392 48470 72408
rect 48377 72326 48470 72392
rect 48377 72224 48470 72290
tri 48377 72208 48393 72224 ne
rect 48393 72208 48470 72224
rect 48210 72109 48358 72191
rect 48098 72076 48175 72092
tri 48175 72076 48191 72092 sw
rect 48098 72010 48191 72076
rect 48227 71951 48341 72109
tri 48377 72076 48393 72092 se
rect 48393 72076 48470 72092
rect 48377 72010 48470 72076
rect 48098 71875 48470 71951
rect 48098 71750 48191 71816
rect 48098 71734 48175 71750
tri 48175 71734 48191 71750 nw
rect 48227 71717 48341 71875
rect 48377 71750 48470 71816
tri 48377 71734 48393 71750 ne
rect 48393 71734 48470 71750
rect 48210 71635 48358 71717
rect 48098 71602 48175 71618
tri 48175 71602 48191 71618 sw
rect 48098 71536 48191 71602
rect 48098 71434 48191 71500
rect 48098 71418 48175 71434
tri 48175 71418 48191 71434 nw
rect 48227 71401 48341 71635
tri 48377 71602 48393 71618 se
rect 48393 71602 48470 71618
rect 48377 71536 48470 71602
rect 48377 71434 48470 71500
tri 48377 71418 48393 71434 ne
rect 48393 71418 48470 71434
rect 48210 71319 48358 71401
rect 48098 71286 48175 71302
tri 48175 71286 48191 71302 sw
rect 48098 71220 48191 71286
rect 48227 71161 48341 71319
tri 48377 71286 48393 71302 se
rect 48393 71286 48470 71302
rect 48377 71220 48470 71286
rect 48098 71085 48470 71161
rect 48098 70960 48191 71026
rect 48098 70944 48175 70960
tri 48175 70944 48191 70960 nw
rect 48227 70927 48341 71085
rect 48377 70960 48470 71026
tri 48377 70944 48393 70960 ne
rect 48393 70944 48470 70960
rect 48210 70845 48358 70927
rect 48098 70812 48175 70828
tri 48175 70812 48191 70828 sw
rect 48098 70746 48191 70812
rect 48098 70644 48191 70710
rect 48098 70628 48175 70644
tri 48175 70628 48191 70644 nw
rect 48227 70611 48341 70845
tri 48377 70812 48393 70828 se
rect 48393 70812 48470 70828
rect 48377 70746 48470 70812
rect 48377 70644 48470 70710
tri 48377 70628 48393 70644 ne
rect 48393 70628 48470 70644
rect 48210 70529 48358 70611
rect 48098 70496 48175 70512
tri 48175 70496 48191 70512 sw
rect 48098 70430 48191 70496
rect 48227 70371 48341 70529
tri 48377 70496 48393 70512 se
rect 48393 70496 48470 70512
rect 48377 70430 48470 70496
rect 48098 70295 48470 70371
rect 48098 70170 48191 70236
rect 48098 70154 48175 70170
tri 48175 70154 48191 70170 nw
rect 48227 70137 48341 70295
rect 48377 70170 48470 70236
tri 48377 70154 48393 70170 ne
rect 48393 70154 48470 70170
rect 48210 70055 48358 70137
rect 48098 70022 48175 70038
tri 48175 70022 48191 70038 sw
rect 48098 69956 48191 70022
rect 48098 69854 48191 69920
rect 48098 69838 48175 69854
tri 48175 69838 48191 69854 nw
rect 48227 69821 48341 70055
tri 48377 70022 48393 70038 se
rect 48393 70022 48470 70038
rect 48377 69956 48470 70022
rect 48377 69854 48470 69920
tri 48377 69838 48393 69854 ne
rect 48393 69838 48470 69854
rect 48210 69739 48358 69821
rect 48098 69706 48175 69722
tri 48175 69706 48191 69722 sw
rect 48098 69640 48191 69706
rect 48227 69581 48341 69739
tri 48377 69706 48393 69722 se
rect 48393 69706 48470 69722
rect 48377 69640 48470 69706
rect 48098 69505 48470 69581
rect 48098 69380 48191 69446
rect 48098 69364 48175 69380
tri 48175 69364 48191 69380 nw
rect 48227 69347 48341 69505
rect 48377 69380 48470 69446
tri 48377 69364 48393 69380 ne
rect 48393 69364 48470 69380
rect 48210 69265 48358 69347
rect 48098 69232 48175 69248
tri 48175 69232 48191 69248 sw
rect 48098 69166 48191 69232
rect 48098 69064 48191 69130
rect 48098 69048 48175 69064
tri 48175 69048 48191 69064 nw
rect 48227 69031 48341 69265
tri 48377 69232 48393 69248 se
rect 48393 69232 48470 69248
rect 48377 69166 48470 69232
rect 48377 69064 48470 69130
tri 48377 69048 48393 69064 ne
rect 48393 69048 48470 69064
rect 48210 68949 48358 69031
rect 48098 68916 48175 68932
tri 48175 68916 48191 68932 sw
rect 48098 68850 48191 68916
rect 48227 68791 48341 68949
tri 48377 68916 48393 68932 se
rect 48393 68916 48470 68932
rect 48377 68850 48470 68916
rect 48098 68715 48470 68791
rect 48098 68590 48191 68656
rect 48098 68574 48175 68590
tri 48175 68574 48191 68590 nw
rect 48227 68557 48341 68715
rect 48377 68590 48470 68656
tri 48377 68574 48393 68590 ne
rect 48393 68574 48470 68590
rect 48210 68475 48358 68557
rect 48098 68442 48175 68458
tri 48175 68442 48191 68458 sw
rect 48098 68376 48191 68442
rect 48098 68274 48191 68340
rect 48098 68258 48175 68274
tri 48175 68258 48191 68274 nw
rect 48227 68241 48341 68475
tri 48377 68442 48393 68458 se
rect 48393 68442 48470 68458
rect 48377 68376 48470 68442
rect 48377 68274 48470 68340
tri 48377 68258 48393 68274 ne
rect 48393 68258 48470 68274
rect 48210 68159 48358 68241
rect 48098 68126 48175 68142
tri 48175 68126 48191 68142 sw
rect 48098 68060 48191 68126
rect 48227 68001 48341 68159
tri 48377 68126 48393 68142 se
rect 48393 68126 48470 68142
rect 48377 68060 48470 68126
rect 48098 67925 48470 68001
rect 48098 67800 48191 67866
rect 48098 67784 48175 67800
tri 48175 67784 48191 67800 nw
rect 48227 67767 48341 67925
rect 48377 67800 48470 67866
tri 48377 67784 48393 67800 ne
rect 48393 67784 48470 67800
rect 48210 67685 48358 67767
rect 48098 67652 48175 67668
tri 48175 67652 48191 67668 sw
rect 48098 67586 48191 67652
rect 48098 67484 48191 67550
rect 48098 67468 48175 67484
tri 48175 67468 48191 67484 nw
rect 48227 67451 48341 67685
tri 48377 67652 48393 67668 se
rect 48393 67652 48470 67668
rect 48377 67586 48470 67652
rect 48377 67484 48470 67550
tri 48377 67468 48393 67484 ne
rect 48393 67468 48470 67484
rect 48210 67369 48358 67451
rect 48098 67336 48175 67352
tri 48175 67336 48191 67352 sw
rect 48098 67270 48191 67336
rect 48227 67211 48341 67369
tri 48377 67336 48393 67352 se
rect 48393 67336 48470 67352
rect 48377 67270 48470 67336
rect 48098 67135 48470 67211
rect 48098 67010 48191 67076
rect 48098 66994 48175 67010
tri 48175 66994 48191 67010 nw
rect 48227 66977 48341 67135
rect 48377 67010 48470 67076
tri 48377 66994 48393 67010 ne
rect 48393 66994 48470 67010
rect 48210 66895 48358 66977
rect 48098 66862 48175 66878
tri 48175 66862 48191 66878 sw
rect 48098 66796 48191 66862
rect 48098 66694 48191 66760
rect 48098 66678 48175 66694
tri 48175 66678 48191 66694 nw
rect 48227 66661 48341 66895
tri 48377 66862 48393 66878 se
rect 48393 66862 48470 66878
rect 48377 66796 48470 66862
rect 48377 66694 48470 66760
tri 48377 66678 48393 66694 ne
rect 48393 66678 48470 66694
rect 48210 66579 48358 66661
rect 48098 66546 48175 66562
tri 48175 66546 48191 66562 sw
rect 48098 66480 48191 66546
rect 48227 66421 48341 66579
tri 48377 66546 48393 66562 se
rect 48393 66546 48470 66562
rect 48377 66480 48470 66546
rect 48098 66345 48470 66421
rect 48098 66220 48191 66286
rect 48098 66204 48175 66220
tri 48175 66204 48191 66220 nw
rect 48227 66187 48341 66345
rect 48377 66220 48470 66286
tri 48377 66204 48393 66220 ne
rect 48393 66204 48470 66220
rect 48210 66105 48358 66187
rect 48098 66072 48175 66088
tri 48175 66072 48191 66088 sw
rect 48098 66006 48191 66072
rect 48098 65904 48191 65970
rect 48098 65888 48175 65904
tri 48175 65888 48191 65904 nw
rect 48227 65871 48341 66105
tri 48377 66072 48393 66088 se
rect 48393 66072 48470 66088
rect 48377 66006 48470 66072
rect 48377 65904 48470 65970
tri 48377 65888 48393 65904 ne
rect 48393 65888 48470 65904
rect 48210 65789 48358 65871
rect 48098 65756 48175 65772
tri 48175 65756 48191 65772 sw
rect 48098 65690 48191 65756
rect 48227 65631 48341 65789
tri 48377 65756 48393 65772 se
rect 48393 65756 48470 65772
rect 48377 65690 48470 65756
rect 48098 65555 48470 65631
rect 48098 65430 48191 65496
rect 48098 65414 48175 65430
tri 48175 65414 48191 65430 nw
rect 48227 65397 48341 65555
rect 48377 65430 48470 65496
tri 48377 65414 48393 65430 ne
rect 48393 65414 48470 65430
rect 48210 65315 48358 65397
rect 48098 65282 48175 65298
tri 48175 65282 48191 65298 sw
rect 48098 65216 48191 65282
rect 48098 65114 48191 65180
rect 48098 65098 48175 65114
tri 48175 65098 48191 65114 nw
rect 48227 65081 48341 65315
tri 48377 65282 48393 65298 se
rect 48393 65282 48470 65298
rect 48377 65216 48470 65282
rect 48377 65114 48470 65180
tri 48377 65098 48393 65114 ne
rect 48393 65098 48470 65114
rect 48210 64999 48358 65081
rect 48098 64966 48175 64982
tri 48175 64966 48191 64982 sw
rect 48098 64900 48191 64966
rect 48227 64841 48341 64999
tri 48377 64966 48393 64982 se
rect 48393 64966 48470 64982
rect 48377 64900 48470 64966
rect 48098 64765 48470 64841
rect 48098 64640 48191 64706
rect 48098 64624 48175 64640
tri 48175 64624 48191 64640 nw
rect 48227 64607 48341 64765
rect 48377 64640 48470 64706
tri 48377 64624 48393 64640 ne
rect 48393 64624 48470 64640
rect 48210 64525 48358 64607
rect 48098 64492 48175 64508
tri 48175 64492 48191 64508 sw
rect 48098 64426 48191 64492
rect 48098 64324 48191 64390
rect 48098 64308 48175 64324
tri 48175 64308 48191 64324 nw
rect 48227 64291 48341 64525
tri 48377 64492 48393 64508 se
rect 48393 64492 48470 64508
rect 48377 64426 48470 64492
rect 48377 64324 48470 64390
tri 48377 64308 48393 64324 ne
rect 48393 64308 48470 64324
rect 48210 64209 48358 64291
rect 48098 64176 48175 64192
tri 48175 64176 48191 64192 sw
rect 48098 64110 48191 64176
rect 48227 64051 48341 64209
tri 48377 64176 48393 64192 se
rect 48393 64176 48470 64192
rect 48377 64110 48470 64176
rect 48098 63975 48470 64051
rect 48098 63850 48191 63916
rect 48098 63834 48175 63850
tri 48175 63834 48191 63850 nw
rect 48227 63817 48341 63975
rect 48377 63850 48470 63916
tri 48377 63834 48393 63850 ne
rect 48393 63834 48470 63850
rect 48210 63735 48358 63817
rect 48098 63702 48175 63718
tri 48175 63702 48191 63718 sw
rect 48098 63636 48191 63702
rect 48098 63534 48191 63600
rect 48098 63518 48175 63534
tri 48175 63518 48191 63534 nw
rect 48227 63501 48341 63735
tri 48377 63702 48393 63718 se
rect 48393 63702 48470 63718
rect 48377 63636 48470 63702
rect 48377 63534 48470 63600
tri 48377 63518 48393 63534 ne
rect 48393 63518 48470 63534
rect 48210 63419 48358 63501
rect 48098 63386 48175 63402
tri 48175 63386 48191 63402 sw
rect 48098 63320 48191 63386
rect 48227 63261 48341 63419
tri 48377 63386 48393 63402 se
rect 48393 63386 48470 63402
rect 48377 63320 48470 63386
rect 48098 63185 48470 63261
rect 48098 63060 48191 63126
rect 48098 63044 48175 63060
tri 48175 63044 48191 63060 nw
rect 48227 63027 48341 63185
rect 48377 63060 48470 63126
tri 48377 63044 48393 63060 ne
rect 48393 63044 48470 63060
rect 48210 62945 48358 63027
rect 48098 62912 48175 62928
tri 48175 62912 48191 62928 sw
rect 48098 62846 48191 62912
rect 48098 62744 48191 62810
rect 48098 62728 48175 62744
tri 48175 62728 48191 62744 nw
rect 48227 62711 48341 62945
tri 48377 62912 48393 62928 se
rect 48393 62912 48470 62928
rect 48377 62846 48470 62912
rect 48377 62744 48470 62810
tri 48377 62728 48393 62744 ne
rect 48393 62728 48470 62744
rect 48210 62629 48358 62711
rect 48098 62596 48175 62612
tri 48175 62596 48191 62612 sw
rect 48098 62530 48191 62596
rect 48227 62471 48341 62629
tri 48377 62596 48393 62612 se
rect 48393 62596 48470 62612
rect 48377 62530 48470 62596
rect 48098 62395 48470 62471
rect 48098 62270 48191 62336
rect 48098 62254 48175 62270
tri 48175 62254 48191 62270 nw
rect 48227 62237 48341 62395
rect 48377 62270 48470 62336
tri 48377 62254 48393 62270 ne
rect 48393 62254 48470 62270
rect 48210 62155 48358 62237
rect 48098 62122 48175 62138
tri 48175 62122 48191 62138 sw
rect 48098 62056 48191 62122
rect 48098 61954 48191 62020
rect 48098 61938 48175 61954
tri 48175 61938 48191 61954 nw
rect 48227 61921 48341 62155
tri 48377 62122 48393 62138 se
rect 48393 62122 48470 62138
rect 48377 62056 48470 62122
rect 48377 61954 48470 62020
tri 48377 61938 48393 61954 ne
rect 48393 61938 48470 61954
rect 48210 61839 48358 61921
rect 48098 61806 48175 61822
tri 48175 61806 48191 61822 sw
rect 48098 61740 48191 61806
rect 48227 61681 48341 61839
tri 48377 61806 48393 61822 se
rect 48393 61806 48470 61822
rect 48377 61740 48470 61806
rect 48098 61605 48470 61681
rect 48098 61480 48191 61546
rect 48098 61464 48175 61480
tri 48175 61464 48191 61480 nw
rect 48227 61447 48341 61605
rect 48377 61480 48470 61546
tri 48377 61464 48393 61480 ne
rect 48393 61464 48470 61480
rect 48210 61365 48358 61447
rect 48098 61332 48175 61348
tri 48175 61332 48191 61348 sw
rect 48098 61266 48191 61332
rect 48098 61164 48191 61230
rect 48098 61148 48175 61164
tri 48175 61148 48191 61164 nw
rect 48227 61131 48341 61365
tri 48377 61332 48393 61348 se
rect 48393 61332 48470 61348
rect 48377 61266 48470 61332
rect 48377 61164 48470 61230
tri 48377 61148 48393 61164 ne
rect 48393 61148 48470 61164
rect 48210 61049 48358 61131
rect 48098 61016 48175 61032
tri 48175 61016 48191 61032 sw
rect 48098 60950 48191 61016
rect 48227 60891 48341 61049
tri 48377 61016 48393 61032 se
rect 48393 61016 48470 61032
rect 48377 60950 48470 61016
rect 48098 60815 48470 60891
rect 48098 60690 48191 60756
rect 48098 60674 48175 60690
tri 48175 60674 48191 60690 nw
rect 48227 60657 48341 60815
rect 48377 60690 48470 60756
tri 48377 60674 48393 60690 ne
rect 48393 60674 48470 60690
rect 48210 60575 48358 60657
rect 48098 60542 48175 60558
tri 48175 60542 48191 60558 sw
rect 48098 60476 48191 60542
rect 48098 60374 48191 60440
rect 48098 60358 48175 60374
tri 48175 60358 48191 60374 nw
rect 48227 60341 48341 60575
tri 48377 60542 48393 60558 se
rect 48393 60542 48470 60558
rect 48377 60476 48470 60542
rect 48377 60374 48470 60440
tri 48377 60358 48393 60374 ne
rect 48393 60358 48470 60374
rect 48210 60259 48358 60341
rect 48098 60226 48175 60242
tri 48175 60226 48191 60242 sw
rect 48098 60160 48191 60226
rect 48227 60101 48341 60259
tri 48377 60226 48393 60242 se
rect 48393 60226 48470 60242
rect 48377 60160 48470 60226
rect 48098 60025 48470 60101
rect 48098 59900 48191 59966
rect 48098 59884 48175 59900
tri 48175 59884 48191 59900 nw
rect 48227 59867 48341 60025
rect 48377 59900 48470 59966
tri 48377 59884 48393 59900 ne
rect 48393 59884 48470 59900
rect 48210 59785 48358 59867
rect 48098 59752 48175 59768
tri 48175 59752 48191 59768 sw
rect 48098 59686 48191 59752
rect 48098 59584 48191 59650
rect 48098 59568 48175 59584
tri 48175 59568 48191 59584 nw
rect 48227 59551 48341 59785
tri 48377 59752 48393 59768 se
rect 48393 59752 48470 59768
rect 48377 59686 48470 59752
rect 48377 59584 48470 59650
tri 48377 59568 48393 59584 ne
rect 48393 59568 48470 59584
rect 48210 59469 48358 59551
rect 48098 59436 48175 59452
tri 48175 59436 48191 59452 sw
rect 48098 59370 48191 59436
rect 48227 59311 48341 59469
tri 48377 59436 48393 59452 se
rect 48393 59436 48470 59452
rect 48377 59370 48470 59436
rect 48098 59235 48470 59311
rect 48098 59110 48191 59176
rect 48098 59094 48175 59110
tri 48175 59094 48191 59110 nw
rect 48227 59077 48341 59235
rect 48377 59110 48470 59176
tri 48377 59094 48393 59110 ne
rect 48393 59094 48470 59110
rect 48210 58995 48358 59077
rect 48098 58962 48175 58978
tri 48175 58962 48191 58978 sw
rect 48098 58896 48191 58962
rect 48098 58794 48191 58860
rect 48098 58778 48175 58794
tri 48175 58778 48191 58794 nw
rect 48227 58761 48341 58995
tri 48377 58962 48393 58978 se
rect 48393 58962 48470 58978
rect 48377 58896 48470 58962
rect 48377 58794 48470 58860
tri 48377 58778 48393 58794 ne
rect 48393 58778 48470 58794
rect 48210 58679 48358 58761
rect 48098 58646 48175 58662
tri 48175 58646 48191 58662 sw
rect 48098 58580 48191 58646
rect 48227 58521 48341 58679
tri 48377 58646 48393 58662 se
rect 48393 58646 48470 58662
rect 48377 58580 48470 58646
rect 48098 58445 48470 58521
rect 48098 58320 48191 58386
rect 48098 58304 48175 58320
tri 48175 58304 48191 58320 nw
rect 48227 58287 48341 58445
rect 48377 58320 48470 58386
tri 48377 58304 48393 58320 ne
rect 48393 58304 48470 58320
rect 48210 58205 48358 58287
rect 48098 58172 48175 58188
tri 48175 58172 48191 58188 sw
rect 48098 58106 48191 58172
rect 48098 58004 48191 58070
rect 48098 57988 48175 58004
tri 48175 57988 48191 58004 nw
rect 48227 57971 48341 58205
tri 48377 58172 48393 58188 se
rect 48393 58172 48470 58188
rect 48377 58106 48470 58172
rect 48377 58004 48470 58070
tri 48377 57988 48393 58004 ne
rect 48393 57988 48470 58004
rect 48210 57889 48358 57971
rect 48098 57856 48175 57872
tri 48175 57856 48191 57872 sw
rect 48098 57790 48191 57856
rect 48227 57731 48341 57889
tri 48377 57856 48393 57872 se
rect 48393 57856 48470 57872
rect 48377 57790 48470 57856
rect 48098 57655 48470 57731
rect 48098 57530 48191 57596
rect 48098 57514 48175 57530
tri 48175 57514 48191 57530 nw
rect 48227 57497 48341 57655
rect 48377 57530 48470 57596
tri 48377 57514 48393 57530 ne
rect 48393 57514 48470 57530
rect 48210 57415 48358 57497
rect 48098 57382 48175 57398
tri 48175 57382 48191 57398 sw
rect 48098 57316 48191 57382
rect 48098 57214 48191 57280
rect 48098 57198 48175 57214
tri 48175 57198 48191 57214 nw
rect 48227 57181 48341 57415
tri 48377 57382 48393 57398 se
rect 48393 57382 48470 57398
rect 48377 57316 48470 57382
rect 48377 57214 48470 57280
tri 48377 57198 48393 57214 ne
rect 48393 57198 48470 57214
rect 48210 57099 48358 57181
rect 48098 57066 48175 57082
tri 48175 57066 48191 57082 sw
rect 48098 57000 48191 57066
rect 48227 56941 48341 57099
tri 48377 57066 48393 57082 se
rect 48393 57066 48470 57082
rect 48377 57000 48470 57066
rect 48098 56865 48470 56941
rect 48098 56740 48191 56806
rect 48098 56724 48175 56740
tri 48175 56724 48191 56740 nw
rect 48227 56707 48341 56865
rect 48377 56740 48470 56806
tri 48377 56724 48393 56740 ne
rect 48393 56724 48470 56740
rect 48210 56625 48358 56707
rect 48098 56592 48175 56608
tri 48175 56592 48191 56608 sw
rect 48098 56526 48191 56592
rect 48098 56424 48191 56490
rect 48098 56408 48175 56424
tri 48175 56408 48191 56424 nw
rect 48227 56391 48341 56625
tri 48377 56592 48393 56608 se
rect 48393 56592 48470 56608
rect 48377 56526 48470 56592
rect 48377 56424 48470 56490
tri 48377 56408 48393 56424 ne
rect 48393 56408 48470 56424
rect 48210 56309 48358 56391
rect 48098 56276 48175 56292
tri 48175 56276 48191 56292 sw
rect 48098 56210 48191 56276
rect 48227 56151 48341 56309
tri 48377 56276 48393 56292 se
rect 48393 56276 48470 56292
rect 48377 56210 48470 56276
rect 48098 56075 48470 56151
rect 48098 55950 48191 56016
rect 48098 55934 48175 55950
tri 48175 55934 48191 55950 nw
rect 48227 55917 48341 56075
rect 48377 55950 48470 56016
tri 48377 55934 48393 55950 ne
rect 48393 55934 48470 55950
rect 48210 55835 48358 55917
rect 48098 55802 48175 55818
tri 48175 55802 48191 55818 sw
rect 48098 55736 48191 55802
rect 48098 55634 48191 55700
rect 48098 55618 48175 55634
tri 48175 55618 48191 55634 nw
rect 48227 55601 48341 55835
tri 48377 55802 48393 55818 se
rect 48393 55802 48470 55818
rect 48377 55736 48470 55802
rect 48377 55634 48470 55700
tri 48377 55618 48393 55634 ne
rect 48393 55618 48470 55634
rect 48210 55519 48358 55601
rect 48098 55486 48175 55502
tri 48175 55486 48191 55502 sw
rect 48098 55420 48191 55486
rect 48227 55361 48341 55519
tri 48377 55486 48393 55502 se
rect 48393 55486 48470 55502
rect 48377 55420 48470 55486
rect 48098 55285 48470 55361
rect 48098 55160 48191 55226
rect 48098 55144 48175 55160
tri 48175 55144 48191 55160 nw
rect 48227 55127 48341 55285
rect 48377 55160 48470 55226
tri 48377 55144 48393 55160 ne
rect 48393 55144 48470 55160
rect 48210 55045 48358 55127
rect 48098 55012 48175 55028
tri 48175 55012 48191 55028 sw
rect 48098 54946 48191 55012
rect 48098 54844 48191 54910
rect 48098 54828 48175 54844
tri 48175 54828 48191 54844 nw
rect 48227 54811 48341 55045
tri 48377 55012 48393 55028 se
rect 48393 55012 48470 55028
rect 48377 54946 48470 55012
rect 48377 54844 48470 54910
tri 48377 54828 48393 54844 ne
rect 48393 54828 48470 54844
rect 48210 54729 48358 54811
rect 48098 54696 48175 54712
tri 48175 54696 48191 54712 sw
rect 48098 54630 48191 54696
rect 48227 54571 48341 54729
tri 48377 54696 48393 54712 se
rect 48393 54696 48470 54712
rect 48377 54630 48470 54696
rect 48098 54495 48470 54571
rect 48098 54370 48191 54436
rect 48098 54354 48175 54370
tri 48175 54354 48191 54370 nw
rect 48227 54337 48341 54495
rect 48377 54370 48470 54436
tri 48377 54354 48393 54370 ne
rect 48393 54354 48470 54370
rect 48210 54255 48358 54337
rect 48098 54222 48175 54238
tri 48175 54222 48191 54238 sw
rect 48098 54156 48191 54222
rect 48098 54054 48191 54120
rect 48098 54038 48175 54054
tri 48175 54038 48191 54054 nw
rect 48227 54021 48341 54255
tri 48377 54222 48393 54238 se
rect 48393 54222 48470 54238
rect 48377 54156 48470 54222
rect 48377 54054 48470 54120
tri 48377 54038 48393 54054 ne
rect 48393 54038 48470 54054
rect 48210 53939 48358 54021
rect 48098 53906 48175 53922
tri 48175 53906 48191 53922 sw
rect 48098 53840 48191 53906
rect 48227 53781 48341 53939
tri 48377 53906 48393 53922 se
rect 48393 53906 48470 53922
rect 48377 53840 48470 53906
rect 48098 53705 48470 53781
rect 48098 53580 48191 53646
rect 48098 53564 48175 53580
tri 48175 53564 48191 53580 nw
rect 48227 53547 48341 53705
rect 48377 53580 48470 53646
tri 48377 53564 48393 53580 ne
rect 48393 53564 48470 53580
rect 48210 53465 48358 53547
rect 48098 53432 48175 53448
tri 48175 53432 48191 53448 sw
rect 48098 53366 48191 53432
rect 48098 53264 48191 53330
rect 48098 53248 48175 53264
tri 48175 53248 48191 53264 nw
rect 48227 53231 48341 53465
tri 48377 53432 48393 53448 se
rect 48393 53432 48470 53448
rect 48377 53366 48470 53432
rect 48377 53264 48470 53330
tri 48377 53248 48393 53264 ne
rect 48393 53248 48470 53264
rect 48210 53149 48358 53231
rect 48098 53116 48175 53132
tri 48175 53116 48191 53132 sw
rect 48098 53050 48191 53116
rect 48227 52991 48341 53149
tri 48377 53116 48393 53132 se
rect 48393 53116 48470 53132
rect 48377 53050 48470 53116
rect 48098 52915 48470 52991
rect 48098 52790 48191 52856
rect 48098 52774 48175 52790
tri 48175 52774 48191 52790 nw
rect 48227 52757 48341 52915
rect 48377 52790 48470 52856
tri 48377 52774 48393 52790 ne
rect 48393 52774 48470 52790
rect 48210 52675 48358 52757
rect 48098 52642 48175 52658
tri 48175 52642 48191 52658 sw
rect 48098 52576 48191 52642
rect 48098 52474 48191 52540
rect 48098 52458 48175 52474
tri 48175 52458 48191 52474 nw
rect 48227 52441 48341 52675
tri 48377 52642 48393 52658 se
rect 48393 52642 48470 52658
rect 48377 52576 48470 52642
rect 48377 52474 48470 52540
tri 48377 52458 48393 52474 ne
rect 48393 52458 48470 52474
rect 48210 52359 48358 52441
rect 48098 52326 48175 52342
tri 48175 52326 48191 52342 sw
rect 48098 52260 48191 52326
rect 48227 52201 48341 52359
tri 48377 52326 48393 52342 se
rect 48393 52326 48470 52342
rect 48377 52260 48470 52326
rect 48098 52125 48470 52201
rect 48098 52000 48191 52066
rect 48098 51984 48175 52000
tri 48175 51984 48191 52000 nw
rect 48227 51967 48341 52125
rect 48377 52000 48470 52066
tri 48377 51984 48393 52000 ne
rect 48393 51984 48470 52000
rect 48210 51885 48358 51967
rect 48098 51852 48175 51868
tri 48175 51852 48191 51868 sw
rect 48098 51786 48191 51852
rect 48098 51684 48191 51750
rect 48098 51668 48175 51684
tri 48175 51668 48191 51684 nw
rect 48227 51651 48341 51885
tri 48377 51852 48393 51868 se
rect 48393 51852 48470 51868
rect 48377 51786 48470 51852
rect 48377 51684 48470 51750
tri 48377 51668 48393 51684 ne
rect 48393 51668 48470 51684
rect 48210 51569 48358 51651
rect 48098 51536 48175 51552
tri 48175 51536 48191 51552 sw
rect 48098 51470 48191 51536
rect 48227 51411 48341 51569
tri 48377 51536 48393 51552 se
rect 48393 51536 48470 51552
rect 48377 51470 48470 51536
rect 48098 51335 48470 51411
rect 48098 51210 48191 51276
rect 48098 51194 48175 51210
tri 48175 51194 48191 51210 nw
rect 48227 51177 48341 51335
rect 48377 51210 48470 51276
tri 48377 51194 48393 51210 ne
rect 48393 51194 48470 51210
rect 48210 51095 48358 51177
rect 48098 51062 48175 51078
tri 48175 51062 48191 51078 sw
rect 48098 50996 48191 51062
rect 48098 50894 48191 50960
rect 48098 50878 48175 50894
tri 48175 50878 48191 50894 nw
rect 48227 50861 48341 51095
tri 48377 51062 48393 51078 se
rect 48393 51062 48470 51078
rect 48377 50996 48470 51062
rect 48377 50894 48470 50960
tri 48377 50878 48393 50894 ne
rect 48393 50878 48470 50894
rect 48210 50779 48358 50861
rect 48098 50746 48175 50762
tri 48175 50746 48191 50762 sw
rect 48098 50680 48191 50746
rect 48227 50621 48341 50779
tri 48377 50746 48393 50762 se
rect 48393 50746 48470 50762
rect 48377 50680 48470 50746
rect 48098 50545 48470 50621
rect 48098 50420 48191 50486
rect 48098 50404 48175 50420
tri 48175 50404 48191 50420 nw
rect 48227 50387 48341 50545
rect 48377 50420 48470 50486
tri 48377 50404 48393 50420 ne
rect 48393 50404 48470 50420
rect 48210 50305 48358 50387
rect 48098 50272 48175 50288
tri 48175 50272 48191 50288 sw
rect 48098 50206 48191 50272
rect 48098 50104 48191 50170
rect 48098 50088 48175 50104
tri 48175 50088 48191 50104 nw
rect 48227 50071 48341 50305
tri 48377 50272 48393 50288 se
rect 48393 50272 48470 50288
rect 48377 50206 48470 50272
rect 48377 50104 48470 50170
tri 48377 50088 48393 50104 ne
rect 48393 50088 48470 50104
rect 48210 49989 48358 50071
rect 48098 49956 48175 49972
tri 48175 49956 48191 49972 sw
rect 48098 49890 48191 49956
rect 48227 49831 48341 49989
tri 48377 49956 48393 49972 se
rect 48393 49956 48470 49972
rect 48377 49890 48470 49956
rect 48098 49755 48470 49831
rect 48098 49630 48191 49696
rect 48098 49614 48175 49630
tri 48175 49614 48191 49630 nw
rect 48227 49597 48341 49755
rect 48377 49630 48470 49696
tri 48377 49614 48393 49630 ne
rect 48393 49614 48470 49630
rect 48210 49515 48358 49597
rect 48098 49482 48175 49498
tri 48175 49482 48191 49498 sw
rect 48098 49416 48191 49482
rect 48098 49314 48191 49380
rect 48098 49298 48175 49314
tri 48175 49298 48191 49314 nw
rect 48227 49281 48341 49515
tri 48377 49482 48393 49498 se
rect 48393 49482 48470 49498
rect 48377 49416 48470 49482
rect 48377 49314 48470 49380
tri 48377 49298 48393 49314 ne
rect 48393 49298 48470 49314
rect 48210 49199 48358 49281
rect 48098 49166 48175 49182
tri 48175 49166 48191 49182 sw
rect 48098 49100 48191 49166
rect 48227 49041 48341 49199
tri 48377 49166 48393 49182 se
rect 48393 49166 48470 49182
rect 48377 49100 48470 49166
rect 48098 48965 48470 49041
rect 48098 48840 48191 48906
rect 48098 48824 48175 48840
tri 48175 48824 48191 48840 nw
rect 48227 48807 48341 48965
rect 48377 48840 48470 48906
tri 48377 48824 48393 48840 ne
rect 48393 48824 48470 48840
rect 48210 48725 48358 48807
rect 48098 48692 48175 48708
tri 48175 48692 48191 48708 sw
rect 48098 48626 48191 48692
rect 48098 48524 48191 48590
rect 48098 48508 48175 48524
tri 48175 48508 48191 48524 nw
rect 48227 48491 48341 48725
tri 48377 48692 48393 48708 se
rect 48393 48692 48470 48708
rect 48377 48626 48470 48692
rect 48377 48524 48470 48590
tri 48377 48508 48393 48524 ne
rect 48393 48508 48470 48524
rect 48210 48409 48358 48491
rect 48098 48376 48175 48392
tri 48175 48376 48191 48392 sw
rect 48098 48310 48191 48376
rect 48227 48251 48341 48409
tri 48377 48376 48393 48392 se
rect 48393 48376 48470 48392
rect 48377 48310 48470 48376
rect 48098 48175 48470 48251
rect 48098 48050 48191 48116
rect 48098 48034 48175 48050
tri 48175 48034 48191 48050 nw
rect 48227 48017 48341 48175
rect 48377 48050 48470 48116
tri 48377 48034 48393 48050 ne
rect 48393 48034 48470 48050
rect 48210 47935 48358 48017
rect 48098 47902 48175 47918
tri 48175 47902 48191 47918 sw
rect 48098 47836 48191 47902
rect 48098 47734 48191 47800
rect 48098 47718 48175 47734
tri 48175 47718 48191 47734 nw
rect 48227 47701 48341 47935
tri 48377 47902 48393 47918 se
rect 48393 47902 48470 47918
rect 48377 47836 48470 47902
rect 48377 47734 48470 47800
tri 48377 47718 48393 47734 ne
rect 48393 47718 48470 47734
rect 48210 47619 48358 47701
rect 48098 47586 48175 47602
tri 48175 47586 48191 47602 sw
rect 48098 47520 48191 47586
rect 48227 47461 48341 47619
tri 48377 47586 48393 47602 se
rect 48393 47586 48470 47602
rect 48377 47520 48470 47586
rect 48098 47385 48470 47461
rect 48098 47260 48191 47326
rect 48098 47244 48175 47260
tri 48175 47244 48191 47260 nw
rect 48227 47227 48341 47385
rect 48377 47260 48470 47326
tri 48377 47244 48393 47260 ne
rect 48393 47244 48470 47260
rect 48210 47145 48358 47227
rect 48098 47112 48175 47128
tri 48175 47112 48191 47128 sw
rect 48098 47046 48191 47112
rect 48098 46944 48191 47010
rect 48098 46928 48175 46944
tri 48175 46928 48191 46944 nw
rect 48227 46911 48341 47145
tri 48377 47112 48393 47128 se
rect 48393 47112 48470 47128
rect 48377 47046 48470 47112
rect 48377 46944 48470 47010
tri 48377 46928 48393 46944 ne
rect 48393 46928 48470 46944
rect 48210 46829 48358 46911
rect 48098 46796 48175 46812
tri 48175 46796 48191 46812 sw
rect 48098 46730 48191 46796
rect 48227 46671 48341 46829
tri 48377 46796 48393 46812 se
rect 48393 46796 48470 46812
rect 48377 46730 48470 46796
rect 48098 46595 48470 46671
rect 48098 46470 48191 46536
rect 48098 46454 48175 46470
tri 48175 46454 48191 46470 nw
rect 48227 46437 48341 46595
rect 48377 46470 48470 46536
tri 48377 46454 48393 46470 ne
rect 48393 46454 48470 46470
rect 48210 46355 48358 46437
rect 48098 46322 48175 46338
tri 48175 46322 48191 46338 sw
rect 48098 46256 48191 46322
rect 48098 46154 48191 46220
rect 48098 46138 48175 46154
tri 48175 46138 48191 46154 nw
rect 48227 46121 48341 46355
tri 48377 46322 48393 46338 se
rect 48393 46322 48470 46338
rect 48377 46256 48470 46322
rect 48377 46154 48470 46220
tri 48377 46138 48393 46154 ne
rect 48393 46138 48470 46154
rect 48210 46039 48358 46121
rect 48098 46006 48175 46022
tri 48175 46006 48191 46022 sw
rect 48098 45940 48191 46006
rect 48227 45881 48341 46039
tri 48377 46006 48393 46022 se
rect 48393 46006 48470 46022
rect 48377 45940 48470 46006
rect 48098 45805 48470 45881
rect 48098 45680 48191 45746
rect 48098 45664 48175 45680
tri 48175 45664 48191 45680 nw
rect 48227 45647 48341 45805
rect 48377 45680 48470 45746
tri 48377 45664 48393 45680 ne
rect 48393 45664 48470 45680
rect 48210 45565 48358 45647
rect 48098 45532 48175 45548
tri 48175 45532 48191 45548 sw
rect 48098 45466 48191 45532
rect 48098 45364 48191 45430
rect 48098 45348 48175 45364
tri 48175 45348 48191 45364 nw
rect 48227 45331 48341 45565
tri 48377 45532 48393 45548 se
rect 48393 45532 48470 45548
rect 48377 45466 48470 45532
rect 48377 45364 48470 45430
tri 48377 45348 48393 45364 ne
rect 48393 45348 48470 45364
rect 48210 45249 48358 45331
rect 48098 45216 48175 45232
tri 48175 45216 48191 45232 sw
rect 48098 45150 48191 45216
rect 48227 45091 48341 45249
tri 48377 45216 48393 45232 se
rect 48393 45216 48470 45232
rect 48377 45150 48470 45216
rect 48098 45015 48470 45091
rect 48098 44890 48191 44956
rect 48098 44874 48175 44890
tri 48175 44874 48191 44890 nw
rect 48227 44857 48341 45015
rect 48377 44890 48470 44956
tri 48377 44874 48393 44890 ne
rect 48393 44874 48470 44890
rect 48210 44775 48358 44857
rect 48098 44742 48175 44758
tri 48175 44742 48191 44758 sw
rect 48098 44676 48191 44742
rect 48098 44574 48191 44640
rect 48098 44558 48175 44574
tri 48175 44558 48191 44574 nw
rect 48227 44541 48341 44775
tri 48377 44742 48393 44758 se
rect 48393 44742 48470 44758
rect 48377 44676 48470 44742
rect 48377 44574 48470 44640
tri 48377 44558 48393 44574 ne
rect 48393 44558 48470 44574
rect 48210 44459 48358 44541
rect 48098 44426 48175 44442
tri 48175 44426 48191 44442 sw
rect 48098 44360 48191 44426
rect 48227 44301 48341 44459
tri 48377 44426 48393 44442 se
rect 48393 44426 48470 44442
rect 48377 44360 48470 44426
rect 48098 44225 48470 44301
rect 48098 44100 48191 44166
rect 48098 44084 48175 44100
tri 48175 44084 48191 44100 nw
rect 48227 44067 48341 44225
rect 48377 44100 48470 44166
tri 48377 44084 48393 44100 ne
rect 48393 44084 48470 44100
rect 48210 43985 48358 44067
rect 48098 43952 48175 43968
tri 48175 43952 48191 43968 sw
rect 48098 43886 48191 43952
rect 48098 43784 48191 43850
rect 48098 43768 48175 43784
tri 48175 43768 48191 43784 nw
rect 48227 43751 48341 43985
tri 48377 43952 48393 43968 se
rect 48393 43952 48470 43968
rect 48377 43886 48470 43952
rect 48377 43784 48470 43850
tri 48377 43768 48393 43784 ne
rect 48393 43768 48470 43784
rect 48210 43669 48358 43751
rect 48098 43636 48175 43652
tri 48175 43636 48191 43652 sw
rect 48098 43570 48191 43636
rect 48227 43511 48341 43669
tri 48377 43636 48393 43652 se
rect 48393 43636 48470 43652
rect 48377 43570 48470 43636
rect 48098 43435 48470 43511
rect 48098 43310 48191 43376
rect 48098 43294 48175 43310
tri 48175 43294 48191 43310 nw
rect 48227 43277 48341 43435
rect 48377 43310 48470 43376
tri 48377 43294 48393 43310 ne
rect 48393 43294 48470 43310
rect 48210 43195 48358 43277
rect 48098 43162 48175 43178
tri 48175 43162 48191 43178 sw
rect 48098 43096 48191 43162
rect 48098 42994 48191 43060
rect 48098 42978 48175 42994
tri 48175 42978 48191 42994 nw
rect 48227 42961 48341 43195
tri 48377 43162 48393 43178 se
rect 48393 43162 48470 43178
rect 48377 43096 48470 43162
rect 48377 42994 48470 43060
tri 48377 42978 48393 42994 ne
rect 48393 42978 48470 42994
rect 48210 42879 48358 42961
rect 48098 42846 48175 42862
tri 48175 42846 48191 42862 sw
rect 48098 42780 48191 42846
rect 48227 42721 48341 42879
tri 48377 42846 48393 42862 se
rect 48393 42846 48470 42862
rect 48377 42780 48470 42846
rect 48098 42645 48470 42721
rect 48098 42520 48191 42586
rect 48098 42504 48175 42520
tri 48175 42504 48191 42520 nw
rect 48227 42487 48341 42645
rect 48377 42520 48470 42586
tri 48377 42504 48393 42520 ne
rect 48393 42504 48470 42520
rect 48210 42405 48358 42487
rect 48098 42372 48175 42388
tri 48175 42372 48191 42388 sw
rect 48098 42306 48191 42372
rect 48098 42204 48191 42270
rect 48098 42188 48175 42204
tri 48175 42188 48191 42204 nw
rect 48227 42171 48341 42405
tri 48377 42372 48393 42388 se
rect 48393 42372 48470 42388
rect 48377 42306 48470 42372
rect 48377 42204 48470 42270
tri 48377 42188 48393 42204 ne
rect 48393 42188 48470 42204
rect 48210 42089 48358 42171
rect 48098 42056 48175 42072
tri 48175 42056 48191 42072 sw
rect 48098 41990 48191 42056
rect 48227 41931 48341 42089
tri 48377 42056 48393 42072 se
rect 48393 42056 48470 42072
rect 48377 41990 48470 42056
rect 48098 41855 48470 41931
rect 48098 41730 48191 41796
rect 48098 41714 48175 41730
tri 48175 41714 48191 41730 nw
rect 48227 41697 48341 41855
rect 48377 41730 48470 41796
tri 48377 41714 48393 41730 ne
rect 48393 41714 48470 41730
rect 48210 41615 48358 41697
rect 48098 41582 48175 41598
tri 48175 41582 48191 41598 sw
rect 48098 41516 48191 41582
rect 48098 41414 48191 41480
rect 48098 41398 48175 41414
tri 48175 41398 48191 41414 nw
rect 48227 41381 48341 41615
tri 48377 41582 48393 41598 se
rect 48393 41582 48470 41598
rect 48377 41516 48470 41582
rect 48377 41414 48470 41480
tri 48377 41398 48393 41414 ne
rect 48393 41398 48470 41414
rect 48210 41299 48358 41381
rect 48098 41266 48175 41282
tri 48175 41266 48191 41282 sw
rect 48098 41200 48191 41266
rect 48227 41141 48341 41299
tri 48377 41266 48393 41282 se
rect 48393 41266 48470 41282
rect 48377 41200 48470 41266
rect 48098 41065 48470 41141
rect 48098 40940 48191 41006
rect 48098 40924 48175 40940
tri 48175 40924 48191 40940 nw
rect 48227 40907 48341 41065
rect 48377 40940 48470 41006
tri 48377 40924 48393 40940 ne
rect 48393 40924 48470 40940
rect 48210 40825 48358 40907
rect 48098 40792 48175 40808
tri 48175 40792 48191 40808 sw
rect 48098 40726 48191 40792
rect 48098 40624 48191 40690
rect 48098 40608 48175 40624
tri 48175 40608 48191 40624 nw
rect 48227 40591 48341 40825
tri 48377 40792 48393 40808 se
rect 48393 40792 48470 40808
rect 48377 40726 48470 40792
rect 48377 40624 48470 40690
tri 48377 40608 48393 40624 ne
rect 48393 40608 48470 40624
rect 48210 40509 48358 40591
rect 48098 40476 48175 40492
tri 48175 40476 48191 40492 sw
rect 48098 40410 48191 40476
rect 48227 40351 48341 40509
tri 48377 40476 48393 40492 se
rect 48393 40476 48470 40492
rect 48377 40410 48470 40476
rect 48098 40275 48470 40351
rect 48098 40150 48191 40216
rect 48098 40134 48175 40150
tri 48175 40134 48191 40150 nw
rect 48227 40117 48341 40275
rect 48377 40150 48470 40216
tri 48377 40134 48393 40150 ne
rect 48393 40134 48470 40150
rect 48210 40035 48358 40117
rect 48098 40002 48175 40018
tri 48175 40002 48191 40018 sw
rect 48098 39936 48191 40002
rect 48098 39834 48191 39900
rect 48098 39818 48175 39834
tri 48175 39818 48191 39834 nw
rect 48227 39801 48341 40035
tri 48377 40002 48393 40018 se
rect 48393 40002 48470 40018
rect 48377 39936 48470 40002
rect 48377 39834 48470 39900
tri 48377 39818 48393 39834 ne
rect 48393 39818 48470 39834
rect 48210 39719 48358 39801
rect 48098 39686 48175 39702
tri 48175 39686 48191 39702 sw
rect 48098 39620 48191 39686
rect 48227 39561 48341 39719
tri 48377 39686 48393 39702 se
rect 48393 39686 48470 39702
rect 48377 39620 48470 39686
rect 48098 39485 48470 39561
rect 48098 39360 48191 39426
rect 48098 39344 48175 39360
tri 48175 39344 48191 39360 nw
rect 48227 39327 48341 39485
rect 48377 39360 48470 39426
tri 48377 39344 48393 39360 ne
rect 48393 39344 48470 39360
rect 48210 39245 48358 39327
rect 48098 39212 48175 39228
tri 48175 39212 48191 39228 sw
rect 48098 39146 48191 39212
rect 48098 39044 48191 39110
rect 48098 39028 48175 39044
tri 48175 39028 48191 39044 nw
rect 48227 39011 48341 39245
tri 48377 39212 48393 39228 se
rect 48393 39212 48470 39228
rect 48377 39146 48470 39212
rect 48377 39044 48470 39110
tri 48377 39028 48393 39044 ne
rect 48393 39028 48470 39044
rect 48210 38929 48358 39011
rect 48098 38896 48175 38912
tri 48175 38896 48191 38912 sw
rect 48098 38830 48191 38896
rect 48227 38771 48341 38929
tri 48377 38896 48393 38912 se
rect 48393 38896 48470 38912
rect 48377 38830 48470 38896
rect 48098 38695 48470 38771
rect 48098 38570 48191 38636
rect 48098 38554 48175 38570
tri 48175 38554 48191 38570 nw
rect 48227 38537 48341 38695
rect 48377 38570 48470 38636
tri 48377 38554 48393 38570 ne
rect 48393 38554 48470 38570
rect 48210 38455 48358 38537
rect 48098 38422 48175 38438
tri 48175 38422 48191 38438 sw
rect 48098 38356 48191 38422
rect 48098 38254 48191 38320
rect 48098 38238 48175 38254
tri 48175 38238 48191 38254 nw
rect 48227 38221 48341 38455
tri 48377 38422 48393 38438 se
rect 48393 38422 48470 38438
rect 48377 38356 48470 38422
rect 48377 38254 48470 38320
tri 48377 38238 48393 38254 ne
rect 48393 38238 48470 38254
rect 48210 38139 48358 38221
rect 48098 38106 48175 38122
tri 48175 38106 48191 38122 sw
rect 48098 38040 48191 38106
rect 48227 37981 48341 38139
tri 48377 38106 48393 38122 se
rect 48393 38106 48470 38122
rect 48377 38040 48470 38106
rect 48098 37905 48470 37981
rect 48098 37780 48191 37846
rect 48098 37764 48175 37780
tri 48175 37764 48191 37780 nw
rect 48227 37747 48341 37905
rect 48377 37780 48470 37846
tri 48377 37764 48393 37780 ne
rect 48393 37764 48470 37780
rect 48210 37665 48358 37747
rect 48098 37632 48175 37648
tri 48175 37632 48191 37648 sw
rect 48098 37566 48191 37632
rect 48098 37464 48191 37530
rect 48098 37448 48175 37464
tri 48175 37448 48191 37464 nw
rect 48227 37431 48341 37665
tri 48377 37632 48393 37648 se
rect 48393 37632 48470 37648
rect 48377 37566 48470 37632
rect 48377 37464 48470 37530
tri 48377 37448 48393 37464 ne
rect 48393 37448 48470 37464
rect 48210 37349 48358 37431
rect 48098 37316 48175 37332
tri 48175 37316 48191 37332 sw
rect 48098 37250 48191 37316
rect 48227 37191 48341 37349
tri 48377 37316 48393 37332 se
rect 48393 37316 48470 37332
rect 48377 37250 48470 37316
rect 48098 37115 48470 37191
rect 48098 36990 48191 37056
rect 48098 36974 48175 36990
tri 48175 36974 48191 36990 nw
rect 48227 36957 48341 37115
rect 48377 36990 48470 37056
tri 48377 36974 48393 36990 ne
rect 48393 36974 48470 36990
rect 48210 36875 48358 36957
rect 48098 36842 48175 36858
tri 48175 36842 48191 36858 sw
rect 48098 36776 48191 36842
rect 48098 36674 48191 36740
rect 48098 36658 48175 36674
tri 48175 36658 48191 36674 nw
rect 48227 36641 48341 36875
tri 48377 36842 48393 36858 se
rect 48393 36842 48470 36858
rect 48377 36776 48470 36842
rect 48377 36674 48470 36740
tri 48377 36658 48393 36674 ne
rect 48393 36658 48470 36674
rect 48210 36559 48358 36641
rect 48098 36526 48175 36542
tri 48175 36526 48191 36542 sw
rect 48098 36460 48191 36526
rect 48227 36401 48341 36559
tri 48377 36526 48393 36542 se
rect 48393 36526 48470 36542
rect 48377 36460 48470 36526
rect 48098 36325 48470 36401
rect 48098 36200 48191 36266
rect 48098 36184 48175 36200
tri 48175 36184 48191 36200 nw
rect 48227 36167 48341 36325
rect 48377 36200 48470 36266
tri 48377 36184 48393 36200 ne
rect 48393 36184 48470 36200
rect 48210 36085 48358 36167
rect 48098 36052 48175 36068
tri 48175 36052 48191 36068 sw
rect 48098 35986 48191 36052
rect 48098 35884 48191 35950
rect 48098 35868 48175 35884
tri 48175 35868 48191 35884 nw
rect 48227 35851 48341 36085
tri 48377 36052 48393 36068 se
rect 48393 36052 48470 36068
rect 48377 35986 48470 36052
rect 48377 35884 48470 35950
tri 48377 35868 48393 35884 ne
rect 48393 35868 48470 35884
rect 48210 35769 48358 35851
rect 48098 35736 48175 35752
tri 48175 35736 48191 35752 sw
rect 48098 35670 48191 35736
rect 48227 35611 48341 35769
tri 48377 35736 48393 35752 se
rect 48393 35736 48470 35752
rect 48377 35670 48470 35736
rect 48098 35535 48470 35611
rect 48098 35410 48191 35476
rect 48098 35394 48175 35410
tri 48175 35394 48191 35410 nw
rect 48227 35377 48341 35535
rect 48377 35410 48470 35476
tri 48377 35394 48393 35410 ne
rect 48393 35394 48470 35410
rect 48210 35295 48358 35377
rect 48098 35262 48175 35278
tri 48175 35262 48191 35278 sw
rect 48098 35196 48191 35262
rect 48098 35094 48191 35160
rect 48098 35078 48175 35094
tri 48175 35078 48191 35094 nw
rect 48227 35061 48341 35295
tri 48377 35262 48393 35278 se
rect 48393 35262 48470 35278
rect 48377 35196 48470 35262
rect 48377 35094 48470 35160
tri 48377 35078 48393 35094 ne
rect 48393 35078 48470 35094
rect 48210 34979 48358 35061
rect 48098 34946 48175 34962
tri 48175 34946 48191 34962 sw
rect 48098 34880 48191 34946
rect 48227 34821 48341 34979
tri 48377 34946 48393 34962 se
rect 48393 34946 48470 34962
rect 48377 34880 48470 34946
rect 48098 34745 48470 34821
rect 48098 34620 48191 34686
rect 48098 34604 48175 34620
tri 48175 34604 48191 34620 nw
rect 48227 34587 48341 34745
rect 48377 34620 48470 34686
tri 48377 34604 48393 34620 ne
rect 48393 34604 48470 34620
rect 48210 34505 48358 34587
rect 48098 34472 48175 34488
tri 48175 34472 48191 34488 sw
rect 48098 34406 48191 34472
rect 48098 34304 48191 34370
rect 48098 34288 48175 34304
tri 48175 34288 48191 34304 nw
rect 48227 34271 48341 34505
tri 48377 34472 48393 34488 se
rect 48393 34472 48470 34488
rect 48377 34406 48470 34472
rect 48377 34304 48470 34370
tri 48377 34288 48393 34304 ne
rect 48393 34288 48470 34304
rect 48210 34189 48358 34271
rect 48098 34156 48175 34172
tri 48175 34156 48191 34172 sw
rect 48098 34090 48191 34156
rect 48227 34031 48341 34189
tri 48377 34156 48393 34172 se
rect 48393 34156 48470 34172
rect 48377 34090 48470 34156
rect 48098 33955 48470 34031
rect 48098 33830 48191 33896
rect 48098 33814 48175 33830
tri 48175 33814 48191 33830 nw
rect 48227 33797 48341 33955
rect 48377 33830 48470 33896
tri 48377 33814 48393 33830 ne
rect 48393 33814 48470 33830
rect 48210 33715 48358 33797
rect 48098 33682 48175 33698
tri 48175 33682 48191 33698 sw
rect 48098 33616 48191 33682
rect 48098 33514 48191 33580
rect 48098 33498 48175 33514
tri 48175 33498 48191 33514 nw
rect 48227 33481 48341 33715
tri 48377 33682 48393 33698 se
rect 48393 33682 48470 33698
rect 48377 33616 48470 33682
rect 48377 33514 48470 33580
tri 48377 33498 48393 33514 ne
rect 48393 33498 48470 33514
rect 48210 33399 48358 33481
rect 48098 33366 48175 33382
tri 48175 33366 48191 33382 sw
rect 48098 33300 48191 33366
rect 48227 33241 48341 33399
tri 48377 33366 48393 33382 se
rect 48393 33366 48470 33382
rect 48377 33300 48470 33366
rect 48098 33165 48470 33241
rect 48098 33040 48191 33106
rect 48098 33024 48175 33040
tri 48175 33024 48191 33040 nw
rect 48227 33007 48341 33165
rect 48377 33040 48470 33106
tri 48377 33024 48393 33040 ne
rect 48393 33024 48470 33040
rect 48210 32925 48358 33007
rect 48098 32892 48175 32908
tri 48175 32892 48191 32908 sw
rect 48098 32826 48191 32892
rect 48098 32724 48191 32790
rect 48098 32708 48175 32724
tri 48175 32708 48191 32724 nw
rect 48227 32691 48341 32925
tri 48377 32892 48393 32908 se
rect 48393 32892 48470 32908
rect 48377 32826 48470 32892
rect 48377 32724 48470 32790
tri 48377 32708 48393 32724 ne
rect 48393 32708 48470 32724
rect 48210 32609 48358 32691
rect 48098 32576 48175 32592
tri 48175 32576 48191 32592 sw
rect 48098 32510 48191 32576
rect 48227 32451 48341 32609
tri 48377 32576 48393 32592 se
rect 48393 32576 48470 32592
rect 48377 32510 48470 32576
rect 48098 32375 48470 32451
rect 48098 32250 48191 32316
rect 48098 32234 48175 32250
tri 48175 32234 48191 32250 nw
rect 48227 32217 48341 32375
rect 48377 32250 48470 32316
tri 48377 32234 48393 32250 ne
rect 48393 32234 48470 32250
rect 48210 32135 48358 32217
rect 48098 32102 48175 32118
tri 48175 32102 48191 32118 sw
rect 48098 32036 48191 32102
rect 48098 31934 48191 32000
rect 48098 31918 48175 31934
tri 48175 31918 48191 31934 nw
rect 48227 31901 48341 32135
tri 48377 32102 48393 32118 se
rect 48393 32102 48470 32118
rect 48377 32036 48470 32102
rect 48377 31934 48470 32000
tri 48377 31918 48393 31934 ne
rect 48393 31918 48470 31934
rect 48210 31819 48358 31901
rect 48098 31786 48175 31802
tri 48175 31786 48191 31802 sw
rect 48098 31720 48191 31786
rect 48227 31661 48341 31819
tri 48377 31786 48393 31802 se
rect 48393 31786 48470 31802
rect 48377 31720 48470 31786
rect 48098 31585 48470 31661
rect 48098 31460 48191 31526
rect 48098 31444 48175 31460
tri 48175 31444 48191 31460 nw
rect 48227 31427 48341 31585
rect 48377 31460 48470 31526
tri 48377 31444 48393 31460 ne
rect 48393 31444 48470 31460
rect 48210 31345 48358 31427
rect 48098 31312 48175 31328
tri 48175 31312 48191 31328 sw
rect 48098 31246 48191 31312
rect 48098 31144 48191 31210
rect 48098 31128 48175 31144
tri 48175 31128 48191 31144 nw
rect 48227 31111 48341 31345
tri 48377 31312 48393 31328 se
rect 48393 31312 48470 31328
rect 48377 31246 48470 31312
rect 48377 31144 48470 31210
tri 48377 31128 48393 31144 ne
rect 48393 31128 48470 31144
rect 48210 31029 48358 31111
rect 48098 30996 48175 31012
tri 48175 30996 48191 31012 sw
rect 48098 30930 48191 30996
rect 48227 30871 48341 31029
tri 48377 30996 48393 31012 se
rect 48393 30996 48470 31012
rect 48377 30930 48470 30996
rect 48098 30795 48470 30871
rect 48098 30670 48191 30736
rect 48098 30654 48175 30670
tri 48175 30654 48191 30670 nw
rect 48227 30637 48341 30795
rect 48377 30670 48470 30736
tri 48377 30654 48393 30670 ne
rect 48393 30654 48470 30670
rect 48210 30555 48358 30637
rect 48098 30522 48175 30538
tri 48175 30522 48191 30538 sw
rect 48098 30456 48191 30522
rect 48098 30354 48191 30420
rect 48098 30338 48175 30354
tri 48175 30338 48191 30354 nw
rect 48227 30321 48341 30555
tri 48377 30522 48393 30538 se
rect 48393 30522 48470 30538
rect 48377 30456 48470 30522
rect 48377 30354 48470 30420
tri 48377 30338 48393 30354 ne
rect 48393 30338 48470 30354
rect 48210 30239 48358 30321
rect 48098 30206 48175 30222
tri 48175 30206 48191 30222 sw
rect 48098 30140 48191 30206
rect 48227 30081 48341 30239
tri 48377 30206 48393 30222 se
rect 48393 30206 48470 30222
rect 48377 30140 48470 30206
rect 48098 30005 48470 30081
rect 48098 29880 48191 29946
rect 48098 29864 48175 29880
tri 48175 29864 48191 29880 nw
rect 48227 29847 48341 30005
rect 48377 29880 48470 29946
tri 48377 29864 48393 29880 ne
rect 48393 29864 48470 29880
rect 48210 29765 48358 29847
rect 48098 29732 48175 29748
tri 48175 29732 48191 29748 sw
rect 48098 29666 48191 29732
rect 48098 29564 48191 29630
rect 48098 29548 48175 29564
tri 48175 29548 48191 29564 nw
rect 48227 29531 48341 29765
tri 48377 29732 48393 29748 se
rect 48393 29732 48470 29748
rect 48377 29666 48470 29732
rect 48377 29564 48470 29630
tri 48377 29548 48393 29564 ne
rect 48393 29548 48470 29564
rect 48210 29449 48358 29531
rect 48098 29416 48175 29432
tri 48175 29416 48191 29432 sw
rect 48098 29350 48191 29416
rect 48227 29291 48341 29449
tri 48377 29416 48393 29432 se
rect 48393 29416 48470 29432
rect 48377 29350 48470 29416
rect 48098 29215 48470 29291
rect 48098 29090 48191 29156
rect 48098 29074 48175 29090
tri 48175 29074 48191 29090 nw
rect 48227 29057 48341 29215
rect 48377 29090 48470 29156
tri 48377 29074 48393 29090 ne
rect 48393 29074 48470 29090
rect 48210 28975 48358 29057
rect 48098 28942 48175 28958
tri 48175 28942 48191 28958 sw
rect 48098 28876 48191 28942
rect 48227 28833 48341 28975
tri 48377 28942 48393 28958 se
rect 48393 28942 48470 28958
rect 48377 28876 48470 28942
rect 48506 28463 48542 80603
rect 48578 28463 48614 80603
rect 48650 80445 48686 80603
rect 48642 80303 48694 80445
rect 48650 28763 48686 80303
rect 48642 28621 48694 28763
rect 48650 28463 48686 28621
rect 48722 28463 48758 80603
rect 48794 28463 48830 80603
rect 48866 28833 48950 80233
rect 48986 28463 49022 80603
rect 49058 28463 49094 80603
rect 49130 80445 49166 80603
rect 49122 80303 49174 80445
rect 49130 28763 49166 80303
rect 49122 28621 49174 28763
rect 49130 28463 49166 28621
rect 49202 28463 49238 80603
rect 49274 28463 49310 80603
rect 49346 80124 49439 80190
rect 49346 80108 49423 80124
tri 49423 80108 49439 80124 nw
rect 49475 80091 49589 80233
rect 49625 80124 49718 80190
tri 49625 80108 49641 80124 ne
rect 49641 80108 49718 80124
rect 49458 80009 49606 80091
rect 49346 79976 49423 79992
tri 49423 79976 49439 79992 sw
rect 49346 79910 49439 79976
rect 49475 79851 49589 80009
tri 49625 79976 49641 79992 se
rect 49641 79976 49718 79992
rect 49625 79910 49718 79976
rect 49346 79775 49718 79851
rect 49346 79650 49439 79716
rect 49346 79634 49423 79650
tri 49423 79634 49439 79650 nw
rect 49475 79617 49589 79775
rect 49625 79650 49718 79716
tri 49625 79634 49641 79650 ne
rect 49641 79634 49718 79650
rect 49458 79535 49606 79617
rect 49346 79502 49423 79518
tri 49423 79502 49439 79518 sw
rect 49346 79436 49439 79502
rect 49346 79334 49439 79400
rect 49346 79318 49423 79334
tri 49423 79318 49439 79334 nw
rect 49475 79301 49589 79535
tri 49625 79502 49641 79518 se
rect 49641 79502 49718 79518
rect 49625 79436 49718 79502
rect 49625 79334 49718 79400
tri 49625 79318 49641 79334 ne
rect 49641 79318 49718 79334
rect 49458 79219 49606 79301
rect 49346 79186 49423 79202
tri 49423 79186 49439 79202 sw
rect 49346 79120 49439 79186
rect 49475 79061 49589 79219
tri 49625 79186 49641 79202 se
rect 49641 79186 49718 79202
rect 49625 79120 49718 79186
rect 49346 78985 49718 79061
rect 49346 78860 49439 78926
rect 49346 78844 49423 78860
tri 49423 78844 49439 78860 nw
rect 49475 78827 49589 78985
rect 49625 78860 49718 78926
tri 49625 78844 49641 78860 ne
rect 49641 78844 49718 78860
rect 49458 78745 49606 78827
rect 49346 78712 49423 78728
tri 49423 78712 49439 78728 sw
rect 49346 78646 49439 78712
rect 49346 78544 49439 78610
rect 49346 78528 49423 78544
tri 49423 78528 49439 78544 nw
rect 49475 78511 49589 78745
tri 49625 78712 49641 78728 se
rect 49641 78712 49718 78728
rect 49625 78646 49718 78712
rect 49625 78544 49718 78610
tri 49625 78528 49641 78544 ne
rect 49641 78528 49718 78544
rect 49458 78429 49606 78511
rect 49346 78396 49423 78412
tri 49423 78396 49439 78412 sw
rect 49346 78330 49439 78396
rect 49475 78271 49589 78429
tri 49625 78396 49641 78412 se
rect 49641 78396 49718 78412
rect 49625 78330 49718 78396
rect 49346 78195 49718 78271
rect 49346 78070 49439 78136
rect 49346 78054 49423 78070
tri 49423 78054 49439 78070 nw
rect 49475 78037 49589 78195
rect 49625 78070 49718 78136
tri 49625 78054 49641 78070 ne
rect 49641 78054 49718 78070
rect 49458 77955 49606 78037
rect 49346 77922 49423 77938
tri 49423 77922 49439 77938 sw
rect 49346 77856 49439 77922
rect 49346 77754 49439 77820
rect 49346 77738 49423 77754
tri 49423 77738 49439 77754 nw
rect 49475 77721 49589 77955
tri 49625 77922 49641 77938 se
rect 49641 77922 49718 77938
rect 49625 77856 49718 77922
rect 49625 77754 49718 77820
tri 49625 77738 49641 77754 ne
rect 49641 77738 49718 77754
rect 49458 77639 49606 77721
rect 49346 77606 49423 77622
tri 49423 77606 49439 77622 sw
rect 49346 77540 49439 77606
rect 49475 77481 49589 77639
tri 49625 77606 49641 77622 se
rect 49641 77606 49718 77622
rect 49625 77540 49718 77606
rect 49346 77405 49718 77481
rect 49346 77280 49439 77346
rect 49346 77264 49423 77280
tri 49423 77264 49439 77280 nw
rect 49475 77247 49589 77405
rect 49625 77280 49718 77346
tri 49625 77264 49641 77280 ne
rect 49641 77264 49718 77280
rect 49458 77165 49606 77247
rect 49346 77132 49423 77148
tri 49423 77132 49439 77148 sw
rect 49346 77066 49439 77132
rect 49346 76964 49439 77030
rect 49346 76948 49423 76964
tri 49423 76948 49439 76964 nw
rect 49475 76931 49589 77165
tri 49625 77132 49641 77148 se
rect 49641 77132 49718 77148
rect 49625 77066 49718 77132
rect 49625 76964 49718 77030
tri 49625 76948 49641 76964 ne
rect 49641 76948 49718 76964
rect 49458 76849 49606 76931
rect 49346 76816 49423 76832
tri 49423 76816 49439 76832 sw
rect 49346 76750 49439 76816
rect 49475 76691 49589 76849
tri 49625 76816 49641 76832 se
rect 49641 76816 49718 76832
rect 49625 76750 49718 76816
rect 49346 76615 49718 76691
rect 49346 76490 49439 76556
rect 49346 76474 49423 76490
tri 49423 76474 49439 76490 nw
rect 49475 76457 49589 76615
rect 49625 76490 49718 76556
tri 49625 76474 49641 76490 ne
rect 49641 76474 49718 76490
rect 49458 76375 49606 76457
rect 49346 76342 49423 76358
tri 49423 76342 49439 76358 sw
rect 49346 76276 49439 76342
rect 49346 76174 49439 76240
rect 49346 76158 49423 76174
tri 49423 76158 49439 76174 nw
rect 49475 76141 49589 76375
tri 49625 76342 49641 76358 se
rect 49641 76342 49718 76358
rect 49625 76276 49718 76342
rect 49625 76174 49718 76240
tri 49625 76158 49641 76174 ne
rect 49641 76158 49718 76174
rect 49458 76059 49606 76141
rect 49346 76026 49423 76042
tri 49423 76026 49439 76042 sw
rect 49346 75960 49439 76026
rect 49475 75901 49589 76059
tri 49625 76026 49641 76042 se
rect 49641 76026 49718 76042
rect 49625 75960 49718 76026
rect 49346 75825 49718 75901
rect 49346 75700 49439 75766
rect 49346 75684 49423 75700
tri 49423 75684 49439 75700 nw
rect 49475 75667 49589 75825
rect 49625 75700 49718 75766
tri 49625 75684 49641 75700 ne
rect 49641 75684 49718 75700
rect 49458 75585 49606 75667
rect 49346 75552 49423 75568
tri 49423 75552 49439 75568 sw
rect 49346 75486 49439 75552
rect 49346 75384 49439 75450
rect 49346 75368 49423 75384
tri 49423 75368 49439 75384 nw
rect 49475 75351 49589 75585
tri 49625 75552 49641 75568 se
rect 49641 75552 49718 75568
rect 49625 75486 49718 75552
rect 49625 75384 49718 75450
tri 49625 75368 49641 75384 ne
rect 49641 75368 49718 75384
rect 49458 75269 49606 75351
rect 49346 75236 49423 75252
tri 49423 75236 49439 75252 sw
rect 49346 75170 49439 75236
rect 49475 75111 49589 75269
tri 49625 75236 49641 75252 se
rect 49641 75236 49718 75252
rect 49625 75170 49718 75236
rect 49346 75035 49718 75111
rect 49346 74910 49439 74976
rect 49346 74894 49423 74910
tri 49423 74894 49439 74910 nw
rect 49475 74877 49589 75035
rect 49625 74910 49718 74976
tri 49625 74894 49641 74910 ne
rect 49641 74894 49718 74910
rect 49458 74795 49606 74877
rect 49346 74762 49423 74778
tri 49423 74762 49439 74778 sw
rect 49346 74696 49439 74762
rect 49346 74594 49439 74660
rect 49346 74578 49423 74594
tri 49423 74578 49439 74594 nw
rect 49475 74561 49589 74795
tri 49625 74762 49641 74778 se
rect 49641 74762 49718 74778
rect 49625 74696 49718 74762
rect 49625 74594 49718 74660
tri 49625 74578 49641 74594 ne
rect 49641 74578 49718 74594
rect 49458 74479 49606 74561
rect 49346 74446 49423 74462
tri 49423 74446 49439 74462 sw
rect 49346 74380 49439 74446
rect 49475 74321 49589 74479
tri 49625 74446 49641 74462 se
rect 49641 74446 49718 74462
rect 49625 74380 49718 74446
rect 49346 74245 49718 74321
rect 49346 74120 49439 74186
rect 49346 74104 49423 74120
tri 49423 74104 49439 74120 nw
rect 49475 74087 49589 74245
rect 49625 74120 49718 74186
tri 49625 74104 49641 74120 ne
rect 49641 74104 49718 74120
rect 49458 74005 49606 74087
rect 49346 73972 49423 73988
tri 49423 73972 49439 73988 sw
rect 49346 73906 49439 73972
rect 49346 73804 49439 73870
rect 49346 73788 49423 73804
tri 49423 73788 49439 73804 nw
rect 49475 73771 49589 74005
tri 49625 73972 49641 73988 se
rect 49641 73972 49718 73988
rect 49625 73906 49718 73972
rect 49625 73804 49718 73870
tri 49625 73788 49641 73804 ne
rect 49641 73788 49718 73804
rect 49458 73689 49606 73771
rect 49346 73656 49423 73672
tri 49423 73656 49439 73672 sw
rect 49346 73590 49439 73656
rect 49475 73531 49589 73689
tri 49625 73656 49641 73672 se
rect 49641 73656 49718 73672
rect 49625 73590 49718 73656
rect 49346 73455 49718 73531
rect 49346 73330 49439 73396
rect 49346 73314 49423 73330
tri 49423 73314 49439 73330 nw
rect 49475 73297 49589 73455
rect 49625 73330 49718 73396
tri 49625 73314 49641 73330 ne
rect 49641 73314 49718 73330
rect 49458 73215 49606 73297
rect 49346 73182 49423 73198
tri 49423 73182 49439 73198 sw
rect 49346 73116 49439 73182
rect 49346 73014 49439 73080
rect 49346 72998 49423 73014
tri 49423 72998 49439 73014 nw
rect 49475 72981 49589 73215
tri 49625 73182 49641 73198 se
rect 49641 73182 49718 73198
rect 49625 73116 49718 73182
rect 49625 73014 49718 73080
tri 49625 72998 49641 73014 ne
rect 49641 72998 49718 73014
rect 49458 72899 49606 72981
rect 49346 72866 49423 72882
tri 49423 72866 49439 72882 sw
rect 49346 72800 49439 72866
rect 49475 72741 49589 72899
tri 49625 72866 49641 72882 se
rect 49641 72866 49718 72882
rect 49625 72800 49718 72866
rect 49346 72665 49718 72741
rect 49346 72540 49439 72606
rect 49346 72524 49423 72540
tri 49423 72524 49439 72540 nw
rect 49475 72507 49589 72665
rect 49625 72540 49718 72606
tri 49625 72524 49641 72540 ne
rect 49641 72524 49718 72540
rect 49458 72425 49606 72507
rect 49346 72392 49423 72408
tri 49423 72392 49439 72408 sw
rect 49346 72326 49439 72392
rect 49346 72224 49439 72290
rect 49346 72208 49423 72224
tri 49423 72208 49439 72224 nw
rect 49475 72191 49589 72425
tri 49625 72392 49641 72408 se
rect 49641 72392 49718 72408
rect 49625 72326 49718 72392
rect 49625 72224 49718 72290
tri 49625 72208 49641 72224 ne
rect 49641 72208 49718 72224
rect 49458 72109 49606 72191
rect 49346 72076 49423 72092
tri 49423 72076 49439 72092 sw
rect 49346 72010 49439 72076
rect 49475 71951 49589 72109
tri 49625 72076 49641 72092 se
rect 49641 72076 49718 72092
rect 49625 72010 49718 72076
rect 49346 71875 49718 71951
rect 49346 71750 49439 71816
rect 49346 71734 49423 71750
tri 49423 71734 49439 71750 nw
rect 49475 71717 49589 71875
rect 49625 71750 49718 71816
tri 49625 71734 49641 71750 ne
rect 49641 71734 49718 71750
rect 49458 71635 49606 71717
rect 49346 71602 49423 71618
tri 49423 71602 49439 71618 sw
rect 49346 71536 49439 71602
rect 49346 71434 49439 71500
rect 49346 71418 49423 71434
tri 49423 71418 49439 71434 nw
rect 49475 71401 49589 71635
tri 49625 71602 49641 71618 se
rect 49641 71602 49718 71618
rect 49625 71536 49718 71602
rect 49625 71434 49718 71500
tri 49625 71418 49641 71434 ne
rect 49641 71418 49718 71434
rect 49458 71319 49606 71401
rect 49346 71286 49423 71302
tri 49423 71286 49439 71302 sw
rect 49346 71220 49439 71286
rect 49475 71161 49589 71319
tri 49625 71286 49641 71302 se
rect 49641 71286 49718 71302
rect 49625 71220 49718 71286
rect 49346 71085 49718 71161
rect 49346 70960 49439 71026
rect 49346 70944 49423 70960
tri 49423 70944 49439 70960 nw
rect 49475 70927 49589 71085
rect 49625 70960 49718 71026
tri 49625 70944 49641 70960 ne
rect 49641 70944 49718 70960
rect 49458 70845 49606 70927
rect 49346 70812 49423 70828
tri 49423 70812 49439 70828 sw
rect 49346 70746 49439 70812
rect 49346 70644 49439 70710
rect 49346 70628 49423 70644
tri 49423 70628 49439 70644 nw
rect 49475 70611 49589 70845
tri 49625 70812 49641 70828 se
rect 49641 70812 49718 70828
rect 49625 70746 49718 70812
rect 49625 70644 49718 70710
tri 49625 70628 49641 70644 ne
rect 49641 70628 49718 70644
rect 49458 70529 49606 70611
rect 49346 70496 49423 70512
tri 49423 70496 49439 70512 sw
rect 49346 70430 49439 70496
rect 49475 70371 49589 70529
tri 49625 70496 49641 70512 se
rect 49641 70496 49718 70512
rect 49625 70430 49718 70496
rect 49346 70295 49718 70371
rect 49346 70170 49439 70236
rect 49346 70154 49423 70170
tri 49423 70154 49439 70170 nw
rect 49475 70137 49589 70295
rect 49625 70170 49718 70236
tri 49625 70154 49641 70170 ne
rect 49641 70154 49718 70170
rect 49458 70055 49606 70137
rect 49346 70022 49423 70038
tri 49423 70022 49439 70038 sw
rect 49346 69956 49439 70022
rect 49346 69854 49439 69920
rect 49346 69838 49423 69854
tri 49423 69838 49439 69854 nw
rect 49475 69821 49589 70055
tri 49625 70022 49641 70038 se
rect 49641 70022 49718 70038
rect 49625 69956 49718 70022
rect 49625 69854 49718 69920
tri 49625 69838 49641 69854 ne
rect 49641 69838 49718 69854
rect 49458 69739 49606 69821
rect 49346 69706 49423 69722
tri 49423 69706 49439 69722 sw
rect 49346 69640 49439 69706
rect 49475 69581 49589 69739
tri 49625 69706 49641 69722 se
rect 49641 69706 49718 69722
rect 49625 69640 49718 69706
rect 49346 69505 49718 69581
rect 49346 69380 49439 69446
rect 49346 69364 49423 69380
tri 49423 69364 49439 69380 nw
rect 49475 69347 49589 69505
rect 49625 69380 49718 69446
tri 49625 69364 49641 69380 ne
rect 49641 69364 49718 69380
rect 49458 69265 49606 69347
rect 49346 69232 49423 69248
tri 49423 69232 49439 69248 sw
rect 49346 69166 49439 69232
rect 49346 69064 49439 69130
rect 49346 69048 49423 69064
tri 49423 69048 49439 69064 nw
rect 49475 69031 49589 69265
tri 49625 69232 49641 69248 se
rect 49641 69232 49718 69248
rect 49625 69166 49718 69232
rect 49625 69064 49718 69130
tri 49625 69048 49641 69064 ne
rect 49641 69048 49718 69064
rect 49458 68949 49606 69031
rect 49346 68916 49423 68932
tri 49423 68916 49439 68932 sw
rect 49346 68850 49439 68916
rect 49475 68791 49589 68949
tri 49625 68916 49641 68932 se
rect 49641 68916 49718 68932
rect 49625 68850 49718 68916
rect 49346 68715 49718 68791
rect 49346 68590 49439 68656
rect 49346 68574 49423 68590
tri 49423 68574 49439 68590 nw
rect 49475 68557 49589 68715
rect 49625 68590 49718 68656
tri 49625 68574 49641 68590 ne
rect 49641 68574 49718 68590
rect 49458 68475 49606 68557
rect 49346 68442 49423 68458
tri 49423 68442 49439 68458 sw
rect 49346 68376 49439 68442
rect 49346 68274 49439 68340
rect 49346 68258 49423 68274
tri 49423 68258 49439 68274 nw
rect 49475 68241 49589 68475
tri 49625 68442 49641 68458 se
rect 49641 68442 49718 68458
rect 49625 68376 49718 68442
rect 49625 68274 49718 68340
tri 49625 68258 49641 68274 ne
rect 49641 68258 49718 68274
rect 49458 68159 49606 68241
rect 49346 68126 49423 68142
tri 49423 68126 49439 68142 sw
rect 49346 68060 49439 68126
rect 49475 68001 49589 68159
tri 49625 68126 49641 68142 se
rect 49641 68126 49718 68142
rect 49625 68060 49718 68126
rect 49346 67925 49718 68001
rect 49346 67800 49439 67866
rect 49346 67784 49423 67800
tri 49423 67784 49439 67800 nw
rect 49475 67767 49589 67925
rect 49625 67800 49718 67866
tri 49625 67784 49641 67800 ne
rect 49641 67784 49718 67800
rect 49458 67685 49606 67767
rect 49346 67652 49423 67668
tri 49423 67652 49439 67668 sw
rect 49346 67586 49439 67652
rect 49346 67484 49439 67550
rect 49346 67468 49423 67484
tri 49423 67468 49439 67484 nw
rect 49475 67451 49589 67685
tri 49625 67652 49641 67668 se
rect 49641 67652 49718 67668
rect 49625 67586 49718 67652
rect 49625 67484 49718 67550
tri 49625 67468 49641 67484 ne
rect 49641 67468 49718 67484
rect 49458 67369 49606 67451
rect 49346 67336 49423 67352
tri 49423 67336 49439 67352 sw
rect 49346 67270 49439 67336
rect 49475 67211 49589 67369
tri 49625 67336 49641 67352 se
rect 49641 67336 49718 67352
rect 49625 67270 49718 67336
rect 49346 67135 49718 67211
rect 49346 67010 49439 67076
rect 49346 66994 49423 67010
tri 49423 66994 49439 67010 nw
rect 49475 66977 49589 67135
rect 49625 67010 49718 67076
tri 49625 66994 49641 67010 ne
rect 49641 66994 49718 67010
rect 49458 66895 49606 66977
rect 49346 66862 49423 66878
tri 49423 66862 49439 66878 sw
rect 49346 66796 49439 66862
rect 49346 66694 49439 66760
rect 49346 66678 49423 66694
tri 49423 66678 49439 66694 nw
rect 49475 66661 49589 66895
tri 49625 66862 49641 66878 se
rect 49641 66862 49718 66878
rect 49625 66796 49718 66862
rect 49625 66694 49718 66760
tri 49625 66678 49641 66694 ne
rect 49641 66678 49718 66694
rect 49458 66579 49606 66661
rect 49346 66546 49423 66562
tri 49423 66546 49439 66562 sw
rect 49346 66480 49439 66546
rect 49475 66421 49589 66579
tri 49625 66546 49641 66562 se
rect 49641 66546 49718 66562
rect 49625 66480 49718 66546
rect 49346 66345 49718 66421
rect 49346 66220 49439 66286
rect 49346 66204 49423 66220
tri 49423 66204 49439 66220 nw
rect 49475 66187 49589 66345
rect 49625 66220 49718 66286
tri 49625 66204 49641 66220 ne
rect 49641 66204 49718 66220
rect 49458 66105 49606 66187
rect 49346 66072 49423 66088
tri 49423 66072 49439 66088 sw
rect 49346 66006 49439 66072
rect 49346 65904 49439 65970
rect 49346 65888 49423 65904
tri 49423 65888 49439 65904 nw
rect 49475 65871 49589 66105
tri 49625 66072 49641 66088 se
rect 49641 66072 49718 66088
rect 49625 66006 49718 66072
rect 49625 65904 49718 65970
tri 49625 65888 49641 65904 ne
rect 49641 65888 49718 65904
rect 49458 65789 49606 65871
rect 49346 65756 49423 65772
tri 49423 65756 49439 65772 sw
rect 49346 65690 49439 65756
rect 49475 65631 49589 65789
tri 49625 65756 49641 65772 se
rect 49641 65756 49718 65772
rect 49625 65690 49718 65756
rect 49346 65555 49718 65631
rect 49346 65430 49439 65496
rect 49346 65414 49423 65430
tri 49423 65414 49439 65430 nw
rect 49475 65397 49589 65555
rect 49625 65430 49718 65496
tri 49625 65414 49641 65430 ne
rect 49641 65414 49718 65430
rect 49458 65315 49606 65397
rect 49346 65282 49423 65298
tri 49423 65282 49439 65298 sw
rect 49346 65216 49439 65282
rect 49346 65114 49439 65180
rect 49346 65098 49423 65114
tri 49423 65098 49439 65114 nw
rect 49475 65081 49589 65315
tri 49625 65282 49641 65298 se
rect 49641 65282 49718 65298
rect 49625 65216 49718 65282
rect 49625 65114 49718 65180
tri 49625 65098 49641 65114 ne
rect 49641 65098 49718 65114
rect 49458 64999 49606 65081
rect 49346 64966 49423 64982
tri 49423 64966 49439 64982 sw
rect 49346 64900 49439 64966
rect 49475 64841 49589 64999
tri 49625 64966 49641 64982 se
rect 49641 64966 49718 64982
rect 49625 64900 49718 64966
rect 49346 64765 49718 64841
rect 49346 64640 49439 64706
rect 49346 64624 49423 64640
tri 49423 64624 49439 64640 nw
rect 49475 64607 49589 64765
rect 49625 64640 49718 64706
tri 49625 64624 49641 64640 ne
rect 49641 64624 49718 64640
rect 49458 64525 49606 64607
rect 49346 64492 49423 64508
tri 49423 64492 49439 64508 sw
rect 49346 64426 49439 64492
rect 49346 64324 49439 64390
rect 49346 64308 49423 64324
tri 49423 64308 49439 64324 nw
rect 49475 64291 49589 64525
tri 49625 64492 49641 64508 se
rect 49641 64492 49718 64508
rect 49625 64426 49718 64492
rect 49625 64324 49718 64390
tri 49625 64308 49641 64324 ne
rect 49641 64308 49718 64324
rect 49458 64209 49606 64291
rect 49346 64176 49423 64192
tri 49423 64176 49439 64192 sw
rect 49346 64110 49439 64176
rect 49475 64051 49589 64209
tri 49625 64176 49641 64192 se
rect 49641 64176 49718 64192
rect 49625 64110 49718 64176
rect 49346 63975 49718 64051
rect 49346 63850 49439 63916
rect 49346 63834 49423 63850
tri 49423 63834 49439 63850 nw
rect 49475 63817 49589 63975
rect 49625 63850 49718 63916
tri 49625 63834 49641 63850 ne
rect 49641 63834 49718 63850
rect 49458 63735 49606 63817
rect 49346 63702 49423 63718
tri 49423 63702 49439 63718 sw
rect 49346 63636 49439 63702
rect 49346 63534 49439 63600
rect 49346 63518 49423 63534
tri 49423 63518 49439 63534 nw
rect 49475 63501 49589 63735
tri 49625 63702 49641 63718 se
rect 49641 63702 49718 63718
rect 49625 63636 49718 63702
rect 49625 63534 49718 63600
tri 49625 63518 49641 63534 ne
rect 49641 63518 49718 63534
rect 49458 63419 49606 63501
rect 49346 63386 49423 63402
tri 49423 63386 49439 63402 sw
rect 49346 63320 49439 63386
rect 49475 63261 49589 63419
tri 49625 63386 49641 63402 se
rect 49641 63386 49718 63402
rect 49625 63320 49718 63386
rect 49346 63185 49718 63261
rect 49346 63060 49439 63126
rect 49346 63044 49423 63060
tri 49423 63044 49439 63060 nw
rect 49475 63027 49589 63185
rect 49625 63060 49718 63126
tri 49625 63044 49641 63060 ne
rect 49641 63044 49718 63060
rect 49458 62945 49606 63027
rect 49346 62912 49423 62928
tri 49423 62912 49439 62928 sw
rect 49346 62846 49439 62912
rect 49346 62744 49439 62810
rect 49346 62728 49423 62744
tri 49423 62728 49439 62744 nw
rect 49475 62711 49589 62945
tri 49625 62912 49641 62928 se
rect 49641 62912 49718 62928
rect 49625 62846 49718 62912
rect 49625 62744 49718 62810
tri 49625 62728 49641 62744 ne
rect 49641 62728 49718 62744
rect 49458 62629 49606 62711
rect 49346 62596 49423 62612
tri 49423 62596 49439 62612 sw
rect 49346 62530 49439 62596
rect 49475 62471 49589 62629
tri 49625 62596 49641 62612 se
rect 49641 62596 49718 62612
rect 49625 62530 49718 62596
rect 49346 62395 49718 62471
rect 49346 62270 49439 62336
rect 49346 62254 49423 62270
tri 49423 62254 49439 62270 nw
rect 49475 62237 49589 62395
rect 49625 62270 49718 62336
tri 49625 62254 49641 62270 ne
rect 49641 62254 49718 62270
rect 49458 62155 49606 62237
rect 49346 62122 49423 62138
tri 49423 62122 49439 62138 sw
rect 49346 62056 49439 62122
rect 49346 61954 49439 62020
rect 49346 61938 49423 61954
tri 49423 61938 49439 61954 nw
rect 49475 61921 49589 62155
tri 49625 62122 49641 62138 se
rect 49641 62122 49718 62138
rect 49625 62056 49718 62122
rect 49625 61954 49718 62020
tri 49625 61938 49641 61954 ne
rect 49641 61938 49718 61954
rect 49458 61839 49606 61921
rect 49346 61806 49423 61822
tri 49423 61806 49439 61822 sw
rect 49346 61740 49439 61806
rect 49475 61681 49589 61839
tri 49625 61806 49641 61822 se
rect 49641 61806 49718 61822
rect 49625 61740 49718 61806
rect 49346 61605 49718 61681
rect 49346 61480 49439 61546
rect 49346 61464 49423 61480
tri 49423 61464 49439 61480 nw
rect 49475 61447 49589 61605
rect 49625 61480 49718 61546
tri 49625 61464 49641 61480 ne
rect 49641 61464 49718 61480
rect 49458 61365 49606 61447
rect 49346 61332 49423 61348
tri 49423 61332 49439 61348 sw
rect 49346 61266 49439 61332
rect 49346 61164 49439 61230
rect 49346 61148 49423 61164
tri 49423 61148 49439 61164 nw
rect 49475 61131 49589 61365
tri 49625 61332 49641 61348 se
rect 49641 61332 49718 61348
rect 49625 61266 49718 61332
rect 49625 61164 49718 61230
tri 49625 61148 49641 61164 ne
rect 49641 61148 49718 61164
rect 49458 61049 49606 61131
rect 49346 61016 49423 61032
tri 49423 61016 49439 61032 sw
rect 49346 60950 49439 61016
rect 49475 60891 49589 61049
tri 49625 61016 49641 61032 se
rect 49641 61016 49718 61032
rect 49625 60950 49718 61016
rect 49346 60815 49718 60891
rect 49346 60690 49439 60756
rect 49346 60674 49423 60690
tri 49423 60674 49439 60690 nw
rect 49475 60657 49589 60815
rect 49625 60690 49718 60756
tri 49625 60674 49641 60690 ne
rect 49641 60674 49718 60690
rect 49458 60575 49606 60657
rect 49346 60542 49423 60558
tri 49423 60542 49439 60558 sw
rect 49346 60476 49439 60542
rect 49346 60374 49439 60440
rect 49346 60358 49423 60374
tri 49423 60358 49439 60374 nw
rect 49475 60341 49589 60575
tri 49625 60542 49641 60558 se
rect 49641 60542 49718 60558
rect 49625 60476 49718 60542
rect 49625 60374 49718 60440
tri 49625 60358 49641 60374 ne
rect 49641 60358 49718 60374
rect 49458 60259 49606 60341
rect 49346 60226 49423 60242
tri 49423 60226 49439 60242 sw
rect 49346 60160 49439 60226
rect 49475 60101 49589 60259
tri 49625 60226 49641 60242 se
rect 49641 60226 49718 60242
rect 49625 60160 49718 60226
rect 49346 60025 49718 60101
rect 49346 59900 49439 59966
rect 49346 59884 49423 59900
tri 49423 59884 49439 59900 nw
rect 49475 59867 49589 60025
rect 49625 59900 49718 59966
tri 49625 59884 49641 59900 ne
rect 49641 59884 49718 59900
rect 49458 59785 49606 59867
rect 49346 59752 49423 59768
tri 49423 59752 49439 59768 sw
rect 49346 59686 49439 59752
rect 49346 59584 49439 59650
rect 49346 59568 49423 59584
tri 49423 59568 49439 59584 nw
rect 49475 59551 49589 59785
tri 49625 59752 49641 59768 se
rect 49641 59752 49718 59768
rect 49625 59686 49718 59752
rect 49625 59584 49718 59650
tri 49625 59568 49641 59584 ne
rect 49641 59568 49718 59584
rect 49458 59469 49606 59551
rect 49346 59436 49423 59452
tri 49423 59436 49439 59452 sw
rect 49346 59370 49439 59436
rect 49475 59311 49589 59469
tri 49625 59436 49641 59452 se
rect 49641 59436 49718 59452
rect 49625 59370 49718 59436
rect 49346 59235 49718 59311
rect 49346 59110 49439 59176
rect 49346 59094 49423 59110
tri 49423 59094 49439 59110 nw
rect 49475 59077 49589 59235
rect 49625 59110 49718 59176
tri 49625 59094 49641 59110 ne
rect 49641 59094 49718 59110
rect 49458 58995 49606 59077
rect 49346 58962 49423 58978
tri 49423 58962 49439 58978 sw
rect 49346 58896 49439 58962
rect 49346 58794 49439 58860
rect 49346 58778 49423 58794
tri 49423 58778 49439 58794 nw
rect 49475 58761 49589 58995
tri 49625 58962 49641 58978 se
rect 49641 58962 49718 58978
rect 49625 58896 49718 58962
rect 49625 58794 49718 58860
tri 49625 58778 49641 58794 ne
rect 49641 58778 49718 58794
rect 49458 58679 49606 58761
rect 49346 58646 49423 58662
tri 49423 58646 49439 58662 sw
rect 49346 58580 49439 58646
rect 49475 58521 49589 58679
tri 49625 58646 49641 58662 se
rect 49641 58646 49718 58662
rect 49625 58580 49718 58646
rect 49346 58445 49718 58521
rect 49346 58320 49439 58386
rect 49346 58304 49423 58320
tri 49423 58304 49439 58320 nw
rect 49475 58287 49589 58445
rect 49625 58320 49718 58386
tri 49625 58304 49641 58320 ne
rect 49641 58304 49718 58320
rect 49458 58205 49606 58287
rect 49346 58172 49423 58188
tri 49423 58172 49439 58188 sw
rect 49346 58106 49439 58172
rect 49346 58004 49439 58070
rect 49346 57988 49423 58004
tri 49423 57988 49439 58004 nw
rect 49475 57971 49589 58205
tri 49625 58172 49641 58188 se
rect 49641 58172 49718 58188
rect 49625 58106 49718 58172
rect 49625 58004 49718 58070
tri 49625 57988 49641 58004 ne
rect 49641 57988 49718 58004
rect 49458 57889 49606 57971
rect 49346 57856 49423 57872
tri 49423 57856 49439 57872 sw
rect 49346 57790 49439 57856
rect 49475 57731 49589 57889
tri 49625 57856 49641 57872 se
rect 49641 57856 49718 57872
rect 49625 57790 49718 57856
rect 49346 57655 49718 57731
rect 49346 57530 49439 57596
rect 49346 57514 49423 57530
tri 49423 57514 49439 57530 nw
rect 49475 57497 49589 57655
rect 49625 57530 49718 57596
tri 49625 57514 49641 57530 ne
rect 49641 57514 49718 57530
rect 49458 57415 49606 57497
rect 49346 57382 49423 57398
tri 49423 57382 49439 57398 sw
rect 49346 57316 49439 57382
rect 49346 57214 49439 57280
rect 49346 57198 49423 57214
tri 49423 57198 49439 57214 nw
rect 49475 57181 49589 57415
tri 49625 57382 49641 57398 se
rect 49641 57382 49718 57398
rect 49625 57316 49718 57382
rect 49625 57214 49718 57280
tri 49625 57198 49641 57214 ne
rect 49641 57198 49718 57214
rect 49458 57099 49606 57181
rect 49346 57066 49423 57082
tri 49423 57066 49439 57082 sw
rect 49346 57000 49439 57066
rect 49475 56941 49589 57099
tri 49625 57066 49641 57082 se
rect 49641 57066 49718 57082
rect 49625 57000 49718 57066
rect 49346 56865 49718 56941
rect 49346 56740 49439 56806
rect 49346 56724 49423 56740
tri 49423 56724 49439 56740 nw
rect 49475 56707 49589 56865
rect 49625 56740 49718 56806
tri 49625 56724 49641 56740 ne
rect 49641 56724 49718 56740
rect 49458 56625 49606 56707
rect 49346 56592 49423 56608
tri 49423 56592 49439 56608 sw
rect 49346 56526 49439 56592
rect 49346 56424 49439 56490
rect 49346 56408 49423 56424
tri 49423 56408 49439 56424 nw
rect 49475 56391 49589 56625
tri 49625 56592 49641 56608 se
rect 49641 56592 49718 56608
rect 49625 56526 49718 56592
rect 49625 56424 49718 56490
tri 49625 56408 49641 56424 ne
rect 49641 56408 49718 56424
rect 49458 56309 49606 56391
rect 49346 56276 49423 56292
tri 49423 56276 49439 56292 sw
rect 49346 56210 49439 56276
rect 49475 56151 49589 56309
tri 49625 56276 49641 56292 se
rect 49641 56276 49718 56292
rect 49625 56210 49718 56276
rect 49346 56075 49718 56151
rect 49346 55950 49439 56016
rect 49346 55934 49423 55950
tri 49423 55934 49439 55950 nw
rect 49475 55917 49589 56075
rect 49625 55950 49718 56016
tri 49625 55934 49641 55950 ne
rect 49641 55934 49718 55950
rect 49458 55835 49606 55917
rect 49346 55802 49423 55818
tri 49423 55802 49439 55818 sw
rect 49346 55736 49439 55802
rect 49346 55634 49439 55700
rect 49346 55618 49423 55634
tri 49423 55618 49439 55634 nw
rect 49475 55601 49589 55835
tri 49625 55802 49641 55818 se
rect 49641 55802 49718 55818
rect 49625 55736 49718 55802
rect 49625 55634 49718 55700
tri 49625 55618 49641 55634 ne
rect 49641 55618 49718 55634
rect 49458 55519 49606 55601
rect 49346 55486 49423 55502
tri 49423 55486 49439 55502 sw
rect 49346 55420 49439 55486
rect 49475 55361 49589 55519
tri 49625 55486 49641 55502 se
rect 49641 55486 49718 55502
rect 49625 55420 49718 55486
rect 49346 55285 49718 55361
rect 49346 55160 49439 55226
rect 49346 55144 49423 55160
tri 49423 55144 49439 55160 nw
rect 49475 55127 49589 55285
rect 49625 55160 49718 55226
tri 49625 55144 49641 55160 ne
rect 49641 55144 49718 55160
rect 49458 55045 49606 55127
rect 49346 55012 49423 55028
tri 49423 55012 49439 55028 sw
rect 49346 54946 49439 55012
rect 49346 54844 49439 54910
rect 49346 54828 49423 54844
tri 49423 54828 49439 54844 nw
rect 49475 54811 49589 55045
tri 49625 55012 49641 55028 se
rect 49641 55012 49718 55028
rect 49625 54946 49718 55012
rect 49625 54844 49718 54910
tri 49625 54828 49641 54844 ne
rect 49641 54828 49718 54844
rect 49458 54729 49606 54811
rect 49346 54696 49423 54712
tri 49423 54696 49439 54712 sw
rect 49346 54630 49439 54696
rect 49475 54571 49589 54729
tri 49625 54696 49641 54712 se
rect 49641 54696 49718 54712
rect 49625 54630 49718 54696
rect 49346 54495 49718 54571
rect 49346 54370 49439 54436
rect 49346 54354 49423 54370
tri 49423 54354 49439 54370 nw
rect 49475 54337 49589 54495
rect 49625 54370 49718 54436
tri 49625 54354 49641 54370 ne
rect 49641 54354 49718 54370
rect 49458 54255 49606 54337
rect 49346 54222 49423 54238
tri 49423 54222 49439 54238 sw
rect 49346 54156 49439 54222
rect 49346 54054 49439 54120
rect 49346 54038 49423 54054
tri 49423 54038 49439 54054 nw
rect 49475 54021 49589 54255
tri 49625 54222 49641 54238 se
rect 49641 54222 49718 54238
rect 49625 54156 49718 54222
rect 49625 54054 49718 54120
tri 49625 54038 49641 54054 ne
rect 49641 54038 49718 54054
rect 49458 53939 49606 54021
rect 49346 53906 49423 53922
tri 49423 53906 49439 53922 sw
rect 49346 53840 49439 53906
rect 49475 53781 49589 53939
tri 49625 53906 49641 53922 se
rect 49641 53906 49718 53922
rect 49625 53840 49718 53906
rect 49346 53705 49718 53781
rect 49346 53580 49439 53646
rect 49346 53564 49423 53580
tri 49423 53564 49439 53580 nw
rect 49475 53547 49589 53705
rect 49625 53580 49718 53646
tri 49625 53564 49641 53580 ne
rect 49641 53564 49718 53580
rect 49458 53465 49606 53547
rect 49346 53432 49423 53448
tri 49423 53432 49439 53448 sw
rect 49346 53366 49439 53432
rect 49346 53264 49439 53330
rect 49346 53248 49423 53264
tri 49423 53248 49439 53264 nw
rect 49475 53231 49589 53465
tri 49625 53432 49641 53448 se
rect 49641 53432 49718 53448
rect 49625 53366 49718 53432
rect 49625 53264 49718 53330
tri 49625 53248 49641 53264 ne
rect 49641 53248 49718 53264
rect 49458 53149 49606 53231
rect 49346 53116 49423 53132
tri 49423 53116 49439 53132 sw
rect 49346 53050 49439 53116
rect 49475 52991 49589 53149
tri 49625 53116 49641 53132 se
rect 49641 53116 49718 53132
rect 49625 53050 49718 53116
rect 49346 52915 49718 52991
rect 49346 52790 49439 52856
rect 49346 52774 49423 52790
tri 49423 52774 49439 52790 nw
rect 49475 52757 49589 52915
rect 49625 52790 49718 52856
tri 49625 52774 49641 52790 ne
rect 49641 52774 49718 52790
rect 49458 52675 49606 52757
rect 49346 52642 49423 52658
tri 49423 52642 49439 52658 sw
rect 49346 52576 49439 52642
rect 49346 52474 49439 52540
rect 49346 52458 49423 52474
tri 49423 52458 49439 52474 nw
rect 49475 52441 49589 52675
tri 49625 52642 49641 52658 se
rect 49641 52642 49718 52658
rect 49625 52576 49718 52642
rect 49625 52474 49718 52540
tri 49625 52458 49641 52474 ne
rect 49641 52458 49718 52474
rect 49458 52359 49606 52441
rect 49346 52326 49423 52342
tri 49423 52326 49439 52342 sw
rect 49346 52260 49439 52326
rect 49475 52201 49589 52359
tri 49625 52326 49641 52342 se
rect 49641 52326 49718 52342
rect 49625 52260 49718 52326
rect 49346 52125 49718 52201
rect 49346 52000 49439 52066
rect 49346 51984 49423 52000
tri 49423 51984 49439 52000 nw
rect 49475 51967 49589 52125
rect 49625 52000 49718 52066
tri 49625 51984 49641 52000 ne
rect 49641 51984 49718 52000
rect 49458 51885 49606 51967
rect 49346 51852 49423 51868
tri 49423 51852 49439 51868 sw
rect 49346 51786 49439 51852
rect 49346 51684 49439 51750
rect 49346 51668 49423 51684
tri 49423 51668 49439 51684 nw
rect 49475 51651 49589 51885
tri 49625 51852 49641 51868 se
rect 49641 51852 49718 51868
rect 49625 51786 49718 51852
rect 49625 51684 49718 51750
tri 49625 51668 49641 51684 ne
rect 49641 51668 49718 51684
rect 49458 51569 49606 51651
rect 49346 51536 49423 51552
tri 49423 51536 49439 51552 sw
rect 49346 51470 49439 51536
rect 49475 51411 49589 51569
tri 49625 51536 49641 51552 se
rect 49641 51536 49718 51552
rect 49625 51470 49718 51536
rect 49346 51335 49718 51411
rect 49346 51210 49439 51276
rect 49346 51194 49423 51210
tri 49423 51194 49439 51210 nw
rect 49475 51177 49589 51335
rect 49625 51210 49718 51276
tri 49625 51194 49641 51210 ne
rect 49641 51194 49718 51210
rect 49458 51095 49606 51177
rect 49346 51062 49423 51078
tri 49423 51062 49439 51078 sw
rect 49346 50996 49439 51062
rect 49346 50894 49439 50960
rect 49346 50878 49423 50894
tri 49423 50878 49439 50894 nw
rect 49475 50861 49589 51095
tri 49625 51062 49641 51078 se
rect 49641 51062 49718 51078
rect 49625 50996 49718 51062
rect 49625 50894 49718 50960
tri 49625 50878 49641 50894 ne
rect 49641 50878 49718 50894
rect 49458 50779 49606 50861
rect 49346 50746 49423 50762
tri 49423 50746 49439 50762 sw
rect 49346 50680 49439 50746
rect 49475 50621 49589 50779
tri 49625 50746 49641 50762 se
rect 49641 50746 49718 50762
rect 49625 50680 49718 50746
rect 49346 50545 49718 50621
rect 49346 50420 49439 50486
rect 49346 50404 49423 50420
tri 49423 50404 49439 50420 nw
rect 49475 50387 49589 50545
rect 49625 50420 49718 50486
tri 49625 50404 49641 50420 ne
rect 49641 50404 49718 50420
rect 49458 50305 49606 50387
rect 49346 50272 49423 50288
tri 49423 50272 49439 50288 sw
rect 49346 50206 49439 50272
rect 49346 50104 49439 50170
rect 49346 50088 49423 50104
tri 49423 50088 49439 50104 nw
rect 49475 50071 49589 50305
tri 49625 50272 49641 50288 se
rect 49641 50272 49718 50288
rect 49625 50206 49718 50272
rect 49625 50104 49718 50170
tri 49625 50088 49641 50104 ne
rect 49641 50088 49718 50104
rect 49458 49989 49606 50071
rect 49346 49956 49423 49972
tri 49423 49956 49439 49972 sw
rect 49346 49890 49439 49956
rect 49475 49831 49589 49989
tri 49625 49956 49641 49972 se
rect 49641 49956 49718 49972
rect 49625 49890 49718 49956
rect 49346 49755 49718 49831
rect 49346 49630 49439 49696
rect 49346 49614 49423 49630
tri 49423 49614 49439 49630 nw
rect 49475 49597 49589 49755
rect 49625 49630 49718 49696
tri 49625 49614 49641 49630 ne
rect 49641 49614 49718 49630
rect 49458 49515 49606 49597
rect 49346 49482 49423 49498
tri 49423 49482 49439 49498 sw
rect 49346 49416 49439 49482
rect 49346 49314 49439 49380
rect 49346 49298 49423 49314
tri 49423 49298 49439 49314 nw
rect 49475 49281 49589 49515
tri 49625 49482 49641 49498 se
rect 49641 49482 49718 49498
rect 49625 49416 49718 49482
rect 49625 49314 49718 49380
tri 49625 49298 49641 49314 ne
rect 49641 49298 49718 49314
rect 49458 49199 49606 49281
rect 49346 49166 49423 49182
tri 49423 49166 49439 49182 sw
rect 49346 49100 49439 49166
rect 49475 49041 49589 49199
tri 49625 49166 49641 49182 se
rect 49641 49166 49718 49182
rect 49625 49100 49718 49166
rect 49346 48965 49718 49041
rect 49346 48840 49439 48906
rect 49346 48824 49423 48840
tri 49423 48824 49439 48840 nw
rect 49475 48807 49589 48965
rect 49625 48840 49718 48906
tri 49625 48824 49641 48840 ne
rect 49641 48824 49718 48840
rect 49458 48725 49606 48807
rect 49346 48692 49423 48708
tri 49423 48692 49439 48708 sw
rect 49346 48626 49439 48692
rect 49346 48524 49439 48590
rect 49346 48508 49423 48524
tri 49423 48508 49439 48524 nw
rect 49475 48491 49589 48725
tri 49625 48692 49641 48708 se
rect 49641 48692 49718 48708
rect 49625 48626 49718 48692
rect 49625 48524 49718 48590
tri 49625 48508 49641 48524 ne
rect 49641 48508 49718 48524
rect 49458 48409 49606 48491
rect 49346 48376 49423 48392
tri 49423 48376 49439 48392 sw
rect 49346 48310 49439 48376
rect 49475 48251 49589 48409
tri 49625 48376 49641 48392 se
rect 49641 48376 49718 48392
rect 49625 48310 49718 48376
rect 49346 48175 49718 48251
rect 49346 48050 49439 48116
rect 49346 48034 49423 48050
tri 49423 48034 49439 48050 nw
rect 49475 48017 49589 48175
rect 49625 48050 49718 48116
tri 49625 48034 49641 48050 ne
rect 49641 48034 49718 48050
rect 49458 47935 49606 48017
rect 49346 47902 49423 47918
tri 49423 47902 49439 47918 sw
rect 49346 47836 49439 47902
rect 49346 47734 49439 47800
rect 49346 47718 49423 47734
tri 49423 47718 49439 47734 nw
rect 49475 47701 49589 47935
tri 49625 47902 49641 47918 se
rect 49641 47902 49718 47918
rect 49625 47836 49718 47902
rect 49625 47734 49718 47800
tri 49625 47718 49641 47734 ne
rect 49641 47718 49718 47734
rect 49458 47619 49606 47701
rect 49346 47586 49423 47602
tri 49423 47586 49439 47602 sw
rect 49346 47520 49439 47586
rect 49475 47461 49589 47619
tri 49625 47586 49641 47602 se
rect 49641 47586 49718 47602
rect 49625 47520 49718 47586
rect 49346 47385 49718 47461
rect 49346 47260 49439 47326
rect 49346 47244 49423 47260
tri 49423 47244 49439 47260 nw
rect 49475 47227 49589 47385
rect 49625 47260 49718 47326
tri 49625 47244 49641 47260 ne
rect 49641 47244 49718 47260
rect 49458 47145 49606 47227
rect 49346 47112 49423 47128
tri 49423 47112 49439 47128 sw
rect 49346 47046 49439 47112
rect 49346 46944 49439 47010
rect 49346 46928 49423 46944
tri 49423 46928 49439 46944 nw
rect 49475 46911 49589 47145
tri 49625 47112 49641 47128 se
rect 49641 47112 49718 47128
rect 49625 47046 49718 47112
rect 49625 46944 49718 47010
tri 49625 46928 49641 46944 ne
rect 49641 46928 49718 46944
rect 49458 46829 49606 46911
rect 49346 46796 49423 46812
tri 49423 46796 49439 46812 sw
rect 49346 46730 49439 46796
rect 49475 46671 49589 46829
tri 49625 46796 49641 46812 se
rect 49641 46796 49718 46812
rect 49625 46730 49718 46796
rect 49346 46595 49718 46671
rect 49346 46470 49439 46536
rect 49346 46454 49423 46470
tri 49423 46454 49439 46470 nw
rect 49475 46437 49589 46595
rect 49625 46470 49718 46536
tri 49625 46454 49641 46470 ne
rect 49641 46454 49718 46470
rect 49458 46355 49606 46437
rect 49346 46322 49423 46338
tri 49423 46322 49439 46338 sw
rect 49346 46256 49439 46322
rect 49346 46154 49439 46220
rect 49346 46138 49423 46154
tri 49423 46138 49439 46154 nw
rect 49475 46121 49589 46355
tri 49625 46322 49641 46338 se
rect 49641 46322 49718 46338
rect 49625 46256 49718 46322
rect 49625 46154 49718 46220
tri 49625 46138 49641 46154 ne
rect 49641 46138 49718 46154
rect 49458 46039 49606 46121
rect 49346 46006 49423 46022
tri 49423 46006 49439 46022 sw
rect 49346 45940 49439 46006
rect 49475 45881 49589 46039
tri 49625 46006 49641 46022 se
rect 49641 46006 49718 46022
rect 49625 45940 49718 46006
rect 49346 45805 49718 45881
rect 49346 45680 49439 45746
rect 49346 45664 49423 45680
tri 49423 45664 49439 45680 nw
rect 49475 45647 49589 45805
rect 49625 45680 49718 45746
tri 49625 45664 49641 45680 ne
rect 49641 45664 49718 45680
rect 49458 45565 49606 45647
rect 49346 45532 49423 45548
tri 49423 45532 49439 45548 sw
rect 49346 45466 49439 45532
rect 49346 45364 49439 45430
rect 49346 45348 49423 45364
tri 49423 45348 49439 45364 nw
rect 49475 45331 49589 45565
tri 49625 45532 49641 45548 se
rect 49641 45532 49718 45548
rect 49625 45466 49718 45532
rect 49625 45364 49718 45430
tri 49625 45348 49641 45364 ne
rect 49641 45348 49718 45364
rect 49458 45249 49606 45331
rect 49346 45216 49423 45232
tri 49423 45216 49439 45232 sw
rect 49346 45150 49439 45216
rect 49475 45091 49589 45249
tri 49625 45216 49641 45232 se
rect 49641 45216 49718 45232
rect 49625 45150 49718 45216
rect 49346 45015 49718 45091
rect 49346 44890 49439 44956
rect 49346 44874 49423 44890
tri 49423 44874 49439 44890 nw
rect 49475 44857 49589 45015
rect 49625 44890 49718 44956
tri 49625 44874 49641 44890 ne
rect 49641 44874 49718 44890
rect 49458 44775 49606 44857
rect 49346 44742 49423 44758
tri 49423 44742 49439 44758 sw
rect 49346 44676 49439 44742
rect 49346 44574 49439 44640
rect 49346 44558 49423 44574
tri 49423 44558 49439 44574 nw
rect 49475 44541 49589 44775
tri 49625 44742 49641 44758 se
rect 49641 44742 49718 44758
rect 49625 44676 49718 44742
rect 49625 44574 49718 44640
tri 49625 44558 49641 44574 ne
rect 49641 44558 49718 44574
rect 49458 44459 49606 44541
rect 49346 44426 49423 44442
tri 49423 44426 49439 44442 sw
rect 49346 44360 49439 44426
rect 49475 44301 49589 44459
tri 49625 44426 49641 44442 se
rect 49641 44426 49718 44442
rect 49625 44360 49718 44426
rect 49346 44225 49718 44301
rect 49346 44100 49439 44166
rect 49346 44084 49423 44100
tri 49423 44084 49439 44100 nw
rect 49475 44067 49589 44225
rect 49625 44100 49718 44166
tri 49625 44084 49641 44100 ne
rect 49641 44084 49718 44100
rect 49458 43985 49606 44067
rect 49346 43952 49423 43968
tri 49423 43952 49439 43968 sw
rect 49346 43886 49439 43952
rect 49346 43784 49439 43850
rect 49346 43768 49423 43784
tri 49423 43768 49439 43784 nw
rect 49475 43751 49589 43985
tri 49625 43952 49641 43968 se
rect 49641 43952 49718 43968
rect 49625 43886 49718 43952
rect 49625 43784 49718 43850
tri 49625 43768 49641 43784 ne
rect 49641 43768 49718 43784
rect 49458 43669 49606 43751
rect 49346 43636 49423 43652
tri 49423 43636 49439 43652 sw
rect 49346 43570 49439 43636
rect 49475 43511 49589 43669
tri 49625 43636 49641 43652 se
rect 49641 43636 49718 43652
rect 49625 43570 49718 43636
rect 49346 43435 49718 43511
rect 49346 43310 49439 43376
rect 49346 43294 49423 43310
tri 49423 43294 49439 43310 nw
rect 49475 43277 49589 43435
rect 49625 43310 49718 43376
tri 49625 43294 49641 43310 ne
rect 49641 43294 49718 43310
rect 49458 43195 49606 43277
rect 49346 43162 49423 43178
tri 49423 43162 49439 43178 sw
rect 49346 43096 49439 43162
rect 49346 42994 49439 43060
rect 49346 42978 49423 42994
tri 49423 42978 49439 42994 nw
rect 49475 42961 49589 43195
tri 49625 43162 49641 43178 se
rect 49641 43162 49718 43178
rect 49625 43096 49718 43162
rect 49625 42994 49718 43060
tri 49625 42978 49641 42994 ne
rect 49641 42978 49718 42994
rect 49458 42879 49606 42961
rect 49346 42846 49423 42862
tri 49423 42846 49439 42862 sw
rect 49346 42780 49439 42846
rect 49475 42721 49589 42879
tri 49625 42846 49641 42862 se
rect 49641 42846 49718 42862
rect 49625 42780 49718 42846
rect 49346 42645 49718 42721
rect 49346 42520 49439 42586
rect 49346 42504 49423 42520
tri 49423 42504 49439 42520 nw
rect 49475 42487 49589 42645
rect 49625 42520 49718 42586
tri 49625 42504 49641 42520 ne
rect 49641 42504 49718 42520
rect 49458 42405 49606 42487
rect 49346 42372 49423 42388
tri 49423 42372 49439 42388 sw
rect 49346 42306 49439 42372
rect 49346 42204 49439 42270
rect 49346 42188 49423 42204
tri 49423 42188 49439 42204 nw
rect 49475 42171 49589 42405
tri 49625 42372 49641 42388 se
rect 49641 42372 49718 42388
rect 49625 42306 49718 42372
rect 49625 42204 49718 42270
tri 49625 42188 49641 42204 ne
rect 49641 42188 49718 42204
rect 49458 42089 49606 42171
rect 49346 42056 49423 42072
tri 49423 42056 49439 42072 sw
rect 49346 41990 49439 42056
rect 49475 41931 49589 42089
tri 49625 42056 49641 42072 se
rect 49641 42056 49718 42072
rect 49625 41990 49718 42056
rect 49346 41855 49718 41931
rect 49346 41730 49439 41796
rect 49346 41714 49423 41730
tri 49423 41714 49439 41730 nw
rect 49475 41697 49589 41855
rect 49625 41730 49718 41796
tri 49625 41714 49641 41730 ne
rect 49641 41714 49718 41730
rect 49458 41615 49606 41697
rect 49346 41582 49423 41598
tri 49423 41582 49439 41598 sw
rect 49346 41516 49439 41582
rect 49346 41414 49439 41480
rect 49346 41398 49423 41414
tri 49423 41398 49439 41414 nw
rect 49475 41381 49589 41615
tri 49625 41582 49641 41598 se
rect 49641 41582 49718 41598
rect 49625 41516 49718 41582
rect 49625 41414 49718 41480
tri 49625 41398 49641 41414 ne
rect 49641 41398 49718 41414
rect 49458 41299 49606 41381
rect 49346 41266 49423 41282
tri 49423 41266 49439 41282 sw
rect 49346 41200 49439 41266
rect 49475 41141 49589 41299
tri 49625 41266 49641 41282 se
rect 49641 41266 49718 41282
rect 49625 41200 49718 41266
rect 49346 41065 49718 41141
rect 49346 40940 49439 41006
rect 49346 40924 49423 40940
tri 49423 40924 49439 40940 nw
rect 49475 40907 49589 41065
rect 49625 40940 49718 41006
tri 49625 40924 49641 40940 ne
rect 49641 40924 49718 40940
rect 49458 40825 49606 40907
rect 49346 40792 49423 40808
tri 49423 40792 49439 40808 sw
rect 49346 40726 49439 40792
rect 49346 40624 49439 40690
rect 49346 40608 49423 40624
tri 49423 40608 49439 40624 nw
rect 49475 40591 49589 40825
tri 49625 40792 49641 40808 se
rect 49641 40792 49718 40808
rect 49625 40726 49718 40792
rect 49625 40624 49718 40690
tri 49625 40608 49641 40624 ne
rect 49641 40608 49718 40624
rect 49458 40509 49606 40591
rect 49346 40476 49423 40492
tri 49423 40476 49439 40492 sw
rect 49346 40410 49439 40476
rect 49475 40351 49589 40509
tri 49625 40476 49641 40492 se
rect 49641 40476 49718 40492
rect 49625 40410 49718 40476
rect 49346 40275 49718 40351
rect 49346 40150 49439 40216
rect 49346 40134 49423 40150
tri 49423 40134 49439 40150 nw
rect 49475 40117 49589 40275
rect 49625 40150 49718 40216
tri 49625 40134 49641 40150 ne
rect 49641 40134 49718 40150
rect 49458 40035 49606 40117
rect 49346 40002 49423 40018
tri 49423 40002 49439 40018 sw
rect 49346 39936 49439 40002
rect 49346 39834 49439 39900
rect 49346 39818 49423 39834
tri 49423 39818 49439 39834 nw
rect 49475 39801 49589 40035
tri 49625 40002 49641 40018 se
rect 49641 40002 49718 40018
rect 49625 39936 49718 40002
rect 49625 39834 49718 39900
tri 49625 39818 49641 39834 ne
rect 49641 39818 49718 39834
rect 49458 39719 49606 39801
rect 49346 39686 49423 39702
tri 49423 39686 49439 39702 sw
rect 49346 39620 49439 39686
rect 49475 39561 49589 39719
tri 49625 39686 49641 39702 se
rect 49641 39686 49718 39702
rect 49625 39620 49718 39686
rect 49346 39485 49718 39561
rect 49346 39360 49439 39426
rect 49346 39344 49423 39360
tri 49423 39344 49439 39360 nw
rect 49475 39327 49589 39485
rect 49625 39360 49718 39426
tri 49625 39344 49641 39360 ne
rect 49641 39344 49718 39360
rect 49458 39245 49606 39327
rect 49346 39212 49423 39228
tri 49423 39212 49439 39228 sw
rect 49346 39146 49439 39212
rect 49346 39044 49439 39110
rect 49346 39028 49423 39044
tri 49423 39028 49439 39044 nw
rect 49475 39011 49589 39245
tri 49625 39212 49641 39228 se
rect 49641 39212 49718 39228
rect 49625 39146 49718 39212
rect 49625 39044 49718 39110
tri 49625 39028 49641 39044 ne
rect 49641 39028 49718 39044
rect 49458 38929 49606 39011
rect 49346 38896 49423 38912
tri 49423 38896 49439 38912 sw
rect 49346 38830 49439 38896
rect 49475 38771 49589 38929
tri 49625 38896 49641 38912 se
rect 49641 38896 49718 38912
rect 49625 38830 49718 38896
rect 49346 38695 49718 38771
rect 49346 38570 49439 38636
rect 49346 38554 49423 38570
tri 49423 38554 49439 38570 nw
rect 49475 38537 49589 38695
rect 49625 38570 49718 38636
tri 49625 38554 49641 38570 ne
rect 49641 38554 49718 38570
rect 49458 38455 49606 38537
rect 49346 38422 49423 38438
tri 49423 38422 49439 38438 sw
rect 49346 38356 49439 38422
rect 49346 38254 49439 38320
rect 49346 38238 49423 38254
tri 49423 38238 49439 38254 nw
rect 49475 38221 49589 38455
tri 49625 38422 49641 38438 se
rect 49641 38422 49718 38438
rect 49625 38356 49718 38422
rect 49625 38254 49718 38320
tri 49625 38238 49641 38254 ne
rect 49641 38238 49718 38254
rect 49458 38139 49606 38221
rect 49346 38106 49423 38122
tri 49423 38106 49439 38122 sw
rect 49346 38040 49439 38106
rect 49475 37981 49589 38139
tri 49625 38106 49641 38122 se
rect 49641 38106 49718 38122
rect 49625 38040 49718 38106
rect 49346 37905 49718 37981
rect 49346 37780 49439 37846
rect 49346 37764 49423 37780
tri 49423 37764 49439 37780 nw
rect 49475 37747 49589 37905
rect 49625 37780 49718 37846
tri 49625 37764 49641 37780 ne
rect 49641 37764 49718 37780
rect 49458 37665 49606 37747
rect 49346 37632 49423 37648
tri 49423 37632 49439 37648 sw
rect 49346 37566 49439 37632
rect 49346 37464 49439 37530
rect 49346 37448 49423 37464
tri 49423 37448 49439 37464 nw
rect 49475 37431 49589 37665
tri 49625 37632 49641 37648 se
rect 49641 37632 49718 37648
rect 49625 37566 49718 37632
rect 49625 37464 49718 37530
tri 49625 37448 49641 37464 ne
rect 49641 37448 49718 37464
rect 49458 37349 49606 37431
rect 49346 37316 49423 37332
tri 49423 37316 49439 37332 sw
rect 49346 37250 49439 37316
rect 49475 37191 49589 37349
tri 49625 37316 49641 37332 se
rect 49641 37316 49718 37332
rect 49625 37250 49718 37316
rect 49346 37115 49718 37191
rect 49346 36990 49439 37056
rect 49346 36974 49423 36990
tri 49423 36974 49439 36990 nw
rect 49475 36957 49589 37115
rect 49625 36990 49718 37056
tri 49625 36974 49641 36990 ne
rect 49641 36974 49718 36990
rect 49458 36875 49606 36957
rect 49346 36842 49423 36858
tri 49423 36842 49439 36858 sw
rect 49346 36776 49439 36842
rect 49346 36674 49439 36740
rect 49346 36658 49423 36674
tri 49423 36658 49439 36674 nw
rect 49475 36641 49589 36875
tri 49625 36842 49641 36858 se
rect 49641 36842 49718 36858
rect 49625 36776 49718 36842
rect 49625 36674 49718 36740
tri 49625 36658 49641 36674 ne
rect 49641 36658 49718 36674
rect 49458 36559 49606 36641
rect 49346 36526 49423 36542
tri 49423 36526 49439 36542 sw
rect 49346 36460 49439 36526
rect 49475 36401 49589 36559
tri 49625 36526 49641 36542 se
rect 49641 36526 49718 36542
rect 49625 36460 49718 36526
rect 49346 36325 49718 36401
rect 49346 36200 49439 36266
rect 49346 36184 49423 36200
tri 49423 36184 49439 36200 nw
rect 49475 36167 49589 36325
rect 49625 36200 49718 36266
tri 49625 36184 49641 36200 ne
rect 49641 36184 49718 36200
rect 49458 36085 49606 36167
rect 49346 36052 49423 36068
tri 49423 36052 49439 36068 sw
rect 49346 35986 49439 36052
rect 49346 35884 49439 35950
rect 49346 35868 49423 35884
tri 49423 35868 49439 35884 nw
rect 49475 35851 49589 36085
tri 49625 36052 49641 36068 se
rect 49641 36052 49718 36068
rect 49625 35986 49718 36052
rect 49625 35884 49718 35950
tri 49625 35868 49641 35884 ne
rect 49641 35868 49718 35884
rect 49458 35769 49606 35851
rect 49346 35736 49423 35752
tri 49423 35736 49439 35752 sw
rect 49346 35670 49439 35736
rect 49475 35611 49589 35769
tri 49625 35736 49641 35752 se
rect 49641 35736 49718 35752
rect 49625 35670 49718 35736
rect 49346 35535 49718 35611
rect 49346 35410 49439 35476
rect 49346 35394 49423 35410
tri 49423 35394 49439 35410 nw
rect 49475 35377 49589 35535
rect 49625 35410 49718 35476
tri 49625 35394 49641 35410 ne
rect 49641 35394 49718 35410
rect 49458 35295 49606 35377
rect 49346 35262 49423 35278
tri 49423 35262 49439 35278 sw
rect 49346 35196 49439 35262
rect 49346 35094 49439 35160
rect 49346 35078 49423 35094
tri 49423 35078 49439 35094 nw
rect 49475 35061 49589 35295
tri 49625 35262 49641 35278 se
rect 49641 35262 49718 35278
rect 49625 35196 49718 35262
rect 49625 35094 49718 35160
tri 49625 35078 49641 35094 ne
rect 49641 35078 49718 35094
rect 49458 34979 49606 35061
rect 49346 34946 49423 34962
tri 49423 34946 49439 34962 sw
rect 49346 34880 49439 34946
rect 49475 34821 49589 34979
tri 49625 34946 49641 34962 se
rect 49641 34946 49718 34962
rect 49625 34880 49718 34946
rect 49346 34745 49718 34821
rect 49346 34620 49439 34686
rect 49346 34604 49423 34620
tri 49423 34604 49439 34620 nw
rect 49475 34587 49589 34745
rect 49625 34620 49718 34686
tri 49625 34604 49641 34620 ne
rect 49641 34604 49718 34620
rect 49458 34505 49606 34587
rect 49346 34472 49423 34488
tri 49423 34472 49439 34488 sw
rect 49346 34406 49439 34472
rect 49346 34304 49439 34370
rect 49346 34288 49423 34304
tri 49423 34288 49439 34304 nw
rect 49475 34271 49589 34505
tri 49625 34472 49641 34488 se
rect 49641 34472 49718 34488
rect 49625 34406 49718 34472
rect 49625 34304 49718 34370
tri 49625 34288 49641 34304 ne
rect 49641 34288 49718 34304
rect 49458 34189 49606 34271
rect 49346 34156 49423 34172
tri 49423 34156 49439 34172 sw
rect 49346 34090 49439 34156
rect 49475 34031 49589 34189
tri 49625 34156 49641 34172 se
rect 49641 34156 49718 34172
rect 49625 34090 49718 34156
rect 49346 33955 49718 34031
rect 49346 33830 49439 33896
rect 49346 33814 49423 33830
tri 49423 33814 49439 33830 nw
rect 49475 33797 49589 33955
rect 49625 33830 49718 33896
tri 49625 33814 49641 33830 ne
rect 49641 33814 49718 33830
rect 49458 33715 49606 33797
rect 49346 33682 49423 33698
tri 49423 33682 49439 33698 sw
rect 49346 33616 49439 33682
rect 49346 33514 49439 33580
rect 49346 33498 49423 33514
tri 49423 33498 49439 33514 nw
rect 49475 33481 49589 33715
tri 49625 33682 49641 33698 se
rect 49641 33682 49718 33698
rect 49625 33616 49718 33682
rect 49625 33514 49718 33580
tri 49625 33498 49641 33514 ne
rect 49641 33498 49718 33514
rect 49458 33399 49606 33481
rect 49346 33366 49423 33382
tri 49423 33366 49439 33382 sw
rect 49346 33300 49439 33366
rect 49475 33241 49589 33399
tri 49625 33366 49641 33382 se
rect 49641 33366 49718 33382
rect 49625 33300 49718 33366
rect 49346 33165 49718 33241
rect 49346 33040 49439 33106
rect 49346 33024 49423 33040
tri 49423 33024 49439 33040 nw
rect 49475 33007 49589 33165
rect 49625 33040 49718 33106
tri 49625 33024 49641 33040 ne
rect 49641 33024 49718 33040
rect 49458 32925 49606 33007
rect 49346 32892 49423 32908
tri 49423 32892 49439 32908 sw
rect 49346 32826 49439 32892
rect 49346 32724 49439 32790
rect 49346 32708 49423 32724
tri 49423 32708 49439 32724 nw
rect 49475 32691 49589 32925
tri 49625 32892 49641 32908 se
rect 49641 32892 49718 32908
rect 49625 32826 49718 32892
rect 49625 32724 49718 32790
tri 49625 32708 49641 32724 ne
rect 49641 32708 49718 32724
rect 49458 32609 49606 32691
rect 49346 32576 49423 32592
tri 49423 32576 49439 32592 sw
rect 49346 32510 49439 32576
rect 49475 32451 49589 32609
tri 49625 32576 49641 32592 se
rect 49641 32576 49718 32592
rect 49625 32510 49718 32576
rect 49346 32375 49718 32451
rect 49346 32250 49439 32316
rect 49346 32234 49423 32250
tri 49423 32234 49439 32250 nw
rect 49475 32217 49589 32375
rect 49625 32250 49718 32316
tri 49625 32234 49641 32250 ne
rect 49641 32234 49718 32250
rect 49458 32135 49606 32217
rect 49346 32102 49423 32118
tri 49423 32102 49439 32118 sw
rect 49346 32036 49439 32102
rect 49346 31934 49439 32000
rect 49346 31918 49423 31934
tri 49423 31918 49439 31934 nw
rect 49475 31901 49589 32135
tri 49625 32102 49641 32118 se
rect 49641 32102 49718 32118
rect 49625 32036 49718 32102
rect 49625 31934 49718 32000
tri 49625 31918 49641 31934 ne
rect 49641 31918 49718 31934
rect 49458 31819 49606 31901
rect 49346 31786 49423 31802
tri 49423 31786 49439 31802 sw
rect 49346 31720 49439 31786
rect 49475 31661 49589 31819
tri 49625 31786 49641 31802 se
rect 49641 31786 49718 31802
rect 49625 31720 49718 31786
rect 49346 31585 49718 31661
rect 49346 31460 49439 31526
rect 49346 31444 49423 31460
tri 49423 31444 49439 31460 nw
rect 49475 31427 49589 31585
rect 49625 31460 49718 31526
tri 49625 31444 49641 31460 ne
rect 49641 31444 49718 31460
rect 49458 31345 49606 31427
rect 49346 31312 49423 31328
tri 49423 31312 49439 31328 sw
rect 49346 31246 49439 31312
rect 49346 31144 49439 31210
rect 49346 31128 49423 31144
tri 49423 31128 49439 31144 nw
rect 49475 31111 49589 31345
tri 49625 31312 49641 31328 se
rect 49641 31312 49718 31328
rect 49625 31246 49718 31312
rect 49625 31144 49718 31210
tri 49625 31128 49641 31144 ne
rect 49641 31128 49718 31144
rect 49458 31029 49606 31111
rect 49346 30996 49423 31012
tri 49423 30996 49439 31012 sw
rect 49346 30930 49439 30996
rect 49475 30871 49589 31029
tri 49625 30996 49641 31012 se
rect 49641 30996 49718 31012
rect 49625 30930 49718 30996
rect 49346 30795 49718 30871
rect 49346 30670 49439 30736
rect 49346 30654 49423 30670
tri 49423 30654 49439 30670 nw
rect 49475 30637 49589 30795
rect 49625 30670 49718 30736
tri 49625 30654 49641 30670 ne
rect 49641 30654 49718 30670
rect 49458 30555 49606 30637
rect 49346 30522 49423 30538
tri 49423 30522 49439 30538 sw
rect 49346 30456 49439 30522
rect 49346 30354 49439 30420
rect 49346 30338 49423 30354
tri 49423 30338 49439 30354 nw
rect 49475 30321 49589 30555
tri 49625 30522 49641 30538 se
rect 49641 30522 49718 30538
rect 49625 30456 49718 30522
rect 49625 30354 49718 30420
tri 49625 30338 49641 30354 ne
rect 49641 30338 49718 30354
rect 49458 30239 49606 30321
rect 49346 30206 49423 30222
tri 49423 30206 49439 30222 sw
rect 49346 30140 49439 30206
rect 49475 30081 49589 30239
tri 49625 30206 49641 30222 se
rect 49641 30206 49718 30222
rect 49625 30140 49718 30206
rect 49346 30005 49718 30081
rect 49346 29880 49439 29946
rect 49346 29864 49423 29880
tri 49423 29864 49439 29880 nw
rect 49475 29847 49589 30005
rect 49625 29880 49718 29946
tri 49625 29864 49641 29880 ne
rect 49641 29864 49718 29880
rect 49458 29765 49606 29847
rect 49346 29732 49423 29748
tri 49423 29732 49439 29748 sw
rect 49346 29666 49439 29732
rect 49346 29564 49439 29630
rect 49346 29548 49423 29564
tri 49423 29548 49439 29564 nw
rect 49475 29531 49589 29765
tri 49625 29732 49641 29748 se
rect 49641 29732 49718 29748
rect 49625 29666 49718 29732
rect 49625 29564 49718 29630
tri 49625 29548 49641 29564 ne
rect 49641 29548 49718 29564
rect 49458 29449 49606 29531
rect 49346 29416 49423 29432
tri 49423 29416 49439 29432 sw
rect 49346 29350 49439 29416
rect 49475 29291 49589 29449
tri 49625 29416 49641 29432 se
rect 49641 29416 49718 29432
rect 49625 29350 49718 29416
rect 49346 29215 49718 29291
rect 49346 29090 49439 29156
rect 49346 29074 49423 29090
tri 49423 29074 49439 29090 nw
rect 49475 29057 49589 29215
rect 49625 29090 49718 29156
tri 49625 29074 49641 29090 ne
rect 49641 29074 49718 29090
rect 49458 28975 49606 29057
rect 49346 28942 49423 28958
tri 49423 28942 49439 28958 sw
rect 49346 28876 49439 28942
rect 49475 28833 49589 28975
tri 49625 28942 49641 28958 se
rect 49641 28942 49718 28958
rect 49625 28876 49718 28942
rect 49754 28463 49790 80603
rect 49826 28463 49862 80603
rect 49898 80445 49934 80603
rect 49890 80303 49942 80445
rect 49898 28763 49934 80303
rect 49890 28621 49942 28763
rect 49898 28463 49934 28621
rect 49970 28463 50006 80603
rect 50042 28463 50078 80603
rect 50114 28833 50198 80233
rect 50234 28463 50270 80603
rect 50306 28463 50342 80603
rect 50378 80445 50414 80603
rect 50370 80303 50422 80445
rect 50378 28763 50414 80303
rect 50370 28621 50422 28763
rect 50378 28463 50414 28621
rect 50450 28463 50486 80603
rect 50522 28463 50558 80603
rect 50594 80124 50687 80190
rect 50594 80108 50671 80124
tri 50671 80108 50687 80124 nw
rect 50723 80091 50837 80233
rect 50873 80124 50966 80190
tri 50873 80108 50889 80124 ne
rect 50889 80108 50966 80124
rect 50706 80009 50854 80091
rect 50594 79976 50671 79992
tri 50671 79976 50687 79992 sw
rect 50594 79910 50687 79976
rect 50723 79851 50837 80009
tri 50873 79976 50889 79992 se
rect 50889 79976 50966 79992
rect 50873 79910 50966 79976
rect 50594 79775 50966 79851
rect 50594 79650 50687 79716
rect 50594 79634 50671 79650
tri 50671 79634 50687 79650 nw
rect 50723 79617 50837 79775
rect 50873 79650 50966 79716
tri 50873 79634 50889 79650 ne
rect 50889 79634 50966 79650
rect 50706 79535 50854 79617
rect 50594 79502 50671 79518
tri 50671 79502 50687 79518 sw
rect 50594 79436 50687 79502
rect 50594 79334 50687 79400
rect 50594 79318 50671 79334
tri 50671 79318 50687 79334 nw
rect 50723 79301 50837 79535
tri 50873 79502 50889 79518 se
rect 50889 79502 50966 79518
rect 50873 79436 50966 79502
rect 50873 79334 50966 79400
tri 50873 79318 50889 79334 ne
rect 50889 79318 50966 79334
rect 50706 79219 50854 79301
rect 50594 79186 50671 79202
tri 50671 79186 50687 79202 sw
rect 50594 79120 50687 79186
rect 50723 79061 50837 79219
tri 50873 79186 50889 79202 se
rect 50889 79186 50966 79202
rect 50873 79120 50966 79186
rect 50594 78985 50966 79061
rect 50594 78860 50687 78926
rect 50594 78844 50671 78860
tri 50671 78844 50687 78860 nw
rect 50723 78827 50837 78985
rect 50873 78860 50966 78926
tri 50873 78844 50889 78860 ne
rect 50889 78844 50966 78860
rect 50706 78745 50854 78827
rect 50594 78712 50671 78728
tri 50671 78712 50687 78728 sw
rect 50594 78646 50687 78712
rect 50594 78544 50687 78610
rect 50594 78528 50671 78544
tri 50671 78528 50687 78544 nw
rect 50723 78511 50837 78745
tri 50873 78712 50889 78728 se
rect 50889 78712 50966 78728
rect 50873 78646 50966 78712
rect 50873 78544 50966 78610
tri 50873 78528 50889 78544 ne
rect 50889 78528 50966 78544
rect 50706 78429 50854 78511
rect 50594 78396 50671 78412
tri 50671 78396 50687 78412 sw
rect 50594 78330 50687 78396
rect 50723 78271 50837 78429
tri 50873 78396 50889 78412 se
rect 50889 78396 50966 78412
rect 50873 78330 50966 78396
rect 50594 78195 50966 78271
rect 50594 78070 50687 78136
rect 50594 78054 50671 78070
tri 50671 78054 50687 78070 nw
rect 50723 78037 50837 78195
rect 50873 78070 50966 78136
tri 50873 78054 50889 78070 ne
rect 50889 78054 50966 78070
rect 50706 77955 50854 78037
rect 50594 77922 50671 77938
tri 50671 77922 50687 77938 sw
rect 50594 77856 50687 77922
rect 50594 77754 50687 77820
rect 50594 77738 50671 77754
tri 50671 77738 50687 77754 nw
rect 50723 77721 50837 77955
tri 50873 77922 50889 77938 se
rect 50889 77922 50966 77938
rect 50873 77856 50966 77922
rect 50873 77754 50966 77820
tri 50873 77738 50889 77754 ne
rect 50889 77738 50966 77754
rect 50706 77639 50854 77721
rect 50594 77606 50671 77622
tri 50671 77606 50687 77622 sw
rect 50594 77540 50687 77606
rect 50723 77481 50837 77639
tri 50873 77606 50889 77622 se
rect 50889 77606 50966 77622
rect 50873 77540 50966 77606
rect 50594 77405 50966 77481
rect 50594 77280 50687 77346
rect 50594 77264 50671 77280
tri 50671 77264 50687 77280 nw
rect 50723 77247 50837 77405
rect 50873 77280 50966 77346
tri 50873 77264 50889 77280 ne
rect 50889 77264 50966 77280
rect 50706 77165 50854 77247
rect 50594 77132 50671 77148
tri 50671 77132 50687 77148 sw
rect 50594 77066 50687 77132
rect 50594 76964 50687 77030
rect 50594 76948 50671 76964
tri 50671 76948 50687 76964 nw
rect 50723 76931 50837 77165
tri 50873 77132 50889 77148 se
rect 50889 77132 50966 77148
rect 50873 77066 50966 77132
rect 50873 76964 50966 77030
tri 50873 76948 50889 76964 ne
rect 50889 76948 50966 76964
rect 50706 76849 50854 76931
rect 50594 76816 50671 76832
tri 50671 76816 50687 76832 sw
rect 50594 76750 50687 76816
rect 50723 76691 50837 76849
tri 50873 76816 50889 76832 se
rect 50889 76816 50966 76832
rect 50873 76750 50966 76816
rect 50594 76615 50966 76691
rect 50594 76490 50687 76556
rect 50594 76474 50671 76490
tri 50671 76474 50687 76490 nw
rect 50723 76457 50837 76615
rect 50873 76490 50966 76556
tri 50873 76474 50889 76490 ne
rect 50889 76474 50966 76490
rect 50706 76375 50854 76457
rect 50594 76342 50671 76358
tri 50671 76342 50687 76358 sw
rect 50594 76276 50687 76342
rect 50594 76174 50687 76240
rect 50594 76158 50671 76174
tri 50671 76158 50687 76174 nw
rect 50723 76141 50837 76375
tri 50873 76342 50889 76358 se
rect 50889 76342 50966 76358
rect 50873 76276 50966 76342
rect 50873 76174 50966 76240
tri 50873 76158 50889 76174 ne
rect 50889 76158 50966 76174
rect 50706 76059 50854 76141
rect 50594 76026 50671 76042
tri 50671 76026 50687 76042 sw
rect 50594 75960 50687 76026
rect 50723 75901 50837 76059
tri 50873 76026 50889 76042 se
rect 50889 76026 50966 76042
rect 50873 75960 50966 76026
rect 50594 75825 50966 75901
rect 50594 75700 50687 75766
rect 50594 75684 50671 75700
tri 50671 75684 50687 75700 nw
rect 50723 75667 50837 75825
rect 50873 75700 50966 75766
tri 50873 75684 50889 75700 ne
rect 50889 75684 50966 75700
rect 50706 75585 50854 75667
rect 50594 75552 50671 75568
tri 50671 75552 50687 75568 sw
rect 50594 75486 50687 75552
rect 50594 75384 50687 75450
rect 50594 75368 50671 75384
tri 50671 75368 50687 75384 nw
rect 50723 75351 50837 75585
tri 50873 75552 50889 75568 se
rect 50889 75552 50966 75568
rect 50873 75486 50966 75552
rect 50873 75384 50966 75450
tri 50873 75368 50889 75384 ne
rect 50889 75368 50966 75384
rect 50706 75269 50854 75351
rect 50594 75236 50671 75252
tri 50671 75236 50687 75252 sw
rect 50594 75170 50687 75236
rect 50723 75111 50837 75269
tri 50873 75236 50889 75252 se
rect 50889 75236 50966 75252
rect 50873 75170 50966 75236
rect 50594 75035 50966 75111
rect 50594 74910 50687 74976
rect 50594 74894 50671 74910
tri 50671 74894 50687 74910 nw
rect 50723 74877 50837 75035
rect 50873 74910 50966 74976
tri 50873 74894 50889 74910 ne
rect 50889 74894 50966 74910
rect 50706 74795 50854 74877
rect 50594 74762 50671 74778
tri 50671 74762 50687 74778 sw
rect 50594 74696 50687 74762
rect 50594 74594 50687 74660
rect 50594 74578 50671 74594
tri 50671 74578 50687 74594 nw
rect 50723 74561 50837 74795
tri 50873 74762 50889 74778 se
rect 50889 74762 50966 74778
rect 50873 74696 50966 74762
rect 50873 74594 50966 74660
tri 50873 74578 50889 74594 ne
rect 50889 74578 50966 74594
rect 50706 74479 50854 74561
rect 50594 74446 50671 74462
tri 50671 74446 50687 74462 sw
rect 50594 74380 50687 74446
rect 50723 74321 50837 74479
tri 50873 74446 50889 74462 se
rect 50889 74446 50966 74462
rect 50873 74380 50966 74446
rect 50594 74245 50966 74321
rect 50594 74120 50687 74186
rect 50594 74104 50671 74120
tri 50671 74104 50687 74120 nw
rect 50723 74087 50837 74245
rect 50873 74120 50966 74186
tri 50873 74104 50889 74120 ne
rect 50889 74104 50966 74120
rect 50706 74005 50854 74087
rect 50594 73972 50671 73988
tri 50671 73972 50687 73988 sw
rect 50594 73906 50687 73972
rect 50594 73804 50687 73870
rect 50594 73788 50671 73804
tri 50671 73788 50687 73804 nw
rect 50723 73771 50837 74005
tri 50873 73972 50889 73988 se
rect 50889 73972 50966 73988
rect 50873 73906 50966 73972
rect 50873 73804 50966 73870
tri 50873 73788 50889 73804 ne
rect 50889 73788 50966 73804
rect 50706 73689 50854 73771
rect 50594 73656 50671 73672
tri 50671 73656 50687 73672 sw
rect 50594 73590 50687 73656
rect 50723 73531 50837 73689
tri 50873 73656 50889 73672 se
rect 50889 73656 50966 73672
rect 50873 73590 50966 73656
rect 50594 73455 50966 73531
rect 50594 73330 50687 73396
rect 50594 73314 50671 73330
tri 50671 73314 50687 73330 nw
rect 50723 73297 50837 73455
rect 50873 73330 50966 73396
tri 50873 73314 50889 73330 ne
rect 50889 73314 50966 73330
rect 50706 73215 50854 73297
rect 50594 73182 50671 73198
tri 50671 73182 50687 73198 sw
rect 50594 73116 50687 73182
rect 50594 73014 50687 73080
rect 50594 72998 50671 73014
tri 50671 72998 50687 73014 nw
rect 50723 72981 50837 73215
tri 50873 73182 50889 73198 se
rect 50889 73182 50966 73198
rect 50873 73116 50966 73182
rect 50873 73014 50966 73080
tri 50873 72998 50889 73014 ne
rect 50889 72998 50966 73014
rect 50706 72899 50854 72981
rect 50594 72866 50671 72882
tri 50671 72866 50687 72882 sw
rect 50594 72800 50687 72866
rect 50723 72741 50837 72899
tri 50873 72866 50889 72882 se
rect 50889 72866 50966 72882
rect 50873 72800 50966 72866
rect 50594 72665 50966 72741
rect 50594 72540 50687 72606
rect 50594 72524 50671 72540
tri 50671 72524 50687 72540 nw
rect 50723 72507 50837 72665
rect 50873 72540 50966 72606
tri 50873 72524 50889 72540 ne
rect 50889 72524 50966 72540
rect 50706 72425 50854 72507
rect 50594 72392 50671 72408
tri 50671 72392 50687 72408 sw
rect 50594 72326 50687 72392
rect 50594 72224 50687 72290
rect 50594 72208 50671 72224
tri 50671 72208 50687 72224 nw
rect 50723 72191 50837 72425
tri 50873 72392 50889 72408 se
rect 50889 72392 50966 72408
rect 50873 72326 50966 72392
rect 50873 72224 50966 72290
tri 50873 72208 50889 72224 ne
rect 50889 72208 50966 72224
rect 50706 72109 50854 72191
rect 50594 72076 50671 72092
tri 50671 72076 50687 72092 sw
rect 50594 72010 50687 72076
rect 50723 71951 50837 72109
tri 50873 72076 50889 72092 se
rect 50889 72076 50966 72092
rect 50873 72010 50966 72076
rect 50594 71875 50966 71951
rect 50594 71750 50687 71816
rect 50594 71734 50671 71750
tri 50671 71734 50687 71750 nw
rect 50723 71717 50837 71875
rect 50873 71750 50966 71816
tri 50873 71734 50889 71750 ne
rect 50889 71734 50966 71750
rect 50706 71635 50854 71717
rect 50594 71602 50671 71618
tri 50671 71602 50687 71618 sw
rect 50594 71536 50687 71602
rect 50594 71434 50687 71500
rect 50594 71418 50671 71434
tri 50671 71418 50687 71434 nw
rect 50723 71401 50837 71635
tri 50873 71602 50889 71618 se
rect 50889 71602 50966 71618
rect 50873 71536 50966 71602
rect 50873 71434 50966 71500
tri 50873 71418 50889 71434 ne
rect 50889 71418 50966 71434
rect 50706 71319 50854 71401
rect 50594 71286 50671 71302
tri 50671 71286 50687 71302 sw
rect 50594 71220 50687 71286
rect 50723 71161 50837 71319
tri 50873 71286 50889 71302 se
rect 50889 71286 50966 71302
rect 50873 71220 50966 71286
rect 50594 71085 50966 71161
rect 50594 70960 50687 71026
rect 50594 70944 50671 70960
tri 50671 70944 50687 70960 nw
rect 50723 70927 50837 71085
rect 50873 70960 50966 71026
tri 50873 70944 50889 70960 ne
rect 50889 70944 50966 70960
rect 50706 70845 50854 70927
rect 50594 70812 50671 70828
tri 50671 70812 50687 70828 sw
rect 50594 70746 50687 70812
rect 50594 70644 50687 70710
rect 50594 70628 50671 70644
tri 50671 70628 50687 70644 nw
rect 50723 70611 50837 70845
tri 50873 70812 50889 70828 se
rect 50889 70812 50966 70828
rect 50873 70746 50966 70812
rect 50873 70644 50966 70710
tri 50873 70628 50889 70644 ne
rect 50889 70628 50966 70644
rect 50706 70529 50854 70611
rect 50594 70496 50671 70512
tri 50671 70496 50687 70512 sw
rect 50594 70430 50687 70496
rect 50723 70371 50837 70529
tri 50873 70496 50889 70512 se
rect 50889 70496 50966 70512
rect 50873 70430 50966 70496
rect 50594 70295 50966 70371
rect 50594 70170 50687 70236
rect 50594 70154 50671 70170
tri 50671 70154 50687 70170 nw
rect 50723 70137 50837 70295
rect 50873 70170 50966 70236
tri 50873 70154 50889 70170 ne
rect 50889 70154 50966 70170
rect 50706 70055 50854 70137
rect 50594 70022 50671 70038
tri 50671 70022 50687 70038 sw
rect 50594 69956 50687 70022
rect 50594 69854 50687 69920
rect 50594 69838 50671 69854
tri 50671 69838 50687 69854 nw
rect 50723 69821 50837 70055
tri 50873 70022 50889 70038 se
rect 50889 70022 50966 70038
rect 50873 69956 50966 70022
rect 50873 69854 50966 69920
tri 50873 69838 50889 69854 ne
rect 50889 69838 50966 69854
rect 50706 69739 50854 69821
rect 50594 69706 50671 69722
tri 50671 69706 50687 69722 sw
rect 50594 69640 50687 69706
rect 50723 69581 50837 69739
tri 50873 69706 50889 69722 se
rect 50889 69706 50966 69722
rect 50873 69640 50966 69706
rect 50594 69505 50966 69581
rect 50594 69380 50687 69446
rect 50594 69364 50671 69380
tri 50671 69364 50687 69380 nw
rect 50723 69347 50837 69505
rect 50873 69380 50966 69446
tri 50873 69364 50889 69380 ne
rect 50889 69364 50966 69380
rect 50706 69265 50854 69347
rect 50594 69232 50671 69248
tri 50671 69232 50687 69248 sw
rect 50594 69166 50687 69232
rect 50594 69064 50687 69130
rect 50594 69048 50671 69064
tri 50671 69048 50687 69064 nw
rect 50723 69031 50837 69265
tri 50873 69232 50889 69248 se
rect 50889 69232 50966 69248
rect 50873 69166 50966 69232
rect 50873 69064 50966 69130
tri 50873 69048 50889 69064 ne
rect 50889 69048 50966 69064
rect 50706 68949 50854 69031
rect 50594 68916 50671 68932
tri 50671 68916 50687 68932 sw
rect 50594 68850 50687 68916
rect 50723 68791 50837 68949
tri 50873 68916 50889 68932 se
rect 50889 68916 50966 68932
rect 50873 68850 50966 68916
rect 50594 68715 50966 68791
rect 50594 68590 50687 68656
rect 50594 68574 50671 68590
tri 50671 68574 50687 68590 nw
rect 50723 68557 50837 68715
rect 50873 68590 50966 68656
tri 50873 68574 50889 68590 ne
rect 50889 68574 50966 68590
rect 50706 68475 50854 68557
rect 50594 68442 50671 68458
tri 50671 68442 50687 68458 sw
rect 50594 68376 50687 68442
rect 50594 68274 50687 68340
rect 50594 68258 50671 68274
tri 50671 68258 50687 68274 nw
rect 50723 68241 50837 68475
tri 50873 68442 50889 68458 se
rect 50889 68442 50966 68458
rect 50873 68376 50966 68442
rect 50873 68274 50966 68340
tri 50873 68258 50889 68274 ne
rect 50889 68258 50966 68274
rect 50706 68159 50854 68241
rect 50594 68126 50671 68142
tri 50671 68126 50687 68142 sw
rect 50594 68060 50687 68126
rect 50723 68001 50837 68159
tri 50873 68126 50889 68142 se
rect 50889 68126 50966 68142
rect 50873 68060 50966 68126
rect 50594 67925 50966 68001
rect 50594 67800 50687 67866
rect 50594 67784 50671 67800
tri 50671 67784 50687 67800 nw
rect 50723 67767 50837 67925
rect 50873 67800 50966 67866
tri 50873 67784 50889 67800 ne
rect 50889 67784 50966 67800
rect 50706 67685 50854 67767
rect 50594 67652 50671 67668
tri 50671 67652 50687 67668 sw
rect 50594 67586 50687 67652
rect 50594 67484 50687 67550
rect 50594 67468 50671 67484
tri 50671 67468 50687 67484 nw
rect 50723 67451 50837 67685
tri 50873 67652 50889 67668 se
rect 50889 67652 50966 67668
rect 50873 67586 50966 67652
rect 50873 67484 50966 67550
tri 50873 67468 50889 67484 ne
rect 50889 67468 50966 67484
rect 50706 67369 50854 67451
rect 50594 67336 50671 67352
tri 50671 67336 50687 67352 sw
rect 50594 67270 50687 67336
rect 50723 67211 50837 67369
tri 50873 67336 50889 67352 se
rect 50889 67336 50966 67352
rect 50873 67270 50966 67336
rect 50594 67135 50966 67211
rect 50594 67010 50687 67076
rect 50594 66994 50671 67010
tri 50671 66994 50687 67010 nw
rect 50723 66977 50837 67135
rect 50873 67010 50966 67076
tri 50873 66994 50889 67010 ne
rect 50889 66994 50966 67010
rect 50706 66895 50854 66977
rect 50594 66862 50671 66878
tri 50671 66862 50687 66878 sw
rect 50594 66796 50687 66862
rect 50594 66694 50687 66760
rect 50594 66678 50671 66694
tri 50671 66678 50687 66694 nw
rect 50723 66661 50837 66895
tri 50873 66862 50889 66878 se
rect 50889 66862 50966 66878
rect 50873 66796 50966 66862
rect 50873 66694 50966 66760
tri 50873 66678 50889 66694 ne
rect 50889 66678 50966 66694
rect 50706 66579 50854 66661
rect 50594 66546 50671 66562
tri 50671 66546 50687 66562 sw
rect 50594 66480 50687 66546
rect 50723 66421 50837 66579
tri 50873 66546 50889 66562 se
rect 50889 66546 50966 66562
rect 50873 66480 50966 66546
rect 50594 66345 50966 66421
rect 50594 66220 50687 66286
rect 50594 66204 50671 66220
tri 50671 66204 50687 66220 nw
rect 50723 66187 50837 66345
rect 50873 66220 50966 66286
tri 50873 66204 50889 66220 ne
rect 50889 66204 50966 66220
rect 50706 66105 50854 66187
rect 50594 66072 50671 66088
tri 50671 66072 50687 66088 sw
rect 50594 66006 50687 66072
rect 50594 65904 50687 65970
rect 50594 65888 50671 65904
tri 50671 65888 50687 65904 nw
rect 50723 65871 50837 66105
tri 50873 66072 50889 66088 se
rect 50889 66072 50966 66088
rect 50873 66006 50966 66072
rect 50873 65904 50966 65970
tri 50873 65888 50889 65904 ne
rect 50889 65888 50966 65904
rect 50706 65789 50854 65871
rect 50594 65756 50671 65772
tri 50671 65756 50687 65772 sw
rect 50594 65690 50687 65756
rect 50723 65631 50837 65789
tri 50873 65756 50889 65772 se
rect 50889 65756 50966 65772
rect 50873 65690 50966 65756
rect 50594 65555 50966 65631
rect 50594 65430 50687 65496
rect 50594 65414 50671 65430
tri 50671 65414 50687 65430 nw
rect 50723 65397 50837 65555
rect 50873 65430 50966 65496
tri 50873 65414 50889 65430 ne
rect 50889 65414 50966 65430
rect 50706 65315 50854 65397
rect 50594 65282 50671 65298
tri 50671 65282 50687 65298 sw
rect 50594 65216 50687 65282
rect 50594 65114 50687 65180
rect 50594 65098 50671 65114
tri 50671 65098 50687 65114 nw
rect 50723 65081 50837 65315
tri 50873 65282 50889 65298 se
rect 50889 65282 50966 65298
rect 50873 65216 50966 65282
rect 50873 65114 50966 65180
tri 50873 65098 50889 65114 ne
rect 50889 65098 50966 65114
rect 50706 64999 50854 65081
rect 50594 64966 50671 64982
tri 50671 64966 50687 64982 sw
rect 50594 64900 50687 64966
rect 50723 64841 50837 64999
tri 50873 64966 50889 64982 se
rect 50889 64966 50966 64982
rect 50873 64900 50966 64966
rect 50594 64765 50966 64841
rect 50594 64640 50687 64706
rect 50594 64624 50671 64640
tri 50671 64624 50687 64640 nw
rect 50723 64607 50837 64765
rect 50873 64640 50966 64706
tri 50873 64624 50889 64640 ne
rect 50889 64624 50966 64640
rect 50706 64525 50854 64607
rect 50594 64492 50671 64508
tri 50671 64492 50687 64508 sw
rect 50594 64426 50687 64492
rect 50594 64324 50687 64390
rect 50594 64308 50671 64324
tri 50671 64308 50687 64324 nw
rect 50723 64291 50837 64525
tri 50873 64492 50889 64508 se
rect 50889 64492 50966 64508
rect 50873 64426 50966 64492
rect 50873 64324 50966 64390
tri 50873 64308 50889 64324 ne
rect 50889 64308 50966 64324
rect 50706 64209 50854 64291
rect 50594 64176 50671 64192
tri 50671 64176 50687 64192 sw
rect 50594 64110 50687 64176
rect 50723 64051 50837 64209
tri 50873 64176 50889 64192 se
rect 50889 64176 50966 64192
rect 50873 64110 50966 64176
rect 50594 63975 50966 64051
rect 50594 63850 50687 63916
rect 50594 63834 50671 63850
tri 50671 63834 50687 63850 nw
rect 50723 63817 50837 63975
rect 50873 63850 50966 63916
tri 50873 63834 50889 63850 ne
rect 50889 63834 50966 63850
rect 50706 63735 50854 63817
rect 50594 63702 50671 63718
tri 50671 63702 50687 63718 sw
rect 50594 63636 50687 63702
rect 50594 63534 50687 63600
rect 50594 63518 50671 63534
tri 50671 63518 50687 63534 nw
rect 50723 63501 50837 63735
tri 50873 63702 50889 63718 se
rect 50889 63702 50966 63718
rect 50873 63636 50966 63702
rect 50873 63534 50966 63600
tri 50873 63518 50889 63534 ne
rect 50889 63518 50966 63534
rect 50706 63419 50854 63501
rect 50594 63386 50671 63402
tri 50671 63386 50687 63402 sw
rect 50594 63320 50687 63386
rect 50723 63261 50837 63419
tri 50873 63386 50889 63402 se
rect 50889 63386 50966 63402
rect 50873 63320 50966 63386
rect 50594 63185 50966 63261
rect 50594 63060 50687 63126
rect 50594 63044 50671 63060
tri 50671 63044 50687 63060 nw
rect 50723 63027 50837 63185
rect 50873 63060 50966 63126
tri 50873 63044 50889 63060 ne
rect 50889 63044 50966 63060
rect 50706 62945 50854 63027
rect 50594 62912 50671 62928
tri 50671 62912 50687 62928 sw
rect 50594 62846 50687 62912
rect 50594 62744 50687 62810
rect 50594 62728 50671 62744
tri 50671 62728 50687 62744 nw
rect 50723 62711 50837 62945
tri 50873 62912 50889 62928 se
rect 50889 62912 50966 62928
rect 50873 62846 50966 62912
rect 50873 62744 50966 62810
tri 50873 62728 50889 62744 ne
rect 50889 62728 50966 62744
rect 50706 62629 50854 62711
rect 50594 62596 50671 62612
tri 50671 62596 50687 62612 sw
rect 50594 62530 50687 62596
rect 50723 62471 50837 62629
tri 50873 62596 50889 62612 se
rect 50889 62596 50966 62612
rect 50873 62530 50966 62596
rect 50594 62395 50966 62471
rect 50594 62270 50687 62336
rect 50594 62254 50671 62270
tri 50671 62254 50687 62270 nw
rect 50723 62237 50837 62395
rect 50873 62270 50966 62336
tri 50873 62254 50889 62270 ne
rect 50889 62254 50966 62270
rect 50706 62155 50854 62237
rect 50594 62122 50671 62138
tri 50671 62122 50687 62138 sw
rect 50594 62056 50687 62122
rect 50594 61954 50687 62020
rect 50594 61938 50671 61954
tri 50671 61938 50687 61954 nw
rect 50723 61921 50837 62155
tri 50873 62122 50889 62138 se
rect 50889 62122 50966 62138
rect 50873 62056 50966 62122
rect 50873 61954 50966 62020
tri 50873 61938 50889 61954 ne
rect 50889 61938 50966 61954
rect 50706 61839 50854 61921
rect 50594 61806 50671 61822
tri 50671 61806 50687 61822 sw
rect 50594 61740 50687 61806
rect 50723 61681 50837 61839
tri 50873 61806 50889 61822 se
rect 50889 61806 50966 61822
rect 50873 61740 50966 61806
rect 50594 61605 50966 61681
rect 50594 61480 50687 61546
rect 50594 61464 50671 61480
tri 50671 61464 50687 61480 nw
rect 50723 61447 50837 61605
rect 50873 61480 50966 61546
tri 50873 61464 50889 61480 ne
rect 50889 61464 50966 61480
rect 50706 61365 50854 61447
rect 50594 61332 50671 61348
tri 50671 61332 50687 61348 sw
rect 50594 61266 50687 61332
rect 50594 61164 50687 61230
rect 50594 61148 50671 61164
tri 50671 61148 50687 61164 nw
rect 50723 61131 50837 61365
tri 50873 61332 50889 61348 se
rect 50889 61332 50966 61348
rect 50873 61266 50966 61332
rect 50873 61164 50966 61230
tri 50873 61148 50889 61164 ne
rect 50889 61148 50966 61164
rect 50706 61049 50854 61131
rect 50594 61016 50671 61032
tri 50671 61016 50687 61032 sw
rect 50594 60950 50687 61016
rect 50723 60891 50837 61049
tri 50873 61016 50889 61032 se
rect 50889 61016 50966 61032
rect 50873 60950 50966 61016
rect 50594 60815 50966 60891
rect 50594 60690 50687 60756
rect 50594 60674 50671 60690
tri 50671 60674 50687 60690 nw
rect 50723 60657 50837 60815
rect 50873 60690 50966 60756
tri 50873 60674 50889 60690 ne
rect 50889 60674 50966 60690
rect 50706 60575 50854 60657
rect 50594 60542 50671 60558
tri 50671 60542 50687 60558 sw
rect 50594 60476 50687 60542
rect 50594 60374 50687 60440
rect 50594 60358 50671 60374
tri 50671 60358 50687 60374 nw
rect 50723 60341 50837 60575
tri 50873 60542 50889 60558 se
rect 50889 60542 50966 60558
rect 50873 60476 50966 60542
rect 50873 60374 50966 60440
tri 50873 60358 50889 60374 ne
rect 50889 60358 50966 60374
rect 50706 60259 50854 60341
rect 50594 60226 50671 60242
tri 50671 60226 50687 60242 sw
rect 50594 60160 50687 60226
rect 50723 60101 50837 60259
tri 50873 60226 50889 60242 se
rect 50889 60226 50966 60242
rect 50873 60160 50966 60226
rect 50594 60025 50966 60101
rect 50594 59900 50687 59966
rect 50594 59884 50671 59900
tri 50671 59884 50687 59900 nw
rect 50723 59867 50837 60025
rect 50873 59900 50966 59966
tri 50873 59884 50889 59900 ne
rect 50889 59884 50966 59900
rect 50706 59785 50854 59867
rect 50594 59752 50671 59768
tri 50671 59752 50687 59768 sw
rect 50594 59686 50687 59752
rect 50594 59584 50687 59650
rect 50594 59568 50671 59584
tri 50671 59568 50687 59584 nw
rect 50723 59551 50837 59785
tri 50873 59752 50889 59768 se
rect 50889 59752 50966 59768
rect 50873 59686 50966 59752
rect 50873 59584 50966 59650
tri 50873 59568 50889 59584 ne
rect 50889 59568 50966 59584
rect 50706 59469 50854 59551
rect 50594 59436 50671 59452
tri 50671 59436 50687 59452 sw
rect 50594 59370 50687 59436
rect 50723 59311 50837 59469
tri 50873 59436 50889 59452 se
rect 50889 59436 50966 59452
rect 50873 59370 50966 59436
rect 50594 59235 50966 59311
rect 50594 59110 50687 59176
rect 50594 59094 50671 59110
tri 50671 59094 50687 59110 nw
rect 50723 59077 50837 59235
rect 50873 59110 50966 59176
tri 50873 59094 50889 59110 ne
rect 50889 59094 50966 59110
rect 50706 58995 50854 59077
rect 50594 58962 50671 58978
tri 50671 58962 50687 58978 sw
rect 50594 58896 50687 58962
rect 50594 58794 50687 58860
rect 50594 58778 50671 58794
tri 50671 58778 50687 58794 nw
rect 50723 58761 50837 58995
tri 50873 58962 50889 58978 se
rect 50889 58962 50966 58978
rect 50873 58896 50966 58962
rect 50873 58794 50966 58860
tri 50873 58778 50889 58794 ne
rect 50889 58778 50966 58794
rect 50706 58679 50854 58761
rect 50594 58646 50671 58662
tri 50671 58646 50687 58662 sw
rect 50594 58580 50687 58646
rect 50723 58521 50837 58679
tri 50873 58646 50889 58662 se
rect 50889 58646 50966 58662
rect 50873 58580 50966 58646
rect 50594 58445 50966 58521
rect 50594 58320 50687 58386
rect 50594 58304 50671 58320
tri 50671 58304 50687 58320 nw
rect 50723 58287 50837 58445
rect 50873 58320 50966 58386
tri 50873 58304 50889 58320 ne
rect 50889 58304 50966 58320
rect 50706 58205 50854 58287
rect 50594 58172 50671 58188
tri 50671 58172 50687 58188 sw
rect 50594 58106 50687 58172
rect 50594 58004 50687 58070
rect 50594 57988 50671 58004
tri 50671 57988 50687 58004 nw
rect 50723 57971 50837 58205
tri 50873 58172 50889 58188 se
rect 50889 58172 50966 58188
rect 50873 58106 50966 58172
rect 50873 58004 50966 58070
tri 50873 57988 50889 58004 ne
rect 50889 57988 50966 58004
rect 50706 57889 50854 57971
rect 50594 57856 50671 57872
tri 50671 57856 50687 57872 sw
rect 50594 57790 50687 57856
rect 50723 57731 50837 57889
tri 50873 57856 50889 57872 se
rect 50889 57856 50966 57872
rect 50873 57790 50966 57856
rect 50594 57655 50966 57731
rect 50594 57530 50687 57596
rect 50594 57514 50671 57530
tri 50671 57514 50687 57530 nw
rect 50723 57497 50837 57655
rect 50873 57530 50966 57596
tri 50873 57514 50889 57530 ne
rect 50889 57514 50966 57530
rect 50706 57415 50854 57497
rect 50594 57382 50671 57398
tri 50671 57382 50687 57398 sw
rect 50594 57316 50687 57382
rect 50594 57214 50687 57280
rect 50594 57198 50671 57214
tri 50671 57198 50687 57214 nw
rect 50723 57181 50837 57415
tri 50873 57382 50889 57398 se
rect 50889 57382 50966 57398
rect 50873 57316 50966 57382
rect 50873 57214 50966 57280
tri 50873 57198 50889 57214 ne
rect 50889 57198 50966 57214
rect 50706 57099 50854 57181
rect 50594 57066 50671 57082
tri 50671 57066 50687 57082 sw
rect 50594 57000 50687 57066
rect 50723 56941 50837 57099
tri 50873 57066 50889 57082 se
rect 50889 57066 50966 57082
rect 50873 57000 50966 57066
rect 50594 56865 50966 56941
rect 50594 56740 50687 56806
rect 50594 56724 50671 56740
tri 50671 56724 50687 56740 nw
rect 50723 56707 50837 56865
rect 50873 56740 50966 56806
tri 50873 56724 50889 56740 ne
rect 50889 56724 50966 56740
rect 50706 56625 50854 56707
rect 50594 56592 50671 56608
tri 50671 56592 50687 56608 sw
rect 50594 56526 50687 56592
rect 50594 56424 50687 56490
rect 50594 56408 50671 56424
tri 50671 56408 50687 56424 nw
rect 50723 56391 50837 56625
tri 50873 56592 50889 56608 se
rect 50889 56592 50966 56608
rect 50873 56526 50966 56592
rect 50873 56424 50966 56490
tri 50873 56408 50889 56424 ne
rect 50889 56408 50966 56424
rect 50706 56309 50854 56391
rect 50594 56276 50671 56292
tri 50671 56276 50687 56292 sw
rect 50594 56210 50687 56276
rect 50723 56151 50837 56309
tri 50873 56276 50889 56292 se
rect 50889 56276 50966 56292
rect 50873 56210 50966 56276
rect 50594 56075 50966 56151
rect 50594 55950 50687 56016
rect 50594 55934 50671 55950
tri 50671 55934 50687 55950 nw
rect 50723 55917 50837 56075
rect 50873 55950 50966 56016
tri 50873 55934 50889 55950 ne
rect 50889 55934 50966 55950
rect 50706 55835 50854 55917
rect 50594 55802 50671 55818
tri 50671 55802 50687 55818 sw
rect 50594 55736 50687 55802
rect 50594 55634 50687 55700
rect 50594 55618 50671 55634
tri 50671 55618 50687 55634 nw
rect 50723 55601 50837 55835
tri 50873 55802 50889 55818 se
rect 50889 55802 50966 55818
rect 50873 55736 50966 55802
rect 50873 55634 50966 55700
tri 50873 55618 50889 55634 ne
rect 50889 55618 50966 55634
rect 50706 55519 50854 55601
rect 50594 55486 50671 55502
tri 50671 55486 50687 55502 sw
rect 50594 55420 50687 55486
rect 50723 55361 50837 55519
tri 50873 55486 50889 55502 se
rect 50889 55486 50966 55502
rect 50873 55420 50966 55486
rect 50594 55285 50966 55361
rect 50594 55160 50687 55226
rect 50594 55144 50671 55160
tri 50671 55144 50687 55160 nw
rect 50723 55127 50837 55285
rect 50873 55160 50966 55226
tri 50873 55144 50889 55160 ne
rect 50889 55144 50966 55160
rect 50706 55045 50854 55127
rect 50594 55012 50671 55028
tri 50671 55012 50687 55028 sw
rect 50594 54946 50687 55012
rect 50594 54844 50687 54910
rect 50594 54828 50671 54844
tri 50671 54828 50687 54844 nw
rect 50723 54811 50837 55045
tri 50873 55012 50889 55028 se
rect 50889 55012 50966 55028
rect 50873 54946 50966 55012
rect 50873 54844 50966 54910
tri 50873 54828 50889 54844 ne
rect 50889 54828 50966 54844
rect 50706 54729 50854 54811
rect 50594 54696 50671 54712
tri 50671 54696 50687 54712 sw
rect 50594 54630 50687 54696
rect 50723 54571 50837 54729
tri 50873 54696 50889 54712 se
rect 50889 54696 50966 54712
rect 50873 54630 50966 54696
rect 50594 54495 50966 54571
rect 50594 54370 50687 54436
rect 50594 54354 50671 54370
tri 50671 54354 50687 54370 nw
rect 50723 54337 50837 54495
rect 50873 54370 50966 54436
tri 50873 54354 50889 54370 ne
rect 50889 54354 50966 54370
rect 50706 54255 50854 54337
rect 50594 54222 50671 54238
tri 50671 54222 50687 54238 sw
rect 50594 54156 50687 54222
rect 50594 54054 50687 54120
rect 50594 54038 50671 54054
tri 50671 54038 50687 54054 nw
rect 50723 54021 50837 54255
tri 50873 54222 50889 54238 se
rect 50889 54222 50966 54238
rect 50873 54156 50966 54222
rect 50873 54054 50966 54120
tri 50873 54038 50889 54054 ne
rect 50889 54038 50966 54054
rect 50706 53939 50854 54021
rect 50594 53906 50671 53922
tri 50671 53906 50687 53922 sw
rect 50594 53840 50687 53906
rect 50723 53781 50837 53939
tri 50873 53906 50889 53922 se
rect 50889 53906 50966 53922
rect 50873 53840 50966 53906
rect 50594 53705 50966 53781
rect 50594 53580 50687 53646
rect 50594 53564 50671 53580
tri 50671 53564 50687 53580 nw
rect 50723 53547 50837 53705
rect 50873 53580 50966 53646
tri 50873 53564 50889 53580 ne
rect 50889 53564 50966 53580
rect 50706 53465 50854 53547
rect 50594 53432 50671 53448
tri 50671 53432 50687 53448 sw
rect 50594 53366 50687 53432
rect 50594 53264 50687 53330
rect 50594 53248 50671 53264
tri 50671 53248 50687 53264 nw
rect 50723 53231 50837 53465
tri 50873 53432 50889 53448 se
rect 50889 53432 50966 53448
rect 50873 53366 50966 53432
rect 50873 53264 50966 53330
tri 50873 53248 50889 53264 ne
rect 50889 53248 50966 53264
rect 50706 53149 50854 53231
rect 50594 53116 50671 53132
tri 50671 53116 50687 53132 sw
rect 50594 53050 50687 53116
rect 50723 52991 50837 53149
tri 50873 53116 50889 53132 se
rect 50889 53116 50966 53132
rect 50873 53050 50966 53116
rect 50594 52915 50966 52991
rect 50594 52790 50687 52856
rect 50594 52774 50671 52790
tri 50671 52774 50687 52790 nw
rect 50723 52757 50837 52915
rect 50873 52790 50966 52856
tri 50873 52774 50889 52790 ne
rect 50889 52774 50966 52790
rect 50706 52675 50854 52757
rect 50594 52642 50671 52658
tri 50671 52642 50687 52658 sw
rect 50594 52576 50687 52642
rect 50594 52474 50687 52540
rect 50594 52458 50671 52474
tri 50671 52458 50687 52474 nw
rect 50723 52441 50837 52675
tri 50873 52642 50889 52658 se
rect 50889 52642 50966 52658
rect 50873 52576 50966 52642
rect 50873 52474 50966 52540
tri 50873 52458 50889 52474 ne
rect 50889 52458 50966 52474
rect 50706 52359 50854 52441
rect 50594 52326 50671 52342
tri 50671 52326 50687 52342 sw
rect 50594 52260 50687 52326
rect 50723 52201 50837 52359
tri 50873 52326 50889 52342 se
rect 50889 52326 50966 52342
rect 50873 52260 50966 52326
rect 50594 52125 50966 52201
rect 50594 52000 50687 52066
rect 50594 51984 50671 52000
tri 50671 51984 50687 52000 nw
rect 50723 51967 50837 52125
rect 50873 52000 50966 52066
tri 50873 51984 50889 52000 ne
rect 50889 51984 50966 52000
rect 50706 51885 50854 51967
rect 50594 51852 50671 51868
tri 50671 51852 50687 51868 sw
rect 50594 51786 50687 51852
rect 50594 51684 50687 51750
rect 50594 51668 50671 51684
tri 50671 51668 50687 51684 nw
rect 50723 51651 50837 51885
tri 50873 51852 50889 51868 se
rect 50889 51852 50966 51868
rect 50873 51786 50966 51852
rect 50873 51684 50966 51750
tri 50873 51668 50889 51684 ne
rect 50889 51668 50966 51684
rect 50706 51569 50854 51651
rect 50594 51536 50671 51552
tri 50671 51536 50687 51552 sw
rect 50594 51470 50687 51536
rect 50723 51411 50837 51569
tri 50873 51536 50889 51552 se
rect 50889 51536 50966 51552
rect 50873 51470 50966 51536
rect 50594 51335 50966 51411
rect 50594 51210 50687 51276
rect 50594 51194 50671 51210
tri 50671 51194 50687 51210 nw
rect 50723 51177 50837 51335
rect 50873 51210 50966 51276
tri 50873 51194 50889 51210 ne
rect 50889 51194 50966 51210
rect 50706 51095 50854 51177
rect 50594 51062 50671 51078
tri 50671 51062 50687 51078 sw
rect 50594 50996 50687 51062
rect 50594 50894 50687 50960
rect 50594 50878 50671 50894
tri 50671 50878 50687 50894 nw
rect 50723 50861 50837 51095
tri 50873 51062 50889 51078 se
rect 50889 51062 50966 51078
rect 50873 50996 50966 51062
rect 50873 50894 50966 50960
tri 50873 50878 50889 50894 ne
rect 50889 50878 50966 50894
rect 50706 50779 50854 50861
rect 50594 50746 50671 50762
tri 50671 50746 50687 50762 sw
rect 50594 50680 50687 50746
rect 50723 50621 50837 50779
tri 50873 50746 50889 50762 se
rect 50889 50746 50966 50762
rect 50873 50680 50966 50746
rect 50594 50545 50966 50621
rect 50594 50420 50687 50486
rect 50594 50404 50671 50420
tri 50671 50404 50687 50420 nw
rect 50723 50387 50837 50545
rect 50873 50420 50966 50486
tri 50873 50404 50889 50420 ne
rect 50889 50404 50966 50420
rect 50706 50305 50854 50387
rect 50594 50272 50671 50288
tri 50671 50272 50687 50288 sw
rect 50594 50206 50687 50272
rect 50594 50104 50687 50170
rect 50594 50088 50671 50104
tri 50671 50088 50687 50104 nw
rect 50723 50071 50837 50305
tri 50873 50272 50889 50288 se
rect 50889 50272 50966 50288
rect 50873 50206 50966 50272
rect 50873 50104 50966 50170
tri 50873 50088 50889 50104 ne
rect 50889 50088 50966 50104
rect 50706 49989 50854 50071
rect 50594 49956 50671 49972
tri 50671 49956 50687 49972 sw
rect 50594 49890 50687 49956
rect 50723 49831 50837 49989
tri 50873 49956 50889 49972 se
rect 50889 49956 50966 49972
rect 50873 49890 50966 49956
rect 50594 49755 50966 49831
rect 50594 49630 50687 49696
rect 50594 49614 50671 49630
tri 50671 49614 50687 49630 nw
rect 50723 49597 50837 49755
rect 50873 49630 50966 49696
tri 50873 49614 50889 49630 ne
rect 50889 49614 50966 49630
rect 50706 49515 50854 49597
rect 50594 49482 50671 49498
tri 50671 49482 50687 49498 sw
rect 50594 49416 50687 49482
rect 50594 49314 50687 49380
rect 50594 49298 50671 49314
tri 50671 49298 50687 49314 nw
rect 50723 49281 50837 49515
tri 50873 49482 50889 49498 se
rect 50889 49482 50966 49498
rect 50873 49416 50966 49482
rect 50873 49314 50966 49380
tri 50873 49298 50889 49314 ne
rect 50889 49298 50966 49314
rect 50706 49199 50854 49281
rect 50594 49166 50671 49182
tri 50671 49166 50687 49182 sw
rect 50594 49100 50687 49166
rect 50723 49041 50837 49199
tri 50873 49166 50889 49182 se
rect 50889 49166 50966 49182
rect 50873 49100 50966 49166
rect 50594 48965 50966 49041
rect 50594 48840 50687 48906
rect 50594 48824 50671 48840
tri 50671 48824 50687 48840 nw
rect 50723 48807 50837 48965
rect 50873 48840 50966 48906
tri 50873 48824 50889 48840 ne
rect 50889 48824 50966 48840
rect 50706 48725 50854 48807
rect 50594 48692 50671 48708
tri 50671 48692 50687 48708 sw
rect 50594 48626 50687 48692
rect 50594 48524 50687 48590
rect 50594 48508 50671 48524
tri 50671 48508 50687 48524 nw
rect 50723 48491 50837 48725
tri 50873 48692 50889 48708 se
rect 50889 48692 50966 48708
rect 50873 48626 50966 48692
rect 50873 48524 50966 48590
tri 50873 48508 50889 48524 ne
rect 50889 48508 50966 48524
rect 50706 48409 50854 48491
rect 50594 48376 50671 48392
tri 50671 48376 50687 48392 sw
rect 50594 48310 50687 48376
rect 50723 48251 50837 48409
tri 50873 48376 50889 48392 se
rect 50889 48376 50966 48392
rect 50873 48310 50966 48376
rect 50594 48175 50966 48251
rect 50594 48050 50687 48116
rect 50594 48034 50671 48050
tri 50671 48034 50687 48050 nw
rect 50723 48017 50837 48175
rect 50873 48050 50966 48116
tri 50873 48034 50889 48050 ne
rect 50889 48034 50966 48050
rect 50706 47935 50854 48017
rect 50594 47902 50671 47918
tri 50671 47902 50687 47918 sw
rect 50594 47836 50687 47902
rect 50594 47734 50687 47800
rect 50594 47718 50671 47734
tri 50671 47718 50687 47734 nw
rect 50723 47701 50837 47935
tri 50873 47902 50889 47918 se
rect 50889 47902 50966 47918
rect 50873 47836 50966 47902
rect 50873 47734 50966 47800
tri 50873 47718 50889 47734 ne
rect 50889 47718 50966 47734
rect 50706 47619 50854 47701
rect 50594 47586 50671 47602
tri 50671 47586 50687 47602 sw
rect 50594 47520 50687 47586
rect 50723 47461 50837 47619
tri 50873 47586 50889 47602 se
rect 50889 47586 50966 47602
rect 50873 47520 50966 47586
rect 50594 47385 50966 47461
rect 50594 47260 50687 47326
rect 50594 47244 50671 47260
tri 50671 47244 50687 47260 nw
rect 50723 47227 50837 47385
rect 50873 47260 50966 47326
tri 50873 47244 50889 47260 ne
rect 50889 47244 50966 47260
rect 50706 47145 50854 47227
rect 50594 47112 50671 47128
tri 50671 47112 50687 47128 sw
rect 50594 47046 50687 47112
rect 50594 46944 50687 47010
rect 50594 46928 50671 46944
tri 50671 46928 50687 46944 nw
rect 50723 46911 50837 47145
tri 50873 47112 50889 47128 se
rect 50889 47112 50966 47128
rect 50873 47046 50966 47112
rect 50873 46944 50966 47010
tri 50873 46928 50889 46944 ne
rect 50889 46928 50966 46944
rect 50706 46829 50854 46911
rect 50594 46796 50671 46812
tri 50671 46796 50687 46812 sw
rect 50594 46730 50687 46796
rect 50723 46671 50837 46829
tri 50873 46796 50889 46812 se
rect 50889 46796 50966 46812
rect 50873 46730 50966 46796
rect 50594 46595 50966 46671
rect 50594 46470 50687 46536
rect 50594 46454 50671 46470
tri 50671 46454 50687 46470 nw
rect 50723 46437 50837 46595
rect 50873 46470 50966 46536
tri 50873 46454 50889 46470 ne
rect 50889 46454 50966 46470
rect 50706 46355 50854 46437
rect 50594 46322 50671 46338
tri 50671 46322 50687 46338 sw
rect 50594 46256 50687 46322
rect 50594 46154 50687 46220
rect 50594 46138 50671 46154
tri 50671 46138 50687 46154 nw
rect 50723 46121 50837 46355
tri 50873 46322 50889 46338 se
rect 50889 46322 50966 46338
rect 50873 46256 50966 46322
rect 50873 46154 50966 46220
tri 50873 46138 50889 46154 ne
rect 50889 46138 50966 46154
rect 50706 46039 50854 46121
rect 50594 46006 50671 46022
tri 50671 46006 50687 46022 sw
rect 50594 45940 50687 46006
rect 50723 45881 50837 46039
tri 50873 46006 50889 46022 se
rect 50889 46006 50966 46022
rect 50873 45940 50966 46006
rect 50594 45805 50966 45881
rect 50594 45680 50687 45746
rect 50594 45664 50671 45680
tri 50671 45664 50687 45680 nw
rect 50723 45647 50837 45805
rect 50873 45680 50966 45746
tri 50873 45664 50889 45680 ne
rect 50889 45664 50966 45680
rect 50706 45565 50854 45647
rect 50594 45532 50671 45548
tri 50671 45532 50687 45548 sw
rect 50594 45466 50687 45532
rect 50594 45364 50687 45430
rect 50594 45348 50671 45364
tri 50671 45348 50687 45364 nw
rect 50723 45331 50837 45565
tri 50873 45532 50889 45548 se
rect 50889 45532 50966 45548
rect 50873 45466 50966 45532
rect 50873 45364 50966 45430
tri 50873 45348 50889 45364 ne
rect 50889 45348 50966 45364
rect 50706 45249 50854 45331
rect 50594 45216 50671 45232
tri 50671 45216 50687 45232 sw
rect 50594 45150 50687 45216
rect 50723 45091 50837 45249
tri 50873 45216 50889 45232 se
rect 50889 45216 50966 45232
rect 50873 45150 50966 45216
rect 50594 45015 50966 45091
rect 50594 44890 50687 44956
rect 50594 44874 50671 44890
tri 50671 44874 50687 44890 nw
rect 50723 44857 50837 45015
rect 50873 44890 50966 44956
tri 50873 44874 50889 44890 ne
rect 50889 44874 50966 44890
rect 50706 44775 50854 44857
rect 50594 44742 50671 44758
tri 50671 44742 50687 44758 sw
rect 50594 44676 50687 44742
rect 50594 44574 50687 44640
rect 50594 44558 50671 44574
tri 50671 44558 50687 44574 nw
rect 50723 44541 50837 44775
tri 50873 44742 50889 44758 se
rect 50889 44742 50966 44758
rect 50873 44676 50966 44742
rect 50873 44574 50966 44640
tri 50873 44558 50889 44574 ne
rect 50889 44558 50966 44574
rect 50706 44459 50854 44541
rect 50594 44426 50671 44442
tri 50671 44426 50687 44442 sw
rect 50594 44360 50687 44426
rect 50723 44301 50837 44459
tri 50873 44426 50889 44442 se
rect 50889 44426 50966 44442
rect 50873 44360 50966 44426
rect 50594 44225 50966 44301
rect 50594 44100 50687 44166
rect 50594 44084 50671 44100
tri 50671 44084 50687 44100 nw
rect 50723 44067 50837 44225
rect 50873 44100 50966 44166
tri 50873 44084 50889 44100 ne
rect 50889 44084 50966 44100
rect 50706 43985 50854 44067
rect 50594 43952 50671 43968
tri 50671 43952 50687 43968 sw
rect 50594 43886 50687 43952
rect 50594 43784 50687 43850
rect 50594 43768 50671 43784
tri 50671 43768 50687 43784 nw
rect 50723 43751 50837 43985
tri 50873 43952 50889 43968 se
rect 50889 43952 50966 43968
rect 50873 43886 50966 43952
rect 50873 43784 50966 43850
tri 50873 43768 50889 43784 ne
rect 50889 43768 50966 43784
rect 50706 43669 50854 43751
rect 50594 43636 50671 43652
tri 50671 43636 50687 43652 sw
rect 50594 43570 50687 43636
rect 50723 43511 50837 43669
tri 50873 43636 50889 43652 se
rect 50889 43636 50966 43652
rect 50873 43570 50966 43636
rect 50594 43435 50966 43511
rect 50594 43310 50687 43376
rect 50594 43294 50671 43310
tri 50671 43294 50687 43310 nw
rect 50723 43277 50837 43435
rect 50873 43310 50966 43376
tri 50873 43294 50889 43310 ne
rect 50889 43294 50966 43310
rect 50706 43195 50854 43277
rect 50594 43162 50671 43178
tri 50671 43162 50687 43178 sw
rect 50594 43096 50687 43162
rect 50594 42994 50687 43060
rect 50594 42978 50671 42994
tri 50671 42978 50687 42994 nw
rect 50723 42961 50837 43195
tri 50873 43162 50889 43178 se
rect 50889 43162 50966 43178
rect 50873 43096 50966 43162
rect 50873 42994 50966 43060
tri 50873 42978 50889 42994 ne
rect 50889 42978 50966 42994
rect 50706 42879 50854 42961
rect 50594 42846 50671 42862
tri 50671 42846 50687 42862 sw
rect 50594 42780 50687 42846
rect 50723 42721 50837 42879
tri 50873 42846 50889 42862 se
rect 50889 42846 50966 42862
rect 50873 42780 50966 42846
rect 50594 42645 50966 42721
rect 50594 42520 50687 42586
rect 50594 42504 50671 42520
tri 50671 42504 50687 42520 nw
rect 50723 42487 50837 42645
rect 50873 42520 50966 42586
tri 50873 42504 50889 42520 ne
rect 50889 42504 50966 42520
rect 50706 42405 50854 42487
rect 50594 42372 50671 42388
tri 50671 42372 50687 42388 sw
rect 50594 42306 50687 42372
rect 50594 42204 50687 42270
rect 50594 42188 50671 42204
tri 50671 42188 50687 42204 nw
rect 50723 42171 50837 42405
tri 50873 42372 50889 42388 se
rect 50889 42372 50966 42388
rect 50873 42306 50966 42372
rect 50873 42204 50966 42270
tri 50873 42188 50889 42204 ne
rect 50889 42188 50966 42204
rect 50706 42089 50854 42171
rect 50594 42056 50671 42072
tri 50671 42056 50687 42072 sw
rect 50594 41990 50687 42056
rect 50723 41931 50837 42089
tri 50873 42056 50889 42072 se
rect 50889 42056 50966 42072
rect 50873 41990 50966 42056
rect 50594 41855 50966 41931
rect 50594 41730 50687 41796
rect 50594 41714 50671 41730
tri 50671 41714 50687 41730 nw
rect 50723 41697 50837 41855
rect 50873 41730 50966 41796
tri 50873 41714 50889 41730 ne
rect 50889 41714 50966 41730
rect 50706 41615 50854 41697
rect 50594 41582 50671 41598
tri 50671 41582 50687 41598 sw
rect 50594 41516 50687 41582
rect 50594 41414 50687 41480
rect 50594 41398 50671 41414
tri 50671 41398 50687 41414 nw
rect 50723 41381 50837 41615
tri 50873 41582 50889 41598 se
rect 50889 41582 50966 41598
rect 50873 41516 50966 41582
rect 50873 41414 50966 41480
tri 50873 41398 50889 41414 ne
rect 50889 41398 50966 41414
rect 50706 41299 50854 41381
rect 50594 41266 50671 41282
tri 50671 41266 50687 41282 sw
rect 50594 41200 50687 41266
rect 50723 41141 50837 41299
tri 50873 41266 50889 41282 se
rect 50889 41266 50966 41282
rect 50873 41200 50966 41266
rect 50594 41065 50966 41141
rect 50594 40940 50687 41006
rect 50594 40924 50671 40940
tri 50671 40924 50687 40940 nw
rect 50723 40907 50837 41065
rect 50873 40940 50966 41006
tri 50873 40924 50889 40940 ne
rect 50889 40924 50966 40940
rect 50706 40825 50854 40907
rect 50594 40792 50671 40808
tri 50671 40792 50687 40808 sw
rect 50594 40726 50687 40792
rect 50594 40624 50687 40690
rect 50594 40608 50671 40624
tri 50671 40608 50687 40624 nw
rect 50723 40591 50837 40825
tri 50873 40792 50889 40808 se
rect 50889 40792 50966 40808
rect 50873 40726 50966 40792
rect 50873 40624 50966 40690
tri 50873 40608 50889 40624 ne
rect 50889 40608 50966 40624
rect 50706 40509 50854 40591
rect 50594 40476 50671 40492
tri 50671 40476 50687 40492 sw
rect 50594 40410 50687 40476
rect 50723 40351 50837 40509
tri 50873 40476 50889 40492 se
rect 50889 40476 50966 40492
rect 50873 40410 50966 40476
rect 50594 40275 50966 40351
rect 50594 40150 50687 40216
rect 50594 40134 50671 40150
tri 50671 40134 50687 40150 nw
rect 50723 40117 50837 40275
rect 50873 40150 50966 40216
tri 50873 40134 50889 40150 ne
rect 50889 40134 50966 40150
rect 50706 40035 50854 40117
rect 50594 40002 50671 40018
tri 50671 40002 50687 40018 sw
rect 50594 39936 50687 40002
rect 50594 39834 50687 39900
rect 50594 39818 50671 39834
tri 50671 39818 50687 39834 nw
rect 50723 39801 50837 40035
tri 50873 40002 50889 40018 se
rect 50889 40002 50966 40018
rect 50873 39936 50966 40002
rect 50873 39834 50966 39900
tri 50873 39818 50889 39834 ne
rect 50889 39818 50966 39834
rect 50706 39719 50854 39801
rect 50594 39686 50671 39702
tri 50671 39686 50687 39702 sw
rect 50594 39620 50687 39686
rect 50723 39561 50837 39719
tri 50873 39686 50889 39702 se
rect 50889 39686 50966 39702
rect 50873 39620 50966 39686
rect 50594 39485 50966 39561
rect 50594 39360 50687 39426
rect 50594 39344 50671 39360
tri 50671 39344 50687 39360 nw
rect 50723 39327 50837 39485
rect 50873 39360 50966 39426
tri 50873 39344 50889 39360 ne
rect 50889 39344 50966 39360
rect 50706 39245 50854 39327
rect 50594 39212 50671 39228
tri 50671 39212 50687 39228 sw
rect 50594 39146 50687 39212
rect 50594 39044 50687 39110
rect 50594 39028 50671 39044
tri 50671 39028 50687 39044 nw
rect 50723 39011 50837 39245
tri 50873 39212 50889 39228 se
rect 50889 39212 50966 39228
rect 50873 39146 50966 39212
rect 50873 39044 50966 39110
tri 50873 39028 50889 39044 ne
rect 50889 39028 50966 39044
rect 50706 38929 50854 39011
rect 50594 38896 50671 38912
tri 50671 38896 50687 38912 sw
rect 50594 38830 50687 38896
rect 50723 38771 50837 38929
tri 50873 38896 50889 38912 se
rect 50889 38896 50966 38912
rect 50873 38830 50966 38896
rect 50594 38695 50966 38771
rect 50594 38570 50687 38636
rect 50594 38554 50671 38570
tri 50671 38554 50687 38570 nw
rect 50723 38537 50837 38695
rect 50873 38570 50966 38636
tri 50873 38554 50889 38570 ne
rect 50889 38554 50966 38570
rect 50706 38455 50854 38537
rect 50594 38422 50671 38438
tri 50671 38422 50687 38438 sw
rect 50594 38356 50687 38422
rect 50594 38254 50687 38320
rect 50594 38238 50671 38254
tri 50671 38238 50687 38254 nw
rect 50723 38221 50837 38455
tri 50873 38422 50889 38438 se
rect 50889 38422 50966 38438
rect 50873 38356 50966 38422
rect 50873 38254 50966 38320
tri 50873 38238 50889 38254 ne
rect 50889 38238 50966 38254
rect 50706 38139 50854 38221
rect 50594 38106 50671 38122
tri 50671 38106 50687 38122 sw
rect 50594 38040 50687 38106
rect 50723 37981 50837 38139
tri 50873 38106 50889 38122 se
rect 50889 38106 50966 38122
rect 50873 38040 50966 38106
rect 50594 37905 50966 37981
rect 50594 37780 50687 37846
rect 50594 37764 50671 37780
tri 50671 37764 50687 37780 nw
rect 50723 37747 50837 37905
rect 50873 37780 50966 37846
tri 50873 37764 50889 37780 ne
rect 50889 37764 50966 37780
rect 50706 37665 50854 37747
rect 50594 37632 50671 37648
tri 50671 37632 50687 37648 sw
rect 50594 37566 50687 37632
rect 50594 37464 50687 37530
rect 50594 37448 50671 37464
tri 50671 37448 50687 37464 nw
rect 50723 37431 50837 37665
tri 50873 37632 50889 37648 se
rect 50889 37632 50966 37648
rect 50873 37566 50966 37632
rect 50873 37464 50966 37530
tri 50873 37448 50889 37464 ne
rect 50889 37448 50966 37464
rect 50706 37349 50854 37431
rect 50594 37316 50671 37332
tri 50671 37316 50687 37332 sw
rect 50594 37250 50687 37316
rect 50723 37191 50837 37349
tri 50873 37316 50889 37332 se
rect 50889 37316 50966 37332
rect 50873 37250 50966 37316
rect 50594 37115 50966 37191
rect 50594 36990 50687 37056
rect 50594 36974 50671 36990
tri 50671 36974 50687 36990 nw
rect 50723 36957 50837 37115
rect 50873 36990 50966 37056
tri 50873 36974 50889 36990 ne
rect 50889 36974 50966 36990
rect 50706 36875 50854 36957
rect 50594 36842 50671 36858
tri 50671 36842 50687 36858 sw
rect 50594 36776 50687 36842
rect 50594 36674 50687 36740
rect 50594 36658 50671 36674
tri 50671 36658 50687 36674 nw
rect 50723 36641 50837 36875
tri 50873 36842 50889 36858 se
rect 50889 36842 50966 36858
rect 50873 36776 50966 36842
rect 50873 36674 50966 36740
tri 50873 36658 50889 36674 ne
rect 50889 36658 50966 36674
rect 50706 36559 50854 36641
rect 50594 36526 50671 36542
tri 50671 36526 50687 36542 sw
rect 50594 36460 50687 36526
rect 50723 36401 50837 36559
tri 50873 36526 50889 36542 se
rect 50889 36526 50966 36542
rect 50873 36460 50966 36526
rect 50594 36325 50966 36401
rect 50594 36200 50687 36266
rect 50594 36184 50671 36200
tri 50671 36184 50687 36200 nw
rect 50723 36167 50837 36325
rect 50873 36200 50966 36266
tri 50873 36184 50889 36200 ne
rect 50889 36184 50966 36200
rect 50706 36085 50854 36167
rect 50594 36052 50671 36068
tri 50671 36052 50687 36068 sw
rect 50594 35986 50687 36052
rect 50594 35884 50687 35950
rect 50594 35868 50671 35884
tri 50671 35868 50687 35884 nw
rect 50723 35851 50837 36085
tri 50873 36052 50889 36068 se
rect 50889 36052 50966 36068
rect 50873 35986 50966 36052
rect 50873 35884 50966 35950
tri 50873 35868 50889 35884 ne
rect 50889 35868 50966 35884
rect 50706 35769 50854 35851
rect 50594 35736 50671 35752
tri 50671 35736 50687 35752 sw
rect 50594 35670 50687 35736
rect 50723 35611 50837 35769
tri 50873 35736 50889 35752 se
rect 50889 35736 50966 35752
rect 50873 35670 50966 35736
rect 50594 35535 50966 35611
rect 50594 35410 50687 35476
rect 50594 35394 50671 35410
tri 50671 35394 50687 35410 nw
rect 50723 35377 50837 35535
rect 50873 35410 50966 35476
tri 50873 35394 50889 35410 ne
rect 50889 35394 50966 35410
rect 50706 35295 50854 35377
rect 50594 35262 50671 35278
tri 50671 35262 50687 35278 sw
rect 50594 35196 50687 35262
rect 50594 35094 50687 35160
rect 50594 35078 50671 35094
tri 50671 35078 50687 35094 nw
rect 50723 35061 50837 35295
tri 50873 35262 50889 35278 se
rect 50889 35262 50966 35278
rect 50873 35196 50966 35262
rect 50873 35094 50966 35160
tri 50873 35078 50889 35094 ne
rect 50889 35078 50966 35094
rect 50706 34979 50854 35061
rect 50594 34946 50671 34962
tri 50671 34946 50687 34962 sw
rect 50594 34880 50687 34946
rect 50723 34821 50837 34979
tri 50873 34946 50889 34962 se
rect 50889 34946 50966 34962
rect 50873 34880 50966 34946
rect 50594 34745 50966 34821
rect 50594 34620 50687 34686
rect 50594 34604 50671 34620
tri 50671 34604 50687 34620 nw
rect 50723 34587 50837 34745
rect 50873 34620 50966 34686
tri 50873 34604 50889 34620 ne
rect 50889 34604 50966 34620
rect 50706 34505 50854 34587
rect 50594 34472 50671 34488
tri 50671 34472 50687 34488 sw
rect 50594 34406 50687 34472
rect 50594 34304 50687 34370
rect 50594 34288 50671 34304
tri 50671 34288 50687 34304 nw
rect 50723 34271 50837 34505
tri 50873 34472 50889 34488 se
rect 50889 34472 50966 34488
rect 50873 34406 50966 34472
rect 50873 34304 50966 34370
tri 50873 34288 50889 34304 ne
rect 50889 34288 50966 34304
rect 50706 34189 50854 34271
rect 50594 34156 50671 34172
tri 50671 34156 50687 34172 sw
rect 50594 34090 50687 34156
rect 50723 34031 50837 34189
tri 50873 34156 50889 34172 se
rect 50889 34156 50966 34172
rect 50873 34090 50966 34156
rect 50594 33955 50966 34031
rect 50594 33830 50687 33896
rect 50594 33814 50671 33830
tri 50671 33814 50687 33830 nw
rect 50723 33797 50837 33955
rect 50873 33830 50966 33896
tri 50873 33814 50889 33830 ne
rect 50889 33814 50966 33830
rect 50706 33715 50854 33797
rect 50594 33682 50671 33698
tri 50671 33682 50687 33698 sw
rect 50594 33616 50687 33682
rect 50594 33514 50687 33580
rect 50594 33498 50671 33514
tri 50671 33498 50687 33514 nw
rect 50723 33481 50837 33715
tri 50873 33682 50889 33698 se
rect 50889 33682 50966 33698
rect 50873 33616 50966 33682
rect 50873 33514 50966 33580
tri 50873 33498 50889 33514 ne
rect 50889 33498 50966 33514
rect 50706 33399 50854 33481
rect 50594 33366 50671 33382
tri 50671 33366 50687 33382 sw
rect 50594 33300 50687 33366
rect 50723 33241 50837 33399
tri 50873 33366 50889 33382 se
rect 50889 33366 50966 33382
rect 50873 33300 50966 33366
rect 50594 33165 50966 33241
rect 50594 33040 50687 33106
rect 50594 33024 50671 33040
tri 50671 33024 50687 33040 nw
rect 50723 33007 50837 33165
rect 50873 33040 50966 33106
tri 50873 33024 50889 33040 ne
rect 50889 33024 50966 33040
rect 50706 32925 50854 33007
rect 50594 32892 50671 32908
tri 50671 32892 50687 32908 sw
rect 50594 32826 50687 32892
rect 50594 32724 50687 32790
rect 50594 32708 50671 32724
tri 50671 32708 50687 32724 nw
rect 50723 32691 50837 32925
tri 50873 32892 50889 32908 se
rect 50889 32892 50966 32908
rect 50873 32826 50966 32892
rect 50873 32724 50966 32790
tri 50873 32708 50889 32724 ne
rect 50889 32708 50966 32724
rect 50706 32609 50854 32691
rect 50594 32576 50671 32592
tri 50671 32576 50687 32592 sw
rect 50594 32510 50687 32576
rect 50723 32451 50837 32609
tri 50873 32576 50889 32592 se
rect 50889 32576 50966 32592
rect 50873 32510 50966 32576
rect 50594 32375 50966 32451
rect 50594 32250 50687 32316
rect 50594 32234 50671 32250
tri 50671 32234 50687 32250 nw
rect 50723 32217 50837 32375
rect 50873 32250 50966 32316
tri 50873 32234 50889 32250 ne
rect 50889 32234 50966 32250
rect 50706 32135 50854 32217
rect 50594 32102 50671 32118
tri 50671 32102 50687 32118 sw
rect 50594 32036 50687 32102
rect 50594 31934 50687 32000
rect 50594 31918 50671 31934
tri 50671 31918 50687 31934 nw
rect 50723 31901 50837 32135
tri 50873 32102 50889 32118 se
rect 50889 32102 50966 32118
rect 50873 32036 50966 32102
rect 50873 31934 50966 32000
tri 50873 31918 50889 31934 ne
rect 50889 31918 50966 31934
rect 50706 31819 50854 31901
rect 50594 31786 50671 31802
tri 50671 31786 50687 31802 sw
rect 50594 31720 50687 31786
rect 50723 31661 50837 31819
tri 50873 31786 50889 31802 se
rect 50889 31786 50966 31802
rect 50873 31720 50966 31786
rect 50594 31585 50966 31661
rect 50594 31460 50687 31526
rect 50594 31444 50671 31460
tri 50671 31444 50687 31460 nw
rect 50723 31427 50837 31585
rect 50873 31460 50966 31526
tri 50873 31444 50889 31460 ne
rect 50889 31444 50966 31460
rect 50706 31345 50854 31427
rect 50594 31312 50671 31328
tri 50671 31312 50687 31328 sw
rect 50594 31246 50687 31312
rect 50594 31144 50687 31210
rect 50594 31128 50671 31144
tri 50671 31128 50687 31144 nw
rect 50723 31111 50837 31345
tri 50873 31312 50889 31328 se
rect 50889 31312 50966 31328
rect 50873 31246 50966 31312
rect 50873 31144 50966 31210
tri 50873 31128 50889 31144 ne
rect 50889 31128 50966 31144
rect 50706 31029 50854 31111
rect 50594 30996 50671 31012
tri 50671 30996 50687 31012 sw
rect 50594 30930 50687 30996
rect 50723 30871 50837 31029
tri 50873 30996 50889 31012 se
rect 50889 30996 50966 31012
rect 50873 30930 50966 30996
rect 50594 30795 50966 30871
rect 50594 30670 50687 30736
rect 50594 30654 50671 30670
tri 50671 30654 50687 30670 nw
rect 50723 30637 50837 30795
rect 50873 30670 50966 30736
tri 50873 30654 50889 30670 ne
rect 50889 30654 50966 30670
rect 50706 30555 50854 30637
rect 50594 30522 50671 30538
tri 50671 30522 50687 30538 sw
rect 50594 30456 50687 30522
rect 50594 30354 50687 30420
rect 50594 30338 50671 30354
tri 50671 30338 50687 30354 nw
rect 50723 30321 50837 30555
tri 50873 30522 50889 30538 se
rect 50889 30522 50966 30538
rect 50873 30456 50966 30522
rect 50873 30354 50966 30420
tri 50873 30338 50889 30354 ne
rect 50889 30338 50966 30354
rect 50706 30239 50854 30321
rect 50594 30206 50671 30222
tri 50671 30206 50687 30222 sw
rect 50594 30140 50687 30206
rect 50723 30081 50837 30239
tri 50873 30206 50889 30222 se
rect 50889 30206 50966 30222
rect 50873 30140 50966 30206
rect 50594 30005 50966 30081
rect 50594 29880 50687 29946
rect 50594 29864 50671 29880
tri 50671 29864 50687 29880 nw
rect 50723 29847 50837 30005
rect 50873 29880 50966 29946
tri 50873 29864 50889 29880 ne
rect 50889 29864 50966 29880
rect 50706 29765 50854 29847
rect 50594 29732 50671 29748
tri 50671 29732 50687 29748 sw
rect 50594 29666 50687 29732
rect 50594 29564 50687 29630
rect 50594 29548 50671 29564
tri 50671 29548 50687 29564 nw
rect 50723 29531 50837 29765
tri 50873 29732 50889 29748 se
rect 50889 29732 50966 29748
rect 50873 29666 50966 29732
rect 50873 29564 50966 29630
tri 50873 29548 50889 29564 ne
rect 50889 29548 50966 29564
rect 50706 29449 50854 29531
rect 50594 29416 50671 29432
tri 50671 29416 50687 29432 sw
rect 50594 29350 50687 29416
rect 50723 29291 50837 29449
tri 50873 29416 50889 29432 se
rect 50889 29416 50966 29432
rect 50873 29350 50966 29416
rect 50594 29215 50966 29291
rect 50594 29090 50687 29156
rect 50594 29074 50671 29090
tri 50671 29074 50687 29090 nw
rect 50723 29057 50837 29215
rect 50873 29090 50966 29156
tri 50873 29074 50889 29090 ne
rect 50889 29074 50966 29090
rect 50706 28975 50854 29057
rect 50594 28942 50671 28958
tri 50671 28942 50687 28958 sw
rect 50594 28876 50687 28942
rect 50723 28833 50837 28975
tri 50873 28942 50889 28958 se
rect 50889 28942 50966 28958
rect 50873 28876 50966 28942
rect 51002 28463 51038 80603
rect 51074 28463 51110 80603
rect 51146 80445 51182 80603
rect 51138 80303 51190 80445
rect 51146 28763 51182 80303
rect 51138 28621 51190 28763
rect 51146 28463 51182 28621
rect 51218 28463 51254 80603
rect 51290 28463 51326 80603
rect 51362 28833 51446 80233
rect 51482 28463 51518 80603
rect 51554 28463 51590 80603
rect 51626 80445 51662 80603
rect 51618 80303 51670 80445
rect 51626 28763 51662 80303
rect 51618 28621 51670 28763
rect 51626 28463 51662 28621
rect 51698 28463 51734 80603
rect 51770 28463 51806 80603
rect 51842 80124 51935 80190
rect 51842 80108 51919 80124
tri 51919 80108 51935 80124 nw
rect 51971 80091 52085 80233
rect 52121 80124 52214 80190
tri 52121 80108 52137 80124 ne
rect 52137 80108 52214 80124
rect 51954 80009 52102 80091
rect 51842 79976 51919 79992
tri 51919 79976 51935 79992 sw
rect 51842 79910 51935 79976
rect 51971 79851 52085 80009
tri 52121 79976 52137 79992 se
rect 52137 79976 52214 79992
rect 52121 79910 52214 79976
rect 51842 79775 52214 79851
rect 51842 79650 51935 79716
rect 51842 79634 51919 79650
tri 51919 79634 51935 79650 nw
rect 51971 79617 52085 79775
rect 52121 79650 52214 79716
tri 52121 79634 52137 79650 ne
rect 52137 79634 52214 79650
rect 51954 79535 52102 79617
rect 51842 79502 51919 79518
tri 51919 79502 51935 79518 sw
rect 51842 79436 51935 79502
rect 51842 79334 51935 79400
rect 51842 79318 51919 79334
tri 51919 79318 51935 79334 nw
rect 51971 79301 52085 79535
tri 52121 79502 52137 79518 se
rect 52137 79502 52214 79518
rect 52121 79436 52214 79502
rect 52121 79334 52214 79400
tri 52121 79318 52137 79334 ne
rect 52137 79318 52214 79334
rect 51954 79219 52102 79301
rect 51842 79186 51919 79202
tri 51919 79186 51935 79202 sw
rect 51842 79120 51935 79186
rect 51971 79061 52085 79219
tri 52121 79186 52137 79202 se
rect 52137 79186 52214 79202
rect 52121 79120 52214 79186
rect 51842 78985 52214 79061
rect 51842 78860 51935 78926
rect 51842 78844 51919 78860
tri 51919 78844 51935 78860 nw
rect 51971 78827 52085 78985
rect 52121 78860 52214 78926
tri 52121 78844 52137 78860 ne
rect 52137 78844 52214 78860
rect 51954 78745 52102 78827
rect 51842 78712 51919 78728
tri 51919 78712 51935 78728 sw
rect 51842 78646 51935 78712
rect 51842 78544 51935 78610
rect 51842 78528 51919 78544
tri 51919 78528 51935 78544 nw
rect 51971 78511 52085 78745
tri 52121 78712 52137 78728 se
rect 52137 78712 52214 78728
rect 52121 78646 52214 78712
rect 52121 78544 52214 78610
tri 52121 78528 52137 78544 ne
rect 52137 78528 52214 78544
rect 51954 78429 52102 78511
rect 51842 78396 51919 78412
tri 51919 78396 51935 78412 sw
rect 51842 78330 51935 78396
rect 51971 78271 52085 78429
tri 52121 78396 52137 78412 se
rect 52137 78396 52214 78412
rect 52121 78330 52214 78396
rect 51842 78195 52214 78271
rect 51842 78070 51935 78136
rect 51842 78054 51919 78070
tri 51919 78054 51935 78070 nw
rect 51971 78037 52085 78195
rect 52121 78070 52214 78136
tri 52121 78054 52137 78070 ne
rect 52137 78054 52214 78070
rect 51954 77955 52102 78037
rect 51842 77922 51919 77938
tri 51919 77922 51935 77938 sw
rect 51842 77856 51935 77922
rect 51842 77754 51935 77820
rect 51842 77738 51919 77754
tri 51919 77738 51935 77754 nw
rect 51971 77721 52085 77955
tri 52121 77922 52137 77938 se
rect 52137 77922 52214 77938
rect 52121 77856 52214 77922
rect 52121 77754 52214 77820
tri 52121 77738 52137 77754 ne
rect 52137 77738 52214 77754
rect 51954 77639 52102 77721
rect 51842 77606 51919 77622
tri 51919 77606 51935 77622 sw
rect 51842 77540 51935 77606
rect 51971 77481 52085 77639
tri 52121 77606 52137 77622 se
rect 52137 77606 52214 77622
rect 52121 77540 52214 77606
rect 51842 77405 52214 77481
rect 51842 77280 51935 77346
rect 51842 77264 51919 77280
tri 51919 77264 51935 77280 nw
rect 51971 77247 52085 77405
rect 52121 77280 52214 77346
tri 52121 77264 52137 77280 ne
rect 52137 77264 52214 77280
rect 51954 77165 52102 77247
rect 51842 77132 51919 77148
tri 51919 77132 51935 77148 sw
rect 51842 77066 51935 77132
rect 51842 76964 51935 77030
rect 51842 76948 51919 76964
tri 51919 76948 51935 76964 nw
rect 51971 76931 52085 77165
tri 52121 77132 52137 77148 se
rect 52137 77132 52214 77148
rect 52121 77066 52214 77132
rect 52121 76964 52214 77030
tri 52121 76948 52137 76964 ne
rect 52137 76948 52214 76964
rect 51954 76849 52102 76931
rect 51842 76816 51919 76832
tri 51919 76816 51935 76832 sw
rect 51842 76750 51935 76816
rect 51971 76691 52085 76849
tri 52121 76816 52137 76832 se
rect 52137 76816 52214 76832
rect 52121 76750 52214 76816
rect 51842 76615 52214 76691
rect 51842 76490 51935 76556
rect 51842 76474 51919 76490
tri 51919 76474 51935 76490 nw
rect 51971 76457 52085 76615
rect 52121 76490 52214 76556
tri 52121 76474 52137 76490 ne
rect 52137 76474 52214 76490
rect 51954 76375 52102 76457
rect 51842 76342 51919 76358
tri 51919 76342 51935 76358 sw
rect 51842 76276 51935 76342
rect 51842 76174 51935 76240
rect 51842 76158 51919 76174
tri 51919 76158 51935 76174 nw
rect 51971 76141 52085 76375
tri 52121 76342 52137 76358 se
rect 52137 76342 52214 76358
rect 52121 76276 52214 76342
rect 52121 76174 52214 76240
tri 52121 76158 52137 76174 ne
rect 52137 76158 52214 76174
rect 51954 76059 52102 76141
rect 51842 76026 51919 76042
tri 51919 76026 51935 76042 sw
rect 51842 75960 51935 76026
rect 51971 75901 52085 76059
tri 52121 76026 52137 76042 se
rect 52137 76026 52214 76042
rect 52121 75960 52214 76026
rect 51842 75825 52214 75901
rect 51842 75700 51935 75766
rect 51842 75684 51919 75700
tri 51919 75684 51935 75700 nw
rect 51971 75667 52085 75825
rect 52121 75700 52214 75766
tri 52121 75684 52137 75700 ne
rect 52137 75684 52214 75700
rect 51954 75585 52102 75667
rect 51842 75552 51919 75568
tri 51919 75552 51935 75568 sw
rect 51842 75486 51935 75552
rect 51842 75384 51935 75450
rect 51842 75368 51919 75384
tri 51919 75368 51935 75384 nw
rect 51971 75351 52085 75585
tri 52121 75552 52137 75568 se
rect 52137 75552 52214 75568
rect 52121 75486 52214 75552
rect 52121 75384 52214 75450
tri 52121 75368 52137 75384 ne
rect 52137 75368 52214 75384
rect 51954 75269 52102 75351
rect 51842 75236 51919 75252
tri 51919 75236 51935 75252 sw
rect 51842 75170 51935 75236
rect 51971 75111 52085 75269
tri 52121 75236 52137 75252 se
rect 52137 75236 52214 75252
rect 52121 75170 52214 75236
rect 51842 75035 52214 75111
rect 51842 74910 51935 74976
rect 51842 74894 51919 74910
tri 51919 74894 51935 74910 nw
rect 51971 74877 52085 75035
rect 52121 74910 52214 74976
tri 52121 74894 52137 74910 ne
rect 52137 74894 52214 74910
rect 51954 74795 52102 74877
rect 51842 74762 51919 74778
tri 51919 74762 51935 74778 sw
rect 51842 74696 51935 74762
rect 51842 74594 51935 74660
rect 51842 74578 51919 74594
tri 51919 74578 51935 74594 nw
rect 51971 74561 52085 74795
tri 52121 74762 52137 74778 se
rect 52137 74762 52214 74778
rect 52121 74696 52214 74762
rect 52121 74594 52214 74660
tri 52121 74578 52137 74594 ne
rect 52137 74578 52214 74594
rect 51954 74479 52102 74561
rect 51842 74446 51919 74462
tri 51919 74446 51935 74462 sw
rect 51842 74380 51935 74446
rect 51971 74321 52085 74479
tri 52121 74446 52137 74462 se
rect 52137 74446 52214 74462
rect 52121 74380 52214 74446
rect 51842 74245 52214 74321
rect 51842 74120 51935 74186
rect 51842 74104 51919 74120
tri 51919 74104 51935 74120 nw
rect 51971 74087 52085 74245
rect 52121 74120 52214 74186
tri 52121 74104 52137 74120 ne
rect 52137 74104 52214 74120
rect 51954 74005 52102 74087
rect 51842 73972 51919 73988
tri 51919 73972 51935 73988 sw
rect 51842 73906 51935 73972
rect 51842 73804 51935 73870
rect 51842 73788 51919 73804
tri 51919 73788 51935 73804 nw
rect 51971 73771 52085 74005
tri 52121 73972 52137 73988 se
rect 52137 73972 52214 73988
rect 52121 73906 52214 73972
rect 52121 73804 52214 73870
tri 52121 73788 52137 73804 ne
rect 52137 73788 52214 73804
rect 51954 73689 52102 73771
rect 51842 73656 51919 73672
tri 51919 73656 51935 73672 sw
rect 51842 73590 51935 73656
rect 51971 73531 52085 73689
tri 52121 73656 52137 73672 se
rect 52137 73656 52214 73672
rect 52121 73590 52214 73656
rect 51842 73455 52214 73531
rect 51842 73330 51935 73396
rect 51842 73314 51919 73330
tri 51919 73314 51935 73330 nw
rect 51971 73297 52085 73455
rect 52121 73330 52214 73396
tri 52121 73314 52137 73330 ne
rect 52137 73314 52214 73330
rect 51954 73215 52102 73297
rect 51842 73182 51919 73198
tri 51919 73182 51935 73198 sw
rect 51842 73116 51935 73182
rect 51842 73014 51935 73080
rect 51842 72998 51919 73014
tri 51919 72998 51935 73014 nw
rect 51971 72981 52085 73215
tri 52121 73182 52137 73198 se
rect 52137 73182 52214 73198
rect 52121 73116 52214 73182
rect 52121 73014 52214 73080
tri 52121 72998 52137 73014 ne
rect 52137 72998 52214 73014
rect 51954 72899 52102 72981
rect 51842 72866 51919 72882
tri 51919 72866 51935 72882 sw
rect 51842 72800 51935 72866
rect 51971 72741 52085 72899
tri 52121 72866 52137 72882 se
rect 52137 72866 52214 72882
rect 52121 72800 52214 72866
rect 51842 72665 52214 72741
rect 51842 72540 51935 72606
rect 51842 72524 51919 72540
tri 51919 72524 51935 72540 nw
rect 51971 72507 52085 72665
rect 52121 72540 52214 72606
tri 52121 72524 52137 72540 ne
rect 52137 72524 52214 72540
rect 51954 72425 52102 72507
rect 51842 72392 51919 72408
tri 51919 72392 51935 72408 sw
rect 51842 72326 51935 72392
rect 51842 72224 51935 72290
rect 51842 72208 51919 72224
tri 51919 72208 51935 72224 nw
rect 51971 72191 52085 72425
tri 52121 72392 52137 72408 se
rect 52137 72392 52214 72408
rect 52121 72326 52214 72392
rect 52121 72224 52214 72290
tri 52121 72208 52137 72224 ne
rect 52137 72208 52214 72224
rect 51954 72109 52102 72191
rect 51842 72076 51919 72092
tri 51919 72076 51935 72092 sw
rect 51842 72010 51935 72076
rect 51971 71951 52085 72109
tri 52121 72076 52137 72092 se
rect 52137 72076 52214 72092
rect 52121 72010 52214 72076
rect 51842 71875 52214 71951
rect 51842 71750 51935 71816
rect 51842 71734 51919 71750
tri 51919 71734 51935 71750 nw
rect 51971 71717 52085 71875
rect 52121 71750 52214 71816
tri 52121 71734 52137 71750 ne
rect 52137 71734 52214 71750
rect 51954 71635 52102 71717
rect 51842 71602 51919 71618
tri 51919 71602 51935 71618 sw
rect 51842 71536 51935 71602
rect 51842 71434 51935 71500
rect 51842 71418 51919 71434
tri 51919 71418 51935 71434 nw
rect 51971 71401 52085 71635
tri 52121 71602 52137 71618 se
rect 52137 71602 52214 71618
rect 52121 71536 52214 71602
rect 52121 71434 52214 71500
tri 52121 71418 52137 71434 ne
rect 52137 71418 52214 71434
rect 51954 71319 52102 71401
rect 51842 71286 51919 71302
tri 51919 71286 51935 71302 sw
rect 51842 71220 51935 71286
rect 51971 71161 52085 71319
tri 52121 71286 52137 71302 se
rect 52137 71286 52214 71302
rect 52121 71220 52214 71286
rect 51842 71085 52214 71161
rect 51842 70960 51935 71026
rect 51842 70944 51919 70960
tri 51919 70944 51935 70960 nw
rect 51971 70927 52085 71085
rect 52121 70960 52214 71026
tri 52121 70944 52137 70960 ne
rect 52137 70944 52214 70960
rect 51954 70845 52102 70927
rect 51842 70812 51919 70828
tri 51919 70812 51935 70828 sw
rect 51842 70746 51935 70812
rect 51842 70644 51935 70710
rect 51842 70628 51919 70644
tri 51919 70628 51935 70644 nw
rect 51971 70611 52085 70845
tri 52121 70812 52137 70828 se
rect 52137 70812 52214 70828
rect 52121 70746 52214 70812
rect 52121 70644 52214 70710
tri 52121 70628 52137 70644 ne
rect 52137 70628 52214 70644
rect 51954 70529 52102 70611
rect 51842 70496 51919 70512
tri 51919 70496 51935 70512 sw
rect 51842 70430 51935 70496
rect 51971 70371 52085 70529
tri 52121 70496 52137 70512 se
rect 52137 70496 52214 70512
rect 52121 70430 52214 70496
rect 51842 70295 52214 70371
rect 51842 70170 51935 70236
rect 51842 70154 51919 70170
tri 51919 70154 51935 70170 nw
rect 51971 70137 52085 70295
rect 52121 70170 52214 70236
tri 52121 70154 52137 70170 ne
rect 52137 70154 52214 70170
rect 51954 70055 52102 70137
rect 51842 70022 51919 70038
tri 51919 70022 51935 70038 sw
rect 51842 69956 51935 70022
rect 51842 69854 51935 69920
rect 51842 69838 51919 69854
tri 51919 69838 51935 69854 nw
rect 51971 69821 52085 70055
tri 52121 70022 52137 70038 se
rect 52137 70022 52214 70038
rect 52121 69956 52214 70022
rect 52121 69854 52214 69920
tri 52121 69838 52137 69854 ne
rect 52137 69838 52214 69854
rect 51954 69739 52102 69821
rect 51842 69706 51919 69722
tri 51919 69706 51935 69722 sw
rect 51842 69640 51935 69706
rect 51971 69581 52085 69739
tri 52121 69706 52137 69722 se
rect 52137 69706 52214 69722
rect 52121 69640 52214 69706
rect 51842 69505 52214 69581
rect 51842 69380 51935 69446
rect 51842 69364 51919 69380
tri 51919 69364 51935 69380 nw
rect 51971 69347 52085 69505
rect 52121 69380 52214 69446
tri 52121 69364 52137 69380 ne
rect 52137 69364 52214 69380
rect 51954 69265 52102 69347
rect 51842 69232 51919 69248
tri 51919 69232 51935 69248 sw
rect 51842 69166 51935 69232
rect 51842 69064 51935 69130
rect 51842 69048 51919 69064
tri 51919 69048 51935 69064 nw
rect 51971 69031 52085 69265
tri 52121 69232 52137 69248 se
rect 52137 69232 52214 69248
rect 52121 69166 52214 69232
rect 52121 69064 52214 69130
tri 52121 69048 52137 69064 ne
rect 52137 69048 52214 69064
rect 51954 68949 52102 69031
rect 51842 68916 51919 68932
tri 51919 68916 51935 68932 sw
rect 51842 68850 51935 68916
rect 51971 68791 52085 68949
tri 52121 68916 52137 68932 se
rect 52137 68916 52214 68932
rect 52121 68850 52214 68916
rect 51842 68715 52214 68791
rect 51842 68590 51935 68656
rect 51842 68574 51919 68590
tri 51919 68574 51935 68590 nw
rect 51971 68557 52085 68715
rect 52121 68590 52214 68656
tri 52121 68574 52137 68590 ne
rect 52137 68574 52214 68590
rect 51954 68475 52102 68557
rect 51842 68442 51919 68458
tri 51919 68442 51935 68458 sw
rect 51842 68376 51935 68442
rect 51842 68274 51935 68340
rect 51842 68258 51919 68274
tri 51919 68258 51935 68274 nw
rect 51971 68241 52085 68475
tri 52121 68442 52137 68458 se
rect 52137 68442 52214 68458
rect 52121 68376 52214 68442
rect 52121 68274 52214 68340
tri 52121 68258 52137 68274 ne
rect 52137 68258 52214 68274
rect 51954 68159 52102 68241
rect 51842 68126 51919 68142
tri 51919 68126 51935 68142 sw
rect 51842 68060 51935 68126
rect 51971 68001 52085 68159
tri 52121 68126 52137 68142 se
rect 52137 68126 52214 68142
rect 52121 68060 52214 68126
rect 51842 67925 52214 68001
rect 51842 67800 51935 67866
rect 51842 67784 51919 67800
tri 51919 67784 51935 67800 nw
rect 51971 67767 52085 67925
rect 52121 67800 52214 67866
tri 52121 67784 52137 67800 ne
rect 52137 67784 52214 67800
rect 51954 67685 52102 67767
rect 51842 67652 51919 67668
tri 51919 67652 51935 67668 sw
rect 51842 67586 51935 67652
rect 51842 67484 51935 67550
rect 51842 67468 51919 67484
tri 51919 67468 51935 67484 nw
rect 51971 67451 52085 67685
tri 52121 67652 52137 67668 se
rect 52137 67652 52214 67668
rect 52121 67586 52214 67652
rect 52121 67484 52214 67550
tri 52121 67468 52137 67484 ne
rect 52137 67468 52214 67484
rect 51954 67369 52102 67451
rect 51842 67336 51919 67352
tri 51919 67336 51935 67352 sw
rect 51842 67270 51935 67336
rect 51971 67211 52085 67369
tri 52121 67336 52137 67352 se
rect 52137 67336 52214 67352
rect 52121 67270 52214 67336
rect 51842 67135 52214 67211
rect 51842 67010 51935 67076
rect 51842 66994 51919 67010
tri 51919 66994 51935 67010 nw
rect 51971 66977 52085 67135
rect 52121 67010 52214 67076
tri 52121 66994 52137 67010 ne
rect 52137 66994 52214 67010
rect 51954 66895 52102 66977
rect 51842 66862 51919 66878
tri 51919 66862 51935 66878 sw
rect 51842 66796 51935 66862
rect 51842 66694 51935 66760
rect 51842 66678 51919 66694
tri 51919 66678 51935 66694 nw
rect 51971 66661 52085 66895
tri 52121 66862 52137 66878 se
rect 52137 66862 52214 66878
rect 52121 66796 52214 66862
rect 52121 66694 52214 66760
tri 52121 66678 52137 66694 ne
rect 52137 66678 52214 66694
rect 51954 66579 52102 66661
rect 51842 66546 51919 66562
tri 51919 66546 51935 66562 sw
rect 51842 66480 51935 66546
rect 51971 66421 52085 66579
tri 52121 66546 52137 66562 se
rect 52137 66546 52214 66562
rect 52121 66480 52214 66546
rect 51842 66345 52214 66421
rect 51842 66220 51935 66286
rect 51842 66204 51919 66220
tri 51919 66204 51935 66220 nw
rect 51971 66187 52085 66345
rect 52121 66220 52214 66286
tri 52121 66204 52137 66220 ne
rect 52137 66204 52214 66220
rect 51954 66105 52102 66187
rect 51842 66072 51919 66088
tri 51919 66072 51935 66088 sw
rect 51842 66006 51935 66072
rect 51842 65904 51935 65970
rect 51842 65888 51919 65904
tri 51919 65888 51935 65904 nw
rect 51971 65871 52085 66105
tri 52121 66072 52137 66088 se
rect 52137 66072 52214 66088
rect 52121 66006 52214 66072
rect 52121 65904 52214 65970
tri 52121 65888 52137 65904 ne
rect 52137 65888 52214 65904
rect 51954 65789 52102 65871
rect 51842 65756 51919 65772
tri 51919 65756 51935 65772 sw
rect 51842 65690 51935 65756
rect 51971 65631 52085 65789
tri 52121 65756 52137 65772 se
rect 52137 65756 52214 65772
rect 52121 65690 52214 65756
rect 51842 65555 52214 65631
rect 51842 65430 51935 65496
rect 51842 65414 51919 65430
tri 51919 65414 51935 65430 nw
rect 51971 65397 52085 65555
rect 52121 65430 52214 65496
tri 52121 65414 52137 65430 ne
rect 52137 65414 52214 65430
rect 51954 65315 52102 65397
rect 51842 65282 51919 65298
tri 51919 65282 51935 65298 sw
rect 51842 65216 51935 65282
rect 51842 65114 51935 65180
rect 51842 65098 51919 65114
tri 51919 65098 51935 65114 nw
rect 51971 65081 52085 65315
tri 52121 65282 52137 65298 se
rect 52137 65282 52214 65298
rect 52121 65216 52214 65282
rect 52121 65114 52214 65180
tri 52121 65098 52137 65114 ne
rect 52137 65098 52214 65114
rect 51954 64999 52102 65081
rect 51842 64966 51919 64982
tri 51919 64966 51935 64982 sw
rect 51842 64900 51935 64966
rect 51971 64841 52085 64999
tri 52121 64966 52137 64982 se
rect 52137 64966 52214 64982
rect 52121 64900 52214 64966
rect 51842 64765 52214 64841
rect 51842 64640 51935 64706
rect 51842 64624 51919 64640
tri 51919 64624 51935 64640 nw
rect 51971 64607 52085 64765
rect 52121 64640 52214 64706
tri 52121 64624 52137 64640 ne
rect 52137 64624 52214 64640
rect 51954 64525 52102 64607
rect 51842 64492 51919 64508
tri 51919 64492 51935 64508 sw
rect 51842 64426 51935 64492
rect 51842 64324 51935 64390
rect 51842 64308 51919 64324
tri 51919 64308 51935 64324 nw
rect 51971 64291 52085 64525
tri 52121 64492 52137 64508 se
rect 52137 64492 52214 64508
rect 52121 64426 52214 64492
rect 52121 64324 52214 64390
tri 52121 64308 52137 64324 ne
rect 52137 64308 52214 64324
rect 51954 64209 52102 64291
rect 51842 64176 51919 64192
tri 51919 64176 51935 64192 sw
rect 51842 64110 51935 64176
rect 51971 64051 52085 64209
tri 52121 64176 52137 64192 se
rect 52137 64176 52214 64192
rect 52121 64110 52214 64176
rect 51842 63975 52214 64051
rect 51842 63850 51935 63916
rect 51842 63834 51919 63850
tri 51919 63834 51935 63850 nw
rect 51971 63817 52085 63975
rect 52121 63850 52214 63916
tri 52121 63834 52137 63850 ne
rect 52137 63834 52214 63850
rect 51954 63735 52102 63817
rect 51842 63702 51919 63718
tri 51919 63702 51935 63718 sw
rect 51842 63636 51935 63702
rect 51842 63534 51935 63600
rect 51842 63518 51919 63534
tri 51919 63518 51935 63534 nw
rect 51971 63501 52085 63735
tri 52121 63702 52137 63718 se
rect 52137 63702 52214 63718
rect 52121 63636 52214 63702
rect 52121 63534 52214 63600
tri 52121 63518 52137 63534 ne
rect 52137 63518 52214 63534
rect 51954 63419 52102 63501
rect 51842 63386 51919 63402
tri 51919 63386 51935 63402 sw
rect 51842 63320 51935 63386
rect 51971 63261 52085 63419
tri 52121 63386 52137 63402 se
rect 52137 63386 52214 63402
rect 52121 63320 52214 63386
rect 51842 63185 52214 63261
rect 51842 63060 51935 63126
rect 51842 63044 51919 63060
tri 51919 63044 51935 63060 nw
rect 51971 63027 52085 63185
rect 52121 63060 52214 63126
tri 52121 63044 52137 63060 ne
rect 52137 63044 52214 63060
rect 51954 62945 52102 63027
rect 51842 62912 51919 62928
tri 51919 62912 51935 62928 sw
rect 51842 62846 51935 62912
rect 51842 62744 51935 62810
rect 51842 62728 51919 62744
tri 51919 62728 51935 62744 nw
rect 51971 62711 52085 62945
tri 52121 62912 52137 62928 se
rect 52137 62912 52214 62928
rect 52121 62846 52214 62912
rect 52121 62744 52214 62810
tri 52121 62728 52137 62744 ne
rect 52137 62728 52214 62744
rect 51954 62629 52102 62711
rect 51842 62596 51919 62612
tri 51919 62596 51935 62612 sw
rect 51842 62530 51935 62596
rect 51971 62471 52085 62629
tri 52121 62596 52137 62612 se
rect 52137 62596 52214 62612
rect 52121 62530 52214 62596
rect 51842 62395 52214 62471
rect 51842 62270 51935 62336
rect 51842 62254 51919 62270
tri 51919 62254 51935 62270 nw
rect 51971 62237 52085 62395
rect 52121 62270 52214 62336
tri 52121 62254 52137 62270 ne
rect 52137 62254 52214 62270
rect 51954 62155 52102 62237
rect 51842 62122 51919 62138
tri 51919 62122 51935 62138 sw
rect 51842 62056 51935 62122
rect 51842 61954 51935 62020
rect 51842 61938 51919 61954
tri 51919 61938 51935 61954 nw
rect 51971 61921 52085 62155
tri 52121 62122 52137 62138 se
rect 52137 62122 52214 62138
rect 52121 62056 52214 62122
rect 52121 61954 52214 62020
tri 52121 61938 52137 61954 ne
rect 52137 61938 52214 61954
rect 51954 61839 52102 61921
rect 51842 61806 51919 61822
tri 51919 61806 51935 61822 sw
rect 51842 61740 51935 61806
rect 51971 61681 52085 61839
tri 52121 61806 52137 61822 se
rect 52137 61806 52214 61822
rect 52121 61740 52214 61806
rect 51842 61605 52214 61681
rect 51842 61480 51935 61546
rect 51842 61464 51919 61480
tri 51919 61464 51935 61480 nw
rect 51971 61447 52085 61605
rect 52121 61480 52214 61546
tri 52121 61464 52137 61480 ne
rect 52137 61464 52214 61480
rect 51954 61365 52102 61447
rect 51842 61332 51919 61348
tri 51919 61332 51935 61348 sw
rect 51842 61266 51935 61332
rect 51842 61164 51935 61230
rect 51842 61148 51919 61164
tri 51919 61148 51935 61164 nw
rect 51971 61131 52085 61365
tri 52121 61332 52137 61348 se
rect 52137 61332 52214 61348
rect 52121 61266 52214 61332
rect 52121 61164 52214 61230
tri 52121 61148 52137 61164 ne
rect 52137 61148 52214 61164
rect 51954 61049 52102 61131
rect 51842 61016 51919 61032
tri 51919 61016 51935 61032 sw
rect 51842 60950 51935 61016
rect 51971 60891 52085 61049
tri 52121 61016 52137 61032 se
rect 52137 61016 52214 61032
rect 52121 60950 52214 61016
rect 51842 60815 52214 60891
rect 51842 60690 51935 60756
rect 51842 60674 51919 60690
tri 51919 60674 51935 60690 nw
rect 51971 60657 52085 60815
rect 52121 60690 52214 60756
tri 52121 60674 52137 60690 ne
rect 52137 60674 52214 60690
rect 51954 60575 52102 60657
rect 51842 60542 51919 60558
tri 51919 60542 51935 60558 sw
rect 51842 60476 51935 60542
rect 51842 60374 51935 60440
rect 51842 60358 51919 60374
tri 51919 60358 51935 60374 nw
rect 51971 60341 52085 60575
tri 52121 60542 52137 60558 se
rect 52137 60542 52214 60558
rect 52121 60476 52214 60542
rect 52121 60374 52214 60440
tri 52121 60358 52137 60374 ne
rect 52137 60358 52214 60374
rect 51954 60259 52102 60341
rect 51842 60226 51919 60242
tri 51919 60226 51935 60242 sw
rect 51842 60160 51935 60226
rect 51971 60101 52085 60259
tri 52121 60226 52137 60242 se
rect 52137 60226 52214 60242
rect 52121 60160 52214 60226
rect 51842 60025 52214 60101
rect 51842 59900 51935 59966
rect 51842 59884 51919 59900
tri 51919 59884 51935 59900 nw
rect 51971 59867 52085 60025
rect 52121 59900 52214 59966
tri 52121 59884 52137 59900 ne
rect 52137 59884 52214 59900
rect 51954 59785 52102 59867
rect 51842 59752 51919 59768
tri 51919 59752 51935 59768 sw
rect 51842 59686 51935 59752
rect 51842 59584 51935 59650
rect 51842 59568 51919 59584
tri 51919 59568 51935 59584 nw
rect 51971 59551 52085 59785
tri 52121 59752 52137 59768 se
rect 52137 59752 52214 59768
rect 52121 59686 52214 59752
rect 52121 59584 52214 59650
tri 52121 59568 52137 59584 ne
rect 52137 59568 52214 59584
rect 51954 59469 52102 59551
rect 51842 59436 51919 59452
tri 51919 59436 51935 59452 sw
rect 51842 59370 51935 59436
rect 51971 59311 52085 59469
tri 52121 59436 52137 59452 se
rect 52137 59436 52214 59452
rect 52121 59370 52214 59436
rect 51842 59235 52214 59311
rect 51842 59110 51935 59176
rect 51842 59094 51919 59110
tri 51919 59094 51935 59110 nw
rect 51971 59077 52085 59235
rect 52121 59110 52214 59176
tri 52121 59094 52137 59110 ne
rect 52137 59094 52214 59110
rect 51954 58995 52102 59077
rect 51842 58962 51919 58978
tri 51919 58962 51935 58978 sw
rect 51842 58896 51935 58962
rect 51842 58794 51935 58860
rect 51842 58778 51919 58794
tri 51919 58778 51935 58794 nw
rect 51971 58761 52085 58995
tri 52121 58962 52137 58978 se
rect 52137 58962 52214 58978
rect 52121 58896 52214 58962
rect 52121 58794 52214 58860
tri 52121 58778 52137 58794 ne
rect 52137 58778 52214 58794
rect 51954 58679 52102 58761
rect 51842 58646 51919 58662
tri 51919 58646 51935 58662 sw
rect 51842 58580 51935 58646
rect 51971 58521 52085 58679
tri 52121 58646 52137 58662 se
rect 52137 58646 52214 58662
rect 52121 58580 52214 58646
rect 51842 58445 52214 58521
rect 51842 58320 51935 58386
rect 51842 58304 51919 58320
tri 51919 58304 51935 58320 nw
rect 51971 58287 52085 58445
rect 52121 58320 52214 58386
tri 52121 58304 52137 58320 ne
rect 52137 58304 52214 58320
rect 51954 58205 52102 58287
rect 51842 58172 51919 58188
tri 51919 58172 51935 58188 sw
rect 51842 58106 51935 58172
rect 51842 58004 51935 58070
rect 51842 57988 51919 58004
tri 51919 57988 51935 58004 nw
rect 51971 57971 52085 58205
tri 52121 58172 52137 58188 se
rect 52137 58172 52214 58188
rect 52121 58106 52214 58172
rect 52121 58004 52214 58070
tri 52121 57988 52137 58004 ne
rect 52137 57988 52214 58004
rect 51954 57889 52102 57971
rect 51842 57856 51919 57872
tri 51919 57856 51935 57872 sw
rect 51842 57790 51935 57856
rect 51971 57731 52085 57889
tri 52121 57856 52137 57872 se
rect 52137 57856 52214 57872
rect 52121 57790 52214 57856
rect 51842 57655 52214 57731
rect 51842 57530 51935 57596
rect 51842 57514 51919 57530
tri 51919 57514 51935 57530 nw
rect 51971 57497 52085 57655
rect 52121 57530 52214 57596
tri 52121 57514 52137 57530 ne
rect 52137 57514 52214 57530
rect 51954 57415 52102 57497
rect 51842 57382 51919 57398
tri 51919 57382 51935 57398 sw
rect 51842 57316 51935 57382
rect 51842 57214 51935 57280
rect 51842 57198 51919 57214
tri 51919 57198 51935 57214 nw
rect 51971 57181 52085 57415
tri 52121 57382 52137 57398 se
rect 52137 57382 52214 57398
rect 52121 57316 52214 57382
rect 52121 57214 52214 57280
tri 52121 57198 52137 57214 ne
rect 52137 57198 52214 57214
rect 51954 57099 52102 57181
rect 51842 57066 51919 57082
tri 51919 57066 51935 57082 sw
rect 51842 57000 51935 57066
rect 51971 56941 52085 57099
tri 52121 57066 52137 57082 se
rect 52137 57066 52214 57082
rect 52121 57000 52214 57066
rect 51842 56865 52214 56941
rect 51842 56740 51935 56806
rect 51842 56724 51919 56740
tri 51919 56724 51935 56740 nw
rect 51971 56707 52085 56865
rect 52121 56740 52214 56806
tri 52121 56724 52137 56740 ne
rect 52137 56724 52214 56740
rect 51954 56625 52102 56707
rect 51842 56592 51919 56608
tri 51919 56592 51935 56608 sw
rect 51842 56526 51935 56592
rect 51842 56424 51935 56490
rect 51842 56408 51919 56424
tri 51919 56408 51935 56424 nw
rect 51971 56391 52085 56625
tri 52121 56592 52137 56608 se
rect 52137 56592 52214 56608
rect 52121 56526 52214 56592
rect 52121 56424 52214 56490
tri 52121 56408 52137 56424 ne
rect 52137 56408 52214 56424
rect 51954 56309 52102 56391
rect 51842 56276 51919 56292
tri 51919 56276 51935 56292 sw
rect 51842 56210 51935 56276
rect 51971 56151 52085 56309
tri 52121 56276 52137 56292 se
rect 52137 56276 52214 56292
rect 52121 56210 52214 56276
rect 51842 56075 52214 56151
rect 51842 55950 51935 56016
rect 51842 55934 51919 55950
tri 51919 55934 51935 55950 nw
rect 51971 55917 52085 56075
rect 52121 55950 52214 56016
tri 52121 55934 52137 55950 ne
rect 52137 55934 52214 55950
rect 51954 55835 52102 55917
rect 51842 55802 51919 55818
tri 51919 55802 51935 55818 sw
rect 51842 55736 51935 55802
rect 51842 55634 51935 55700
rect 51842 55618 51919 55634
tri 51919 55618 51935 55634 nw
rect 51971 55601 52085 55835
tri 52121 55802 52137 55818 se
rect 52137 55802 52214 55818
rect 52121 55736 52214 55802
rect 52121 55634 52214 55700
tri 52121 55618 52137 55634 ne
rect 52137 55618 52214 55634
rect 51954 55519 52102 55601
rect 51842 55486 51919 55502
tri 51919 55486 51935 55502 sw
rect 51842 55420 51935 55486
rect 51971 55361 52085 55519
tri 52121 55486 52137 55502 se
rect 52137 55486 52214 55502
rect 52121 55420 52214 55486
rect 51842 55285 52214 55361
rect 51842 55160 51935 55226
rect 51842 55144 51919 55160
tri 51919 55144 51935 55160 nw
rect 51971 55127 52085 55285
rect 52121 55160 52214 55226
tri 52121 55144 52137 55160 ne
rect 52137 55144 52214 55160
rect 51954 55045 52102 55127
rect 51842 55012 51919 55028
tri 51919 55012 51935 55028 sw
rect 51842 54946 51935 55012
rect 51842 54844 51935 54910
rect 51842 54828 51919 54844
tri 51919 54828 51935 54844 nw
rect 51971 54811 52085 55045
tri 52121 55012 52137 55028 se
rect 52137 55012 52214 55028
rect 52121 54946 52214 55012
rect 52121 54844 52214 54910
tri 52121 54828 52137 54844 ne
rect 52137 54828 52214 54844
rect 51954 54729 52102 54811
rect 51842 54696 51919 54712
tri 51919 54696 51935 54712 sw
rect 51842 54630 51935 54696
rect 51971 54571 52085 54729
tri 52121 54696 52137 54712 se
rect 52137 54696 52214 54712
rect 52121 54630 52214 54696
rect 51842 54495 52214 54571
rect 51842 54370 51935 54436
rect 51842 54354 51919 54370
tri 51919 54354 51935 54370 nw
rect 51971 54337 52085 54495
rect 52121 54370 52214 54436
tri 52121 54354 52137 54370 ne
rect 52137 54354 52214 54370
rect 51954 54255 52102 54337
rect 51842 54222 51919 54238
tri 51919 54222 51935 54238 sw
rect 51842 54156 51935 54222
rect 51842 54054 51935 54120
rect 51842 54038 51919 54054
tri 51919 54038 51935 54054 nw
rect 51971 54021 52085 54255
tri 52121 54222 52137 54238 se
rect 52137 54222 52214 54238
rect 52121 54156 52214 54222
rect 52121 54054 52214 54120
tri 52121 54038 52137 54054 ne
rect 52137 54038 52214 54054
rect 51954 53939 52102 54021
rect 51842 53906 51919 53922
tri 51919 53906 51935 53922 sw
rect 51842 53840 51935 53906
rect 51971 53781 52085 53939
tri 52121 53906 52137 53922 se
rect 52137 53906 52214 53922
rect 52121 53840 52214 53906
rect 51842 53705 52214 53781
rect 51842 53580 51935 53646
rect 51842 53564 51919 53580
tri 51919 53564 51935 53580 nw
rect 51971 53547 52085 53705
rect 52121 53580 52214 53646
tri 52121 53564 52137 53580 ne
rect 52137 53564 52214 53580
rect 51954 53465 52102 53547
rect 51842 53432 51919 53448
tri 51919 53432 51935 53448 sw
rect 51842 53366 51935 53432
rect 51842 53264 51935 53330
rect 51842 53248 51919 53264
tri 51919 53248 51935 53264 nw
rect 51971 53231 52085 53465
tri 52121 53432 52137 53448 se
rect 52137 53432 52214 53448
rect 52121 53366 52214 53432
rect 52121 53264 52214 53330
tri 52121 53248 52137 53264 ne
rect 52137 53248 52214 53264
rect 51954 53149 52102 53231
rect 51842 53116 51919 53132
tri 51919 53116 51935 53132 sw
rect 51842 53050 51935 53116
rect 51971 52991 52085 53149
tri 52121 53116 52137 53132 se
rect 52137 53116 52214 53132
rect 52121 53050 52214 53116
rect 51842 52915 52214 52991
rect 51842 52790 51935 52856
rect 51842 52774 51919 52790
tri 51919 52774 51935 52790 nw
rect 51971 52757 52085 52915
rect 52121 52790 52214 52856
tri 52121 52774 52137 52790 ne
rect 52137 52774 52214 52790
rect 51954 52675 52102 52757
rect 51842 52642 51919 52658
tri 51919 52642 51935 52658 sw
rect 51842 52576 51935 52642
rect 51842 52474 51935 52540
rect 51842 52458 51919 52474
tri 51919 52458 51935 52474 nw
rect 51971 52441 52085 52675
tri 52121 52642 52137 52658 se
rect 52137 52642 52214 52658
rect 52121 52576 52214 52642
rect 52121 52474 52214 52540
tri 52121 52458 52137 52474 ne
rect 52137 52458 52214 52474
rect 51954 52359 52102 52441
rect 51842 52326 51919 52342
tri 51919 52326 51935 52342 sw
rect 51842 52260 51935 52326
rect 51971 52201 52085 52359
tri 52121 52326 52137 52342 se
rect 52137 52326 52214 52342
rect 52121 52260 52214 52326
rect 51842 52125 52214 52201
rect 51842 52000 51935 52066
rect 51842 51984 51919 52000
tri 51919 51984 51935 52000 nw
rect 51971 51967 52085 52125
rect 52121 52000 52214 52066
tri 52121 51984 52137 52000 ne
rect 52137 51984 52214 52000
rect 51954 51885 52102 51967
rect 51842 51852 51919 51868
tri 51919 51852 51935 51868 sw
rect 51842 51786 51935 51852
rect 51842 51684 51935 51750
rect 51842 51668 51919 51684
tri 51919 51668 51935 51684 nw
rect 51971 51651 52085 51885
tri 52121 51852 52137 51868 se
rect 52137 51852 52214 51868
rect 52121 51786 52214 51852
rect 52121 51684 52214 51750
tri 52121 51668 52137 51684 ne
rect 52137 51668 52214 51684
rect 51954 51569 52102 51651
rect 51842 51536 51919 51552
tri 51919 51536 51935 51552 sw
rect 51842 51470 51935 51536
rect 51971 51411 52085 51569
tri 52121 51536 52137 51552 se
rect 52137 51536 52214 51552
rect 52121 51470 52214 51536
rect 51842 51335 52214 51411
rect 51842 51210 51935 51276
rect 51842 51194 51919 51210
tri 51919 51194 51935 51210 nw
rect 51971 51177 52085 51335
rect 52121 51210 52214 51276
tri 52121 51194 52137 51210 ne
rect 52137 51194 52214 51210
rect 51954 51095 52102 51177
rect 51842 51062 51919 51078
tri 51919 51062 51935 51078 sw
rect 51842 50996 51935 51062
rect 51842 50894 51935 50960
rect 51842 50878 51919 50894
tri 51919 50878 51935 50894 nw
rect 51971 50861 52085 51095
tri 52121 51062 52137 51078 se
rect 52137 51062 52214 51078
rect 52121 50996 52214 51062
rect 52121 50894 52214 50960
tri 52121 50878 52137 50894 ne
rect 52137 50878 52214 50894
rect 51954 50779 52102 50861
rect 51842 50746 51919 50762
tri 51919 50746 51935 50762 sw
rect 51842 50680 51935 50746
rect 51971 50621 52085 50779
tri 52121 50746 52137 50762 se
rect 52137 50746 52214 50762
rect 52121 50680 52214 50746
rect 51842 50545 52214 50621
rect 51842 50420 51935 50486
rect 51842 50404 51919 50420
tri 51919 50404 51935 50420 nw
rect 51971 50387 52085 50545
rect 52121 50420 52214 50486
tri 52121 50404 52137 50420 ne
rect 52137 50404 52214 50420
rect 51954 50305 52102 50387
rect 51842 50272 51919 50288
tri 51919 50272 51935 50288 sw
rect 51842 50206 51935 50272
rect 51842 50104 51935 50170
rect 51842 50088 51919 50104
tri 51919 50088 51935 50104 nw
rect 51971 50071 52085 50305
tri 52121 50272 52137 50288 se
rect 52137 50272 52214 50288
rect 52121 50206 52214 50272
rect 52121 50104 52214 50170
tri 52121 50088 52137 50104 ne
rect 52137 50088 52214 50104
rect 51954 49989 52102 50071
rect 51842 49956 51919 49972
tri 51919 49956 51935 49972 sw
rect 51842 49890 51935 49956
rect 51971 49831 52085 49989
tri 52121 49956 52137 49972 se
rect 52137 49956 52214 49972
rect 52121 49890 52214 49956
rect 51842 49755 52214 49831
rect 51842 49630 51935 49696
rect 51842 49614 51919 49630
tri 51919 49614 51935 49630 nw
rect 51971 49597 52085 49755
rect 52121 49630 52214 49696
tri 52121 49614 52137 49630 ne
rect 52137 49614 52214 49630
rect 51954 49515 52102 49597
rect 51842 49482 51919 49498
tri 51919 49482 51935 49498 sw
rect 51842 49416 51935 49482
rect 51842 49314 51935 49380
rect 51842 49298 51919 49314
tri 51919 49298 51935 49314 nw
rect 51971 49281 52085 49515
tri 52121 49482 52137 49498 se
rect 52137 49482 52214 49498
rect 52121 49416 52214 49482
rect 52121 49314 52214 49380
tri 52121 49298 52137 49314 ne
rect 52137 49298 52214 49314
rect 51954 49199 52102 49281
rect 51842 49166 51919 49182
tri 51919 49166 51935 49182 sw
rect 51842 49100 51935 49166
rect 51971 49041 52085 49199
tri 52121 49166 52137 49182 se
rect 52137 49166 52214 49182
rect 52121 49100 52214 49166
rect 51842 48965 52214 49041
rect 51842 48840 51935 48906
rect 51842 48824 51919 48840
tri 51919 48824 51935 48840 nw
rect 51971 48807 52085 48965
rect 52121 48840 52214 48906
tri 52121 48824 52137 48840 ne
rect 52137 48824 52214 48840
rect 51954 48725 52102 48807
rect 51842 48692 51919 48708
tri 51919 48692 51935 48708 sw
rect 51842 48626 51935 48692
rect 51842 48524 51935 48590
rect 51842 48508 51919 48524
tri 51919 48508 51935 48524 nw
rect 51971 48491 52085 48725
tri 52121 48692 52137 48708 se
rect 52137 48692 52214 48708
rect 52121 48626 52214 48692
rect 52121 48524 52214 48590
tri 52121 48508 52137 48524 ne
rect 52137 48508 52214 48524
rect 51954 48409 52102 48491
rect 51842 48376 51919 48392
tri 51919 48376 51935 48392 sw
rect 51842 48310 51935 48376
rect 51971 48251 52085 48409
tri 52121 48376 52137 48392 se
rect 52137 48376 52214 48392
rect 52121 48310 52214 48376
rect 51842 48175 52214 48251
rect 51842 48050 51935 48116
rect 51842 48034 51919 48050
tri 51919 48034 51935 48050 nw
rect 51971 48017 52085 48175
rect 52121 48050 52214 48116
tri 52121 48034 52137 48050 ne
rect 52137 48034 52214 48050
rect 51954 47935 52102 48017
rect 51842 47902 51919 47918
tri 51919 47902 51935 47918 sw
rect 51842 47836 51935 47902
rect 51842 47734 51935 47800
rect 51842 47718 51919 47734
tri 51919 47718 51935 47734 nw
rect 51971 47701 52085 47935
tri 52121 47902 52137 47918 se
rect 52137 47902 52214 47918
rect 52121 47836 52214 47902
rect 52121 47734 52214 47800
tri 52121 47718 52137 47734 ne
rect 52137 47718 52214 47734
rect 51954 47619 52102 47701
rect 51842 47586 51919 47602
tri 51919 47586 51935 47602 sw
rect 51842 47520 51935 47586
rect 51971 47461 52085 47619
tri 52121 47586 52137 47602 se
rect 52137 47586 52214 47602
rect 52121 47520 52214 47586
rect 51842 47385 52214 47461
rect 51842 47260 51935 47326
rect 51842 47244 51919 47260
tri 51919 47244 51935 47260 nw
rect 51971 47227 52085 47385
rect 52121 47260 52214 47326
tri 52121 47244 52137 47260 ne
rect 52137 47244 52214 47260
rect 51954 47145 52102 47227
rect 51842 47112 51919 47128
tri 51919 47112 51935 47128 sw
rect 51842 47046 51935 47112
rect 51842 46944 51935 47010
rect 51842 46928 51919 46944
tri 51919 46928 51935 46944 nw
rect 51971 46911 52085 47145
tri 52121 47112 52137 47128 se
rect 52137 47112 52214 47128
rect 52121 47046 52214 47112
rect 52121 46944 52214 47010
tri 52121 46928 52137 46944 ne
rect 52137 46928 52214 46944
rect 51954 46829 52102 46911
rect 51842 46796 51919 46812
tri 51919 46796 51935 46812 sw
rect 51842 46730 51935 46796
rect 51971 46671 52085 46829
tri 52121 46796 52137 46812 se
rect 52137 46796 52214 46812
rect 52121 46730 52214 46796
rect 51842 46595 52214 46671
rect 51842 46470 51935 46536
rect 51842 46454 51919 46470
tri 51919 46454 51935 46470 nw
rect 51971 46437 52085 46595
rect 52121 46470 52214 46536
tri 52121 46454 52137 46470 ne
rect 52137 46454 52214 46470
rect 51954 46355 52102 46437
rect 51842 46322 51919 46338
tri 51919 46322 51935 46338 sw
rect 51842 46256 51935 46322
rect 51842 46154 51935 46220
rect 51842 46138 51919 46154
tri 51919 46138 51935 46154 nw
rect 51971 46121 52085 46355
tri 52121 46322 52137 46338 se
rect 52137 46322 52214 46338
rect 52121 46256 52214 46322
rect 52121 46154 52214 46220
tri 52121 46138 52137 46154 ne
rect 52137 46138 52214 46154
rect 51954 46039 52102 46121
rect 51842 46006 51919 46022
tri 51919 46006 51935 46022 sw
rect 51842 45940 51935 46006
rect 51971 45881 52085 46039
tri 52121 46006 52137 46022 se
rect 52137 46006 52214 46022
rect 52121 45940 52214 46006
rect 51842 45805 52214 45881
rect 51842 45680 51935 45746
rect 51842 45664 51919 45680
tri 51919 45664 51935 45680 nw
rect 51971 45647 52085 45805
rect 52121 45680 52214 45746
tri 52121 45664 52137 45680 ne
rect 52137 45664 52214 45680
rect 51954 45565 52102 45647
rect 51842 45532 51919 45548
tri 51919 45532 51935 45548 sw
rect 51842 45466 51935 45532
rect 51842 45364 51935 45430
rect 51842 45348 51919 45364
tri 51919 45348 51935 45364 nw
rect 51971 45331 52085 45565
tri 52121 45532 52137 45548 se
rect 52137 45532 52214 45548
rect 52121 45466 52214 45532
rect 52121 45364 52214 45430
tri 52121 45348 52137 45364 ne
rect 52137 45348 52214 45364
rect 51954 45249 52102 45331
rect 51842 45216 51919 45232
tri 51919 45216 51935 45232 sw
rect 51842 45150 51935 45216
rect 51971 45091 52085 45249
tri 52121 45216 52137 45232 se
rect 52137 45216 52214 45232
rect 52121 45150 52214 45216
rect 51842 45015 52214 45091
rect 51842 44890 51935 44956
rect 51842 44874 51919 44890
tri 51919 44874 51935 44890 nw
rect 51971 44857 52085 45015
rect 52121 44890 52214 44956
tri 52121 44874 52137 44890 ne
rect 52137 44874 52214 44890
rect 51954 44775 52102 44857
rect 51842 44742 51919 44758
tri 51919 44742 51935 44758 sw
rect 51842 44676 51935 44742
rect 51842 44574 51935 44640
rect 51842 44558 51919 44574
tri 51919 44558 51935 44574 nw
rect 51971 44541 52085 44775
tri 52121 44742 52137 44758 se
rect 52137 44742 52214 44758
rect 52121 44676 52214 44742
rect 52121 44574 52214 44640
tri 52121 44558 52137 44574 ne
rect 52137 44558 52214 44574
rect 51954 44459 52102 44541
rect 51842 44426 51919 44442
tri 51919 44426 51935 44442 sw
rect 51842 44360 51935 44426
rect 51971 44301 52085 44459
tri 52121 44426 52137 44442 se
rect 52137 44426 52214 44442
rect 52121 44360 52214 44426
rect 51842 44225 52214 44301
rect 51842 44100 51935 44166
rect 51842 44084 51919 44100
tri 51919 44084 51935 44100 nw
rect 51971 44067 52085 44225
rect 52121 44100 52214 44166
tri 52121 44084 52137 44100 ne
rect 52137 44084 52214 44100
rect 51954 43985 52102 44067
rect 51842 43952 51919 43968
tri 51919 43952 51935 43968 sw
rect 51842 43886 51935 43952
rect 51842 43784 51935 43850
rect 51842 43768 51919 43784
tri 51919 43768 51935 43784 nw
rect 51971 43751 52085 43985
tri 52121 43952 52137 43968 se
rect 52137 43952 52214 43968
rect 52121 43886 52214 43952
rect 52121 43784 52214 43850
tri 52121 43768 52137 43784 ne
rect 52137 43768 52214 43784
rect 51954 43669 52102 43751
rect 51842 43636 51919 43652
tri 51919 43636 51935 43652 sw
rect 51842 43570 51935 43636
rect 51971 43511 52085 43669
tri 52121 43636 52137 43652 se
rect 52137 43636 52214 43652
rect 52121 43570 52214 43636
rect 51842 43435 52214 43511
rect 51842 43310 51935 43376
rect 51842 43294 51919 43310
tri 51919 43294 51935 43310 nw
rect 51971 43277 52085 43435
rect 52121 43310 52214 43376
tri 52121 43294 52137 43310 ne
rect 52137 43294 52214 43310
rect 51954 43195 52102 43277
rect 51842 43162 51919 43178
tri 51919 43162 51935 43178 sw
rect 51842 43096 51935 43162
rect 51842 42994 51935 43060
rect 51842 42978 51919 42994
tri 51919 42978 51935 42994 nw
rect 51971 42961 52085 43195
tri 52121 43162 52137 43178 se
rect 52137 43162 52214 43178
rect 52121 43096 52214 43162
rect 52121 42994 52214 43060
tri 52121 42978 52137 42994 ne
rect 52137 42978 52214 42994
rect 51954 42879 52102 42961
rect 51842 42846 51919 42862
tri 51919 42846 51935 42862 sw
rect 51842 42780 51935 42846
rect 51971 42721 52085 42879
tri 52121 42846 52137 42862 se
rect 52137 42846 52214 42862
rect 52121 42780 52214 42846
rect 51842 42645 52214 42721
rect 51842 42520 51935 42586
rect 51842 42504 51919 42520
tri 51919 42504 51935 42520 nw
rect 51971 42487 52085 42645
rect 52121 42520 52214 42586
tri 52121 42504 52137 42520 ne
rect 52137 42504 52214 42520
rect 51954 42405 52102 42487
rect 51842 42372 51919 42388
tri 51919 42372 51935 42388 sw
rect 51842 42306 51935 42372
rect 51842 42204 51935 42270
rect 51842 42188 51919 42204
tri 51919 42188 51935 42204 nw
rect 51971 42171 52085 42405
tri 52121 42372 52137 42388 se
rect 52137 42372 52214 42388
rect 52121 42306 52214 42372
rect 52121 42204 52214 42270
tri 52121 42188 52137 42204 ne
rect 52137 42188 52214 42204
rect 51954 42089 52102 42171
rect 51842 42056 51919 42072
tri 51919 42056 51935 42072 sw
rect 51842 41990 51935 42056
rect 51971 41931 52085 42089
tri 52121 42056 52137 42072 se
rect 52137 42056 52214 42072
rect 52121 41990 52214 42056
rect 51842 41855 52214 41931
rect 51842 41730 51935 41796
rect 51842 41714 51919 41730
tri 51919 41714 51935 41730 nw
rect 51971 41697 52085 41855
rect 52121 41730 52214 41796
tri 52121 41714 52137 41730 ne
rect 52137 41714 52214 41730
rect 51954 41615 52102 41697
rect 51842 41582 51919 41598
tri 51919 41582 51935 41598 sw
rect 51842 41516 51935 41582
rect 51842 41414 51935 41480
rect 51842 41398 51919 41414
tri 51919 41398 51935 41414 nw
rect 51971 41381 52085 41615
tri 52121 41582 52137 41598 se
rect 52137 41582 52214 41598
rect 52121 41516 52214 41582
rect 52121 41414 52214 41480
tri 52121 41398 52137 41414 ne
rect 52137 41398 52214 41414
rect 51954 41299 52102 41381
rect 51842 41266 51919 41282
tri 51919 41266 51935 41282 sw
rect 51842 41200 51935 41266
rect 51971 41141 52085 41299
tri 52121 41266 52137 41282 se
rect 52137 41266 52214 41282
rect 52121 41200 52214 41266
rect 51842 41065 52214 41141
rect 51842 40940 51935 41006
rect 51842 40924 51919 40940
tri 51919 40924 51935 40940 nw
rect 51971 40907 52085 41065
rect 52121 40940 52214 41006
tri 52121 40924 52137 40940 ne
rect 52137 40924 52214 40940
rect 51954 40825 52102 40907
rect 51842 40792 51919 40808
tri 51919 40792 51935 40808 sw
rect 51842 40726 51935 40792
rect 51842 40624 51935 40690
rect 51842 40608 51919 40624
tri 51919 40608 51935 40624 nw
rect 51971 40591 52085 40825
tri 52121 40792 52137 40808 se
rect 52137 40792 52214 40808
rect 52121 40726 52214 40792
rect 52121 40624 52214 40690
tri 52121 40608 52137 40624 ne
rect 52137 40608 52214 40624
rect 51954 40509 52102 40591
rect 51842 40476 51919 40492
tri 51919 40476 51935 40492 sw
rect 51842 40410 51935 40476
rect 51971 40351 52085 40509
tri 52121 40476 52137 40492 se
rect 52137 40476 52214 40492
rect 52121 40410 52214 40476
rect 51842 40275 52214 40351
rect 51842 40150 51935 40216
rect 51842 40134 51919 40150
tri 51919 40134 51935 40150 nw
rect 51971 40117 52085 40275
rect 52121 40150 52214 40216
tri 52121 40134 52137 40150 ne
rect 52137 40134 52214 40150
rect 51954 40035 52102 40117
rect 51842 40002 51919 40018
tri 51919 40002 51935 40018 sw
rect 51842 39936 51935 40002
rect 51842 39834 51935 39900
rect 51842 39818 51919 39834
tri 51919 39818 51935 39834 nw
rect 51971 39801 52085 40035
tri 52121 40002 52137 40018 se
rect 52137 40002 52214 40018
rect 52121 39936 52214 40002
rect 52121 39834 52214 39900
tri 52121 39818 52137 39834 ne
rect 52137 39818 52214 39834
rect 51954 39719 52102 39801
rect 51842 39686 51919 39702
tri 51919 39686 51935 39702 sw
rect 51842 39620 51935 39686
rect 51971 39561 52085 39719
tri 52121 39686 52137 39702 se
rect 52137 39686 52214 39702
rect 52121 39620 52214 39686
rect 51842 39485 52214 39561
rect 51842 39360 51935 39426
rect 51842 39344 51919 39360
tri 51919 39344 51935 39360 nw
rect 51971 39327 52085 39485
rect 52121 39360 52214 39426
tri 52121 39344 52137 39360 ne
rect 52137 39344 52214 39360
rect 51954 39245 52102 39327
rect 51842 39212 51919 39228
tri 51919 39212 51935 39228 sw
rect 51842 39146 51935 39212
rect 51842 39044 51935 39110
rect 51842 39028 51919 39044
tri 51919 39028 51935 39044 nw
rect 51971 39011 52085 39245
tri 52121 39212 52137 39228 se
rect 52137 39212 52214 39228
rect 52121 39146 52214 39212
rect 52121 39044 52214 39110
tri 52121 39028 52137 39044 ne
rect 52137 39028 52214 39044
rect 51954 38929 52102 39011
rect 51842 38896 51919 38912
tri 51919 38896 51935 38912 sw
rect 51842 38830 51935 38896
rect 51971 38771 52085 38929
tri 52121 38896 52137 38912 se
rect 52137 38896 52214 38912
rect 52121 38830 52214 38896
rect 51842 38695 52214 38771
rect 51842 38570 51935 38636
rect 51842 38554 51919 38570
tri 51919 38554 51935 38570 nw
rect 51971 38537 52085 38695
rect 52121 38570 52214 38636
tri 52121 38554 52137 38570 ne
rect 52137 38554 52214 38570
rect 51954 38455 52102 38537
rect 51842 38422 51919 38438
tri 51919 38422 51935 38438 sw
rect 51842 38356 51935 38422
rect 51842 38254 51935 38320
rect 51842 38238 51919 38254
tri 51919 38238 51935 38254 nw
rect 51971 38221 52085 38455
tri 52121 38422 52137 38438 se
rect 52137 38422 52214 38438
rect 52121 38356 52214 38422
rect 52121 38254 52214 38320
tri 52121 38238 52137 38254 ne
rect 52137 38238 52214 38254
rect 51954 38139 52102 38221
rect 51842 38106 51919 38122
tri 51919 38106 51935 38122 sw
rect 51842 38040 51935 38106
rect 51971 37981 52085 38139
tri 52121 38106 52137 38122 se
rect 52137 38106 52214 38122
rect 52121 38040 52214 38106
rect 51842 37905 52214 37981
rect 51842 37780 51935 37846
rect 51842 37764 51919 37780
tri 51919 37764 51935 37780 nw
rect 51971 37747 52085 37905
rect 52121 37780 52214 37846
tri 52121 37764 52137 37780 ne
rect 52137 37764 52214 37780
rect 51954 37665 52102 37747
rect 51842 37632 51919 37648
tri 51919 37632 51935 37648 sw
rect 51842 37566 51935 37632
rect 51842 37464 51935 37530
rect 51842 37448 51919 37464
tri 51919 37448 51935 37464 nw
rect 51971 37431 52085 37665
tri 52121 37632 52137 37648 se
rect 52137 37632 52214 37648
rect 52121 37566 52214 37632
rect 52121 37464 52214 37530
tri 52121 37448 52137 37464 ne
rect 52137 37448 52214 37464
rect 51954 37349 52102 37431
rect 51842 37316 51919 37332
tri 51919 37316 51935 37332 sw
rect 51842 37250 51935 37316
rect 51971 37191 52085 37349
tri 52121 37316 52137 37332 se
rect 52137 37316 52214 37332
rect 52121 37250 52214 37316
rect 51842 37115 52214 37191
rect 51842 36990 51935 37056
rect 51842 36974 51919 36990
tri 51919 36974 51935 36990 nw
rect 51971 36957 52085 37115
rect 52121 36990 52214 37056
tri 52121 36974 52137 36990 ne
rect 52137 36974 52214 36990
rect 51954 36875 52102 36957
rect 51842 36842 51919 36858
tri 51919 36842 51935 36858 sw
rect 51842 36776 51935 36842
rect 51842 36674 51935 36740
rect 51842 36658 51919 36674
tri 51919 36658 51935 36674 nw
rect 51971 36641 52085 36875
tri 52121 36842 52137 36858 se
rect 52137 36842 52214 36858
rect 52121 36776 52214 36842
rect 52121 36674 52214 36740
tri 52121 36658 52137 36674 ne
rect 52137 36658 52214 36674
rect 51954 36559 52102 36641
rect 51842 36526 51919 36542
tri 51919 36526 51935 36542 sw
rect 51842 36460 51935 36526
rect 51971 36401 52085 36559
tri 52121 36526 52137 36542 se
rect 52137 36526 52214 36542
rect 52121 36460 52214 36526
rect 51842 36325 52214 36401
rect 51842 36200 51935 36266
rect 51842 36184 51919 36200
tri 51919 36184 51935 36200 nw
rect 51971 36167 52085 36325
rect 52121 36200 52214 36266
tri 52121 36184 52137 36200 ne
rect 52137 36184 52214 36200
rect 51954 36085 52102 36167
rect 51842 36052 51919 36068
tri 51919 36052 51935 36068 sw
rect 51842 35986 51935 36052
rect 51842 35884 51935 35950
rect 51842 35868 51919 35884
tri 51919 35868 51935 35884 nw
rect 51971 35851 52085 36085
tri 52121 36052 52137 36068 se
rect 52137 36052 52214 36068
rect 52121 35986 52214 36052
rect 52121 35884 52214 35950
tri 52121 35868 52137 35884 ne
rect 52137 35868 52214 35884
rect 51954 35769 52102 35851
rect 51842 35736 51919 35752
tri 51919 35736 51935 35752 sw
rect 51842 35670 51935 35736
rect 51971 35611 52085 35769
tri 52121 35736 52137 35752 se
rect 52137 35736 52214 35752
rect 52121 35670 52214 35736
rect 51842 35535 52214 35611
rect 51842 35410 51935 35476
rect 51842 35394 51919 35410
tri 51919 35394 51935 35410 nw
rect 51971 35377 52085 35535
rect 52121 35410 52214 35476
tri 52121 35394 52137 35410 ne
rect 52137 35394 52214 35410
rect 51954 35295 52102 35377
rect 51842 35262 51919 35278
tri 51919 35262 51935 35278 sw
rect 51842 35196 51935 35262
rect 51842 35094 51935 35160
rect 51842 35078 51919 35094
tri 51919 35078 51935 35094 nw
rect 51971 35061 52085 35295
tri 52121 35262 52137 35278 se
rect 52137 35262 52214 35278
rect 52121 35196 52214 35262
rect 52121 35094 52214 35160
tri 52121 35078 52137 35094 ne
rect 52137 35078 52214 35094
rect 51954 34979 52102 35061
rect 51842 34946 51919 34962
tri 51919 34946 51935 34962 sw
rect 51842 34880 51935 34946
rect 51971 34821 52085 34979
tri 52121 34946 52137 34962 se
rect 52137 34946 52214 34962
rect 52121 34880 52214 34946
rect 51842 34745 52214 34821
rect 51842 34620 51935 34686
rect 51842 34604 51919 34620
tri 51919 34604 51935 34620 nw
rect 51971 34587 52085 34745
rect 52121 34620 52214 34686
tri 52121 34604 52137 34620 ne
rect 52137 34604 52214 34620
rect 51954 34505 52102 34587
rect 51842 34472 51919 34488
tri 51919 34472 51935 34488 sw
rect 51842 34406 51935 34472
rect 51842 34304 51935 34370
rect 51842 34288 51919 34304
tri 51919 34288 51935 34304 nw
rect 51971 34271 52085 34505
tri 52121 34472 52137 34488 se
rect 52137 34472 52214 34488
rect 52121 34406 52214 34472
rect 52121 34304 52214 34370
tri 52121 34288 52137 34304 ne
rect 52137 34288 52214 34304
rect 51954 34189 52102 34271
rect 51842 34156 51919 34172
tri 51919 34156 51935 34172 sw
rect 51842 34090 51935 34156
rect 51971 34031 52085 34189
tri 52121 34156 52137 34172 se
rect 52137 34156 52214 34172
rect 52121 34090 52214 34156
rect 51842 33955 52214 34031
rect 51842 33830 51935 33896
rect 51842 33814 51919 33830
tri 51919 33814 51935 33830 nw
rect 51971 33797 52085 33955
rect 52121 33830 52214 33896
tri 52121 33814 52137 33830 ne
rect 52137 33814 52214 33830
rect 51954 33715 52102 33797
rect 51842 33682 51919 33698
tri 51919 33682 51935 33698 sw
rect 51842 33616 51935 33682
rect 51842 33514 51935 33580
rect 51842 33498 51919 33514
tri 51919 33498 51935 33514 nw
rect 51971 33481 52085 33715
tri 52121 33682 52137 33698 se
rect 52137 33682 52214 33698
rect 52121 33616 52214 33682
rect 52121 33514 52214 33580
tri 52121 33498 52137 33514 ne
rect 52137 33498 52214 33514
rect 51954 33399 52102 33481
rect 51842 33366 51919 33382
tri 51919 33366 51935 33382 sw
rect 51842 33300 51935 33366
rect 51971 33241 52085 33399
tri 52121 33366 52137 33382 se
rect 52137 33366 52214 33382
rect 52121 33300 52214 33366
rect 51842 33165 52214 33241
rect 51842 33040 51935 33106
rect 51842 33024 51919 33040
tri 51919 33024 51935 33040 nw
rect 51971 33007 52085 33165
rect 52121 33040 52214 33106
tri 52121 33024 52137 33040 ne
rect 52137 33024 52214 33040
rect 51954 32925 52102 33007
rect 51842 32892 51919 32908
tri 51919 32892 51935 32908 sw
rect 51842 32826 51935 32892
rect 51842 32724 51935 32790
rect 51842 32708 51919 32724
tri 51919 32708 51935 32724 nw
rect 51971 32691 52085 32925
tri 52121 32892 52137 32908 se
rect 52137 32892 52214 32908
rect 52121 32826 52214 32892
rect 52121 32724 52214 32790
tri 52121 32708 52137 32724 ne
rect 52137 32708 52214 32724
rect 51954 32609 52102 32691
rect 51842 32576 51919 32592
tri 51919 32576 51935 32592 sw
rect 51842 32510 51935 32576
rect 51971 32451 52085 32609
tri 52121 32576 52137 32592 se
rect 52137 32576 52214 32592
rect 52121 32510 52214 32576
rect 51842 32375 52214 32451
rect 51842 32250 51935 32316
rect 51842 32234 51919 32250
tri 51919 32234 51935 32250 nw
rect 51971 32217 52085 32375
rect 52121 32250 52214 32316
tri 52121 32234 52137 32250 ne
rect 52137 32234 52214 32250
rect 51954 32135 52102 32217
rect 51842 32102 51919 32118
tri 51919 32102 51935 32118 sw
rect 51842 32036 51935 32102
rect 51842 31934 51935 32000
rect 51842 31918 51919 31934
tri 51919 31918 51935 31934 nw
rect 51971 31901 52085 32135
tri 52121 32102 52137 32118 se
rect 52137 32102 52214 32118
rect 52121 32036 52214 32102
rect 52121 31934 52214 32000
tri 52121 31918 52137 31934 ne
rect 52137 31918 52214 31934
rect 51954 31819 52102 31901
rect 51842 31786 51919 31802
tri 51919 31786 51935 31802 sw
rect 51842 31720 51935 31786
rect 51971 31661 52085 31819
tri 52121 31786 52137 31802 se
rect 52137 31786 52214 31802
rect 52121 31720 52214 31786
rect 51842 31585 52214 31661
rect 51842 31460 51935 31526
rect 51842 31444 51919 31460
tri 51919 31444 51935 31460 nw
rect 51971 31427 52085 31585
rect 52121 31460 52214 31526
tri 52121 31444 52137 31460 ne
rect 52137 31444 52214 31460
rect 51954 31345 52102 31427
rect 51842 31312 51919 31328
tri 51919 31312 51935 31328 sw
rect 51842 31246 51935 31312
rect 51842 31144 51935 31210
rect 51842 31128 51919 31144
tri 51919 31128 51935 31144 nw
rect 51971 31111 52085 31345
tri 52121 31312 52137 31328 se
rect 52137 31312 52214 31328
rect 52121 31246 52214 31312
rect 52121 31144 52214 31210
tri 52121 31128 52137 31144 ne
rect 52137 31128 52214 31144
rect 51954 31029 52102 31111
rect 51842 30996 51919 31012
tri 51919 30996 51935 31012 sw
rect 51842 30930 51935 30996
rect 51971 30871 52085 31029
tri 52121 30996 52137 31012 se
rect 52137 30996 52214 31012
rect 52121 30930 52214 30996
rect 51842 30795 52214 30871
rect 51842 30670 51935 30736
rect 51842 30654 51919 30670
tri 51919 30654 51935 30670 nw
rect 51971 30637 52085 30795
rect 52121 30670 52214 30736
tri 52121 30654 52137 30670 ne
rect 52137 30654 52214 30670
rect 51954 30555 52102 30637
rect 51842 30522 51919 30538
tri 51919 30522 51935 30538 sw
rect 51842 30456 51935 30522
rect 51842 30354 51935 30420
rect 51842 30338 51919 30354
tri 51919 30338 51935 30354 nw
rect 51971 30321 52085 30555
tri 52121 30522 52137 30538 se
rect 52137 30522 52214 30538
rect 52121 30456 52214 30522
rect 52121 30354 52214 30420
tri 52121 30338 52137 30354 ne
rect 52137 30338 52214 30354
rect 51954 30239 52102 30321
rect 51842 30206 51919 30222
tri 51919 30206 51935 30222 sw
rect 51842 30140 51935 30206
rect 51971 30081 52085 30239
tri 52121 30206 52137 30222 se
rect 52137 30206 52214 30222
rect 52121 30140 52214 30206
rect 51842 30005 52214 30081
rect 51842 29880 51935 29946
rect 51842 29864 51919 29880
tri 51919 29864 51935 29880 nw
rect 51971 29847 52085 30005
rect 52121 29880 52214 29946
tri 52121 29864 52137 29880 ne
rect 52137 29864 52214 29880
rect 51954 29765 52102 29847
rect 51842 29732 51919 29748
tri 51919 29732 51935 29748 sw
rect 51842 29666 51935 29732
rect 51842 29564 51935 29630
rect 51842 29548 51919 29564
tri 51919 29548 51935 29564 nw
rect 51971 29531 52085 29765
tri 52121 29732 52137 29748 se
rect 52137 29732 52214 29748
rect 52121 29666 52214 29732
rect 52121 29564 52214 29630
tri 52121 29548 52137 29564 ne
rect 52137 29548 52214 29564
rect 51954 29449 52102 29531
rect 51842 29416 51919 29432
tri 51919 29416 51935 29432 sw
rect 51842 29350 51935 29416
rect 51971 29291 52085 29449
tri 52121 29416 52137 29432 se
rect 52137 29416 52214 29432
rect 52121 29350 52214 29416
rect 51842 29215 52214 29291
rect 51842 29090 51935 29156
rect 51842 29074 51919 29090
tri 51919 29074 51935 29090 nw
rect 51971 29057 52085 29215
rect 52121 29090 52214 29156
tri 52121 29074 52137 29090 ne
rect 52137 29074 52214 29090
rect 51954 28975 52102 29057
rect 51842 28942 51919 28958
tri 51919 28942 51935 28958 sw
rect 51842 28876 51935 28942
rect 51971 28833 52085 28975
tri 52121 28942 52137 28958 se
rect 52137 28942 52214 28958
rect 52121 28876 52214 28942
rect 52250 28463 52286 80603
rect 52322 28463 52358 80603
rect 52394 80445 52430 80603
rect 52386 80303 52438 80445
rect 52394 28763 52430 80303
rect 52386 28621 52438 28763
rect 52394 28463 52430 28621
rect 52466 28463 52502 80603
rect 52538 28463 52574 80603
rect 52610 28833 52694 80233
rect 52730 28463 52766 80603
rect 52802 28463 52838 80603
rect 52874 80445 52910 80603
rect 52866 80303 52918 80445
rect 52874 28763 52910 80303
rect 52866 28621 52918 28763
rect 52874 28463 52910 28621
rect 52946 28463 52982 80603
rect 53018 28463 53054 80603
rect 53090 80124 53183 80190
rect 53090 80108 53167 80124
tri 53167 80108 53183 80124 nw
rect 53219 80091 53333 80233
rect 53369 80124 53462 80190
tri 53369 80108 53385 80124 ne
rect 53385 80108 53462 80124
rect 53202 80009 53350 80091
rect 53090 79976 53167 79992
tri 53167 79976 53183 79992 sw
rect 53090 79910 53183 79976
rect 53219 79851 53333 80009
tri 53369 79976 53385 79992 se
rect 53385 79976 53462 79992
rect 53369 79910 53462 79976
rect 53090 79775 53462 79851
rect 53090 79650 53183 79716
rect 53090 79634 53167 79650
tri 53167 79634 53183 79650 nw
rect 53219 79617 53333 79775
rect 53369 79650 53462 79716
tri 53369 79634 53385 79650 ne
rect 53385 79634 53462 79650
rect 53202 79535 53350 79617
rect 53090 79502 53167 79518
tri 53167 79502 53183 79518 sw
rect 53090 79436 53183 79502
rect 53090 79334 53183 79400
rect 53090 79318 53167 79334
tri 53167 79318 53183 79334 nw
rect 53219 79301 53333 79535
tri 53369 79502 53385 79518 se
rect 53385 79502 53462 79518
rect 53369 79436 53462 79502
rect 53369 79334 53462 79400
tri 53369 79318 53385 79334 ne
rect 53385 79318 53462 79334
rect 53202 79219 53350 79301
rect 53090 79186 53167 79202
tri 53167 79186 53183 79202 sw
rect 53090 79120 53183 79186
rect 53219 79061 53333 79219
tri 53369 79186 53385 79202 se
rect 53385 79186 53462 79202
rect 53369 79120 53462 79186
rect 53090 78985 53462 79061
rect 53090 78860 53183 78926
rect 53090 78844 53167 78860
tri 53167 78844 53183 78860 nw
rect 53219 78827 53333 78985
rect 53369 78860 53462 78926
tri 53369 78844 53385 78860 ne
rect 53385 78844 53462 78860
rect 53202 78745 53350 78827
rect 53090 78712 53167 78728
tri 53167 78712 53183 78728 sw
rect 53090 78646 53183 78712
rect 53090 78544 53183 78610
rect 53090 78528 53167 78544
tri 53167 78528 53183 78544 nw
rect 53219 78511 53333 78745
tri 53369 78712 53385 78728 se
rect 53385 78712 53462 78728
rect 53369 78646 53462 78712
rect 53369 78544 53462 78610
tri 53369 78528 53385 78544 ne
rect 53385 78528 53462 78544
rect 53202 78429 53350 78511
rect 53090 78396 53167 78412
tri 53167 78396 53183 78412 sw
rect 53090 78330 53183 78396
rect 53219 78271 53333 78429
tri 53369 78396 53385 78412 se
rect 53385 78396 53462 78412
rect 53369 78330 53462 78396
rect 53090 78195 53462 78271
rect 53090 78070 53183 78136
rect 53090 78054 53167 78070
tri 53167 78054 53183 78070 nw
rect 53219 78037 53333 78195
rect 53369 78070 53462 78136
tri 53369 78054 53385 78070 ne
rect 53385 78054 53462 78070
rect 53202 77955 53350 78037
rect 53090 77922 53167 77938
tri 53167 77922 53183 77938 sw
rect 53090 77856 53183 77922
rect 53090 77754 53183 77820
rect 53090 77738 53167 77754
tri 53167 77738 53183 77754 nw
rect 53219 77721 53333 77955
tri 53369 77922 53385 77938 se
rect 53385 77922 53462 77938
rect 53369 77856 53462 77922
rect 53369 77754 53462 77820
tri 53369 77738 53385 77754 ne
rect 53385 77738 53462 77754
rect 53202 77639 53350 77721
rect 53090 77606 53167 77622
tri 53167 77606 53183 77622 sw
rect 53090 77540 53183 77606
rect 53219 77481 53333 77639
tri 53369 77606 53385 77622 se
rect 53385 77606 53462 77622
rect 53369 77540 53462 77606
rect 53090 77405 53462 77481
rect 53090 77280 53183 77346
rect 53090 77264 53167 77280
tri 53167 77264 53183 77280 nw
rect 53219 77247 53333 77405
rect 53369 77280 53462 77346
tri 53369 77264 53385 77280 ne
rect 53385 77264 53462 77280
rect 53202 77165 53350 77247
rect 53090 77132 53167 77148
tri 53167 77132 53183 77148 sw
rect 53090 77066 53183 77132
rect 53090 76964 53183 77030
rect 53090 76948 53167 76964
tri 53167 76948 53183 76964 nw
rect 53219 76931 53333 77165
tri 53369 77132 53385 77148 se
rect 53385 77132 53462 77148
rect 53369 77066 53462 77132
rect 53369 76964 53462 77030
tri 53369 76948 53385 76964 ne
rect 53385 76948 53462 76964
rect 53202 76849 53350 76931
rect 53090 76816 53167 76832
tri 53167 76816 53183 76832 sw
rect 53090 76750 53183 76816
rect 53219 76691 53333 76849
tri 53369 76816 53385 76832 se
rect 53385 76816 53462 76832
rect 53369 76750 53462 76816
rect 53090 76615 53462 76691
rect 53090 76490 53183 76556
rect 53090 76474 53167 76490
tri 53167 76474 53183 76490 nw
rect 53219 76457 53333 76615
rect 53369 76490 53462 76556
tri 53369 76474 53385 76490 ne
rect 53385 76474 53462 76490
rect 53202 76375 53350 76457
rect 53090 76342 53167 76358
tri 53167 76342 53183 76358 sw
rect 53090 76276 53183 76342
rect 53090 76174 53183 76240
rect 53090 76158 53167 76174
tri 53167 76158 53183 76174 nw
rect 53219 76141 53333 76375
tri 53369 76342 53385 76358 se
rect 53385 76342 53462 76358
rect 53369 76276 53462 76342
rect 53369 76174 53462 76240
tri 53369 76158 53385 76174 ne
rect 53385 76158 53462 76174
rect 53202 76059 53350 76141
rect 53090 76026 53167 76042
tri 53167 76026 53183 76042 sw
rect 53090 75960 53183 76026
rect 53219 75901 53333 76059
tri 53369 76026 53385 76042 se
rect 53385 76026 53462 76042
rect 53369 75960 53462 76026
rect 53090 75825 53462 75901
rect 53090 75700 53183 75766
rect 53090 75684 53167 75700
tri 53167 75684 53183 75700 nw
rect 53219 75667 53333 75825
rect 53369 75700 53462 75766
tri 53369 75684 53385 75700 ne
rect 53385 75684 53462 75700
rect 53202 75585 53350 75667
rect 53090 75552 53167 75568
tri 53167 75552 53183 75568 sw
rect 53090 75486 53183 75552
rect 53090 75384 53183 75450
rect 53090 75368 53167 75384
tri 53167 75368 53183 75384 nw
rect 53219 75351 53333 75585
tri 53369 75552 53385 75568 se
rect 53385 75552 53462 75568
rect 53369 75486 53462 75552
rect 53369 75384 53462 75450
tri 53369 75368 53385 75384 ne
rect 53385 75368 53462 75384
rect 53202 75269 53350 75351
rect 53090 75236 53167 75252
tri 53167 75236 53183 75252 sw
rect 53090 75170 53183 75236
rect 53219 75111 53333 75269
tri 53369 75236 53385 75252 se
rect 53385 75236 53462 75252
rect 53369 75170 53462 75236
rect 53090 75035 53462 75111
rect 53090 74910 53183 74976
rect 53090 74894 53167 74910
tri 53167 74894 53183 74910 nw
rect 53219 74877 53333 75035
rect 53369 74910 53462 74976
tri 53369 74894 53385 74910 ne
rect 53385 74894 53462 74910
rect 53202 74795 53350 74877
rect 53090 74762 53167 74778
tri 53167 74762 53183 74778 sw
rect 53090 74696 53183 74762
rect 53090 74594 53183 74660
rect 53090 74578 53167 74594
tri 53167 74578 53183 74594 nw
rect 53219 74561 53333 74795
tri 53369 74762 53385 74778 se
rect 53385 74762 53462 74778
rect 53369 74696 53462 74762
rect 53369 74594 53462 74660
tri 53369 74578 53385 74594 ne
rect 53385 74578 53462 74594
rect 53202 74479 53350 74561
rect 53090 74446 53167 74462
tri 53167 74446 53183 74462 sw
rect 53090 74380 53183 74446
rect 53219 74321 53333 74479
tri 53369 74446 53385 74462 se
rect 53385 74446 53462 74462
rect 53369 74380 53462 74446
rect 53090 74245 53462 74321
rect 53090 74120 53183 74186
rect 53090 74104 53167 74120
tri 53167 74104 53183 74120 nw
rect 53219 74087 53333 74245
rect 53369 74120 53462 74186
tri 53369 74104 53385 74120 ne
rect 53385 74104 53462 74120
rect 53202 74005 53350 74087
rect 53090 73972 53167 73988
tri 53167 73972 53183 73988 sw
rect 53090 73906 53183 73972
rect 53090 73804 53183 73870
rect 53090 73788 53167 73804
tri 53167 73788 53183 73804 nw
rect 53219 73771 53333 74005
tri 53369 73972 53385 73988 se
rect 53385 73972 53462 73988
rect 53369 73906 53462 73972
rect 53369 73804 53462 73870
tri 53369 73788 53385 73804 ne
rect 53385 73788 53462 73804
rect 53202 73689 53350 73771
rect 53090 73656 53167 73672
tri 53167 73656 53183 73672 sw
rect 53090 73590 53183 73656
rect 53219 73531 53333 73689
tri 53369 73656 53385 73672 se
rect 53385 73656 53462 73672
rect 53369 73590 53462 73656
rect 53090 73455 53462 73531
rect 53090 73330 53183 73396
rect 53090 73314 53167 73330
tri 53167 73314 53183 73330 nw
rect 53219 73297 53333 73455
rect 53369 73330 53462 73396
tri 53369 73314 53385 73330 ne
rect 53385 73314 53462 73330
rect 53202 73215 53350 73297
rect 53090 73182 53167 73198
tri 53167 73182 53183 73198 sw
rect 53090 73116 53183 73182
rect 53090 73014 53183 73080
rect 53090 72998 53167 73014
tri 53167 72998 53183 73014 nw
rect 53219 72981 53333 73215
tri 53369 73182 53385 73198 se
rect 53385 73182 53462 73198
rect 53369 73116 53462 73182
rect 53369 73014 53462 73080
tri 53369 72998 53385 73014 ne
rect 53385 72998 53462 73014
rect 53202 72899 53350 72981
rect 53090 72866 53167 72882
tri 53167 72866 53183 72882 sw
rect 53090 72800 53183 72866
rect 53219 72741 53333 72899
tri 53369 72866 53385 72882 se
rect 53385 72866 53462 72882
rect 53369 72800 53462 72866
rect 53090 72665 53462 72741
rect 53090 72540 53183 72606
rect 53090 72524 53167 72540
tri 53167 72524 53183 72540 nw
rect 53219 72507 53333 72665
rect 53369 72540 53462 72606
tri 53369 72524 53385 72540 ne
rect 53385 72524 53462 72540
rect 53202 72425 53350 72507
rect 53090 72392 53167 72408
tri 53167 72392 53183 72408 sw
rect 53090 72326 53183 72392
rect 53090 72224 53183 72290
rect 53090 72208 53167 72224
tri 53167 72208 53183 72224 nw
rect 53219 72191 53333 72425
tri 53369 72392 53385 72408 se
rect 53385 72392 53462 72408
rect 53369 72326 53462 72392
rect 53369 72224 53462 72290
tri 53369 72208 53385 72224 ne
rect 53385 72208 53462 72224
rect 53202 72109 53350 72191
rect 53090 72076 53167 72092
tri 53167 72076 53183 72092 sw
rect 53090 72010 53183 72076
rect 53219 71951 53333 72109
tri 53369 72076 53385 72092 se
rect 53385 72076 53462 72092
rect 53369 72010 53462 72076
rect 53090 71875 53462 71951
rect 53090 71750 53183 71816
rect 53090 71734 53167 71750
tri 53167 71734 53183 71750 nw
rect 53219 71717 53333 71875
rect 53369 71750 53462 71816
tri 53369 71734 53385 71750 ne
rect 53385 71734 53462 71750
rect 53202 71635 53350 71717
rect 53090 71602 53167 71618
tri 53167 71602 53183 71618 sw
rect 53090 71536 53183 71602
rect 53090 71434 53183 71500
rect 53090 71418 53167 71434
tri 53167 71418 53183 71434 nw
rect 53219 71401 53333 71635
tri 53369 71602 53385 71618 se
rect 53385 71602 53462 71618
rect 53369 71536 53462 71602
rect 53369 71434 53462 71500
tri 53369 71418 53385 71434 ne
rect 53385 71418 53462 71434
rect 53202 71319 53350 71401
rect 53090 71286 53167 71302
tri 53167 71286 53183 71302 sw
rect 53090 71220 53183 71286
rect 53219 71161 53333 71319
tri 53369 71286 53385 71302 se
rect 53385 71286 53462 71302
rect 53369 71220 53462 71286
rect 53090 71085 53462 71161
rect 53090 70960 53183 71026
rect 53090 70944 53167 70960
tri 53167 70944 53183 70960 nw
rect 53219 70927 53333 71085
rect 53369 70960 53462 71026
tri 53369 70944 53385 70960 ne
rect 53385 70944 53462 70960
rect 53202 70845 53350 70927
rect 53090 70812 53167 70828
tri 53167 70812 53183 70828 sw
rect 53090 70746 53183 70812
rect 53090 70644 53183 70710
rect 53090 70628 53167 70644
tri 53167 70628 53183 70644 nw
rect 53219 70611 53333 70845
tri 53369 70812 53385 70828 se
rect 53385 70812 53462 70828
rect 53369 70746 53462 70812
rect 53369 70644 53462 70710
tri 53369 70628 53385 70644 ne
rect 53385 70628 53462 70644
rect 53202 70529 53350 70611
rect 53090 70496 53167 70512
tri 53167 70496 53183 70512 sw
rect 53090 70430 53183 70496
rect 53219 70371 53333 70529
tri 53369 70496 53385 70512 se
rect 53385 70496 53462 70512
rect 53369 70430 53462 70496
rect 53090 70295 53462 70371
rect 53090 70170 53183 70236
rect 53090 70154 53167 70170
tri 53167 70154 53183 70170 nw
rect 53219 70137 53333 70295
rect 53369 70170 53462 70236
tri 53369 70154 53385 70170 ne
rect 53385 70154 53462 70170
rect 53202 70055 53350 70137
rect 53090 70022 53167 70038
tri 53167 70022 53183 70038 sw
rect 53090 69956 53183 70022
rect 53090 69854 53183 69920
rect 53090 69838 53167 69854
tri 53167 69838 53183 69854 nw
rect 53219 69821 53333 70055
tri 53369 70022 53385 70038 se
rect 53385 70022 53462 70038
rect 53369 69956 53462 70022
rect 53369 69854 53462 69920
tri 53369 69838 53385 69854 ne
rect 53385 69838 53462 69854
rect 53202 69739 53350 69821
rect 53090 69706 53167 69722
tri 53167 69706 53183 69722 sw
rect 53090 69640 53183 69706
rect 53219 69581 53333 69739
tri 53369 69706 53385 69722 se
rect 53385 69706 53462 69722
rect 53369 69640 53462 69706
rect 53090 69505 53462 69581
rect 53090 69380 53183 69446
rect 53090 69364 53167 69380
tri 53167 69364 53183 69380 nw
rect 53219 69347 53333 69505
rect 53369 69380 53462 69446
tri 53369 69364 53385 69380 ne
rect 53385 69364 53462 69380
rect 53202 69265 53350 69347
rect 53090 69232 53167 69248
tri 53167 69232 53183 69248 sw
rect 53090 69166 53183 69232
rect 53090 69064 53183 69130
rect 53090 69048 53167 69064
tri 53167 69048 53183 69064 nw
rect 53219 69031 53333 69265
tri 53369 69232 53385 69248 se
rect 53385 69232 53462 69248
rect 53369 69166 53462 69232
rect 53369 69064 53462 69130
tri 53369 69048 53385 69064 ne
rect 53385 69048 53462 69064
rect 53202 68949 53350 69031
rect 53090 68916 53167 68932
tri 53167 68916 53183 68932 sw
rect 53090 68850 53183 68916
rect 53219 68791 53333 68949
tri 53369 68916 53385 68932 se
rect 53385 68916 53462 68932
rect 53369 68850 53462 68916
rect 53090 68715 53462 68791
rect 53090 68590 53183 68656
rect 53090 68574 53167 68590
tri 53167 68574 53183 68590 nw
rect 53219 68557 53333 68715
rect 53369 68590 53462 68656
tri 53369 68574 53385 68590 ne
rect 53385 68574 53462 68590
rect 53202 68475 53350 68557
rect 53090 68442 53167 68458
tri 53167 68442 53183 68458 sw
rect 53090 68376 53183 68442
rect 53090 68274 53183 68340
rect 53090 68258 53167 68274
tri 53167 68258 53183 68274 nw
rect 53219 68241 53333 68475
tri 53369 68442 53385 68458 se
rect 53385 68442 53462 68458
rect 53369 68376 53462 68442
rect 53369 68274 53462 68340
tri 53369 68258 53385 68274 ne
rect 53385 68258 53462 68274
rect 53202 68159 53350 68241
rect 53090 68126 53167 68142
tri 53167 68126 53183 68142 sw
rect 53090 68060 53183 68126
rect 53219 68001 53333 68159
tri 53369 68126 53385 68142 se
rect 53385 68126 53462 68142
rect 53369 68060 53462 68126
rect 53090 67925 53462 68001
rect 53090 67800 53183 67866
rect 53090 67784 53167 67800
tri 53167 67784 53183 67800 nw
rect 53219 67767 53333 67925
rect 53369 67800 53462 67866
tri 53369 67784 53385 67800 ne
rect 53385 67784 53462 67800
rect 53202 67685 53350 67767
rect 53090 67652 53167 67668
tri 53167 67652 53183 67668 sw
rect 53090 67586 53183 67652
rect 53090 67484 53183 67550
rect 53090 67468 53167 67484
tri 53167 67468 53183 67484 nw
rect 53219 67451 53333 67685
tri 53369 67652 53385 67668 se
rect 53385 67652 53462 67668
rect 53369 67586 53462 67652
rect 53369 67484 53462 67550
tri 53369 67468 53385 67484 ne
rect 53385 67468 53462 67484
rect 53202 67369 53350 67451
rect 53090 67336 53167 67352
tri 53167 67336 53183 67352 sw
rect 53090 67270 53183 67336
rect 53219 67211 53333 67369
tri 53369 67336 53385 67352 se
rect 53385 67336 53462 67352
rect 53369 67270 53462 67336
rect 53090 67135 53462 67211
rect 53090 67010 53183 67076
rect 53090 66994 53167 67010
tri 53167 66994 53183 67010 nw
rect 53219 66977 53333 67135
rect 53369 67010 53462 67076
tri 53369 66994 53385 67010 ne
rect 53385 66994 53462 67010
rect 53202 66895 53350 66977
rect 53090 66862 53167 66878
tri 53167 66862 53183 66878 sw
rect 53090 66796 53183 66862
rect 53090 66694 53183 66760
rect 53090 66678 53167 66694
tri 53167 66678 53183 66694 nw
rect 53219 66661 53333 66895
tri 53369 66862 53385 66878 se
rect 53385 66862 53462 66878
rect 53369 66796 53462 66862
rect 53369 66694 53462 66760
tri 53369 66678 53385 66694 ne
rect 53385 66678 53462 66694
rect 53202 66579 53350 66661
rect 53090 66546 53167 66562
tri 53167 66546 53183 66562 sw
rect 53090 66480 53183 66546
rect 53219 66421 53333 66579
tri 53369 66546 53385 66562 se
rect 53385 66546 53462 66562
rect 53369 66480 53462 66546
rect 53090 66345 53462 66421
rect 53090 66220 53183 66286
rect 53090 66204 53167 66220
tri 53167 66204 53183 66220 nw
rect 53219 66187 53333 66345
rect 53369 66220 53462 66286
tri 53369 66204 53385 66220 ne
rect 53385 66204 53462 66220
rect 53202 66105 53350 66187
rect 53090 66072 53167 66088
tri 53167 66072 53183 66088 sw
rect 53090 66006 53183 66072
rect 53090 65904 53183 65970
rect 53090 65888 53167 65904
tri 53167 65888 53183 65904 nw
rect 53219 65871 53333 66105
tri 53369 66072 53385 66088 se
rect 53385 66072 53462 66088
rect 53369 66006 53462 66072
rect 53369 65904 53462 65970
tri 53369 65888 53385 65904 ne
rect 53385 65888 53462 65904
rect 53202 65789 53350 65871
rect 53090 65756 53167 65772
tri 53167 65756 53183 65772 sw
rect 53090 65690 53183 65756
rect 53219 65631 53333 65789
tri 53369 65756 53385 65772 se
rect 53385 65756 53462 65772
rect 53369 65690 53462 65756
rect 53090 65555 53462 65631
rect 53090 65430 53183 65496
rect 53090 65414 53167 65430
tri 53167 65414 53183 65430 nw
rect 53219 65397 53333 65555
rect 53369 65430 53462 65496
tri 53369 65414 53385 65430 ne
rect 53385 65414 53462 65430
rect 53202 65315 53350 65397
rect 53090 65282 53167 65298
tri 53167 65282 53183 65298 sw
rect 53090 65216 53183 65282
rect 53090 65114 53183 65180
rect 53090 65098 53167 65114
tri 53167 65098 53183 65114 nw
rect 53219 65081 53333 65315
tri 53369 65282 53385 65298 se
rect 53385 65282 53462 65298
rect 53369 65216 53462 65282
rect 53369 65114 53462 65180
tri 53369 65098 53385 65114 ne
rect 53385 65098 53462 65114
rect 53202 64999 53350 65081
rect 53090 64966 53167 64982
tri 53167 64966 53183 64982 sw
rect 53090 64900 53183 64966
rect 53219 64841 53333 64999
tri 53369 64966 53385 64982 se
rect 53385 64966 53462 64982
rect 53369 64900 53462 64966
rect 53090 64765 53462 64841
rect 53090 64640 53183 64706
rect 53090 64624 53167 64640
tri 53167 64624 53183 64640 nw
rect 53219 64607 53333 64765
rect 53369 64640 53462 64706
tri 53369 64624 53385 64640 ne
rect 53385 64624 53462 64640
rect 53202 64525 53350 64607
rect 53090 64492 53167 64508
tri 53167 64492 53183 64508 sw
rect 53090 64426 53183 64492
rect 53090 64324 53183 64390
rect 53090 64308 53167 64324
tri 53167 64308 53183 64324 nw
rect 53219 64291 53333 64525
tri 53369 64492 53385 64508 se
rect 53385 64492 53462 64508
rect 53369 64426 53462 64492
rect 53369 64324 53462 64390
tri 53369 64308 53385 64324 ne
rect 53385 64308 53462 64324
rect 53202 64209 53350 64291
rect 53090 64176 53167 64192
tri 53167 64176 53183 64192 sw
rect 53090 64110 53183 64176
rect 53219 64051 53333 64209
tri 53369 64176 53385 64192 se
rect 53385 64176 53462 64192
rect 53369 64110 53462 64176
rect 53090 63975 53462 64051
rect 53090 63850 53183 63916
rect 53090 63834 53167 63850
tri 53167 63834 53183 63850 nw
rect 53219 63817 53333 63975
rect 53369 63850 53462 63916
tri 53369 63834 53385 63850 ne
rect 53385 63834 53462 63850
rect 53202 63735 53350 63817
rect 53090 63702 53167 63718
tri 53167 63702 53183 63718 sw
rect 53090 63636 53183 63702
rect 53090 63534 53183 63600
rect 53090 63518 53167 63534
tri 53167 63518 53183 63534 nw
rect 53219 63501 53333 63735
tri 53369 63702 53385 63718 se
rect 53385 63702 53462 63718
rect 53369 63636 53462 63702
rect 53369 63534 53462 63600
tri 53369 63518 53385 63534 ne
rect 53385 63518 53462 63534
rect 53202 63419 53350 63501
rect 53090 63386 53167 63402
tri 53167 63386 53183 63402 sw
rect 53090 63320 53183 63386
rect 53219 63261 53333 63419
tri 53369 63386 53385 63402 se
rect 53385 63386 53462 63402
rect 53369 63320 53462 63386
rect 53090 63185 53462 63261
rect 53090 63060 53183 63126
rect 53090 63044 53167 63060
tri 53167 63044 53183 63060 nw
rect 53219 63027 53333 63185
rect 53369 63060 53462 63126
tri 53369 63044 53385 63060 ne
rect 53385 63044 53462 63060
rect 53202 62945 53350 63027
rect 53090 62912 53167 62928
tri 53167 62912 53183 62928 sw
rect 53090 62846 53183 62912
rect 53090 62744 53183 62810
rect 53090 62728 53167 62744
tri 53167 62728 53183 62744 nw
rect 53219 62711 53333 62945
tri 53369 62912 53385 62928 se
rect 53385 62912 53462 62928
rect 53369 62846 53462 62912
rect 53369 62744 53462 62810
tri 53369 62728 53385 62744 ne
rect 53385 62728 53462 62744
rect 53202 62629 53350 62711
rect 53090 62596 53167 62612
tri 53167 62596 53183 62612 sw
rect 53090 62530 53183 62596
rect 53219 62471 53333 62629
tri 53369 62596 53385 62612 se
rect 53385 62596 53462 62612
rect 53369 62530 53462 62596
rect 53090 62395 53462 62471
rect 53090 62270 53183 62336
rect 53090 62254 53167 62270
tri 53167 62254 53183 62270 nw
rect 53219 62237 53333 62395
rect 53369 62270 53462 62336
tri 53369 62254 53385 62270 ne
rect 53385 62254 53462 62270
rect 53202 62155 53350 62237
rect 53090 62122 53167 62138
tri 53167 62122 53183 62138 sw
rect 53090 62056 53183 62122
rect 53090 61954 53183 62020
rect 53090 61938 53167 61954
tri 53167 61938 53183 61954 nw
rect 53219 61921 53333 62155
tri 53369 62122 53385 62138 se
rect 53385 62122 53462 62138
rect 53369 62056 53462 62122
rect 53369 61954 53462 62020
tri 53369 61938 53385 61954 ne
rect 53385 61938 53462 61954
rect 53202 61839 53350 61921
rect 53090 61806 53167 61822
tri 53167 61806 53183 61822 sw
rect 53090 61740 53183 61806
rect 53219 61681 53333 61839
tri 53369 61806 53385 61822 se
rect 53385 61806 53462 61822
rect 53369 61740 53462 61806
rect 53090 61605 53462 61681
rect 53090 61480 53183 61546
rect 53090 61464 53167 61480
tri 53167 61464 53183 61480 nw
rect 53219 61447 53333 61605
rect 53369 61480 53462 61546
tri 53369 61464 53385 61480 ne
rect 53385 61464 53462 61480
rect 53202 61365 53350 61447
rect 53090 61332 53167 61348
tri 53167 61332 53183 61348 sw
rect 53090 61266 53183 61332
rect 53090 61164 53183 61230
rect 53090 61148 53167 61164
tri 53167 61148 53183 61164 nw
rect 53219 61131 53333 61365
tri 53369 61332 53385 61348 se
rect 53385 61332 53462 61348
rect 53369 61266 53462 61332
rect 53369 61164 53462 61230
tri 53369 61148 53385 61164 ne
rect 53385 61148 53462 61164
rect 53202 61049 53350 61131
rect 53090 61016 53167 61032
tri 53167 61016 53183 61032 sw
rect 53090 60950 53183 61016
rect 53219 60891 53333 61049
tri 53369 61016 53385 61032 se
rect 53385 61016 53462 61032
rect 53369 60950 53462 61016
rect 53090 60815 53462 60891
rect 53090 60690 53183 60756
rect 53090 60674 53167 60690
tri 53167 60674 53183 60690 nw
rect 53219 60657 53333 60815
rect 53369 60690 53462 60756
tri 53369 60674 53385 60690 ne
rect 53385 60674 53462 60690
rect 53202 60575 53350 60657
rect 53090 60542 53167 60558
tri 53167 60542 53183 60558 sw
rect 53090 60476 53183 60542
rect 53090 60374 53183 60440
rect 53090 60358 53167 60374
tri 53167 60358 53183 60374 nw
rect 53219 60341 53333 60575
tri 53369 60542 53385 60558 se
rect 53385 60542 53462 60558
rect 53369 60476 53462 60542
rect 53369 60374 53462 60440
tri 53369 60358 53385 60374 ne
rect 53385 60358 53462 60374
rect 53202 60259 53350 60341
rect 53090 60226 53167 60242
tri 53167 60226 53183 60242 sw
rect 53090 60160 53183 60226
rect 53219 60101 53333 60259
tri 53369 60226 53385 60242 se
rect 53385 60226 53462 60242
rect 53369 60160 53462 60226
rect 53090 60025 53462 60101
rect 53090 59900 53183 59966
rect 53090 59884 53167 59900
tri 53167 59884 53183 59900 nw
rect 53219 59867 53333 60025
rect 53369 59900 53462 59966
tri 53369 59884 53385 59900 ne
rect 53385 59884 53462 59900
rect 53202 59785 53350 59867
rect 53090 59752 53167 59768
tri 53167 59752 53183 59768 sw
rect 53090 59686 53183 59752
rect 53090 59584 53183 59650
rect 53090 59568 53167 59584
tri 53167 59568 53183 59584 nw
rect 53219 59551 53333 59785
tri 53369 59752 53385 59768 se
rect 53385 59752 53462 59768
rect 53369 59686 53462 59752
rect 53369 59584 53462 59650
tri 53369 59568 53385 59584 ne
rect 53385 59568 53462 59584
rect 53202 59469 53350 59551
rect 53090 59436 53167 59452
tri 53167 59436 53183 59452 sw
rect 53090 59370 53183 59436
rect 53219 59311 53333 59469
tri 53369 59436 53385 59452 se
rect 53385 59436 53462 59452
rect 53369 59370 53462 59436
rect 53090 59235 53462 59311
rect 53090 59110 53183 59176
rect 53090 59094 53167 59110
tri 53167 59094 53183 59110 nw
rect 53219 59077 53333 59235
rect 53369 59110 53462 59176
tri 53369 59094 53385 59110 ne
rect 53385 59094 53462 59110
rect 53202 58995 53350 59077
rect 53090 58962 53167 58978
tri 53167 58962 53183 58978 sw
rect 53090 58896 53183 58962
rect 53090 58794 53183 58860
rect 53090 58778 53167 58794
tri 53167 58778 53183 58794 nw
rect 53219 58761 53333 58995
tri 53369 58962 53385 58978 se
rect 53385 58962 53462 58978
rect 53369 58896 53462 58962
rect 53369 58794 53462 58860
tri 53369 58778 53385 58794 ne
rect 53385 58778 53462 58794
rect 53202 58679 53350 58761
rect 53090 58646 53167 58662
tri 53167 58646 53183 58662 sw
rect 53090 58580 53183 58646
rect 53219 58521 53333 58679
tri 53369 58646 53385 58662 se
rect 53385 58646 53462 58662
rect 53369 58580 53462 58646
rect 53090 58445 53462 58521
rect 53090 58320 53183 58386
rect 53090 58304 53167 58320
tri 53167 58304 53183 58320 nw
rect 53219 58287 53333 58445
rect 53369 58320 53462 58386
tri 53369 58304 53385 58320 ne
rect 53385 58304 53462 58320
rect 53202 58205 53350 58287
rect 53090 58172 53167 58188
tri 53167 58172 53183 58188 sw
rect 53090 58106 53183 58172
rect 53090 58004 53183 58070
rect 53090 57988 53167 58004
tri 53167 57988 53183 58004 nw
rect 53219 57971 53333 58205
tri 53369 58172 53385 58188 se
rect 53385 58172 53462 58188
rect 53369 58106 53462 58172
rect 53369 58004 53462 58070
tri 53369 57988 53385 58004 ne
rect 53385 57988 53462 58004
rect 53202 57889 53350 57971
rect 53090 57856 53167 57872
tri 53167 57856 53183 57872 sw
rect 53090 57790 53183 57856
rect 53219 57731 53333 57889
tri 53369 57856 53385 57872 se
rect 53385 57856 53462 57872
rect 53369 57790 53462 57856
rect 53090 57655 53462 57731
rect 53090 57530 53183 57596
rect 53090 57514 53167 57530
tri 53167 57514 53183 57530 nw
rect 53219 57497 53333 57655
rect 53369 57530 53462 57596
tri 53369 57514 53385 57530 ne
rect 53385 57514 53462 57530
rect 53202 57415 53350 57497
rect 53090 57382 53167 57398
tri 53167 57382 53183 57398 sw
rect 53090 57316 53183 57382
rect 53090 57214 53183 57280
rect 53090 57198 53167 57214
tri 53167 57198 53183 57214 nw
rect 53219 57181 53333 57415
tri 53369 57382 53385 57398 se
rect 53385 57382 53462 57398
rect 53369 57316 53462 57382
rect 53369 57214 53462 57280
tri 53369 57198 53385 57214 ne
rect 53385 57198 53462 57214
rect 53202 57099 53350 57181
rect 53090 57066 53167 57082
tri 53167 57066 53183 57082 sw
rect 53090 57000 53183 57066
rect 53219 56941 53333 57099
tri 53369 57066 53385 57082 se
rect 53385 57066 53462 57082
rect 53369 57000 53462 57066
rect 53090 56865 53462 56941
rect 53090 56740 53183 56806
rect 53090 56724 53167 56740
tri 53167 56724 53183 56740 nw
rect 53219 56707 53333 56865
rect 53369 56740 53462 56806
tri 53369 56724 53385 56740 ne
rect 53385 56724 53462 56740
rect 53202 56625 53350 56707
rect 53090 56592 53167 56608
tri 53167 56592 53183 56608 sw
rect 53090 56526 53183 56592
rect 53090 56424 53183 56490
rect 53090 56408 53167 56424
tri 53167 56408 53183 56424 nw
rect 53219 56391 53333 56625
tri 53369 56592 53385 56608 se
rect 53385 56592 53462 56608
rect 53369 56526 53462 56592
rect 53369 56424 53462 56490
tri 53369 56408 53385 56424 ne
rect 53385 56408 53462 56424
rect 53202 56309 53350 56391
rect 53090 56276 53167 56292
tri 53167 56276 53183 56292 sw
rect 53090 56210 53183 56276
rect 53219 56151 53333 56309
tri 53369 56276 53385 56292 se
rect 53385 56276 53462 56292
rect 53369 56210 53462 56276
rect 53090 56075 53462 56151
rect 53090 55950 53183 56016
rect 53090 55934 53167 55950
tri 53167 55934 53183 55950 nw
rect 53219 55917 53333 56075
rect 53369 55950 53462 56016
tri 53369 55934 53385 55950 ne
rect 53385 55934 53462 55950
rect 53202 55835 53350 55917
rect 53090 55802 53167 55818
tri 53167 55802 53183 55818 sw
rect 53090 55736 53183 55802
rect 53090 55634 53183 55700
rect 53090 55618 53167 55634
tri 53167 55618 53183 55634 nw
rect 53219 55601 53333 55835
tri 53369 55802 53385 55818 se
rect 53385 55802 53462 55818
rect 53369 55736 53462 55802
rect 53369 55634 53462 55700
tri 53369 55618 53385 55634 ne
rect 53385 55618 53462 55634
rect 53202 55519 53350 55601
rect 53090 55486 53167 55502
tri 53167 55486 53183 55502 sw
rect 53090 55420 53183 55486
rect 53219 55361 53333 55519
tri 53369 55486 53385 55502 se
rect 53385 55486 53462 55502
rect 53369 55420 53462 55486
rect 53090 55285 53462 55361
rect 53090 55160 53183 55226
rect 53090 55144 53167 55160
tri 53167 55144 53183 55160 nw
rect 53219 55127 53333 55285
rect 53369 55160 53462 55226
tri 53369 55144 53385 55160 ne
rect 53385 55144 53462 55160
rect 53202 55045 53350 55127
rect 53090 55012 53167 55028
tri 53167 55012 53183 55028 sw
rect 53090 54946 53183 55012
rect 53090 54844 53183 54910
rect 53090 54828 53167 54844
tri 53167 54828 53183 54844 nw
rect 53219 54811 53333 55045
tri 53369 55012 53385 55028 se
rect 53385 55012 53462 55028
rect 53369 54946 53462 55012
rect 53369 54844 53462 54910
tri 53369 54828 53385 54844 ne
rect 53385 54828 53462 54844
rect 53202 54729 53350 54811
rect 53090 54696 53167 54712
tri 53167 54696 53183 54712 sw
rect 53090 54630 53183 54696
rect 53219 54571 53333 54729
tri 53369 54696 53385 54712 se
rect 53385 54696 53462 54712
rect 53369 54630 53462 54696
rect 53090 54495 53462 54571
rect 53090 54370 53183 54436
rect 53090 54354 53167 54370
tri 53167 54354 53183 54370 nw
rect 53219 54337 53333 54495
rect 53369 54370 53462 54436
tri 53369 54354 53385 54370 ne
rect 53385 54354 53462 54370
rect 53202 54255 53350 54337
rect 53090 54222 53167 54238
tri 53167 54222 53183 54238 sw
rect 53090 54156 53183 54222
rect 53090 54054 53183 54120
rect 53090 54038 53167 54054
tri 53167 54038 53183 54054 nw
rect 53219 54021 53333 54255
tri 53369 54222 53385 54238 se
rect 53385 54222 53462 54238
rect 53369 54156 53462 54222
rect 53369 54054 53462 54120
tri 53369 54038 53385 54054 ne
rect 53385 54038 53462 54054
rect 53202 53939 53350 54021
rect 53090 53906 53167 53922
tri 53167 53906 53183 53922 sw
rect 53090 53840 53183 53906
rect 53219 53781 53333 53939
tri 53369 53906 53385 53922 se
rect 53385 53906 53462 53922
rect 53369 53840 53462 53906
rect 53090 53705 53462 53781
rect 53090 53580 53183 53646
rect 53090 53564 53167 53580
tri 53167 53564 53183 53580 nw
rect 53219 53547 53333 53705
rect 53369 53580 53462 53646
tri 53369 53564 53385 53580 ne
rect 53385 53564 53462 53580
rect 53202 53465 53350 53547
rect 53090 53432 53167 53448
tri 53167 53432 53183 53448 sw
rect 53090 53366 53183 53432
rect 53090 53264 53183 53330
rect 53090 53248 53167 53264
tri 53167 53248 53183 53264 nw
rect 53219 53231 53333 53465
tri 53369 53432 53385 53448 se
rect 53385 53432 53462 53448
rect 53369 53366 53462 53432
rect 53369 53264 53462 53330
tri 53369 53248 53385 53264 ne
rect 53385 53248 53462 53264
rect 53202 53149 53350 53231
rect 53090 53116 53167 53132
tri 53167 53116 53183 53132 sw
rect 53090 53050 53183 53116
rect 53219 52991 53333 53149
tri 53369 53116 53385 53132 se
rect 53385 53116 53462 53132
rect 53369 53050 53462 53116
rect 53090 52915 53462 52991
rect 53090 52790 53183 52856
rect 53090 52774 53167 52790
tri 53167 52774 53183 52790 nw
rect 53219 52757 53333 52915
rect 53369 52790 53462 52856
tri 53369 52774 53385 52790 ne
rect 53385 52774 53462 52790
rect 53202 52675 53350 52757
rect 53090 52642 53167 52658
tri 53167 52642 53183 52658 sw
rect 53090 52576 53183 52642
rect 53090 52474 53183 52540
rect 53090 52458 53167 52474
tri 53167 52458 53183 52474 nw
rect 53219 52441 53333 52675
tri 53369 52642 53385 52658 se
rect 53385 52642 53462 52658
rect 53369 52576 53462 52642
rect 53369 52474 53462 52540
tri 53369 52458 53385 52474 ne
rect 53385 52458 53462 52474
rect 53202 52359 53350 52441
rect 53090 52326 53167 52342
tri 53167 52326 53183 52342 sw
rect 53090 52260 53183 52326
rect 53219 52201 53333 52359
tri 53369 52326 53385 52342 se
rect 53385 52326 53462 52342
rect 53369 52260 53462 52326
rect 53090 52125 53462 52201
rect 53090 52000 53183 52066
rect 53090 51984 53167 52000
tri 53167 51984 53183 52000 nw
rect 53219 51967 53333 52125
rect 53369 52000 53462 52066
tri 53369 51984 53385 52000 ne
rect 53385 51984 53462 52000
rect 53202 51885 53350 51967
rect 53090 51852 53167 51868
tri 53167 51852 53183 51868 sw
rect 53090 51786 53183 51852
rect 53090 51684 53183 51750
rect 53090 51668 53167 51684
tri 53167 51668 53183 51684 nw
rect 53219 51651 53333 51885
tri 53369 51852 53385 51868 se
rect 53385 51852 53462 51868
rect 53369 51786 53462 51852
rect 53369 51684 53462 51750
tri 53369 51668 53385 51684 ne
rect 53385 51668 53462 51684
rect 53202 51569 53350 51651
rect 53090 51536 53167 51552
tri 53167 51536 53183 51552 sw
rect 53090 51470 53183 51536
rect 53219 51411 53333 51569
tri 53369 51536 53385 51552 se
rect 53385 51536 53462 51552
rect 53369 51470 53462 51536
rect 53090 51335 53462 51411
rect 53090 51210 53183 51276
rect 53090 51194 53167 51210
tri 53167 51194 53183 51210 nw
rect 53219 51177 53333 51335
rect 53369 51210 53462 51276
tri 53369 51194 53385 51210 ne
rect 53385 51194 53462 51210
rect 53202 51095 53350 51177
rect 53090 51062 53167 51078
tri 53167 51062 53183 51078 sw
rect 53090 50996 53183 51062
rect 53090 50894 53183 50960
rect 53090 50878 53167 50894
tri 53167 50878 53183 50894 nw
rect 53219 50861 53333 51095
tri 53369 51062 53385 51078 se
rect 53385 51062 53462 51078
rect 53369 50996 53462 51062
rect 53369 50894 53462 50960
tri 53369 50878 53385 50894 ne
rect 53385 50878 53462 50894
rect 53202 50779 53350 50861
rect 53090 50746 53167 50762
tri 53167 50746 53183 50762 sw
rect 53090 50680 53183 50746
rect 53219 50621 53333 50779
tri 53369 50746 53385 50762 se
rect 53385 50746 53462 50762
rect 53369 50680 53462 50746
rect 53090 50545 53462 50621
rect 53090 50420 53183 50486
rect 53090 50404 53167 50420
tri 53167 50404 53183 50420 nw
rect 53219 50387 53333 50545
rect 53369 50420 53462 50486
tri 53369 50404 53385 50420 ne
rect 53385 50404 53462 50420
rect 53202 50305 53350 50387
rect 53090 50272 53167 50288
tri 53167 50272 53183 50288 sw
rect 53090 50206 53183 50272
rect 53090 50104 53183 50170
rect 53090 50088 53167 50104
tri 53167 50088 53183 50104 nw
rect 53219 50071 53333 50305
tri 53369 50272 53385 50288 se
rect 53385 50272 53462 50288
rect 53369 50206 53462 50272
rect 53369 50104 53462 50170
tri 53369 50088 53385 50104 ne
rect 53385 50088 53462 50104
rect 53202 49989 53350 50071
rect 53090 49956 53167 49972
tri 53167 49956 53183 49972 sw
rect 53090 49890 53183 49956
rect 53219 49831 53333 49989
tri 53369 49956 53385 49972 se
rect 53385 49956 53462 49972
rect 53369 49890 53462 49956
rect 53090 49755 53462 49831
rect 53090 49630 53183 49696
rect 53090 49614 53167 49630
tri 53167 49614 53183 49630 nw
rect 53219 49597 53333 49755
rect 53369 49630 53462 49696
tri 53369 49614 53385 49630 ne
rect 53385 49614 53462 49630
rect 53202 49515 53350 49597
rect 53090 49482 53167 49498
tri 53167 49482 53183 49498 sw
rect 53090 49416 53183 49482
rect 53090 49314 53183 49380
rect 53090 49298 53167 49314
tri 53167 49298 53183 49314 nw
rect 53219 49281 53333 49515
tri 53369 49482 53385 49498 se
rect 53385 49482 53462 49498
rect 53369 49416 53462 49482
rect 53369 49314 53462 49380
tri 53369 49298 53385 49314 ne
rect 53385 49298 53462 49314
rect 53202 49199 53350 49281
rect 53090 49166 53167 49182
tri 53167 49166 53183 49182 sw
rect 53090 49100 53183 49166
rect 53219 49041 53333 49199
tri 53369 49166 53385 49182 se
rect 53385 49166 53462 49182
rect 53369 49100 53462 49166
rect 53090 48965 53462 49041
rect 53090 48840 53183 48906
rect 53090 48824 53167 48840
tri 53167 48824 53183 48840 nw
rect 53219 48807 53333 48965
rect 53369 48840 53462 48906
tri 53369 48824 53385 48840 ne
rect 53385 48824 53462 48840
rect 53202 48725 53350 48807
rect 53090 48692 53167 48708
tri 53167 48692 53183 48708 sw
rect 53090 48626 53183 48692
rect 53090 48524 53183 48590
rect 53090 48508 53167 48524
tri 53167 48508 53183 48524 nw
rect 53219 48491 53333 48725
tri 53369 48692 53385 48708 se
rect 53385 48692 53462 48708
rect 53369 48626 53462 48692
rect 53369 48524 53462 48590
tri 53369 48508 53385 48524 ne
rect 53385 48508 53462 48524
rect 53202 48409 53350 48491
rect 53090 48376 53167 48392
tri 53167 48376 53183 48392 sw
rect 53090 48310 53183 48376
rect 53219 48251 53333 48409
tri 53369 48376 53385 48392 se
rect 53385 48376 53462 48392
rect 53369 48310 53462 48376
rect 53090 48175 53462 48251
rect 53090 48050 53183 48116
rect 53090 48034 53167 48050
tri 53167 48034 53183 48050 nw
rect 53219 48017 53333 48175
rect 53369 48050 53462 48116
tri 53369 48034 53385 48050 ne
rect 53385 48034 53462 48050
rect 53202 47935 53350 48017
rect 53090 47902 53167 47918
tri 53167 47902 53183 47918 sw
rect 53090 47836 53183 47902
rect 53090 47734 53183 47800
rect 53090 47718 53167 47734
tri 53167 47718 53183 47734 nw
rect 53219 47701 53333 47935
tri 53369 47902 53385 47918 se
rect 53385 47902 53462 47918
rect 53369 47836 53462 47902
rect 53369 47734 53462 47800
tri 53369 47718 53385 47734 ne
rect 53385 47718 53462 47734
rect 53202 47619 53350 47701
rect 53090 47586 53167 47602
tri 53167 47586 53183 47602 sw
rect 53090 47520 53183 47586
rect 53219 47461 53333 47619
tri 53369 47586 53385 47602 se
rect 53385 47586 53462 47602
rect 53369 47520 53462 47586
rect 53090 47385 53462 47461
rect 53090 47260 53183 47326
rect 53090 47244 53167 47260
tri 53167 47244 53183 47260 nw
rect 53219 47227 53333 47385
rect 53369 47260 53462 47326
tri 53369 47244 53385 47260 ne
rect 53385 47244 53462 47260
rect 53202 47145 53350 47227
rect 53090 47112 53167 47128
tri 53167 47112 53183 47128 sw
rect 53090 47046 53183 47112
rect 53090 46944 53183 47010
rect 53090 46928 53167 46944
tri 53167 46928 53183 46944 nw
rect 53219 46911 53333 47145
tri 53369 47112 53385 47128 se
rect 53385 47112 53462 47128
rect 53369 47046 53462 47112
rect 53369 46944 53462 47010
tri 53369 46928 53385 46944 ne
rect 53385 46928 53462 46944
rect 53202 46829 53350 46911
rect 53090 46796 53167 46812
tri 53167 46796 53183 46812 sw
rect 53090 46730 53183 46796
rect 53219 46671 53333 46829
tri 53369 46796 53385 46812 se
rect 53385 46796 53462 46812
rect 53369 46730 53462 46796
rect 53090 46595 53462 46671
rect 53090 46470 53183 46536
rect 53090 46454 53167 46470
tri 53167 46454 53183 46470 nw
rect 53219 46437 53333 46595
rect 53369 46470 53462 46536
tri 53369 46454 53385 46470 ne
rect 53385 46454 53462 46470
rect 53202 46355 53350 46437
rect 53090 46322 53167 46338
tri 53167 46322 53183 46338 sw
rect 53090 46256 53183 46322
rect 53090 46154 53183 46220
rect 53090 46138 53167 46154
tri 53167 46138 53183 46154 nw
rect 53219 46121 53333 46355
tri 53369 46322 53385 46338 se
rect 53385 46322 53462 46338
rect 53369 46256 53462 46322
rect 53369 46154 53462 46220
tri 53369 46138 53385 46154 ne
rect 53385 46138 53462 46154
rect 53202 46039 53350 46121
rect 53090 46006 53167 46022
tri 53167 46006 53183 46022 sw
rect 53090 45940 53183 46006
rect 53219 45881 53333 46039
tri 53369 46006 53385 46022 se
rect 53385 46006 53462 46022
rect 53369 45940 53462 46006
rect 53090 45805 53462 45881
rect 53090 45680 53183 45746
rect 53090 45664 53167 45680
tri 53167 45664 53183 45680 nw
rect 53219 45647 53333 45805
rect 53369 45680 53462 45746
tri 53369 45664 53385 45680 ne
rect 53385 45664 53462 45680
rect 53202 45565 53350 45647
rect 53090 45532 53167 45548
tri 53167 45532 53183 45548 sw
rect 53090 45466 53183 45532
rect 53090 45364 53183 45430
rect 53090 45348 53167 45364
tri 53167 45348 53183 45364 nw
rect 53219 45331 53333 45565
tri 53369 45532 53385 45548 se
rect 53385 45532 53462 45548
rect 53369 45466 53462 45532
rect 53369 45364 53462 45430
tri 53369 45348 53385 45364 ne
rect 53385 45348 53462 45364
rect 53202 45249 53350 45331
rect 53090 45216 53167 45232
tri 53167 45216 53183 45232 sw
rect 53090 45150 53183 45216
rect 53219 45091 53333 45249
tri 53369 45216 53385 45232 se
rect 53385 45216 53462 45232
rect 53369 45150 53462 45216
rect 53090 45015 53462 45091
rect 53090 44890 53183 44956
rect 53090 44874 53167 44890
tri 53167 44874 53183 44890 nw
rect 53219 44857 53333 45015
rect 53369 44890 53462 44956
tri 53369 44874 53385 44890 ne
rect 53385 44874 53462 44890
rect 53202 44775 53350 44857
rect 53090 44742 53167 44758
tri 53167 44742 53183 44758 sw
rect 53090 44676 53183 44742
rect 53090 44574 53183 44640
rect 53090 44558 53167 44574
tri 53167 44558 53183 44574 nw
rect 53219 44541 53333 44775
tri 53369 44742 53385 44758 se
rect 53385 44742 53462 44758
rect 53369 44676 53462 44742
rect 53369 44574 53462 44640
tri 53369 44558 53385 44574 ne
rect 53385 44558 53462 44574
rect 53202 44459 53350 44541
rect 53090 44426 53167 44442
tri 53167 44426 53183 44442 sw
rect 53090 44360 53183 44426
rect 53219 44301 53333 44459
tri 53369 44426 53385 44442 se
rect 53385 44426 53462 44442
rect 53369 44360 53462 44426
rect 53090 44225 53462 44301
rect 53090 44100 53183 44166
rect 53090 44084 53167 44100
tri 53167 44084 53183 44100 nw
rect 53219 44067 53333 44225
rect 53369 44100 53462 44166
tri 53369 44084 53385 44100 ne
rect 53385 44084 53462 44100
rect 53202 43985 53350 44067
rect 53090 43952 53167 43968
tri 53167 43952 53183 43968 sw
rect 53090 43886 53183 43952
rect 53090 43784 53183 43850
rect 53090 43768 53167 43784
tri 53167 43768 53183 43784 nw
rect 53219 43751 53333 43985
tri 53369 43952 53385 43968 se
rect 53385 43952 53462 43968
rect 53369 43886 53462 43952
rect 53369 43784 53462 43850
tri 53369 43768 53385 43784 ne
rect 53385 43768 53462 43784
rect 53202 43669 53350 43751
rect 53090 43636 53167 43652
tri 53167 43636 53183 43652 sw
rect 53090 43570 53183 43636
rect 53219 43511 53333 43669
tri 53369 43636 53385 43652 se
rect 53385 43636 53462 43652
rect 53369 43570 53462 43636
rect 53090 43435 53462 43511
rect 53090 43310 53183 43376
rect 53090 43294 53167 43310
tri 53167 43294 53183 43310 nw
rect 53219 43277 53333 43435
rect 53369 43310 53462 43376
tri 53369 43294 53385 43310 ne
rect 53385 43294 53462 43310
rect 53202 43195 53350 43277
rect 53090 43162 53167 43178
tri 53167 43162 53183 43178 sw
rect 53090 43096 53183 43162
rect 53090 42994 53183 43060
rect 53090 42978 53167 42994
tri 53167 42978 53183 42994 nw
rect 53219 42961 53333 43195
tri 53369 43162 53385 43178 se
rect 53385 43162 53462 43178
rect 53369 43096 53462 43162
rect 53369 42994 53462 43060
tri 53369 42978 53385 42994 ne
rect 53385 42978 53462 42994
rect 53202 42879 53350 42961
rect 53090 42846 53167 42862
tri 53167 42846 53183 42862 sw
rect 53090 42780 53183 42846
rect 53219 42721 53333 42879
tri 53369 42846 53385 42862 se
rect 53385 42846 53462 42862
rect 53369 42780 53462 42846
rect 53090 42645 53462 42721
rect 53090 42520 53183 42586
rect 53090 42504 53167 42520
tri 53167 42504 53183 42520 nw
rect 53219 42487 53333 42645
rect 53369 42520 53462 42586
tri 53369 42504 53385 42520 ne
rect 53385 42504 53462 42520
rect 53202 42405 53350 42487
rect 53090 42372 53167 42388
tri 53167 42372 53183 42388 sw
rect 53090 42306 53183 42372
rect 53090 42204 53183 42270
rect 53090 42188 53167 42204
tri 53167 42188 53183 42204 nw
rect 53219 42171 53333 42405
tri 53369 42372 53385 42388 se
rect 53385 42372 53462 42388
rect 53369 42306 53462 42372
rect 53369 42204 53462 42270
tri 53369 42188 53385 42204 ne
rect 53385 42188 53462 42204
rect 53202 42089 53350 42171
rect 53090 42056 53167 42072
tri 53167 42056 53183 42072 sw
rect 53090 41990 53183 42056
rect 53219 41931 53333 42089
tri 53369 42056 53385 42072 se
rect 53385 42056 53462 42072
rect 53369 41990 53462 42056
rect 53090 41855 53462 41931
rect 53090 41730 53183 41796
rect 53090 41714 53167 41730
tri 53167 41714 53183 41730 nw
rect 53219 41697 53333 41855
rect 53369 41730 53462 41796
tri 53369 41714 53385 41730 ne
rect 53385 41714 53462 41730
rect 53202 41615 53350 41697
rect 53090 41582 53167 41598
tri 53167 41582 53183 41598 sw
rect 53090 41516 53183 41582
rect 53090 41414 53183 41480
rect 53090 41398 53167 41414
tri 53167 41398 53183 41414 nw
rect 53219 41381 53333 41615
tri 53369 41582 53385 41598 se
rect 53385 41582 53462 41598
rect 53369 41516 53462 41582
rect 53369 41414 53462 41480
tri 53369 41398 53385 41414 ne
rect 53385 41398 53462 41414
rect 53202 41299 53350 41381
rect 53090 41266 53167 41282
tri 53167 41266 53183 41282 sw
rect 53090 41200 53183 41266
rect 53219 41141 53333 41299
tri 53369 41266 53385 41282 se
rect 53385 41266 53462 41282
rect 53369 41200 53462 41266
rect 53090 41065 53462 41141
rect 53090 40940 53183 41006
rect 53090 40924 53167 40940
tri 53167 40924 53183 40940 nw
rect 53219 40907 53333 41065
rect 53369 40940 53462 41006
tri 53369 40924 53385 40940 ne
rect 53385 40924 53462 40940
rect 53202 40825 53350 40907
rect 53090 40792 53167 40808
tri 53167 40792 53183 40808 sw
rect 53090 40726 53183 40792
rect 53090 40624 53183 40690
rect 53090 40608 53167 40624
tri 53167 40608 53183 40624 nw
rect 53219 40591 53333 40825
tri 53369 40792 53385 40808 se
rect 53385 40792 53462 40808
rect 53369 40726 53462 40792
rect 53369 40624 53462 40690
tri 53369 40608 53385 40624 ne
rect 53385 40608 53462 40624
rect 53202 40509 53350 40591
rect 53090 40476 53167 40492
tri 53167 40476 53183 40492 sw
rect 53090 40410 53183 40476
rect 53219 40351 53333 40509
tri 53369 40476 53385 40492 se
rect 53385 40476 53462 40492
rect 53369 40410 53462 40476
rect 53090 40275 53462 40351
rect 53090 40150 53183 40216
rect 53090 40134 53167 40150
tri 53167 40134 53183 40150 nw
rect 53219 40117 53333 40275
rect 53369 40150 53462 40216
tri 53369 40134 53385 40150 ne
rect 53385 40134 53462 40150
rect 53202 40035 53350 40117
rect 53090 40002 53167 40018
tri 53167 40002 53183 40018 sw
rect 53090 39936 53183 40002
rect 53090 39834 53183 39900
rect 53090 39818 53167 39834
tri 53167 39818 53183 39834 nw
rect 53219 39801 53333 40035
tri 53369 40002 53385 40018 se
rect 53385 40002 53462 40018
rect 53369 39936 53462 40002
rect 53369 39834 53462 39900
tri 53369 39818 53385 39834 ne
rect 53385 39818 53462 39834
rect 53202 39719 53350 39801
rect 53090 39686 53167 39702
tri 53167 39686 53183 39702 sw
rect 53090 39620 53183 39686
rect 53219 39561 53333 39719
tri 53369 39686 53385 39702 se
rect 53385 39686 53462 39702
rect 53369 39620 53462 39686
rect 53090 39485 53462 39561
rect 53090 39360 53183 39426
rect 53090 39344 53167 39360
tri 53167 39344 53183 39360 nw
rect 53219 39327 53333 39485
rect 53369 39360 53462 39426
tri 53369 39344 53385 39360 ne
rect 53385 39344 53462 39360
rect 53202 39245 53350 39327
rect 53090 39212 53167 39228
tri 53167 39212 53183 39228 sw
rect 53090 39146 53183 39212
rect 53090 39044 53183 39110
rect 53090 39028 53167 39044
tri 53167 39028 53183 39044 nw
rect 53219 39011 53333 39245
tri 53369 39212 53385 39228 se
rect 53385 39212 53462 39228
rect 53369 39146 53462 39212
rect 53369 39044 53462 39110
tri 53369 39028 53385 39044 ne
rect 53385 39028 53462 39044
rect 53202 38929 53350 39011
rect 53090 38896 53167 38912
tri 53167 38896 53183 38912 sw
rect 53090 38830 53183 38896
rect 53219 38771 53333 38929
tri 53369 38896 53385 38912 se
rect 53385 38896 53462 38912
rect 53369 38830 53462 38896
rect 53090 38695 53462 38771
rect 53090 38570 53183 38636
rect 53090 38554 53167 38570
tri 53167 38554 53183 38570 nw
rect 53219 38537 53333 38695
rect 53369 38570 53462 38636
tri 53369 38554 53385 38570 ne
rect 53385 38554 53462 38570
rect 53202 38455 53350 38537
rect 53090 38422 53167 38438
tri 53167 38422 53183 38438 sw
rect 53090 38356 53183 38422
rect 53090 38254 53183 38320
rect 53090 38238 53167 38254
tri 53167 38238 53183 38254 nw
rect 53219 38221 53333 38455
tri 53369 38422 53385 38438 se
rect 53385 38422 53462 38438
rect 53369 38356 53462 38422
rect 53369 38254 53462 38320
tri 53369 38238 53385 38254 ne
rect 53385 38238 53462 38254
rect 53202 38139 53350 38221
rect 53090 38106 53167 38122
tri 53167 38106 53183 38122 sw
rect 53090 38040 53183 38106
rect 53219 37981 53333 38139
tri 53369 38106 53385 38122 se
rect 53385 38106 53462 38122
rect 53369 38040 53462 38106
rect 53090 37905 53462 37981
rect 53090 37780 53183 37846
rect 53090 37764 53167 37780
tri 53167 37764 53183 37780 nw
rect 53219 37747 53333 37905
rect 53369 37780 53462 37846
tri 53369 37764 53385 37780 ne
rect 53385 37764 53462 37780
rect 53202 37665 53350 37747
rect 53090 37632 53167 37648
tri 53167 37632 53183 37648 sw
rect 53090 37566 53183 37632
rect 53090 37464 53183 37530
rect 53090 37448 53167 37464
tri 53167 37448 53183 37464 nw
rect 53219 37431 53333 37665
tri 53369 37632 53385 37648 se
rect 53385 37632 53462 37648
rect 53369 37566 53462 37632
rect 53369 37464 53462 37530
tri 53369 37448 53385 37464 ne
rect 53385 37448 53462 37464
rect 53202 37349 53350 37431
rect 53090 37316 53167 37332
tri 53167 37316 53183 37332 sw
rect 53090 37250 53183 37316
rect 53219 37191 53333 37349
tri 53369 37316 53385 37332 se
rect 53385 37316 53462 37332
rect 53369 37250 53462 37316
rect 53090 37115 53462 37191
rect 53090 36990 53183 37056
rect 53090 36974 53167 36990
tri 53167 36974 53183 36990 nw
rect 53219 36957 53333 37115
rect 53369 36990 53462 37056
tri 53369 36974 53385 36990 ne
rect 53385 36974 53462 36990
rect 53202 36875 53350 36957
rect 53090 36842 53167 36858
tri 53167 36842 53183 36858 sw
rect 53090 36776 53183 36842
rect 53090 36674 53183 36740
rect 53090 36658 53167 36674
tri 53167 36658 53183 36674 nw
rect 53219 36641 53333 36875
tri 53369 36842 53385 36858 se
rect 53385 36842 53462 36858
rect 53369 36776 53462 36842
rect 53369 36674 53462 36740
tri 53369 36658 53385 36674 ne
rect 53385 36658 53462 36674
rect 53202 36559 53350 36641
rect 53090 36526 53167 36542
tri 53167 36526 53183 36542 sw
rect 53090 36460 53183 36526
rect 53219 36401 53333 36559
tri 53369 36526 53385 36542 se
rect 53385 36526 53462 36542
rect 53369 36460 53462 36526
rect 53090 36325 53462 36401
rect 53090 36200 53183 36266
rect 53090 36184 53167 36200
tri 53167 36184 53183 36200 nw
rect 53219 36167 53333 36325
rect 53369 36200 53462 36266
tri 53369 36184 53385 36200 ne
rect 53385 36184 53462 36200
rect 53202 36085 53350 36167
rect 53090 36052 53167 36068
tri 53167 36052 53183 36068 sw
rect 53090 35986 53183 36052
rect 53090 35884 53183 35950
rect 53090 35868 53167 35884
tri 53167 35868 53183 35884 nw
rect 53219 35851 53333 36085
tri 53369 36052 53385 36068 se
rect 53385 36052 53462 36068
rect 53369 35986 53462 36052
rect 53369 35884 53462 35950
tri 53369 35868 53385 35884 ne
rect 53385 35868 53462 35884
rect 53202 35769 53350 35851
rect 53090 35736 53167 35752
tri 53167 35736 53183 35752 sw
rect 53090 35670 53183 35736
rect 53219 35611 53333 35769
tri 53369 35736 53385 35752 se
rect 53385 35736 53462 35752
rect 53369 35670 53462 35736
rect 53090 35535 53462 35611
rect 53090 35410 53183 35476
rect 53090 35394 53167 35410
tri 53167 35394 53183 35410 nw
rect 53219 35377 53333 35535
rect 53369 35410 53462 35476
tri 53369 35394 53385 35410 ne
rect 53385 35394 53462 35410
rect 53202 35295 53350 35377
rect 53090 35262 53167 35278
tri 53167 35262 53183 35278 sw
rect 53090 35196 53183 35262
rect 53090 35094 53183 35160
rect 53090 35078 53167 35094
tri 53167 35078 53183 35094 nw
rect 53219 35061 53333 35295
tri 53369 35262 53385 35278 se
rect 53385 35262 53462 35278
rect 53369 35196 53462 35262
rect 53369 35094 53462 35160
tri 53369 35078 53385 35094 ne
rect 53385 35078 53462 35094
rect 53202 34979 53350 35061
rect 53090 34946 53167 34962
tri 53167 34946 53183 34962 sw
rect 53090 34880 53183 34946
rect 53219 34821 53333 34979
tri 53369 34946 53385 34962 se
rect 53385 34946 53462 34962
rect 53369 34880 53462 34946
rect 53090 34745 53462 34821
rect 53090 34620 53183 34686
rect 53090 34604 53167 34620
tri 53167 34604 53183 34620 nw
rect 53219 34587 53333 34745
rect 53369 34620 53462 34686
tri 53369 34604 53385 34620 ne
rect 53385 34604 53462 34620
rect 53202 34505 53350 34587
rect 53090 34472 53167 34488
tri 53167 34472 53183 34488 sw
rect 53090 34406 53183 34472
rect 53090 34304 53183 34370
rect 53090 34288 53167 34304
tri 53167 34288 53183 34304 nw
rect 53219 34271 53333 34505
tri 53369 34472 53385 34488 se
rect 53385 34472 53462 34488
rect 53369 34406 53462 34472
rect 53369 34304 53462 34370
tri 53369 34288 53385 34304 ne
rect 53385 34288 53462 34304
rect 53202 34189 53350 34271
rect 53090 34156 53167 34172
tri 53167 34156 53183 34172 sw
rect 53090 34090 53183 34156
rect 53219 34031 53333 34189
tri 53369 34156 53385 34172 se
rect 53385 34156 53462 34172
rect 53369 34090 53462 34156
rect 53090 33955 53462 34031
rect 53090 33830 53183 33896
rect 53090 33814 53167 33830
tri 53167 33814 53183 33830 nw
rect 53219 33797 53333 33955
rect 53369 33830 53462 33896
tri 53369 33814 53385 33830 ne
rect 53385 33814 53462 33830
rect 53202 33715 53350 33797
rect 53090 33682 53167 33698
tri 53167 33682 53183 33698 sw
rect 53090 33616 53183 33682
rect 53090 33514 53183 33580
rect 53090 33498 53167 33514
tri 53167 33498 53183 33514 nw
rect 53219 33481 53333 33715
tri 53369 33682 53385 33698 se
rect 53385 33682 53462 33698
rect 53369 33616 53462 33682
rect 53369 33514 53462 33580
tri 53369 33498 53385 33514 ne
rect 53385 33498 53462 33514
rect 53202 33399 53350 33481
rect 53090 33366 53167 33382
tri 53167 33366 53183 33382 sw
rect 53090 33300 53183 33366
rect 53219 33241 53333 33399
tri 53369 33366 53385 33382 se
rect 53385 33366 53462 33382
rect 53369 33300 53462 33366
rect 53090 33165 53462 33241
rect 53090 33040 53183 33106
rect 53090 33024 53167 33040
tri 53167 33024 53183 33040 nw
rect 53219 33007 53333 33165
rect 53369 33040 53462 33106
tri 53369 33024 53385 33040 ne
rect 53385 33024 53462 33040
rect 53202 32925 53350 33007
rect 53090 32892 53167 32908
tri 53167 32892 53183 32908 sw
rect 53090 32826 53183 32892
rect 53090 32724 53183 32790
rect 53090 32708 53167 32724
tri 53167 32708 53183 32724 nw
rect 53219 32691 53333 32925
tri 53369 32892 53385 32908 se
rect 53385 32892 53462 32908
rect 53369 32826 53462 32892
rect 53369 32724 53462 32790
tri 53369 32708 53385 32724 ne
rect 53385 32708 53462 32724
rect 53202 32609 53350 32691
rect 53090 32576 53167 32592
tri 53167 32576 53183 32592 sw
rect 53090 32510 53183 32576
rect 53219 32451 53333 32609
tri 53369 32576 53385 32592 se
rect 53385 32576 53462 32592
rect 53369 32510 53462 32576
rect 53090 32375 53462 32451
rect 53090 32250 53183 32316
rect 53090 32234 53167 32250
tri 53167 32234 53183 32250 nw
rect 53219 32217 53333 32375
rect 53369 32250 53462 32316
tri 53369 32234 53385 32250 ne
rect 53385 32234 53462 32250
rect 53202 32135 53350 32217
rect 53090 32102 53167 32118
tri 53167 32102 53183 32118 sw
rect 53090 32036 53183 32102
rect 53090 31934 53183 32000
rect 53090 31918 53167 31934
tri 53167 31918 53183 31934 nw
rect 53219 31901 53333 32135
tri 53369 32102 53385 32118 se
rect 53385 32102 53462 32118
rect 53369 32036 53462 32102
rect 53369 31934 53462 32000
tri 53369 31918 53385 31934 ne
rect 53385 31918 53462 31934
rect 53202 31819 53350 31901
rect 53090 31786 53167 31802
tri 53167 31786 53183 31802 sw
rect 53090 31720 53183 31786
rect 53219 31661 53333 31819
tri 53369 31786 53385 31802 se
rect 53385 31786 53462 31802
rect 53369 31720 53462 31786
rect 53090 31585 53462 31661
rect 53090 31460 53183 31526
rect 53090 31444 53167 31460
tri 53167 31444 53183 31460 nw
rect 53219 31427 53333 31585
rect 53369 31460 53462 31526
tri 53369 31444 53385 31460 ne
rect 53385 31444 53462 31460
rect 53202 31345 53350 31427
rect 53090 31312 53167 31328
tri 53167 31312 53183 31328 sw
rect 53090 31246 53183 31312
rect 53090 31144 53183 31210
rect 53090 31128 53167 31144
tri 53167 31128 53183 31144 nw
rect 53219 31111 53333 31345
tri 53369 31312 53385 31328 se
rect 53385 31312 53462 31328
rect 53369 31246 53462 31312
rect 53369 31144 53462 31210
tri 53369 31128 53385 31144 ne
rect 53385 31128 53462 31144
rect 53202 31029 53350 31111
rect 53090 30996 53167 31012
tri 53167 30996 53183 31012 sw
rect 53090 30930 53183 30996
rect 53219 30871 53333 31029
tri 53369 30996 53385 31012 se
rect 53385 30996 53462 31012
rect 53369 30930 53462 30996
rect 53090 30795 53462 30871
rect 53090 30670 53183 30736
rect 53090 30654 53167 30670
tri 53167 30654 53183 30670 nw
rect 53219 30637 53333 30795
rect 53369 30670 53462 30736
tri 53369 30654 53385 30670 ne
rect 53385 30654 53462 30670
rect 53202 30555 53350 30637
rect 53090 30522 53167 30538
tri 53167 30522 53183 30538 sw
rect 53090 30456 53183 30522
rect 53090 30354 53183 30420
rect 53090 30338 53167 30354
tri 53167 30338 53183 30354 nw
rect 53219 30321 53333 30555
tri 53369 30522 53385 30538 se
rect 53385 30522 53462 30538
rect 53369 30456 53462 30522
rect 53369 30354 53462 30420
tri 53369 30338 53385 30354 ne
rect 53385 30338 53462 30354
rect 53202 30239 53350 30321
rect 53090 30206 53167 30222
tri 53167 30206 53183 30222 sw
rect 53090 30140 53183 30206
rect 53219 30081 53333 30239
tri 53369 30206 53385 30222 se
rect 53385 30206 53462 30222
rect 53369 30140 53462 30206
rect 53090 30005 53462 30081
rect 53090 29880 53183 29946
rect 53090 29864 53167 29880
tri 53167 29864 53183 29880 nw
rect 53219 29847 53333 30005
rect 53369 29880 53462 29946
tri 53369 29864 53385 29880 ne
rect 53385 29864 53462 29880
rect 53202 29765 53350 29847
rect 53090 29732 53167 29748
tri 53167 29732 53183 29748 sw
rect 53090 29666 53183 29732
rect 53090 29564 53183 29630
rect 53090 29548 53167 29564
tri 53167 29548 53183 29564 nw
rect 53219 29531 53333 29765
tri 53369 29732 53385 29748 se
rect 53385 29732 53462 29748
rect 53369 29666 53462 29732
rect 53369 29564 53462 29630
tri 53369 29548 53385 29564 ne
rect 53385 29548 53462 29564
rect 53202 29449 53350 29531
rect 53090 29416 53167 29432
tri 53167 29416 53183 29432 sw
rect 53090 29350 53183 29416
rect 53219 29291 53333 29449
tri 53369 29416 53385 29432 se
rect 53385 29416 53462 29432
rect 53369 29350 53462 29416
rect 53090 29215 53462 29291
rect 53090 29090 53183 29156
rect 53090 29074 53167 29090
tri 53167 29074 53183 29090 nw
rect 53219 29057 53333 29215
rect 53369 29090 53462 29156
tri 53369 29074 53385 29090 ne
rect 53385 29074 53462 29090
rect 53202 28975 53350 29057
rect 53090 28942 53167 28958
tri 53167 28942 53183 28958 sw
rect 53090 28876 53183 28942
rect 53219 28833 53333 28975
tri 53369 28942 53385 28958 se
rect 53385 28942 53462 28958
rect 53369 28876 53462 28942
rect 53498 28463 53534 80603
rect 53570 28463 53606 80603
rect 53642 80445 53678 80603
rect 53634 80303 53686 80445
rect 53642 28763 53678 80303
rect 53634 28621 53686 28763
rect 53642 28463 53678 28621
rect 53714 28463 53750 80603
rect 53786 28463 53822 80603
rect 53858 28833 53942 80233
rect 53978 28463 54014 80603
rect 54050 28463 54086 80603
rect 54122 80445 54158 80603
rect 54114 80303 54166 80445
rect 54122 28763 54158 80303
rect 54114 28621 54166 28763
rect 54122 28463 54158 28621
rect 54194 28463 54230 80603
rect 54266 28463 54302 80603
rect 54338 80124 54431 80190
rect 54338 80108 54415 80124
tri 54415 80108 54431 80124 nw
rect 54467 80091 54581 80233
rect 54617 80124 54710 80190
tri 54617 80108 54633 80124 ne
rect 54633 80108 54710 80124
rect 54450 80009 54598 80091
rect 54338 79976 54415 79992
tri 54415 79976 54431 79992 sw
rect 54338 79910 54431 79976
rect 54467 79851 54581 80009
tri 54617 79976 54633 79992 se
rect 54633 79976 54710 79992
rect 54617 79910 54710 79976
rect 54338 79775 54710 79851
rect 54338 79650 54431 79716
rect 54338 79634 54415 79650
tri 54415 79634 54431 79650 nw
rect 54467 79617 54581 79775
rect 54617 79650 54710 79716
tri 54617 79634 54633 79650 ne
rect 54633 79634 54710 79650
rect 54450 79535 54598 79617
rect 54338 79502 54415 79518
tri 54415 79502 54431 79518 sw
rect 54338 79436 54431 79502
rect 54338 79334 54431 79400
rect 54338 79318 54415 79334
tri 54415 79318 54431 79334 nw
rect 54467 79301 54581 79535
tri 54617 79502 54633 79518 se
rect 54633 79502 54710 79518
rect 54617 79436 54710 79502
rect 54617 79334 54710 79400
tri 54617 79318 54633 79334 ne
rect 54633 79318 54710 79334
rect 54450 79219 54598 79301
rect 54338 79186 54415 79202
tri 54415 79186 54431 79202 sw
rect 54338 79120 54431 79186
rect 54467 79061 54581 79219
tri 54617 79186 54633 79202 se
rect 54633 79186 54710 79202
rect 54617 79120 54710 79186
rect 54338 78985 54710 79061
rect 54338 78860 54431 78926
rect 54338 78844 54415 78860
tri 54415 78844 54431 78860 nw
rect 54467 78827 54581 78985
rect 54617 78860 54710 78926
tri 54617 78844 54633 78860 ne
rect 54633 78844 54710 78860
rect 54450 78745 54598 78827
rect 54338 78712 54415 78728
tri 54415 78712 54431 78728 sw
rect 54338 78646 54431 78712
rect 54338 78544 54431 78610
rect 54338 78528 54415 78544
tri 54415 78528 54431 78544 nw
rect 54467 78511 54581 78745
tri 54617 78712 54633 78728 se
rect 54633 78712 54710 78728
rect 54617 78646 54710 78712
rect 54617 78544 54710 78610
tri 54617 78528 54633 78544 ne
rect 54633 78528 54710 78544
rect 54450 78429 54598 78511
rect 54338 78396 54415 78412
tri 54415 78396 54431 78412 sw
rect 54338 78330 54431 78396
rect 54467 78271 54581 78429
tri 54617 78396 54633 78412 se
rect 54633 78396 54710 78412
rect 54617 78330 54710 78396
rect 54338 78195 54710 78271
rect 54338 78070 54431 78136
rect 54338 78054 54415 78070
tri 54415 78054 54431 78070 nw
rect 54467 78037 54581 78195
rect 54617 78070 54710 78136
tri 54617 78054 54633 78070 ne
rect 54633 78054 54710 78070
rect 54450 77955 54598 78037
rect 54338 77922 54415 77938
tri 54415 77922 54431 77938 sw
rect 54338 77856 54431 77922
rect 54338 77754 54431 77820
rect 54338 77738 54415 77754
tri 54415 77738 54431 77754 nw
rect 54467 77721 54581 77955
tri 54617 77922 54633 77938 se
rect 54633 77922 54710 77938
rect 54617 77856 54710 77922
rect 54617 77754 54710 77820
tri 54617 77738 54633 77754 ne
rect 54633 77738 54710 77754
rect 54450 77639 54598 77721
rect 54338 77606 54415 77622
tri 54415 77606 54431 77622 sw
rect 54338 77540 54431 77606
rect 54467 77481 54581 77639
tri 54617 77606 54633 77622 se
rect 54633 77606 54710 77622
rect 54617 77540 54710 77606
rect 54338 77405 54710 77481
rect 54338 77280 54431 77346
rect 54338 77264 54415 77280
tri 54415 77264 54431 77280 nw
rect 54467 77247 54581 77405
rect 54617 77280 54710 77346
tri 54617 77264 54633 77280 ne
rect 54633 77264 54710 77280
rect 54450 77165 54598 77247
rect 54338 77132 54415 77148
tri 54415 77132 54431 77148 sw
rect 54338 77066 54431 77132
rect 54338 76964 54431 77030
rect 54338 76948 54415 76964
tri 54415 76948 54431 76964 nw
rect 54467 76931 54581 77165
tri 54617 77132 54633 77148 se
rect 54633 77132 54710 77148
rect 54617 77066 54710 77132
rect 54617 76964 54710 77030
tri 54617 76948 54633 76964 ne
rect 54633 76948 54710 76964
rect 54450 76849 54598 76931
rect 54338 76816 54415 76832
tri 54415 76816 54431 76832 sw
rect 54338 76750 54431 76816
rect 54467 76691 54581 76849
tri 54617 76816 54633 76832 se
rect 54633 76816 54710 76832
rect 54617 76750 54710 76816
rect 54338 76615 54710 76691
rect 54338 76490 54431 76556
rect 54338 76474 54415 76490
tri 54415 76474 54431 76490 nw
rect 54467 76457 54581 76615
rect 54617 76490 54710 76556
tri 54617 76474 54633 76490 ne
rect 54633 76474 54710 76490
rect 54450 76375 54598 76457
rect 54338 76342 54415 76358
tri 54415 76342 54431 76358 sw
rect 54338 76276 54431 76342
rect 54338 76174 54431 76240
rect 54338 76158 54415 76174
tri 54415 76158 54431 76174 nw
rect 54467 76141 54581 76375
tri 54617 76342 54633 76358 se
rect 54633 76342 54710 76358
rect 54617 76276 54710 76342
rect 54617 76174 54710 76240
tri 54617 76158 54633 76174 ne
rect 54633 76158 54710 76174
rect 54450 76059 54598 76141
rect 54338 76026 54415 76042
tri 54415 76026 54431 76042 sw
rect 54338 75960 54431 76026
rect 54467 75901 54581 76059
tri 54617 76026 54633 76042 se
rect 54633 76026 54710 76042
rect 54617 75960 54710 76026
rect 54338 75825 54710 75901
rect 54338 75700 54431 75766
rect 54338 75684 54415 75700
tri 54415 75684 54431 75700 nw
rect 54467 75667 54581 75825
rect 54617 75700 54710 75766
tri 54617 75684 54633 75700 ne
rect 54633 75684 54710 75700
rect 54450 75585 54598 75667
rect 54338 75552 54415 75568
tri 54415 75552 54431 75568 sw
rect 54338 75486 54431 75552
rect 54338 75384 54431 75450
rect 54338 75368 54415 75384
tri 54415 75368 54431 75384 nw
rect 54467 75351 54581 75585
tri 54617 75552 54633 75568 se
rect 54633 75552 54710 75568
rect 54617 75486 54710 75552
rect 54617 75384 54710 75450
tri 54617 75368 54633 75384 ne
rect 54633 75368 54710 75384
rect 54450 75269 54598 75351
rect 54338 75236 54415 75252
tri 54415 75236 54431 75252 sw
rect 54338 75170 54431 75236
rect 54467 75111 54581 75269
tri 54617 75236 54633 75252 se
rect 54633 75236 54710 75252
rect 54617 75170 54710 75236
rect 54338 75035 54710 75111
rect 54338 74910 54431 74976
rect 54338 74894 54415 74910
tri 54415 74894 54431 74910 nw
rect 54467 74877 54581 75035
rect 54617 74910 54710 74976
tri 54617 74894 54633 74910 ne
rect 54633 74894 54710 74910
rect 54450 74795 54598 74877
rect 54338 74762 54415 74778
tri 54415 74762 54431 74778 sw
rect 54338 74696 54431 74762
rect 54338 74594 54431 74660
rect 54338 74578 54415 74594
tri 54415 74578 54431 74594 nw
rect 54467 74561 54581 74795
tri 54617 74762 54633 74778 se
rect 54633 74762 54710 74778
rect 54617 74696 54710 74762
rect 54617 74594 54710 74660
tri 54617 74578 54633 74594 ne
rect 54633 74578 54710 74594
rect 54450 74479 54598 74561
rect 54338 74446 54415 74462
tri 54415 74446 54431 74462 sw
rect 54338 74380 54431 74446
rect 54467 74321 54581 74479
tri 54617 74446 54633 74462 se
rect 54633 74446 54710 74462
rect 54617 74380 54710 74446
rect 54338 74245 54710 74321
rect 54338 74120 54431 74186
rect 54338 74104 54415 74120
tri 54415 74104 54431 74120 nw
rect 54467 74087 54581 74245
rect 54617 74120 54710 74186
tri 54617 74104 54633 74120 ne
rect 54633 74104 54710 74120
rect 54450 74005 54598 74087
rect 54338 73972 54415 73988
tri 54415 73972 54431 73988 sw
rect 54338 73906 54431 73972
rect 54338 73804 54431 73870
rect 54338 73788 54415 73804
tri 54415 73788 54431 73804 nw
rect 54467 73771 54581 74005
tri 54617 73972 54633 73988 se
rect 54633 73972 54710 73988
rect 54617 73906 54710 73972
rect 54617 73804 54710 73870
tri 54617 73788 54633 73804 ne
rect 54633 73788 54710 73804
rect 54450 73689 54598 73771
rect 54338 73656 54415 73672
tri 54415 73656 54431 73672 sw
rect 54338 73590 54431 73656
rect 54467 73531 54581 73689
tri 54617 73656 54633 73672 se
rect 54633 73656 54710 73672
rect 54617 73590 54710 73656
rect 54338 73455 54710 73531
rect 54338 73330 54431 73396
rect 54338 73314 54415 73330
tri 54415 73314 54431 73330 nw
rect 54467 73297 54581 73455
rect 54617 73330 54710 73396
tri 54617 73314 54633 73330 ne
rect 54633 73314 54710 73330
rect 54450 73215 54598 73297
rect 54338 73182 54415 73198
tri 54415 73182 54431 73198 sw
rect 54338 73116 54431 73182
rect 54338 73014 54431 73080
rect 54338 72998 54415 73014
tri 54415 72998 54431 73014 nw
rect 54467 72981 54581 73215
tri 54617 73182 54633 73198 se
rect 54633 73182 54710 73198
rect 54617 73116 54710 73182
rect 54617 73014 54710 73080
tri 54617 72998 54633 73014 ne
rect 54633 72998 54710 73014
rect 54450 72899 54598 72981
rect 54338 72866 54415 72882
tri 54415 72866 54431 72882 sw
rect 54338 72800 54431 72866
rect 54467 72741 54581 72899
tri 54617 72866 54633 72882 se
rect 54633 72866 54710 72882
rect 54617 72800 54710 72866
rect 54338 72665 54710 72741
rect 54338 72540 54431 72606
rect 54338 72524 54415 72540
tri 54415 72524 54431 72540 nw
rect 54467 72507 54581 72665
rect 54617 72540 54710 72606
tri 54617 72524 54633 72540 ne
rect 54633 72524 54710 72540
rect 54450 72425 54598 72507
rect 54338 72392 54415 72408
tri 54415 72392 54431 72408 sw
rect 54338 72326 54431 72392
rect 54338 72224 54431 72290
rect 54338 72208 54415 72224
tri 54415 72208 54431 72224 nw
rect 54467 72191 54581 72425
tri 54617 72392 54633 72408 se
rect 54633 72392 54710 72408
rect 54617 72326 54710 72392
rect 54617 72224 54710 72290
tri 54617 72208 54633 72224 ne
rect 54633 72208 54710 72224
rect 54450 72109 54598 72191
rect 54338 72076 54415 72092
tri 54415 72076 54431 72092 sw
rect 54338 72010 54431 72076
rect 54467 71951 54581 72109
tri 54617 72076 54633 72092 se
rect 54633 72076 54710 72092
rect 54617 72010 54710 72076
rect 54338 71875 54710 71951
rect 54338 71750 54431 71816
rect 54338 71734 54415 71750
tri 54415 71734 54431 71750 nw
rect 54467 71717 54581 71875
rect 54617 71750 54710 71816
tri 54617 71734 54633 71750 ne
rect 54633 71734 54710 71750
rect 54450 71635 54598 71717
rect 54338 71602 54415 71618
tri 54415 71602 54431 71618 sw
rect 54338 71536 54431 71602
rect 54338 71434 54431 71500
rect 54338 71418 54415 71434
tri 54415 71418 54431 71434 nw
rect 54467 71401 54581 71635
tri 54617 71602 54633 71618 se
rect 54633 71602 54710 71618
rect 54617 71536 54710 71602
rect 54617 71434 54710 71500
tri 54617 71418 54633 71434 ne
rect 54633 71418 54710 71434
rect 54450 71319 54598 71401
rect 54338 71286 54415 71302
tri 54415 71286 54431 71302 sw
rect 54338 71220 54431 71286
rect 54467 71161 54581 71319
tri 54617 71286 54633 71302 se
rect 54633 71286 54710 71302
rect 54617 71220 54710 71286
rect 54338 71085 54710 71161
rect 54338 70960 54431 71026
rect 54338 70944 54415 70960
tri 54415 70944 54431 70960 nw
rect 54467 70927 54581 71085
rect 54617 70960 54710 71026
tri 54617 70944 54633 70960 ne
rect 54633 70944 54710 70960
rect 54450 70845 54598 70927
rect 54338 70812 54415 70828
tri 54415 70812 54431 70828 sw
rect 54338 70746 54431 70812
rect 54338 70644 54431 70710
rect 54338 70628 54415 70644
tri 54415 70628 54431 70644 nw
rect 54467 70611 54581 70845
tri 54617 70812 54633 70828 se
rect 54633 70812 54710 70828
rect 54617 70746 54710 70812
rect 54617 70644 54710 70710
tri 54617 70628 54633 70644 ne
rect 54633 70628 54710 70644
rect 54450 70529 54598 70611
rect 54338 70496 54415 70512
tri 54415 70496 54431 70512 sw
rect 54338 70430 54431 70496
rect 54467 70371 54581 70529
tri 54617 70496 54633 70512 se
rect 54633 70496 54710 70512
rect 54617 70430 54710 70496
rect 54338 70295 54710 70371
rect 54338 70170 54431 70236
rect 54338 70154 54415 70170
tri 54415 70154 54431 70170 nw
rect 54467 70137 54581 70295
rect 54617 70170 54710 70236
tri 54617 70154 54633 70170 ne
rect 54633 70154 54710 70170
rect 54450 70055 54598 70137
rect 54338 70022 54415 70038
tri 54415 70022 54431 70038 sw
rect 54338 69956 54431 70022
rect 54338 69854 54431 69920
rect 54338 69838 54415 69854
tri 54415 69838 54431 69854 nw
rect 54467 69821 54581 70055
tri 54617 70022 54633 70038 se
rect 54633 70022 54710 70038
rect 54617 69956 54710 70022
rect 54617 69854 54710 69920
tri 54617 69838 54633 69854 ne
rect 54633 69838 54710 69854
rect 54450 69739 54598 69821
rect 54338 69706 54415 69722
tri 54415 69706 54431 69722 sw
rect 54338 69640 54431 69706
rect 54467 69581 54581 69739
tri 54617 69706 54633 69722 se
rect 54633 69706 54710 69722
rect 54617 69640 54710 69706
rect 54338 69505 54710 69581
rect 54338 69380 54431 69446
rect 54338 69364 54415 69380
tri 54415 69364 54431 69380 nw
rect 54467 69347 54581 69505
rect 54617 69380 54710 69446
tri 54617 69364 54633 69380 ne
rect 54633 69364 54710 69380
rect 54450 69265 54598 69347
rect 54338 69232 54415 69248
tri 54415 69232 54431 69248 sw
rect 54338 69166 54431 69232
rect 54338 69064 54431 69130
rect 54338 69048 54415 69064
tri 54415 69048 54431 69064 nw
rect 54467 69031 54581 69265
tri 54617 69232 54633 69248 se
rect 54633 69232 54710 69248
rect 54617 69166 54710 69232
rect 54617 69064 54710 69130
tri 54617 69048 54633 69064 ne
rect 54633 69048 54710 69064
rect 54450 68949 54598 69031
rect 54338 68916 54415 68932
tri 54415 68916 54431 68932 sw
rect 54338 68850 54431 68916
rect 54467 68791 54581 68949
tri 54617 68916 54633 68932 se
rect 54633 68916 54710 68932
rect 54617 68850 54710 68916
rect 54338 68715 54710 68791
rect 54338 68590 54431 68656
rect 54338 68574 54415 68590
tri 54415 68574 54431 68590 nw
rect 54467 68557 54581 68715
rect 54617 68590 54710 68656
tri 54617 68574 54633 68590 ne
rect 54633 68574 54710 68590
rect 54450 68475 54598 68557
rect 54338 68442 54415 68458
tri 54415 68442 54431 68458 sw
rect 54338 68376 54431 68442
rect 54338 68274 54431 68340
rect 54338 68258 54415 68274
tri 54415 68258 54431 68274 nw
rect 54467 68241 54581 68475
tri 54617 68442 54633 68458 se
rect 54633 68442 54710 68458
rect 54617 68376 54710 68442
rect 54617 68274 54710 68340
tri 54617 68258 54633 68274 ne
rect 54633 68258 54710 68274
rect 54450 68159 54598 68241
rect 54338 68126 54415 68142
tri 54415 68126 54431 68142 sw
rect 54338 68060 54431 68126
rect 54467 68001 54581 68159
tri 54617 68126 54633 68142 se
rect 54633 68126 54710 68142
rect 54617 68060 54710 68126
rect 54338 67925 54710 68001
rect 54338 67800 54431 67866
rect 54338 67784 54415 67800
tri 54415 67784 54431 67800 nw
rect 54467 67767 54581 67925
rect 54617 67800 54710 67866
tri 54617 67784 54633 67800 ne
rect 54633 67784 54710 67800
rect 54450 67685 54598 67767
rect 54338 67652 54415 67668
tri 54415 67652 54431 67668 sw
rect 54338 67586 54431 67652
rect 54338 67484 54431 67550
rect 54338 67468 54415 67484
tri 54415 67468 54431 67484 nw
rect 54467 67451 54581 67685
tri 54617 67652 54633 67668 se
rect 54633 67652 54710 67668
rect 54617 67586 54710 67652
rect 54617 67484 54710 67550
tri 54617 67468 54633 67484 ne
rect 54633 67468 54710 67484
rect 54450 67369 54598 67451
rect 54338 67336 54415 67352
tri 54415 67336 54431 67352 sw
rect 54338 67270 54431 67336
rect 54467 67211 54581 67369
tri 54617 67336 54633 67352 se
rect 54633 67336 54710 67352
rect 54617 67270 54710 67336
rect 54338 67135 54710 67211
rect 54338 67010 54431 67076
rect 54338 66994 54415 67010
tri 54415 66994 54431 67010 nw
rect 54467 66977 54581 67135
rect 54617 67010 54710 67076
tri 54617 66994 54633 67010 ne
rect 54633 66994 54710 67010
rect 54450 66895 54598 66977
rect 54338 66862 54415 66878
tri 54415 66862 54431 66878 sw
rect 54338 66796 54431 66862
rect 54338 66694 54431 66760
rect 54338 66678 54415 66694
tri 54415 66678 54431 66694 nw
rect 54467 66661 54581 66895
tri 54617 66862 54633 66878 se
rect 54633 66862 54710 66878
rect 54617 66796 54710 66862
rect 54617 66694 54710 66760
tri 54617 66678 54633 66694 ne
rect 54633 66678 54710 66694
rect 54450 66579 54598 66661
rect 54338 66546 54415 66562
tri 54415 66546 54431 66562 sw
rect 54338 66480 54431 66546
rect 54467 66421 54581 66579
tri 54617 66546 54633 66562 se
rect 54633 66546 54710 66562
rect 54617 66480 54710 66546
rect 54338 66345 54710 66421
rect 54338 66220 54431 66286
rect 54338 66204 54415 66220
tri 54415 66204 54431 66220 nw
rect 54467 66187 54581 66345
rect 54617 66220 54710 66286
tri 54617 66204 54633 66220 ne
rect 54633 66204 54710 66220
rect 54450 66105 54598 66187
rect 54338 66072 54415 66088
tri 54415 66072 54431 66088 sw
rect 54338 66006 54431 66072
rect 54338 65904 54431 65970
rect 54338 65888 54415 65904
tri 54415 65888 54431 65904 nw
rect 54467 65871 54581 66105
tri 54617 66072 54633 66088 se
rect 54633 66072 54710 66088
rect 54617 66006 54710 66072
rect 54617 65904 54710 65970
tri 54617 65888 54633 65904 ne
rect 54633 65888 54710 65904
rect 54450 65789 54598 65871
rect 54338 65756 54415 65772
tri 54415 65756 54431 65772 sw
rect 54338 65690 54431 65756
rect 54467 65631 54581 65789
tri 54617 65756 54633 65772 se
rect 54633 65756 54710 65772
rect 54617 65690 54710 65756
rect 54338 65555 54710 65631
rect 54338 65430 54431 65496
rect 54338 65414 54415 65430
tri 54415 65414 54431 65430 nw
rect 54467 65397 54581 65555
rect 54617 65430 54710 65496
tri 54617 65414 54633 65430 ne
rect 54633 65414 54710 65430
rect 54450 65315 54598 65397
rect 54338 65282 54415 65298
tri 54415 65282 54431 65298 sw
rect 54338 65216 54431 65282
rect 54338 65114 54431 65180
rect 54338 65098 54415 65114
tri 54415 65098 54431 65114 nw
rect 54467 65081 54581 65315
tri 54617 65282 54633 65298 se
rect 54633 65282 54710 65298
rect 54617 65216 54710 65282
rect 54617 65114 54710 65180
tri 54617 65098 54633 65114 ne
rect 54633 65098 54710 65114
rect 54450 64999 54598 65081
rect 54338 64966 54415 64982
tri 54415 64966 54431 64982 sw
rect 54338 64900 54431 64966
rect 54467 64841 54581 64999
tri 54617 64966 54633 64982 se
rect 54633 64966 54710 64982
rect 54617 64900 54710 64966
rect 54338 64765 54710 64841
rect 54338 64640 54431 64706
rect 54338 64624 54415 64640
tri 54415 64624 54431 64640 nw
rect 54467 64607 54581 64765
rect 54617 64640 54710 64706
tri 54617 64624 54633 64640 ne
rect 54633 64624 54710 64640
rect 54450 64525 54598 64607
rect 54338 64492 54415 64508
tri 54415 64492 54431 64508 sw
rect 54338 64426 54431 64492
rect 54338 64324 54431 64390
rect 54338 64308 54415 64324
tri 54415 64308 54431 64324 nw
rect 54467 64291 54581 64525
tri 54617 64492 54633 64508 se
rect 54633 64492 54710 64508
rect 54617 64426 54710 64492
rect 54617 64324 54710 64390
tri 54617 64308 54633 64324 ne
rect 54633 64308 54710 64324
rect 54450 64209 54598 64291
rect 54338 64176 54415 64192
tri 54415 64176 54431 64192 sw
rect 54338 64110 54431 64176
rect 54467 64051 54581 64209
tri 54617 64176 54633 64192 se
rect 54633 64176 54710 64192
rect 54617 64110 54710 64176
rect 54338 63975 54710 64051
rect 54338 63850 54431 63916
rect 54338 63834 54415 63850
tri 54415 63834 54431 63850 nw
rect 54467 63817 54581 63975
rect 54617 63850 54710 63916
tri 54617 63834 54633 63850 ne
rect 54633 63834 54710 63850
rect 54450 63735 54598 63817
rect 54338 63702 54415 63718
tri 54415 63702 54431 63718 sw
rect 54338 63636 54431 63702
rect 54338 63534 54431 63600
rect 54338 63518 54415 63534
tri 54415 63518 54431 63534 nw
rect 54467 63501 54581 63735
tri 54617 63702 54633 63718 se
rect 54633 63702 54710 63718
rect 54617 63636 54710 63702
rect 54617 63534 54710 63600
tri 54617 63518 54633 63534 ne
rect 54633 63518 54710 63534
rect 54450 63419 54598 63501
rect 54338 63386 54415 63402
tri 54415 63386 54431 63402 sw
rect 54338 63320 54431 63386
rect 54467 63261 54581 63419
tri 54617 63386 54633 63402 se
rect 54633 63386 54710 63402
rect 54617 63320 54710 63386
rect 54338 63185 54710 63261
rect 54338 63060 54431 63126
rect 54338 63044 54415 63060
tri 54415 63044 54431 63060 nw
rect 54467 63027 54581 63185
rect 54617 63060 54710 63126
tri 54617 63044 54633 63060 ne
rect 54633 63044 54710 63060
rect 54450 62945 54598 63027
rect 54338 62912 54415 62928
tri 54415 62912 54431 62928 sw
rect 54338 62846 54431 62912
rect 54338 62744 54431 62810
rect 54338 62728 54415 62744
tri 54415 62728 54431 62744 nw
rect 54467 62711 54581 62945
tri 54617 62912 54633 62928 se
rect 54633 62912 54710 62928
rect 54617 62846 54710 62912
rect 54617 62744 54710 62810
tri 54617 62728 54633 62744 ne
rect 54633 62728 54710 62744
rect 54450 62629 54598 62711
rect 54338 62596 54415 62612
tri 54415 62596 54431 62612 sw
rect 54338 62530 54431 62596
rect 54467 62471 54581 62629
tri 54617 62596 54633 62612 se
rect 54633 62596 54710 62612
rect 54617 62530 54710 62596
rect 54338 62395 54710 62471
rect 54338 62270 54431 62336
rect 54338 62254 54415 62270
tri 54415 62254 54431 62270 nw
rect 54467 62237 54581 62395
rect 54617 62270 54710 62336
tri 54617 62254 54633 62270 ne
rect 54633 62254 54710 62270
rect 54450 62155 54598 62237
rect 54338 62122 54415 62138
tri 54415 62122 54431 62138 sw
rect 54338 62056 54431 62122
rect 54338 61954 54431 62020
rect 54338 61938 54415 61954
tri 54415 61938 54431 61954 nw
rect 54467 61921 54581 62155
tri 54617 62122 54633 62138 se
rect 54633 62122 54710 62138
rect 54617 62056 54710 62122
rect 54617 61954 54710 62020
tri 54617 61938 54633 61954 ne
rect 54633 61938 54710 61954
rect 54450 61839 54598 61921
rect 54338 61806 54415 61822
tri 54415 61806 54431 61822 sw
rect 54338 61740 54431 61806
rect 54467 61681 54581 61839
tri 54617 61806 54633 61822 se
rect 54633 61806 54710 61822
rect 54617 61740 54710 61806
rect 54338 61605 54710 61681
rect 54338 61480 54431 61546
rect 54338 61464 54415 61480
tri 54415 61464 54431 61480 nw
rect 54467 61447 54581 61605
rect 54617 61480 54710 61546
tri 54617 61464 54633 61480 ne
rect 54633 61464 54710 61480
rect 54450 61365 54598 61447
rect 54338 61332 54415 61348
tri 54415 61332 54431 61348 sw
rect 54338 61266 54431 61332
rect 54338 61164 54431 61230
rect 54338 61148 54415 61164
tri 54415 61148 54431 61164 nw
rect 54467 61131 54581 61365
tri 54617 61332 54633 61348 se
rect 54633 61332 54710 61348
rect 54617 61266 54710 61332
rect 54617 61164 54710 61230
tri 54617 61148 54633 61164 ne
rect 54633 61148 54710 61164
rect 54450 61049 54598 61131
rect 54338 61016 54415 61032
tri 54415 61016 54431 61032 sw
rect 54338 60950 54431 61016
rect 54467 60891 54581 61049
tri 54617 61016 54633 61032 se
rect 54633 61016 54710 61032
rect 54617 60950 54710 61016
rect 54338 60815 54710 60891
rect 54338 60690 54431 60756
rect 54338 60674 54415 60690
tri 54415 60674 54431 60690 nw
rect 54467 60657 54581 60815
rect 54617 60690 54710 60756
tri 54617 60674 54633 60690 ne
rect 54633 60674 54710 60690
rect 54450 60575 54598 60657
rect 54338 60542 54415 60558
tri 54415 60542 54431 60558 sw
rect 54338 60476 54431 60542
rect 54338 60374 54431 60440
rect 54338 60358 54415 60374
tri 54415 60358 54431 60374 nw
rect 54467 60341 54581 60575
tri 54617 60542 54633 60558 se
rect 54633 60542 54710 60558
rect 54617 60476 54710 60542
rect 54617 60374 54710 60440
tri 54617 60358 54633 60374 ne
rect 54633 60358 54710 60374
rect 54450 60259 54598 60341
rect 54338 60226 54415 60242
tri 54415 60226 54431 60242 sw
rect 54338 60160 54431 60226
rect 54467 60101 54581 60259
tri 54617 60226 54633 60242 se
rect 54633 60226 54710 60242
rect 54617 60160 54710 60226
rect 54338 60025 54710 60101
rect 54338 59900 54431 59966
rect 54338 59884 54415 59900
tri 54415 59884 54431 59900 nw
rect 54467 59867 54581 60025
rect 54617 59900 54710 59966
tri 54617 59884 54633 59900 ne
rect 54633 59884 54710 59900
rect 54450 59785 54598 59867
rect 54338 59752 54415 59768
tri 54415 59752 54431 59768 sw
rect 54338 59686 54431 59752
rect 54338 59584 54431 59650
rect 54338 59568 54415 59584
tri 54415 59568 54431 59584 nw
rect 54467 59551 54581 59785
tri 54617 59752 54633 59768 se
rect 54633 59752 54710 59768
rect 54617 59686 54710 59752
rect 54617 59584 54710 59650
tri 54617 59568 54633 59584 ne
rect 54633 59568 54710 59584
rect 54450 59469 54598 59551
rect 54338 59436 54415 59452
tri 54415 59436 54431 59452 sw
rect 54338 59370 54431 59436
rect 54467 59311 54581 59469
tri 54617 59436 54633 59452 se
rect 54633 59436 54710 59452
rect 54617 59370 54710 59436
rect 54338 59235 54710 59311
rect 54338 59110 54431 59176
rect 54338 59094 54415 59110
tri 54415 59094 54431 59110 nw
rect 54467 59077 54581 59235
rect 54617 59110 54710 59176
tri 54617 59094 54633 59110 ne
rect 54633 59094 54710 59110
rect 54450 58995 54598 59077
rect 54338 58962 54415 58978
tri 54415 58962 54431 58978 sw
rect 54338 58896 54431 58962
rect 54338 58794 54431 58860
rect 54338 58778 54415 58794
tri 54415 58778 54431 58794 nw
rect 54467 58761 54581 58995
tri 54617 58962 54633 58978 se
rect 54633 58962 54710 58978
rect 54617 58896 54710 58962
rect 54617 58794 54710 58860
tri 54617 58778 54633 58794 ne
rect 54633 58778 54710 58794
rect 54450 58679 54598 58761
rect 54338 58646 54415 58662
tri 54415 58646 54431 58662 sw
rect 54338 58580 54431 58646
rect 54467 58521 54581 58679
tri 54617 58646 54633 58662 se
rect 54633 58646 54710 58662
rect 54617 58580 54710 58646
rect 54338 58445 54710 58521
rect 54338 58320 54431 58386
rect 54338 58304 54415 58320
tri 54415 58304 54431 58320 nw
rect 54467 58287 54581 58445
rect 54617 58320 54710 58386
tri 54617 58304 54633 58320 ne
rect 54633 58304 54710 58320
rect 54450 58205 54598 58287
rect 54338 58172 54415 58188
tri 54415 58172 54431 58188 sw
rect 54338 58106 54431 58172
rect 54338 58004 54431 58070
rect 54338 57988 54415 58004
tri 54415 57988 54431 58004 nw
rect 54467 57971 54581 58205
tri 54617 58172 54633 58188 se
rect 54633 58172 54710 58188
rect 54617 58106 54710 58172
rect 54617 58004 54710 58070
tri 54617 57988 54633 58004 ne
rect 54633 57988 54710 58004
rect 54450 57889 54598 57971
rect 54338 57856 54415 57872
tri 54415 57856 54431 57872 sw
rect 54338 57790 54431 57856
rect 54467 57731 54581 57889
tri 54617 57856 54633 57872 se
rect 54633 57856 54710 57872
rect 54617 57790 54710 57856
rect 54338 57655 54710 57731
rect 54338 57530 54431 57596
rect 54338 57514 54415 57530
tri 54415 57514 54431 57530 nw
rect 54467 57497 54581 57655
rect 54617 57530 54710 57596
tri 54617 57514 54633 57530 ne
rect 54633 57514 54710 57530
rect 54450 57415 54598 57497
rect 54338 57382 54415 57398
tri 54415 57382 54431 57398 sw
rect 54338 57316 54431 57382
rect 54338 57214 54431 57280
rect 54338 57198 54415 57214
tri 54415 57198 54431 57214 nw
rect 54467 57181 54581 57415
tri 54617 57382 54633 57398 se
rect 54633 57382 54710 57398
rect 54617 57316 54710 57382
rect 54617 57214 54710 57280
tri 54617 57198 54633 57214 ne
rect 54633 57198 54710 57214
rect 54450 57099 54598 57181
rect 54338 57066 54415 57082
tri 54415 57066 54431 57082 sw
rect 54338 57000 54431 57066
rect 54467 56941 54581 57099
tri 54617 57066 54633 57082 se
rect 54633 57066 54710 57082
rect 54617 57000 54710 57066
rect 54338 56865 54710 56941
rect 54338 56740 54431 56806
rect 54338 56724 54415 56740
tri 54415 56724 54431 56740 nw
rect 54467 56707 54581 56865
rect 54617 56740 54710 56806
tri 54617 56724 54633 56740 ne
rect 54633 56724 54710 56740
rect 54450 56625 54598 56707
rect 54338 56592 54415 56608
tri 54415 56592 54431 56608 sw
rect 54338 56526 54431 56592
rect 54338 56424 54431 56490
rect 54338 56408 54415 56424
tri 54415 56408 54431 56424 nw
rect 54467 56391 54581 56625
tri 54617 56592 54633 56608 se
rect 54633 56592 54710 56608
rect 54617 56526 54710 56592
rect 54617 56424 54710 56490
tri 54617 56408 54633 56424 ne
rect 54633 56408 54710 56424
rect 54450 56309 54598 56391
rect 54338 56276 54415 56292
tri 54415 56276 54431 56292 sw
rect 54338 56210 54431 56276
rect 54467 56151 54581 56309
tri 54617 56276 54633 56292 se
rect 54633 56276 54710 56292
rect 54617 56210 54710 56276
rect 54338 56075 54710 56151
rect 54338 55950 54431 56016
rect 54338 55934 54415 55950
tri 54415 55934 54431 55950 nw
rect 54467 55917 54581 56075
rect 54617 55950 54710 56016
tri 54617 55934 54633 55950 ne
rect 54633 55934 54710 55950
rect 54450 55835 54598 55917
rect 54338 55802 54415 55818
tri 54415 55802 54431 55818 sw
rect 54338 55736 54431 55802
rect 54338 55634 54431 55700
rect 54338 55618 54415 55634
tri 54415 55618 54431 55634 nw
rect 54467 55601 54581 55835
tri 54617 55802 54633 55818 se
rect 54633 55802 54710 55818
rect 54617 55736 54710 55802
rect 54617 55634 54710 55700
tri 54617 55618 54633 55634 ne
rect 54633 55618 54710 55634
rect 54450 55519 54598 55601
rect 54338 55486 54415 55502
tri 54415 55486 54431 55502 sw
rect 54338 55420 54431 55486
rect 54467 55361 54581 55519
tri 54617 55486 54633 55502 se
rect 54633 55486 54710 55502
rect 54617 55420 54710 55486
rect 54338 55285 54710 55361
rect 54338 55160 54431 55226
rect 54338 55144 54415 55160
tri 54415 55144 54431 55160 nw
rect 54467 55127 54581 55285
rect 54617 55160 54710 55226
tri 54617 55144 54633 55160 ne
rect 54633 55144 54710 55160
rect 54450 55045 54598 55127
rect 54338 55012 54415 55028
tri 54415 55012 54431 55028 sw
rect 54338 54946 54431 55012
rect 54338 54844 54431 54910
rect 54338 54828 54415 54844
tri 54415 54828 54431 54844 nw
rect 54467 54811 54581 55045
tri 54617 55012 54633 55028 se
rect 54633 55012 54710 55028
rect 54617 54946 54710 55012
rect 54617 54844 54710 54910
tri 54617 54828 54633 54844 ne
rect 54633 54828 54710 54844
rect 54450 54729 54598 54811
rect 54338 54696 54415 54712
tri 54415 54696 54431 54712 sw
rect 54338 54630 54431 54696
rect 54467 54571 54581 54729
tri 54617 54696 54633 54712 se
rect 54633 54696 54710 54712
rect 54617 54630 54710 54696
rect 54338 54495 54710 54571
rect 54338 54370 54431 54436
rect 54338 54354 54415 54370
tri 54415 54354 54431 54370 nw
rect 54467 54337 54581 54495
rect 54617 54370 54710 54436
tri 54617 54354 54633 54370 ne
rect 54633 54354 54710 54370
rect 54450 54255 54598 54337
rect 54338 54222 54415 54238
tri 54415 54222 54431 54238 sw
rect 54338 54156 54431 54222
rect 54338 54054 54431 54120
rect 54338 54038 54415 54054
tri 54415 54038 54431 54054 nw
rect 54467 54021 54581 54255
tri 54617 54222 54633 54238 se
rect 54633 54222 54710 54238
rect 54617 54156 54710 54222
rect 54617 54054 54710 54120
tri 54617 54038 54633 54054 ne
rect 54633 54038 54710 54054
rect 54450 53939 54598 54021
rect 54338 53906 54415 53922
tri 54415 53906 54431 53922 sw
rect 54338 53840 54431 53906
rect 54467 53781 54581 53939
tri 54617 53906 54633 53922 se
rect 54633 53906 54710 53922
rect 54617 53840 54710 53906
rect 54338 53705 54710 53781
rect 54338 53580 54431 53646
rect 54338 53564 54415 53580
tri 54415 53564 54431 53580 nw
rect 54467 53547 54581 53705
rect 54617 53580 54710 53646
tri 54617 53564 54633 53580 ne
rect 54633 53564 54710 53580
rect 54450 53465 54598 53547
rect 54338 53432 54415 53448
tri 54415 53432 54431 53448 sw
rect 54338 53366 54431 53432
rect 54338 53264 54431 53330
rect 54338 53248 54415 53264
tri 54415 53248 54431 53264 nw
rect 54467 53231 54581 53465
tri 54617 53432 54633 53448 se
rect 54633 53432 54710 53448
rect 54617 53366 54710 53432
rect 54617 53264 54710 53330
tri 54617 53248 54633 53264 ne
rect 54633 53248 54710 53264
rect 54450 53149 54598 53231
rect 54338 53116 54415 53132
tri 54415 53116 54431 53132 sw
rect 54338 53050 54431 53116
rect 54467 52991 54581 53149
tri 54617 53116 54633 53132 se
rect 54633 53116 54710 53132
rect 54617 53050 54710 53116
rect 54338 52915 54710 52991
rect 54338 52790 54431 52856
rect 54338 52774 54415 52790
tri 54415 52774 54431 52790 nw
rect 54467 52757 54581 52915
rect 54617 52790 54710 52856
tri 54617 52774 54633 52790 ne
rect 54633 52774 54710 52790
rect 54450 52675 54598 52757
rect 54338 52642 54415 52658
tri 54415 52642 54431 52658 sw
rect 54338 52576 54431 52642
rect 54338 52474 54431 52540
rect 54338 52458 54415 52474
tri 54415 52458 54431 52474 nw
rect 54467 52441 54581 52675
tri 54617 52642 54633 52658 se
rect 54633 52642 54710 52658
rect 54617 52576 54710 52642
rect 54617 52474 54710 52540
tri 54617 52458 54633 52474 ne
rect 54633 52458 54710 52474
rect 54450 52359 54598 52441
rect 54338 52326 54415 52342
tri 54415 52326 54431 52342 sw
rect 54338 52260 54431 52326
rect 54467 52201 54581 52359
tri 54617 52326 54633 52342 se
rect 54633 52326 54710 52342
rect 54617 52260 54710 52326
rect 54338 52125 54710 52201
rect 54338 52000 54431 52066
rect 54338 51984 54415 52000
tri 54415 51984 54431 52000 nw
rect 54467 51967 54581 52125
rect 54617 52000 54710 52066
tri 54617 51984 54633 52000 ne
rect 54633 51984 54710 52000
rect 54450 51885 54598 51967
rect 54338 51852 54415 51868
tri 54415 51852 54431 51868 sw
rect 54338 51786 54431 51852
rect 54338 51684 54431 51750
rect 54338 51668 54415 51684
tri 54415 51668 54431 51684 nw
rect 54467 51651 54581 51885
tri 54617 51852 54633 51868 se
rect 54633 51852 54710 51868
rect 54617 51786 54710 51852
rect 54617 51684 54710 51750
tri 54617 51668 54633 51684 ne
rect 54633 51668 54710 51684
rect 54450 51569 54598 51651
rect 54338 51536 54415 51552
tri 54415 51536 54431 51552 sw
rect 54338 51470 54431 51536
rect 54467 51411 54581 51569
tri 54617 51536 54633 51552 se
rect 54633 51536 54710 51552
rect 54617 51470 54710 51536
rect 54338 51335 54710 51411
rect 54338 51210 54431 51276
rect 54338 51194 54415 51210
tri 54415 51194 54431 51210 nw
rect 54467 51177 54581 51335
rect 54617 51210 54710 51276
tri 54617 51194 54633 51210 ne
rect 54633 51194 54710 51210
rect 54450 51095 54598 51177
rect 54338 51062 54415 51078
tri 54415 51062 54431 51078 sw
rect 54338 50996 54431 51062
rect 54338 50894 54431 50960
rect 54338 50878 54415 50894
tri 54415 50878 54431 50894 nw
rect 54467 50861 54581 51095
tri 54617 51062 54633 51078 se
rect 54633 51062 54710 51078
rect 54617 50996 54710 51062
rect 54617 50894 54710 50960
tri 54617 50878 54633 50894 ne
rect 54633 50878 54710 50894
rect 54450 50779 54598 50861
rect 54338 50746 54415 50762
tri 54415 50746 54431 50762 sw
rect 54338 50680 54431 50746
rect 54467 50621 54581 50779
tri 54617 50746 54633 50762 se
rect 54633 50746 54710 50762
rect 54617 50680 54710 50746
rect 54338 50545 54710 50621
rect 54338 50420 54431 50486
rect 54338 50404 54415 50420
tri 54415 50404 54431 50420 nw
rect 54467 50387 54581 50545
rect 54617 50420 54710 50486
tri 54617 50404 54633 50420 ne
rect 54633 50404 54710 50420
rect 54450 50305 54598 50387
rect 54338 50272 54415 50288
tri 54415 50272 54431 50288 sw
rect 54338 50206 54431 50272
rect 54338 50104 54431 50170
rect 54338 50088 54415 50104
tri 54415 50088 54431 50104 nw
rect 54467 50071 54581 50305
tri 54617 50272 54633 50288 se
rect 54633 50272 54710 50288
rect 54617 50206 54710 50272
rect 54617 50104 54710 50170
tri 54617 50088 54633 50104 ne
rect 54633 50088 54710 50104
rect 54450 49989 54598 50071
rect 54338 49956 54415 49972
tri 54415 49956 54431 49972 sw
rect 54338 49890 54431 49956
rect 54467 49831 54581 49989
tri 54617 49956 54633 49972 se
rect 54633 49956 54710 49972
rect 54617 49890 54710 49956
rect 54338 49755 54710 49831
rect 54338 49630 54431 49696
rect 54338 49614 54415 49630
tri 54415 49614 54431 49630 nw
rect 54467 49597 54581 49755
rect 54617 49630 54710 49696
tri 54617 49614 54633 49630 ne
rect 54633 49614 54710 49630
rect 54450 49515 54598 49597
rect 54338 49482 54415 49498
tri 54415 49482 54431 49498 sw
rect 54338 49416 54431 49482
rect 54338 49314 54431 49380
rect 54338 49298 54415 49314
tri 54415 49298 54431 49314 nw
rect 54467 49281 54581 49515
tri 54617 49482 54633 49498 se
rect 54633 49482 54710 49498
rect 54617 49416 54710 49482
rect 54617 49314 54710 49380
tri 54617 49298 54633 49314 ne
rect 54633 49298 54710 49314
rect 54450 49199 54598 49281
rect 54338 49166 54415 49182
tri 54415 49166 54431 49182 sw
rect 54338 49100 54431 49166
rect 54467 49041 54581 49199
tri 54617 49166 54633 49182 se
rect 54633 49166 54710 49182
rect 54617 49100 54710 49166
rect 54338 48965 54710 49041
rect 54338 48840 54431 48906
rect 54338 48824 54415 48840
tri 54415 48824 54431 48840 nw
rect 54467 48807 54581 48965
rect 54617 48840 54710 48906
tri 54617 48824 54633 48840 ne
rect 54633 48824 54710 48840
rect 54450 48725 54598 48807
rect 54338 48692 54415 48708
tri 54415 48692 54431 48708 sw
rect 54338 48626 54431 48692
rect 54338 48524 54431 48590
rect 54338 48508 54415 48524
tri 54415 48508 54431 48524 nw
rect 54467 48491 54581 48725
tri 54617 48692 54633 48708 se
rect 54633 48692 54710 48708
rect 54617 48626 54710 48692
rect 54617 48524 54710 48590
tri 54617 48508 54633 48524 ne
rect 54633 48508 54710 48524
rect 54450 48409 54598 48491
rect 54338 48376 54415 48392
tri 54415 48376 54431 48392 sw
rect 54338 48310 54431 48376
rect 54467 48251 54581 48409
tri 54617 48376 54633 48392 se
rect 54633 48376 54710 48392
rect 54617 48310 54710 48376
rect 54338 48175 54710 48251
rect 54338 48050 54431 48116
rect 54338 48034 54415 48050
tri 54415 48034 54431 48050 nw
rect 54467 48017 54581 48175
rect 54617 48050 54710 48116
tri 54617 48034 54633 48050 ne
rect 54633 48034 54710 48050
rect 54450 47935 54598 48017
rect 54338 47902 54415 47918
tri 54415 47902 54431 47918 sw
rect 54338 47836 54431 47902
rect 54338 47734 54431 47800
rect 54338 47718 54415 47734
tri 54415 47718 54431 47734 nw
rect 54467 47701 54581 47935
tri 54617 47902 54633 47918 se
rect 54633 47902 54710 47918
rect 54617 47836 54710 47902
rect 54617 47734 54710 47800
tri 54617 47718 54633 47734 ne
rect 54633 47718 54710 47734
rect 54450 47619 54598 47701
rect 54338 47586 54415 47602
tri 54415 47586 54431 47602 sw
rect 54338 47520 54431 47586
rect 54467 47461 54581 47619
tri 54617 47586 54633 47602 se
rect 54633 47586 54710 47602
rect 54617 47520 54710 47586
rect 54338 47385 54710 47461
rect 54338 47260 54431 47326
rect 54338 47244 54415 47260
tri 54415 47244 54431 47260 nw
rect 54467 47227 54581 47385
rect 54617 47260 54710 47326
tri 54617 47244 54633 47260 ne
rect 54633 47244 54710 47260
rect 54450 47145 54598 47227
rect 54338 47112 54415 47128
tri 54415 47112 54431 47128 sw
rect 54338 47046 54431 47112
rect 54338 46944 54431 47010
rect 54338 46928 54415 46944
tri 54415 46928 54431 46944 nw
rect 54467 46911 54581 47145
tri 54617 47112 54633 47128 se
rect 54633 47112 54710 47128
rect 54617 47046 54710 47112
rect 54617 46944 54710 47010
tri 54617 46928 54633 46944 ne
rect 54633 46928 54710 46944
rect 54450 46829 54598 46911
rect 54338 46796 54415 46812
tri 54415 46796 54431 46812 sw
rect 54338 46730 54431 46796
rect 54467 46671 54581 46829
tri 54617 46796 54633 46812 se
rect 54633 46796 54710 46812
rect 54617 46730 54710 46796
rect 54338 46595 54710 46671
rect 54338 46470 54431 46536
rect 54338 46454 54415 46470
tri 54415 46454 54431 46470 nw
rect 54467 46437 54581 46595
rect 54617 46470 54710 46536
tri 54617 46454 54633 46470 ne
rect 54633 46454 54710 46470
rect 54450 46355 54598 46437
rect 54338 46322 54415 46338
tri 54415 46322 54431 46338 sw
rect 54338 46256 54431 46322
rect 54338 46154 54431 46220
rect 54338 46138 54415 46154
tri 54415 46138 54431 46154 nw
rect 54467 46121 54581 46355
tri 54617 46322 54633 46338 se
rect 54633 46322 54710 46338
rect 54617 46256 54710 46322
rect 54617 46154 54710 46220
tri 54617 46138 54633 46154 ne
rect 54633 46138 54710 46154
rect 54450 46039 54598 46121
rect 54338 46006 54415 46022
tri 54415 46006 54431 46022 sw
rect 54338 45940 54431 46006
rect 54467 45881 54581 46039
tri 54617 46006 54633 46022 se
rect 54633 46006 54710 46022
rect 54617 45940 54710 46006
rect 54338 45805 54710 45881
rect 54338 45680 54431 45746
rect 54338 45664 54415 45680
tri 54415 45664 54431 45680 nw
rect 54467 45647 54581 45805
rect 54617 45680 54710 45746
tri 54617 45664 54633 45680 ne
rect 54633 45664 54710 45680
rect 54450 45565 54598 45647
rect 54338 45532 54415 45548
tri 54415 45532 54431 45548 sw
rect 54338 45466 54431 45532
rect 54338 45364 54431 45430
rect 54338 45348 54415 45364
tri 54415 45348 54431 45364 nw
rect 54467 45331 54581 45565
tri 54617 45532 54633 45548 se
rect 54633 45532 54710 45548
rect 54617 45466 54710 45532
rect 54617 45364 54710 45430
tri 54617 45348 54633 45364 ne
rect 54633 45348 54710 45364
rect 54450 45249 54598 45331
rect 54338 45216 54415 45232
tri 54415 45216 54431 45232 sw
rect 54338 45150 54431 45216
rect 54467 45091 54581 45249
tri 54617 45216 54633 45232 se
rect 54633 45216 54710 45232
rect 54617 45150 54710 45216
rect 54338 45015 54710 45091
rect 54338 44890 54431 44956
rect 54338 44874 54415 44890
tri 54415 44874 54431 44890 nw
rect 54467 44857 54581 45015
rect 54617 44890 54710 44956
tri 54617 44874 54633 44890 ne
rect 54633 44874 54710 44890
rect 54450 44775 54598 44857
rect 54338 44742 54415 44758
tri 54415 44742 54431 44758 sw
rect 54338 44676 54431 44742
rect 54338 44574 54431 44640
rect 54338 44558 54415 44574
tri 54415 44558 54431 44574 nw
rect 54467 44541 54581 44775
tri 54617 44742 54633 44758 se
rect 54633 44742 54710 44758
rect 54617 44676 54710 44742
rect 54617 44574 54710 44640
tri 54617 44558 54633 44574 ne
rect 54633 44558 54710 44574
rect 54450 44459 54598 44541
rect 54338 44426 54415 44442
tri 54415 44426 54431 44442 sw
rect 54338 44360 54431 44426
rect 54467 44301 54581 44459
tri 54617 44426 54633 44442 se
rect 54633 44426 54710 44442
rect 54617 44360 54710 44426
rect 54338 44225 54710 44301
rect 54338 44100 54431 44166
rect 54338 44084 54415 44100
tri 54415 44084 54431 44100 nw
rect 54467 44067 54581 44225
rect 54617 44100 54710 44166
tri 54617 44084 54633 44100 ne
rect 54633 44084 54710 44100
rect 54450 43985 54598 44067
rect 54338 43952 54415 43968
tri 54415 43952 54431 43968 sw
rect 54338 43886 54431 43952
rect 54338 43784 54431 43850
rect 54338 43768 54415 43784
tri 54415 43768 54431 43784 nw
rect 54467 43751 54581 43985
tri 54617 43952 54633 43968 se
rect 54633 43952 54710 43968
rect 54617 43886 54710 43952
rect 54617 43784 54710 43850
tri 54617 43768 54633 43784 ne
rect 54633 43768 54710 43784
rect 54450 43669 54598 43751
rect 54338 43636 54415 43652
tri 54415 43636 54431 43652 sw
rect 54338 43570 54431 43636
rect 54467 43511 54581 43669
tri 54617 43636 54633 43652 se
rect 54633 43636 54710 43652
rect 54617 43570 54710 43636
rect 54338 43435 54710 43511
rect 54338 43310 54431 43376
rect 54338 43294 54415 43310
tri 54415 43294 54431 43310 nw
rect 54467 43277 54581 43435
rect 54617 43310 54710 43376
tri 54617 43294 54633 43310 ne
rect 54633 43294 54710 43310
rect 54450 43195 54598 43277
rect 54338 43162 54415 43178
tri 54415 43162 54431 43178 sw
rect 54338 43096 54431 43162
rect 54338 42994 54431 43060
rect 54338 42978 54415 42994
tri 54415 42978 54431 42994 nw
rect 54467 42961 54581 43195
tri 54617 43162 54633 43178 se
rect 54633 43162 54710 43178
rect 54617 43096 54710 43162
rect 54617 42994 54710 43060
tri 54617 42978 54633 42994 ne
rect 54633 42978 54710 42994
rect 54450 42879 54598 42961
rect 54338 42846 54415 42862
tri 54415 42846 54431 42862 sw
rect 54338 42780 54431 42846
rect 54467 42721 54581 42879
tri 54617 42846 54633 42862 se
rect 54633 42846 54710 42862
rect 54617 42780 54710 42846
rect 54338 42645 54710 42721
rect 54338 42520 54431 42586
rect 54338 42504 54415 42520
tri 54415 42504 54431 42520 nw
rect 54467 42487 54581 42645
rect 54617 42520 54710 42586
tri 54617 42504 54633 42520 ne
rect 54633 42504 54710 42520
rect 54450 42405 54598 42487
rect 54338 42372 54415 42388
tri 54415 42372 54431 42388 sw
rect 54338 42306 54431 42372
rect 54338 42204 54431 42270
rect 54338 42188 54415 42204
tri 54415 42188 54431 42204 nw
rect 54467 42171 54581 42405
tri 54617 42372 54633 42388 se
rect 54633 42372 54710 42388
rect 54617 42306 54710 42372
rect 54617 42204 54710 42270
tri 54617 42188 54633 42204 ne
rect 54633 42188 54710 42204
rect 54450 42089 54598 42171
rect 54338 42056 54415 42072
tri 54415 42056 54431 42072 sw
rect 54338 41990 54431 42056
rect 54467 41931 54581 42089
tri 54617 42056 54633 42072 se
rect 54633 42056 54710 42072
rect 54617 41990 54710 42056
rect 54338 41855 54710 41931
rect 54338 41730 54431 41796
rect 54338 41714 54415 41730
tri 54415 41714 54431 41730 nw
rect 54467 41697 54581 41855
rect 54617 41730 54710 41796
tri 54617 41714 54633 41730 ne
rect 54633 41714 54710 41730
rect 54450 41615 54598 41697
rect 54338 41582 54415 41598
tri 54415 41582 54431 41598 sw
rect 54338 41516 54431 41582
rect 54338 41414 54431 41480
rect 54338 41398 54415 41414
tri 54415 41398 54431 41414 nw
rect 54467 41381 54581 41615
tri 54617 41582 54633 41598 se
rect 54633 41582 54710 41598
rect 54617 41516 54710 41582
rect 54617 41414 54710 41480
tri 54617 41398 54633 41414 ne
rect 54633 41398 54710 41414
rect 54450 41299 54598 41381
rect 54338 41266 54415 41282
tri 54415 41266 54431 41282 sw
rect 54338 41200 54431 41266
rect 54467 41141 54581 41299
tri 54617 41266 54633 41282 se
rect 54633 41266 54710 41282
rect 54617 41200 54710 41266
rect 54338 41065 54710 41141
rect 54338 40940 54431 41006
rect 54338 40924 54415 40940
tri 54415 40924 54431 40940 nw
rect 54467 40907 54581 41065
rect 54617 40940 54710 41006
tri 54617 40924 54633 40940 ne
rect 54633 40924 54710 40940
rect 54450 40825 54598 40907
rect 54338 40792 54415 40808
tri 54415 40792 54431 40808 sw
rect 54338 40726 54431 40792
rect 54338 40624 54431 40690
rect 54338 40608 54415 40624
tri 54415 40608 54431 40624 nw
rect 54467 40591 54581 40825
tri 54617 40792 54633 40808 se
rect 54633 40792 54710 40808
rect 54617 40726 54710 40792
rect 54617 40624 54710 40690
tri 54617 40608 54633 40624 ne
rect 54633 40608 54710 40624
rect 54450 40509 54598 40591
rect 54338 40476 54415 40492
tri 54415 40476 54431 40492 sw
rect 54338 40410 54431 40476
rect 54467 40351 54581 40509
tri 54617 40476 54633 40492 se
rect 54633 40476 54710 40492
rect 54617 40410 54710 40476
rect 54338 40275 54710 40351
rect 54338 40150 54431 40216
rect 54338 40134 54415 40150
tri 54415 40134 54431 40150 nw
rect 54467 40117 54581 40275
rect 54617 40150 54710 40216
tri 54617 40134 54633 40150 ne
rect 54633 40134 54710 40150
rect 54450 40035 54598 40117
rect 54338 40002 54415 40018
tri 54415 40002 54431 40018 sw
rect 54338 39936 54431 40002
rect 54338 39834 54431 39900
rect 54338 39818 54415 39834
tri 54415 39818 54431 39834 nw
rect 54467 39801 54581 40035
tri 54617 40002 54633 40018 se
rect 54633 40002 54710 40018
rect 54617 39936 54710 40002
rect 54617 39834 54710 39900
tri 54617 39818 54633 39834 ne
rect 54633 39818 54710 39834
rect 54450 39719 54598 39801
rect 54338 39686 54415 39702
tri 54415 39686 54431 39702 sw
rect 54338 39620 54431 39686
rect 54467 39561 54581 39719
tri 54617 39686 54633 39702 se
rect 54633 39686 54710 39702
rect 54617 39620 54710 39686
rect 54338 39485 54710 39561
rect 54338 39360 54431 39426
rect 54338 39344 54415 39360
tri 54415 39344 54431 39360 nw
rect 54467 39327 54581 39485
rect 54617 39360 54710 39426
tri 54617 39344 54633 39360 ne
rect 54633 39344 54710 39360
rect 54450 39245 54598 39327
rect 54338 39212 54415 39228
tri 54415 39212 54431 39228 sw
rect 54338 39146 54431 39212
rect 54338 39044 54431 39110
rect 54338 39028 54415 39044
tri 54415 39028 54431 39044 nw
rect 54467 39011 54581 39245
tri 54617 39212 54633 39228 se
rect 54633 39212 54710 39228
rect 54617 39146 54710 39212
rect 54617 39044 54710 39110
tri 54617 39028 54633 39044 ne
rect 54633 39028 54710 39044
rect 54450 38929 54598 39011
rect 54338 38896 54415 38912
tri 54415 38896 54431 38912 sw
rect 54338 38830 54431 38896
rect 54467 38771 54581 38929
tri 54617 38896 54633 38912 se
rect 54633 38896 54710 38912
rect 54617 38830 54710 38896
rect 54338 38695 54710 38771
rect 54338 38570 54431 38636
rect 54338 38554 54415 38570
tri 54415 38554 54431 38570 nw
rect 54467 38537 54581 38695
rect 54617 38570 54710 38636
tri 54617 38554 54633 38570 ne
rect 54633 38554 54710 38570
rect 54450 38455 54598 38537
rect 54338 38422 54415 38438
tri 54415 38422 54431 38438 sw
rect 54338 38356 54431 38422
rect 54338 38254 54431 38320
rect 54338 38238 54415 38254
tri 54415 38238 54431 38254 nw
rect 54467 38221 54581 38455
tri 54617 38422 54633 38438 se
rect 54633 38422 54710 38438
rect 54617 38356 54710 38422
rect 54617 38254 54710 38320
tri 54617 38238 54633 38254 ne
rect 54633 38238 54710 38254
rect 54450 38139 54598 38221
rect 54338 38106 54415 38122
tri 54415 38106 54431 38122 sw
rect 54338 38040 54431 38106
rect 54467 37981 54581 38139
tri 54617 38106 54633 38122 se
rect 54633 38106 54710 38122
rect 54617 38040 54710 38106
rect 54338 37905 54710 37981
rect 54338 37780 54431 37846
rect 54338 37764 54415 37780
tri 54415 37764 54431 37780 nw
rect 54467 37747 54581 37905
rect 54617 37780 54710 37846
tri 54617 37764 54633 37780 ne
rect 54633 37764 54710 37780
rect 54450 37665 54598 37747
rect 54338 37632 54415 37648
tri 54415 37632 54431 37648 sw
rect 54338 37566 54431 37632
rect 54338 37464 54431 37530
rect 54338 37448 54415 37464
tri 54415 37448 54431 37464 nw
rect 54467 37431 54581 37665
tri 54617 37632 54633 37648 se
rect 54633 37632 54710 37648
rect 54617 37566 54710 37632
rect 54617 37464 54710 37530
tri 54617 37448 54633 37464 ne
rect 54633 37448 54710 37464
rect 54450 37349 54598 37431
rect 54338 37316 54415 37332
tri 54415 37316 54431 37332 sw
rect 54338 37250 54431 37316
rect 54467 37191 54581 37349
tri 54617 37316 54633 37332 se
rect 54633 37316 54710 37332
rect 54617 37250 54710 37316
rect 54338 37115 54710 37191
rect 54338 36990 54431 37056
rect 54338 36974 54415 36990
tri 54415 36974 54431 36990 nw
rect 54467 36957 54581 37115
rect 54617 36990 54710 37056
tri 54617 36974 54633 36990 ne
rect 54633 36974 54710 36990
rect 54450 36875 54598 36957
rect 54338 36842 54415 36858
tri 54415 36842 54431 36858 sw
rect 54338 36776 54431 36842
rect 54338 36674 54431 36740
rect 54338 36658 54415 36674
tri 54415 36658 54431 36674 nw
rect 54467 36641 54581 36875
tri 54617 36842 54633 36858 se
rect 54633 36842 54710 36858
rect 54617 36776 54710 36842
rect 54617 36674 54710 36740
tri 54617 36658 54633 36674 ne
rect 54633 36658 54710 36674
rect 54450 36559 54598 36641
rect 54338 36526 54415 36542
tri 54415 36526 54431 36542 sw
rect 54338 36460 54431 36526
rect 54467 36401 54581 36559
tri 54617 36526 54633 36542 se
rect 54633 36526 54710 36542
rect 54617 36460 54710 36526
rect 54338 36325 54710 36401
rect 54338 36200 54431 36266
rect 54338 36184 54415 36200
tri 54415 36184 54431 36200 nw
rect 54467 36167 54581 36325
rect 54617 36200 54710 36266
tri 54617 36184 54633 36200 ne
rect 54633 36184 54710 36200
rect 54450 36085 54598 36167
rect 54338 36052 54415 36068
tri 54415 36052 54431 36068 sw
rect 54338 35986 54431 36052
rect 54338 35884 54431 35950
rect 54338 35868 54415 35884
tri 54415 35868 54431 35884 nw
rect 54467 35851 54581 36085
tri 54617 36052 54633 36068 se
rect 54633 36052 54710 36068
rect 54617 35986 54710 36052
rect 54617 35884 54710 35950
tri 54617 35868 54633 35884 ne
rect 54633 35868 54710 35884
rect 54450 35769 54598 35851
rect 54338 35736 54415 35752
tri 54415 35736 54431 35752 sw
rect 54338 35670 54431 35736
rect 54467 35611 54581 35769
tri 54617 35736 54633 35752 se
rect 54633 35736 54710 35752
rect 54617 35670 54710 35736
rect 54338 35535 54710 35611
rect 54338 35410 54431 35476
rect 54338 35394 54415 35410
tri 54415 35394 54431 35410 nw
rect 54467 35377 54581 35535
rect 54617 35410 54710 35476
tri 54617 35394 54633 35410 ne
rect 54633 35394 54710 35410
rect 54450 35295 54598 35377
rect 54338 35262 54415 35278
tri 54415 35262 54431 35278 sw
rect 54338 35196 54431 35262
rect 54338 35094 54431 35160
rect 54338 35078 54415 35094
tri 54415 35078 54431 35094 nw
rect 54467 35061 54581 35295
tri 54617 35262 54633 35278 se
rect 54633 35262 54710 35278
rect 54617 35196 54710 35262
rect 54617 35094 54710 35160
tri 54617 35078 54633 35094 ne
rect 54633 35078 54710 35094
rect 54450 34979 54598 35061
rect 54338 34946 54415 34962
tri 54415 34946 54431 34962 sw
rect 54338 34880 54431 34946
rect 54467 34821 54581 34979
tri 54617 34946 54633 34962 se
rect 54633 34946 54710 34962
rect 54617 34880 54710 34946
rect 54338 34745 54710 34821
rect 54338 34620 54431 34686
rect 54338 34604 54415 34620
tri 54415 34604 54431 34620 nw
rect 54467 34587 54581 34745
rect 54617 34620 54710 34686
tri 54617 34604 54633 34620 ne
rect 54633 34604 54710 34620
rect 54450 34505 54598 34587
rect 54338 34472 54415 34488
tri 54415 34472 54431 34488 sw
rect 54338 34406 54431 34472
rect 54338 34304 54431 34370
rect 54338 34288 54415 34304
tri 54415 34288 54431 34304 nw
rect 54467 34271 54581 34505
tri 54617 34472 54633 34488 se
rect 54633 34472 54710 34488
rect 54617 34406 54710 34472
rect 54617 34304 54710 34370
tri 54617 34288 54633 34304 ne
rect 54633 34288 54710 34304
rect 54450 34189 54598 34271
rect 54338 34156 54415 34172
tri 54415 34156 54431 34172 sw
rect 54338 34090 54431 34156
rect 54467 34031 54581 34189
tri 54617 34156 54633 34172 se
rect 54633 34156 54710 34172
rect 54617 34090 54710 34156
rect 54338 33955 54710 34031
rect 54338 33830 54431 33896
rect 54338 33814 54415 33830
tri 54415 33814 54431 33830 nw
rect 54467 33797 54581 33955
rect 54617 33830 54710 33896
tri 54617 33814 54633 33830 ne
rect 54633 33814 54710 33830
rect 54450 33715 54598 33797
rect 54338 33682 54415 33698
tri 54415 33682 54431 33698 sw
rect 54338 33616 54431 33682
rect 54338 33514 54431 33580
rect 54338 33498 54415 33514
tri 54415 33498 54431 33514 nw
rect 54467 33481 54581 33715
tri 54617 33682 54633 33698 se
rect 54633 33682 54710 33698
rect 54617 33616 54710 33682
rect 54617 33514 54710 33580
tri 54617 33498 54633 33514 ne
rect 54633 33498 54710 33514
rect 54450 33399 54598 33481
rect 54338 33366 54415 33382
tri 54415 33366 54431 33382 sw
rect 54338 33300 54431 33366
rect 54467 33241 54581 33399
tri 54617 33366 54633 33382 se
rect 54633 33366 54710 33382
rect 54617 33300 54710 33366
rect 54338 33165 54710 33241
rect 54338 33040 54431 33106
rect 54338 33024 54415 33040
tri 54415 33024 54431 33040 nw
rect 54467 33007 54581 33165
rect 54617 33040 54710 33106
tri 54617 33024 54633 33040 ne
rect 54633 33024 54710 33040
rect 54450 32925 54598 33007
rect 54338 32892 54415 32908
tri 54415 32892 54431 32908 sw
rect 54338 32826 54431 32892
rect 54338 32724 54431 32790
rect 54338 32708 54415 32724
tri 54415 32708 54431 32724 nw
rect 54467 32691 54581 32925
tri 54617 32892 54633 32908 se
rect 54633 32892 54710 32908
rect 54617 32826 54710 32892
rect 54617 32724 54710 32790
tri 54617 32708 54633 32724 ne
rect 54633 32708 54710 32724
rect 54450 32609 54598 32691
rect 54338 32576 54415 32592
tri 54415 32576 54431 32592 sw
rect 54338 32510 54431 32576
rect 54467 32451 54581 32609
tri 54617 32576 54633 32592 se
rect 54633 32576 54710 32592
rect 54617 32510 54710 32576
rect 54338 32375 54710 32451
rect 54338 32250 54431 32316
rect 54338 32234 54415 32250
tri 54415 32234 54431 32250 nw
rect 54467 32217 54581 32375
rect 54617 32250 54710 32316
tri 54617 32234 54633 32250 ne
rect 54633 32234 54710 32250
rect 54450 32135 54598 32217
rect 54338 32102 54415 32118
tri 54415 32102 54431 32118 sw
rect 54338 32036 54431 32102
rect 54338 31934 54431 32000
rect 54338 31918 54415 31934
tri 54415 31918 54431 31934 nw
rect 54467 31901 54581 32135
tri 54617 32102 54633 32118 se
rect 54633 32102 54710 32118
rect 54617 32036 54710 32102
rect 54617 31934 54710 32000
tri 54617 31918 54633 31934 ne
rect 54633 31918 54710 31934
rect 54450 31819 54598 31901
rect 54338 31786 54415 31802
tri 54415 31786 54431 31802 sw
rect 54338 31720 54431 31786
rect 54467 31661 54581 31819
tri 54617 31786 54633 31802 se
rect 54633 31786 54710 31802
rect 54617 31720 54710 31786
rect 54338 31585 54710 31661
rect 54338 31460 54431 31526
rect 54338 31444 54415 31460
tri 54415 31444 54431 31460 nw
rect 54467 31427 54581 31585
rect 54617 31460 54710 31526
tri 54617 31444 54633 31460 ne
rect 54633 31444 54710 31460
rect 54450 31345 54598 31427
rect 54338 31312 54415 31328
tri 54415 31312 54431 31328 sw
rect 54338 31246 54431 31312
rect 54338 31144 54431 31210
rect 54338 31128 54415 31144
tri 54415 31128 54431 31144 nw
rect 54467 31111 54581 31345
tri 54617 31312 54633 31328 se
rect 54633 31312 54710 31328
rect 54617 31246 54710 31312
rect 54617 31144 54710 31210
tri 54617 31128 54633 31144 ne
rect 54633 31128 54710 31144
rect 54450 31029 54598 31111
rect 54338 30996 54415 31012
tri 54415 30996 54431 31012 sw
rect 54338 30930 54431 30996
rect 54467 30871 54581 31029
tri 54617 30996 54633 31012 se
rect 54633 30996 54710 31012
rect 54617 30930 54710 30996
rect 54338 30795 54710 30871
rect 54338 30670 54431 30736
rect 54338 30654 54415 30670
tri 54415 30654 54431 30670 nw
rect 54467 30637 54581 30795
rect 54617 30670 54710 30736
tri 54617 30654 54633 30670 ne
rect 54633 30654 54710 30670
rect 54450 30555 54598 30637
rect 54338 30522 54415 30538
tri 54415 30522 54431 30538 sw
rect 54338 30456 54431 30522
rect 54338 30354 54431 30420
rect 54338 30338 54415 30354
tri 54415 30338 54431 30354 nw
rect 54467 30321 54581 30555
tri 54617 30522 54633 30538 se
rect 54633 30522 54710 30538
rect 54617 30456 54710 30522
rect 54617 30354 54710 30420
tri 54617 30338 54633 30354 ne
rect 54633 30338 54710 30354
rect 54450 30239 54598 30321
rect 54338 30206 54415 30222
tri 54415 30206 54431 30222 sw
rect 54338 30140 54431 30206
rect 54467 30081 54581 30239
tri 54617 30206 54633 30222 se
rect 54633 30206 54710 30222
rect 54617 30140 54710 30206
rect 54338 30005 54710 30081
rect 54338 29880 54431 29946
rect 54338 29864 54415 29880
tri 54415 29864 54431 29880 nw
rect 54467 29847 54581 30005
rect 54617 29880 54710 29946
tri 54617 29864 54633 29880 ne
rect 54633 29864 54710 29880
rect 54450 29765 54598 29847
rect 54338 29732 54415 29748
tri 54415 29732 54431 29748 sw
rect 54338 29666 54431 29732
rect 54338 29564 54431 29630
rect 54338 29548 54415 29564
tri 54415 29548 54431 29564 nw
rect 54467 29531 54581 29765
tri 54617 29732 54633 29748 se
rect 54633 29732 54710 29748
rect 54617 29666 54710 29732
rect 54617 29564 54710 29630
tri 54617 29548 54633 29564 ne
rect 54633 29548 54710 29564
rect 54450 29449 54598 29531
rect 54338 29416 54415 29432
tri 54415 29416 54431 29432 sw
rect 54338 29350 54431 29416
rect 54467 29291 54581 29449
tri 54617 29416 54633 29432 se
rect 54633 29416 54710 29432
rect 54617 29350 54710 29416
rect 54338 29215 54710 29291
rect 54338 29090 54431 29156
rect 54338 29074 54415 29090
tri 54415 29074 54431 29090 nw
rect 54467 29057 54581 29215
rect 54617 29090 54710 29156
tri 54617 29074 54633 29090 ne
rect 54633 29074 54710 29090
rect 54450 28975 54598 29057
rect 54338 28942 54415 28958
tri 54415 28942 54431 28958 sw
rect 54338 28876 54431 28942
rect 54467 28833 54581 28975
tri 54617 28942 54633 28958 se
rect 54633 28942 54710 28958
rect 54617 28876 54710 28942
rect 54746 28463 54782 80603
rect 54818 28463 54854 80603
rect 54890 80445 54926 80603
rect 54882 80303 54934 80445
rect 54890 28763 54926 80303
rect 54882 28621 54934 28763
rect 54890 28463 54926 28621
rect 54962 28463 54998 80603
rect 55034 28463 55070 80603
rect 55106 28833 55190 80233
rect 55226 28463 55262 80603
rect 55298 28463 55334 80603
rect 55370 80445 55406 80603
rect 55362 80303 55414 80445
rect 55370 28763 55406 80303
rect 55362 28621 55414 28763
rect 55370 28463 55406 28621
rect 55442 28463 55478 80603
rect 55514 28463 55550 80603
rect 55586 80124 55679 80190
rect 55586 80108 55663 80124
tri 55663 80108 55679 80124 nw
rect 55715 80091 55829 80233
rect 55865 80124 55958 80190
tri 55865 80108 55881 80124 ne
rect 55881 80108 55958 80124
rect 55698 80009 55846 80091
rect 55586 79976 55663 79992
tri 55663 79976 55679 79992 sw
rect 55586 79910 55679 79976
rect 55715 79851 55829 80009
tri 55865 79976 55881 79992 se
rect 55881 79976 55958 79992
rect 55865 79910 55958 79976
rect 55586 79775 55958 79851
rect 55586 79650 55679 79716
rect 55586 79634 55663 79650
tri 55663 79634 55679 79650 nw
rect 55715 79617 55829 79775
rect 55865 79650 55958 79716
tri 55865 79634 55881 79650 ne
rect 55881 79634 55958 79650
rect 55698 79535 55846 79617
rect 55586 79502 55663 79518
tri 55663 79502 55679 79518 sw
rect 55586 79436 55679 79502
rect 55586 79334 55679 79400
rect 55586 79318 55663 79334
tri 55663 79318 55679 79334 nw
rect 55715 79301 55829 79535
tri 55865 79502 55881 79518 se
rect 55881 79502 55958 79518
rect 55865 79436 55958 79502
rect 55865 79334 55958 79400
tri 55865 79318 55881 79334 ne
rect 55881 79318 55958 79334
rect 55698 79219 55846 79301
rect 55586 79186 55663 79202
tri 55663 79186 55679 79202 sw
rect 55586 79120 55679 79186
rect 55715 79061 55829 79219
tri 55865 79186 55881 79202 se
rect 55881 79186 55958 79202
rect 55865 79120 55958 79186
rect 55586 78985 55958 79061
rect 55586 78860 55679 78926
rect 55586 78844 55663 78860
tri 55663 78844 55679 78860 nw
rect 55715 78827 55829 78985
rect 55865 78860 55958 78926
tri 55865 78844 55881 78860 ne
rect 55881 78844 55958 78860
rect 55698 78745 55846 78827
rect 55586 78712 55663 78728
tri 55663 78712 55679 78728 sw
rect 55586 78646 55679 78712
rect 55586 78544 55679 78610
rect 55586 78528 55663 78544
tri 55663 78528 55679 78544 nw
rect 55715 78511 55829 78745
tri 55865 78712 55881 78728 se
rect 55881 78712 55958 78728
rect 55865 78646 55958 78712
rect 55865 78544 55958 78610
tri 55865 78528 55881 78544 ne
rect 55881 78528 55958 78544
rect 55698 78429 55846 78511
rect 55586 78396 55663 78412
tri 55663 78396 55679 78412 sw
rect 55586 78330 55679 78396
rect 55715 78271 55829 78429
tri 55865 78396 55881 78412 se
rect 55881 78396 55958 78412
rect 55865 78330 55958 78396
rect 55586 78195 55958 78271
rect 55586 78070 55679 78136
rect 55586 78054 55663 78070
tri 55663 78054 55679 78070 nw
rect 55715 78037 55829 78195
rect 55865 78070 55958 78136
tri 55865 78054 55881 78070 ne
rect 55881 78054 55958 78070
rect 55698 77955 55846 78037
rect 55586 77922 55663 77938
tri 55663 77922 55679 77938 sw
rect 55586 77856 55679 77922
rect 55586 77754 55679 77820
rect 55586 77738 55663 77754
tri 55663 77738 55679 77754 nw
rect 55715 77721 55829 77955
tri 55865 77922 55881 77938 se
rect 55881 77922 55958 77938
rect 55865 77856 55958 77922
rect 55865 77754 55958 77820
tri 55865 77738 55881 77754 ne
rect 55881 77738 55958 77754
rect 55698 77639 55846 77721
rect 55586 77606 55663 77622
tri 55663 77606 55679 77622 sw
rect 55586 77540 55679 77606
rect 55715 77481 55829 77639
tri 55865 77606 55881 77622 se
rect 55881 77606 55958 77622
rect 55865 77540 55958 77606
rect 55586 77405 55958 77481
rect 55586 77280 55679 77346
rect 55586 77264 55663 77280
tri 55663 77264 55679 77280 nw
rect 55715 77247 55829 77405
rect 55865 77280 55958 77346
tri 55865 77264 55881 77280 ne
rect 55881 77264 55958 77280
rect 55698 77165 55846 77247
rect 55586 77132 55663 77148
tri 55663 77132 55679 77148 sw
rect 55586 77066 55679 77132
rect 55586 76964 55679 77030
rect 55586 76948 55663 76964
tri 55663 76948 55679 76964 nw
rect 55715 76931 55829 77165
tri 55865 77132 55881 77148 se
rect 55881 77132 55958 77148
rect 55865 77066 55958 77132
rect 55865 76964 55958 77030
tri 55865 76948 55881 76964 ne
rect 55881 76948 55958 76964
rect 55698 76849 55846 76931
rect 55586 76816 55663 76832
tri 55663 76816 55679 76832 sw
rect 55586 76750 55679 76816
rect 55715 76691 55829 76849
tri 55865 76816 55881 76832 se
rect 55881 76816 55958 76832
rect 55865 76750 55958 76816
rect 55586 76615 55958 76691
rect 55586 76490 55679 76556
rect 55586 76474 55663 76490
tri 55663 76474 55679 76490 nw
rect 55715 76457 55829 76615
rect 55865 76490 55958 76556
tri 55865 76474 55881 76490 ne
rect 55881 76474 55958 76490
rect 55698 76375 55846 76457
rect 55586 76342 55663 76358
tri 55663 76342 55679 76358 sw
rect 55586 76276 55679 76342
rect 55586 76174 55679 76240
rect 55586 76158 55663 76174
tri 55663 76158 55679 76174 nw
rect 55715 76141 55829 76375
tri 55865 76342 55881 76358 se
rect 55881 76342 55958 76358
rect 55865 76276 55958 76342
rect 55865 76174 55958 76240
tri 55865 76158 55881 76174 ne
rect 55881 76158 55958 76174
rect 55698 76059 55846 76141
rect 55586 76026 55663 76042
tri 55663 76026 55679 76042 sw
rect 55586 75960 55679 76026
rect 55715 75901 55829 76059
tri 55865 76026 55881 76042 se
rect 55881 76026 55958 76042
rect 55865 75960 55958 76026
rect 55586 75825 55958 75901
rect 55586 75700 55679 75766
rect 55586 75684 55663 75700
tri 55663 75684 55679 75700 nw
rect 55715 75667 55829 75825
rect 55865 75700 55958 75766
tri 55865 75684 55881 75700 ne
rect 55881 75684 55958 75700
rect 55698 75585 55846 75667
rect 55586 75552 55663 75568
tri 55663 75552 55679 75568 sw
rect 55586 75486 55679 75552
rect 55586 75384 55679 75450
rect 55586 75368 55663 75384
tri 55663 75368 55679 75384 nw
rect 55715 75351 55829 75585
tri 55865 75552 55881 75568 se
rect 55881 75552 55958 75568
rect 55865 75486 55958 75552
rect 55865 75384 55958 75450
tri 55865 75368 55881 75384 ne
rect 55881 75368 55958 75384
rect 55698 75269 55846 75351
rect 55586 75236 55663 75252
tri 55663 75236 55679 75252 sw
rect 55586 75170 55679 75236
rect 55715 75111 55829 75269
tri 55865 75236 55881 75252 se
rect 55881 75236 55958 75252
rect 55865 75170 55958 75236
rect 55586 75035 55958 75111
rect 55586 74910 55679 74976
rect 55586 74894 55663 74910
tri 55663 74894 55679 74910 nw
rect 55715 74877 55829 75035
rect 55865 74910 55958 74976
tri 55865 74894 55881 74910 ne
rect 55881 74894 55958 74910
rect 55698 74795 55846 74877
rect 55586 74762 55663 74778
tri 55663 74762 55679 74778 sw
rect 55586 74696 55679 74762
rect 55586 74594 55679 74660
rect 55586 74578 55663 74594
tri 55663 74578 55679 74594 nw
rect 55715 74561 55829 74795
tri 55865 74762 55881 74778 se
rect 55881 74762 55958 74778
rect 55865 74696 55958 74762
rect 55865 74594 55958 74660
tri 55865 74578 55881 74594 ne
rect 55881 74578 55958 74594
rect 55698 74479 55846 74561
rect 55586 74446 55663 74462
tri 55663 74446 55679 74462 sw
rect 55586 74380 55679 74446
rect 55715 74321 55829 74479
tri 55865 74446 55881 74462 se
rect 55881 74446 55958 74462
rect 55865 74380 55958 74446
rect 55586 74245 55958 74321
rect 55586 74120 55679 74186
rect 55586 74104 55663 74120
tri 55663 74104 55679 74120 nw
rect 55715 74087 55829 74245
rect 55865 74120 55958 74186
tri 55865 74104 55881 74120 ne
rect 55881 74104 55958 74120
rect 55698 74005 55846 74087
rect 55586 73972 55663 73988
tri 55663 73972 55679 73988 sw
rect 55586 73906 55679 73972
rect 55586 73804 55679 73870
rect 55586 73788 55663 73804
tri 55663 73788 55679 73804 nw
rect 55715 73771 55829 74005
tri 55865 73972 55881 73988 se
rect 55881 73972 55958 73988
rect 55865 73906 55958 73972
rect 55865 73804 55958 73870
tri 55865 73788 55881 73804 ne
rect 55881 73788 55958 73804
rect 55698 73689 55846 73771
rect 55586 73656 55663 73672
tri 55663 73656 55679 73672 sw
rect 55586 73590 55679 73656
rect 55715 73531 55829 73689
tri 55865 73656 55881 73672 se
rect 55881 73656 55958 73672
rect 55865 73590 55958 73656
rect 55586 73455 55958 73531
rect 55586 73330 55679 73396
rect 55586 73314 55663 73330
tri 55663 73314 55679 73330 nw
rect 55715 73297 55829 73455
rect 55865 73330 55958 73396
tri 55865 73314 55881 73330 ne
rect 55881 73314 55958 73330
rect 55698 73215 55846 73297
rect 55586 73182 55663 73198
tri 55663 73182 55679 73198 sw
rect 55586 73116 55679 73182
rect 55586 73014 55679 73080
rect 55586 72998 55663 73014
tri 55663 72998 55679 73014 nw
rect 55715 72981 55829 73215
tri 55865 73182 55881 73198 se
rect 55881 73182 55958 73198
rect 55865 73116 55958 73182
rect 55865 73014 55958 73080
tri 55865 72998 55881 73014 ne
rect 55881 72998 55958 73014
rect 55698 72899 55846 72981
rect 55586 72866 55663 72882
tri 55663 72866 55679 72882 sw
rect 55586 72800 55679 72866
rect 55715 72741 55829 72899
tri 55865 72866 55881 72882 se
rect 55881 72866 55958 72882
rect 55865 72800 55958 72866
rect 55586 72665 55958 72741
rect 55586 72540 55679 72606
rect 55586 72524 55663 72540
tri 55663 72524 55679 72540 nw
rect 55715 72507 55829 72665
rect 55865 72540 55958 72606
tri 55865 72524 55881 72540 ne
rect 55881 72524 55958 72540
rect 55698 72425 55846 72507
rect 55586 72392 55663 72408
tri 55663 72392 55679 72408 sw
rect 55586 72326 55679 72392
rect 55586 72224 55679 72290
rect 55586 72208 55663 72224
tri 55663 72208 55679 72224 nw
rect 55715 72191 55829 72425
tri 55865 72392 55881 72408 se
rect 55881 72392 55958 72408
rect 55865 72326 55958 72392
rect 55865 72224 55958 72290
tri 55865 72208 55881 72224 ne
rect 55881 72208 55958 72224
rect 55698 72109 55846 72191
rect 55586 72076 55663 72092
tri 55663 72076 55679 72092 sw
rect 55586 72010 55679 72076
rect 55715 71951 55829 72109
tri 55865 72076 55881 72092 se
rect 55881 72076 55958 72092
rect 55865 72010 55958 72076
rect 55586 71875 55958 71951
rect 55586 71750 55679 71816
rect 55586 71734 55663 71750
tri 55663 71734 55679 71750 nw
rect 55715 71717 55829 71875
rect 55865 71750 55958 71816
tri 55865 71734 55881 71750 ne
rect 55881 71734 55958 71750
rect 55698 71635 55846 71717
rect 55586 71602 55663 71618
tri 55663 71602 55679 71618 sw
rect 55586 71536 55679 71602
rect 55586 71434 55679 71500
rect 55586 71418 55663 71434
tri 55663 71418 55679 71434 nw
rect 55715 71401 55829 71635
tri 55865 71602 55881 71618 se
rect 55881 71602 55958 71618
rect 55865 71536 55958 71602
rect 55865 71434 55958 71500
tri 55865 71418 55881 71434 ne
rect 55881 71418 55958 71434
rect 55698 71319 55846 71401
rect 55586 71286 55663 71302
tri 55663 71286 55679 71302 sw
rect 55586 71220 55679 71286
rect 55715 71161 55829 71319
tri 55865 71286 55881 71302 se
rect 55881 71286 55958 71302
rect 55865 71220 55958 71286
rect 55586 71085 55958 71161
rect 55586 70960 55679 71026
rect 55586 70944 55663 70960
tri 55663 70944 55679 70960 nw
rect 55715 70927 55829 71085
rect 55865 70960 55958 71026
tri 55865 70944 55881 70960 ne
rect 55881 70944 55958 70960
rect 55698 70845 55846 70927
rect 55586 70812 55663 70828
tri 55663 70812 55679 70828 sw
rect 55586 70746 55679 70812
rect 55586 70644 55679 70710
rect 55586 70628 55663 70644
tri 55663 70628 55679 70644 nw
rect 55715 70611 55829 70845
tri 55865 70812 55881 70828 se
rect 55881 70812 55958 70828
rect 55865 70746 55958 70812
rect 55865 70644 55958 70710
tri 55865 70628 55881 70644 ne
rect 55881 70628 55958 70644
rect 55698 70529 55846 70611
rect 55586 70496 55663 70512
tri 55663 70496 55679 70512 sw
rect 55586 70430 55679 70496
rect 55715 70371 55829 70529
tri 55865 70496 55881 70512 se
rect 55881 70496 55958 70512
rect 55865 70430 55958 70496
rect 55586 70295 55958 70371
rect 55586 70170 55679 70236
rect 55586 70154 55663 70170
tri 55663 70154 55679 70170 nw
rect 55715 70137 55829 70295
rect 55865 70170 55958 70236
tri 55865 70154 55881 70170 ne
rect 55881 70154 55958 70170
rect 55698 70055 55846 70137
rect 55586 70022 55663 70038
tri 55663 70022 55679 70038 sw
rect 55586 69956 55679 70022
rect 55586 69854 55679 69920
rect 55586 69838 55663 69854
tri 55663 69838 55679 69854 nw
rect 55715 69821 55829 70055
tri 55865 70022 55881 70038 se
rect 55881 70022 55958 70038
rect 55865 69956 55958 70022
rect 55865 69854 55958 69920
tri 55865 69838 55881 69854 ne
rect 55881 69838 55958 69854
rect 55698 69739 55846 69821
rect 55586 69706 55663 69722
tri 55663 69706 55679 69722 sw
rect 55586 69640 55679 69706
rect 55715 69581 55829 69739
tri 55865 69706 55881 69722 se
rect 55881 69706 55958 69722
rect 55865 69640 55958 69706
rect 55586 69505 55958 69581
rect 55586 69380 55679 69446
rect 55586 69364 55663 69380
tri 55663 69364 55679 69380 nw
rect 55715 69347 55829 69505
rect 55865 69380 55958 69446
tri 55865 69364 55881 69380 ne
rect 55881 69364 55958 69380
rect 55698 69265 55846 69347
rect 55586 69232 55663 69248
tri 55663 69232 55679 69248 sw
rect 55586 69166 55679 69232
rect 55586 69064 55679 69130
rect 55586 69048 55663 69064
tri 55663 69048 55679 69064 nw
rect 55715 69031 55829 69265
tri 55865 69232 55881 69248 se
rect 55881 69232 55958 69248
rect 55865 69166 55958 69232
rect 55865 69064 55958 69130
tri 55865 69048 55881 69064 ne
rect 55881 69048 55958 69064
rect 55698 68949 55846 69031
rect 55586 68916 55663 68932
tri 55663 68916 55679 68932 sw
rect 55586 68850 55679 68916
rect 55715 68791 55829 68949
tri 55865 68916 55881 68932 se
rect 55881 68916 55958 68932
rect 55865 68850 55958 68916
rect 55586 68715 55958 68791
rect 55586 68590 55679 68656
rect 55586 68574 55663 68590
tri 55663 68574 55679 68590 nw
rect 55715 68557 55829 68715
rect 55865 68590 55958 68656
tri 55865 68574 55881 68590 ne
rect 55881 68574 55958 68590
rect 55698 68475 55846 68557
rect 55586 68442 55663 68458
tri 55663 68442 55679 68458 sw
rect 55586 68376 55679 68442
rect 55586 68274 55679 68340
rect 55586 68258 55663 68274
tri 55663 68258 55679 68274 nw
rect 55715 68241 55829 68475
tri 55865 68442 55881 68458 se
rect 55881 68442 55958 68458
rect 55865 68376 55958 68442
rect 55865 68274 55958 68340
tri 55865 68258 55881 68274 ne
rect 55881 68258 55958 68274
rect 55698 68159 55846 68241
rect 55586 68126 55663 68142
tri 55663 68126 55679 68142 sw
rect 55586 68060 55679 68126
rect 55715 68001 55829 68159
tri 55865 68126 55881 68142 se
rect 55881 68126 55958 68142
rect 55865 68060 55958 68126
rect 55586 67925 55958 68001
rect 55586 67800 55679 67866
rect 55586 67784 55663 67800
tri 55663 67784 55679 67800 nw
rect 55715 67767 55829 67925
rect 55865 67800 55958 67866
tri 55865 67784 55881 67800 ne
rect 55881 67784 55958 67800
rect 55698 67685 55846 67767
rect 55586 67652 55663 67668
tri 55663 67652 55679 67668 sw
rect 55586 67586 55679 67652
rect 55586 67484 55679 67550
rect 55586 67468 55663 67484
tri 55663 67468 55679 67484 nw
rect 55715 67451 55829 67685
tri 55865 67652 55881 67668 se
rect 55881 67652 55958 67668
rect 55865 67586 55958 67652
rect 55865 67484 55958 67550
tri 55865 67468 55881 67484 ne
rect 55881 67468 55958 67484
rect 55698 67369 55846 67451
rect 55586 67336 55663 67352
tri 55663 67336 55679 67352 sw
rect 55586 67270 55679 67336
rect 55715 67211 55829 67369
tri 55865 67336 55881 67352 se
rect 55881 67336 55958 67352
rect 55865 67270 55958 67336
rect 55586 67135 55958 67211
rect 55586 67010 55679 67076
rect 55586 66994 55663 67010
tri 55663 66994 55679 67010 nw
rect 55715 66977 55829 67135
rect 55865 67010 55958 67076
tri 55865 66994 55881 67010 ne
rect 55881 66994 55958 67010
rect 55698 66895 55846 66977
rect 55586 66862 55663 66878
tri 55663 66862 55679 66878 sw
rect 55586 66796 55679 66862
rect 55586 66694 55679 66760
rect 55586 66678 55663 66694
tri 55663 66678 55679 66694 nw
rect 55715 66661 55829 66895
tri 55865 66862 55881 66878 se
rect 55881 66862 55958 66878
rect 55865 66796 55958 66862
rect 55865 66694 55958 66760
tri 55865 66678 55881 66694 ne
rect 55881 66678 55958 66694
rect 55698 66579 55846 66661
rect 55586 66546 55663 66562
tri 55663 66546 55679 66562 sw
rect 55586 66480 55679 66546
rect 55715 66421 55829 66579
tri 55865 66546 55881 66562 se
rect 55881 66546 55958 66562
rect 55865 66480 55958 66546
rect 55586 66345 55958 66421
rect 55586 66220 55679 66286
rect 55586 66204 55663 66220
tri 55663 66204 55679 66220 nw
rect 55715 66187 55829 66345
rect 55865 66220 55958 66286
tri 55865 66204 55881 66220 ne
rect 55881 66204 55958 66220
rect 55698 66105 55846 66187
rect 55586 66072 55663 66088
tri 55663 66072 55679 66088 sw
rect 55586 66006 55679 66072
rect 55586 65904 55679 65970
rect 55586 65888 55663 65904
tri 55663 65888 55679 65904 nw
rect 55715 65871 55829 66105
tri 55865 66072 55881 66088 se
rect 55881 66072 55958 66088
rect 55865 66006 55958 66072
rect 55865 65904 55958 65970
tri 55865 65888 55881 65904 ne
rect 55881 65888 55958 65904
rect 55698 65789 55846 65871
rect 55586 65756 55663 65772
tri 55663 65756 55679 65772 sw
rect 55586 65690 55679 65756
rect 55715 65631 55829 65789
tri 55865 65756 55881 65772 se
rect 55881 65756 55958 65772
rect 55865 65690 55958 65756
rect 55586 65555 55958 65631
rect 55586 65430 55679 65496
rect 55586 65414 55663 65430
tri 55663 65414 55679 65430 nw
rect 55715 65397 55829 65555
rect 55865 65430 55958 65496
tri 55865 65414 55881 65430 ne
rect 55881 65414 55958 65430
rect 55698 65315 55846 65397
rect 55586 65282 55663 65298
tri 55663 65282 55679 65298 sw
rect 55586 65216 55679 65282
rect 55586 65114 55679 65180
rect 55586 65098 55663 65114
tri 55663 65098 55679 65114 nw
rect 55715 65081 55829 65315
tri 55865 65282 55881 65298 se
rect 55881 65282 55958 65298
rect 55865 65216 55958 65282
rect 55865 65114 55958 65180
tri 55865 65098 55881 65114 ne
rect 55881 65098 55958 65114
rect 55698 64999 55846 65081
rect 55586 64966 55663 64982
tri 55663 64966 55679 64982 sw
rect 55586 64900 55679 64966
rect 55715 64841 55829 64999
tri 55865 64966 55881 64982 se
rect 55881 64966 55958 64982
rect 55865 64900 55958 64966
rect 55586 64765 55958 64841
rect 55586 64640 55679 64706
rect 55586 64624 55663 64640
tri 55663 64624 55679 64640 nw
rect 55715 64607 55829 64765
rect 55865 64640 55958 64706
tri 55865 64624 55881 64640 ne
rect 55881 64624 55958 64640
rect 55698 64525 55846 64607
rect 55586 64492 55663 64508
tri 55663 64492 55679 64508 sw
rect 55586 64426 55679 64492
rect 55586 64324 55679 64390
rect 55586 64308 55663 64324
tri 55663 64308 55679 64324 nw
rect 55715 64291 55829 64525
tri 55865 64492 55881 64508 se
rect 55881 64492 55958 64508
rect 55865 64426 55958 64492
rect 55865 64324 55958 64390
tri 55865 64308 55881 64324 ne
rect 55881 64308 55958 64324
rect 55698 64209 55846 64291
rect 55586 64176 55663 64192
tri 55663 64176 55679 64192 sw
rect 55586 64110 55679 64176
rect 55715 64051 55829 64209
tri 55865 64176 55881 64192 se
rect 55881 64176 55958 64192
rect 55865 64110 55958 64176
rect 55586 63975 55958 64051
rect 55586 63850 55679 63916
rect 55586 63834 55663 63850
tri 55663 63834 55679 63850 nw
rect 55715 63817 55829 63975
rect 55865 63850 55958 63916
tri 55865 63834 55881 63850 ne
rect 55881 63834 55958 63850
rect 55698 63735 55846 63817
rect 55586 63702 55663 63718
tri 55663 63702 55679 63718 sw
rect 55586 63636 55679 63702
rect 55586 63534 55679 63600
rect 55586 63518 55663 63534
tri 55663 63518 55679 63534 nw
rect 55715 63501 55829 63735
tri 55865 63702 55881 63718 se
rect 55881 63702 55958 63718
rect 55865 63636 55958 63702
rect 55865 63534 55958 63600
tri 55865 63518 55881 63534 ne
rect 55881 63518 55958 63534
rect 55698 63419 55846 63501
rect 55586 63386 55663 63402
tri 55663 63386 55679 63402 sw
rect 55586 63320 55679 63386
rect 55715 63261 55829 63419
tri 55865 63386 55881 63402 se
rect 55881 63386 55958 63402
rect 55865 63320 55958 63386
rect 55586 63185 55958 63261
rect 55586 63060 55679 63126
rect 55586 63044 55663 63060
tri 55663 63044 55679 63060 nw
rect 55715 63027 55829 63185
rect 55865 63060 55958 63126
tri 55865 63044 55881 63060 ne
rect 55881 63044 55958 63060
rect 55698 62945 55846 63027
rect 55586 62912 55663 62928
tri 55663 62912 55679 62928 sw
rect 55586 62846 55679 62912
rect 55586 62744 55679 62810
rect 55586 62728 55663 62744
tri 55663 62728 55679 62744 nw
rect 55715 62711 55829 62945
tri 55865 62912 55881 62928 se
rect 55881 62912 55958 62928
rect 55865 62846 55958 62912
rect 55865 62744 55958 62810
tri 55865 62728 55881 62744 ne
rect 55881 62728 55958 62744
rect 55698 62629 55846 62711
rect 55586 62596 55663 62612
tri 55663 62596 55679 62612 sw
rect 55586 62530 55679 62596
rect 55715 62471 55829 62629
tri 55865 62596 55881 62612 se
rect 55881 62596 55958 62612
rect 55865 62530 55958 62596
rect 55586 62395 55958 62471
rect 55586 62270 55679 62336
rect 55586 62254 55663 62270
tri 55663 62254 55679 62270 nw
rect 55715 62237 55829 62395
rect 55865 62270 55958 62336
tri 55865 62254 55881 62270 ne
rect 55881 62254 55958 62270
rect 55698 62155 55846 62237
rect 55586 62122 55663 62138
tri 55663 62122 55679 62138 sw
rect 55586 62056 55679 62122
rect 55586 61954 55679 62020
rect 55586 61938 55663 61954
tri 55663 61938 55679 61954 nw
rect 55715 61921 55829 62155
tri 55865 62122 55881 62138 se
rect 55881 62122 55958 62138
rect 55865 62056 55958 62122
rect 55865 61954 55958 62020
tri 55865 61938 55881 61954 ne
rect 55881 61938 55958 61954
rect 55698 61839 55846 61921
rect 55586 61806 55663 61822
tri 55663 61806 55679 61822 sw
rect 55586 61740 55679 61806
rect 55715 61681 55829 61839
tri 55865 61806 55881 61822 se
rect 55881 61806 55958 61822
rect 55865 61740 55958 61806
rect 55586 61605 55958 61681
rect 55586 61480 55679 61546
rect 55586 61464 55663 61480
tri 55663 61464 55679 61480 nw
rect 55715 61447 55829 61605
rect 55865 61480 55958 61546
tri 55865 61464 55881 61480 ne
rect 55881 61464 55958 61480
rect 55698 61365 55846 61447
rect 55586 61332 55663 61348
tri 55663 61332 55679 61348 sw
rect 55586 61266 55679 61332
rect 55586 61164 55679 61230
rect 55586 61148 55663 61164
tri 55663 61148 55679 61164 nw
rect 55715 61131 55829 61365
tri 55865 61332 55881 61348 se
rect 55881 61332 55958 61348
rect 55865 61266 55958 61332
rect 55865 61164 55958 61230
tri 55865 61148 55881 61164 ne
rect 55881 61148 55958 61164
rect 55698 61049 55846 61131
rect 55586 61016 55663 61032
tri 55663 61016 55679 61032 sw
rect 55586 60950 55679 61016
rect 55715 60891 55829 61049
tri 55865 61016 55881 61032 se
rect 55881 61016 55958 61032
rect 55865 60950 55958 61016
rect 55586 60815 55958 60891
rect 55586 60690 55679 60756
rect 55586 60674 55663 60690
tri 55663 60674 55679 60690 nw
rect 55715 60657 55829 60815
rect 55865 60690 55958 60756
tri 55865 60674 55881 60690 ne
rect 55881 60674 55958 60690
rect 55698 60575 55846 60657
rect 55586 60542 55663 60558
tri 55663 60542 55679 60558 sw
rect 55586 60476 55679 60542
rect 55586 60374 55679 60440
rect 55586 60358 55663 60374
tri 55663 60358 55679 60374 nw
rect 55715 60341 55829 60575
tri 55865 60542 55881 60558 se
rect 55881 60542 55958 60558
rect 55865 60476 55958 60542
rect 55865 60374 55958 60440
tri 55865 60358 55881 60374 ne
rect 55881 60358 55958 60374
rect 55698 60259 55846 60341
rect 55586 60226 55663 60242
tri 55663 60226 55679 60242 sw
rect 55586 60160 55679 60226
rect 55715 60101 55829 60259
tri 55865 60226 55881 60242 se
rect 55881 60226 55958 60242
rect 55865 60160 55958 60226
rect 55586 60025 55958 60101
rect 55586 59900 55679 59966
rect 55586 59884 55663 59900
tri 55663 59884 55679 59900 nw
rect 55715 59867 55829 60025
rect 55865 59900 55958 59966
tri 55865 59884 55881 59900 ne
rect 55881 59884 55958 59900
rect 55698 59785 55846 59867
rect 55586 59752 55663 59768
tri 55663 59752 55679 59768 sw
rect 55586 59686 55679 59752
rect 55586 59584 55679 59650
rect 55586 59568 55663 59584
tri 55663 59568 55679 59584 nw
rect 55715 59551 55829 59785
tri 55865 59752 55881 59768 se
rect 55881 59752 55958 59768
rect 55865 59686 55958 59752
rect 55865 59584 55958 59650
tri 55865 59568 55881 59584 ne
rect 55881 59568 55958 59584
rect 55698 59469 55846 59551
rect 55586 59436 55663 59452
tri 55663 59436 55679 59452 sw
rect 55586 59370 55679 59436
rect 55715 59311 55829 59469
tri 55865 59436 55881 59452 se
rect 55881 59436 55958 59452
rect 55865 59370 55958 59436
rect 55586 59235 55958 59311
rect 55586 59110 55679 59176
rect 55586 59094 55663 59110
tri 55663 59094 55679 59110 nw
rect 55715 59077 55829 59235
rect 55865 59110 55958 59176
tri 55865 59094 55881 59110 ne
rect 55881 59094 55958 59110
rect 55698 58995 55846 59077
rect 55586 58962 55663 58978
tri 55663 58962 55679 58978 sw
rect 55586 58896 55679 58962
rect 55586 58794 55679 58860
rect 55586 58778 55663 58794
tri 55663 58778 55679 58794 nw
rect 55715 58761 55829 58995
tri 55865 58962 55881 58978 se
rect 55881 58962 55958 58978
rect 55865 58896 55958 58962
rect 55865 58794 55958 58860
tri 55865 58778 55881 58794 ne
rect 55881 58778 55958 58794
rect 55698 58679 55846 58761
rect 55586 58646 55663 58662
tri 55663 58646 55679 58662 sw
rect 55586 58580 55679 58646
rect 55715 58521 55829 58679
tri 55865 58646 55881 58662 se
rect 55881 58646 55958 58662
rect 55865 58580 55958 58646
rect 55586 58445 55958 58521
rect 55586 58320 55679 58386
rect 55586 58304 55663 58320
tri 55663 58304 55679 58320 nw
rect 55715 58287 55829 58445
rect 55865 58320 55958 58386
tri 55865 58304 55881 58320 ne
rect 55881 58304 55958 58320
rect 55698 58205 55846 58287
rect 55586 58172 55663 58188
tri 55663 58172 55679 58188 sw
rect 55586 58106 55679 58172
rect 55586 58004 55679 58070
rect 55586 57988 55663 58004
tri 55663 57988 55679 58004 nw
rect 55715 57971 55829 58205
tri 55865 58172 55881 58188 se
rect 55881 58172 55958 58188
rect 55865 58106 55958 58172
rect 55865 58004 55958 58070
tri 55865 57988 55881 58004 ne
rect 55881 57988 55958 58004
rect 55698 57889 55846 57971
rect 55586 57856 55663 57872
tri 55663 57856 55679 57872 sw
rect 55586 57790 55679 57856
rect 55715 57731 55829 57889
tri 55865 57856 55881 57872 se
rect 55881 57856 55958 57872
rect 55865 57790 55958 57856
rect 55586 57655 55958 57731
rect 55586 57530 55679 57596
rect 55586 57514 55663 57530
tri 55663 57514 55679 57530 nw
rect 55715 57497 55829 57655
rect 55865 57530 55958 57596
tri 55865 57514 55881 57530 ne
rect 55881 57514 55958 57530
rect 55698 57415 55846 57497
rect 55586 57382 55663 57398
tri 55663 57382 55679 57398 sw
rect 55586 57316 55679 57382
rect 55586 57214 55679 57280
rect 55586 57198 55663 57214
tri 55663 57198 55679 57214 nw
rect 55715 57181 55829 57415
tri 55865 57382 55881 57398 se
rect 55881 57382 55958 57398
rect 55865 57316 55958 57382
rect 55865 57214 55958 57280
tri 55865 57198 55881 57214 ne
rect 55881 57198 55958 57214
rect 55698 57099 55846 57181
rect 55586 57066 55663 57082
tri 55663 57066 55679 57082 sw
rect 55586 57000 55679 57066
rect 55715 56941 55829 57099
tri 55865 57066 55881 57082 se
rect 55881 57066 55958 57082
rect 55865 57000 55958 57066
rect 55586 56865 55958 56941
rect 55586 56740 55679 56806
rect 55586 56724 55663 56740
tri 55663 56724 55679 56740 nw
rect 55715 56707 55829 56865
rect 55865 56740 55958 56806
tri 55865 56724 55881 56740 ne
rect 55881 56724 55958 56740
rect 55698 56625 55846 56707
rect 55586 56592 55663 56608
tri 55663 56592 55679 56608 sw
rect 55586 56526 55679 56592
rect 55586 56424 55679 56490
rect 55586 56408 55663 56424
tri 55663 56408 55679 56424 nw
rect 55715 56391 55829 56625
tri 55865 56592 55881 56608 se
rect 55881 56592 55958 56608
rect 55865 56526 55958 56592
rect 55865 56424 55958 56490
tri 55865 56408 55881 56424 ne
rect 55881 56408 55958 56424
rect 55698 56309 55846 56391
rect 55586 56276 55663 56292
tri 55663 56276 55679 56292 sw
rect 55586 56210 55679 56276
rect 55715 56151 55829 56309
tri 55865 56276 55881 56292 se
rect 55881 56276 55958 56292
rect 55865 56210 55958 56276
rect 55586 56075 55958 56151
rect 55586 55950 55679 56016
rect 55586 55934 55663 55950
tri 55663 55934 55679 55950 nw
rect 55715 55917 55829 56075
rect 55865 55950 55958 56016
tri 55865 55934 55881 55950 ne
rect 55881 55934 55958 55950
rect 55698 55835 55846 55917
rect 55586 55802 55663 55818
tri 55663 55802 55679 55818 sw
rect 55586 55736 55679 55802
rect 55586 55634 55679 55700
rect 55586 55618 55663 55634
tri 55663 55618 55679 55634 nw
rect 55715 55601 55829 55835
tri 55865 55802 55881 55818 se
rect 55881 55802 55958 55818
rect 55865 55736 55958 55802
rect 55865 55634 55958 55700
tri 55865 55618 55881 55634 ne
rect 55881 55618 55958 55634
rect 55698 55519 55846 55601
rect 55586 55486 55663 55502
tri 55663 55486 55679 55502 sw
rect 55586 55420 55679 55486
rect 55715 55361 55829 55519
tri 55865 55486 55881 55502 se
rect 55881 55486 55958 55502
rect 55865 55420 55958 55486
rect 55586 55285 55958 55361
rect 55586 55160 55679 55226
rect 55586 55144 55663 55160
tri 55663 55144 55679 55160 nw
rect 55715 55127 55829 55285
rect 55865 55160 55958 55226
tri 55865 55144 55881 55160 ne
rect 55881 55144 55958 55160
rect 55698 55045 55846 55127
rect 55586 55012 55663 55028
tri 55663 55012 55679 55028 sw
rect 55586 54946 55679 55012
rect 55586 54844 55679 54910
rect 55586 54828 55663 54844
tri 55663 54828 55679 54844 nw
rect 55715 54811 55829 55045
tri 55865 55012 55881 55028 se
rect 55881 55012 55958 55028
rect 55865 54946 55958 55012
rect 55865 54844 55958 54910
tri 55865 54828 55881 54844 ne
rect 55881 54828 55958 54844
rect 55698 54729 55846 54811
rect 55586 54696 55663 54712
tri 55663 54696 55679 54712 sw
rect 55586 54630 55679 54696
rect 55715 54571 55829 54729
tri 55865 54696 55881 54712 se
rect 55881 54696 55958 54712
rect 55865 54630 55958 54696
rect 55586 54495 55958 54571
rect 55586 54370 55679 54436
rect 55586 54354 55663 54370
tri 55663 54354 55679 54370 nw
rect 55715 54337 55829 54495
rect 55865 54370 55958 54436
tri 55865 54354 55881 54370 ne
rect 55881 54354 55958 54370
rect 55698 54255 55846 54337
rect 55586 54222 55663 54238
tri 55663 54222 55679 54238 sw
rect 55586 54156 55679 54222
rect 55586 54054 55679 54120
rect 55586 54038 55663 54054
tri 55663 54038 55679 54054 nw
rect 55715 54021 55829 54255
tri 55865 54222 55881 54238 se
rect 55881 54222 55958 54238
rect 55865 54156 55958 54222
rect 55865 54054 55958 54120
tri 55865 54038 55881 54054 ne
rect 55881 54038 55958 54054
rect 55698 53939 55846 54021
rect 55586 53906 55663 53922
tri 55663 53906 55679 53922 sw
rect 55586 53840 55679 53906
rect 55715 53781 55829 53939
tri 55865 53906 55881 53922 se
rect 55881 53906 55958 53922
rect 55865 53840 55958 53906
rect 55586 53705 55958 53781
rect 55586 53580 55679 53646
rect 55586 53564 55663 53580
tri 55663 53564 55679 53580 nw
rect 55715 53547 55829 53705
rect 55865 53580 55958 53646
tri 55865 53564 55881 53580 ne
rect 55881 53564 55958 53580
rect 55698 53465 55846 53547
rect 55586 53432 55663 53448
tri 55663 53432 55679 53448 sw
rect 55586 53366 55679 53432
rect 55586 53264 55679 53330
rect 55586 53248 55663 53264
tri 55663 53248 55679 53264 nw
rect 55715 53231 55829 53465
tri 55865 53432 55881 53448 se
rect 55881 53432 55958 53448
rect 55865 53366 55958 53432
rect 55865 53264 55958 53330
tri 55865 53248 55881 53264 ne
rect 55881 53248 55958 53264
rect 55698 53149 55846 53231
rect 55586 53116 55663 53132
tri 55663 53116 55679 53132 sw
rect 55586 53050 55679 53116
rect 55715 52991 55829 53149
tri 55865 53116 55881 53132 se
rect 55881 53116 55958 53132
rect 55865 53050 55958 53116
rect 55586 52915 55958 52991
rect 55586 52790 55679 52856
rect 55586 52774 55663 52790
tri 55663 52774 55679 52790 nw
rect 55715 52757 55829 52915
rect 55865 52790 55958 52856
tri 55865 52774 55881 52790 ne
rect 55881 52774 55958 52790
rect 55698 52675 55846 52757
rect 55586 52642 55663 52658
tri 55663 52642 55679 52658 sw
rect 55586 52576 55679 52642
rect 55586 52474 55679 52540
rect 55586 52458 55663 52474
tri 55663 52458 55679 52474 nw
rect 55715 52441 55829 52675
tri 55865 52642 55881 52658 se
rect 55881 52642 55958 52658
rect 55865 52576 55958 52642
rect 55865 52474 55958 52540
tri 55865 52458 55881 52474 ne
rect 55881 52458 55958 52474
rect 55698 52359 55846 52441
rect 55586 52326 55663 52342
tri 55663 52326 55679 52342 sw
rect 55586 52260 55679 52326
rect 55715 52201 55829 52359
tri 55865 52326 55881 52342 se
rect 55881 52326 55958 52342
rect 55865 52260 55958 52326
rect 55586 52125 55958 52201
rect 55586 52000 55679 52066
rect 55586 51984 55663 52000
tri 55663 51984 55679 52000 nw
rect 55715 51967 55829 52125
rect 55865 52000 55958 52066
tri 55865 51984 55881 52000 ne
rect 55881 51984 55958 52000
rect 55698 51885 55846 51967
rect 55586 51852 55663 51868
tri 55663 51852 55679 51868 sw
rect 55586 51786 55679 51852
rect 55586 51684 55679 51750
rect 55586 51668 55663 51684
tri 55663 51668 55679 51684 nw
rect 55715 51651 55829 51885
tri 55865 51852 55881 51868 se
rect 55881 51852 55958 51868
rect 55865 51786 55958 51852
rect 55865 51684 55958 51750
tri 55865 51668 55881 51684 ne
rect 55881 51668 55958 51684
rect 55698 51569 55846 51651
rect 55586 51536 55663 51552
tri 55663 51536 55679 51552 sw
rect 55586 51470 55679 51536
rect 55715 51411 55829 51569
tri 55865 51536 55881 51552 se
rect 55881 51536 55958 51552
rect 55865 51470 55958 51536
rect 55586 51335 55958 51411
rect 55586 51210 55679 51276
rect 55586 51194 55663 51210
tri 55663 51194 55679 51210 nw
rect 55715 51177 55829 51335
rect 55865 51210 55958 51276
tri 55865 51194 55881 51210 ne
rect 55881 51194 55958 51210
rect 55698 51095 55846 51177
rect 55586 51062 55663 51078
tri 55663 51062 55679 51078 sw
rect 55586 50996 55679 51062
rect 55586 50894 55679 50960
rect 55586 50878 55663 50894
tri 55663 50878 55679 50894 nw
rect 55715 50861 55829 51095
tri 55865 51062 55881 51078 se
rect 55881 51062 55958 51078
rect 55865 50996 55958 51062
rect 55865 50894 55958 50960
tri 55865 50878 55881 50894 ne
rect 55881 50878 55958 50894
rect 55698 50779 55846 50861
rect 55586 50746 55663 50762
tri 55663 50746 55679 50762 sw
rect 55586 50680 55679 50746
rect 55715 50621 55829 50779
tri 55865 50746 55881 50762 se
rect 55881 50746 55958 50762
rect 55865 50680 55958 50746
rect 55586 50545 55958 50621
rect 55586 50420 55679 50486
rect 55586 50404 55663 50420
tri 55663 50404 55679 50420 nw
rect 55715 50387 55829 50545
rect 55865 50420 55958 50486
tri 55865 50404 55881 50420 ne
rect 55881 50404 55958 50420
rect 55698 50305 55846 50387
rect 55586 50272 55663 50288
tri 55663 50272 55679 50288 sw
rect 55586 50206 55679 50272
rect 55586 50104 55679 50170
rect 55586 50088 55663 50104
tri 55663 50088 55679 50104 nw
rect 55715 50071 55829 50305
tri 55865 50272 55881 50288 se
rect 55881 50272 55958 50288
rect 55865 50206 55958 50272
rect 55865 50104 55958 50170
tri 55865 50088 55881 50104 ne
rect 55881 50088 55958 50104
rect 55698 49989 55846 50071
rect 55586 49956 55663 49972
tri 55663 49956 55679 49972 sw
rect 55586 49890 55679 49956
rect 55715 49831 55829 49989
tri 55865 49956 55881 49972 se
rect 55881 49956 55958 49972
rect 55865 49890 55958 49956
rect 55586 49755 55958 49831
rect 55586 49630 55679 49696
rect 55586 49614 55663 49630
tri 55663 49614 55679 49630 nw
rect 55715 49597 55829 49755
rect 55865 49630 55958 49696
tri 55865 49614 55881 49630 ne
rect 55881 49614 55958 49630
rect 55698 49515 55846 49597
rect 55586 49482 55663 49498
tri 55663 49482 55679 49498 sw
rect 55586 49416 55679 49482
rect 55586 49314 55679 49380
rect 55586 49298 55663 49314
tri 55663 49298 55679 49314 nw
rect 55715 49281 55829 49515
tri 55865 49482 55881 49498 se
rect 55881 49482 55958 49498
rect 55865 49416 55958 49482
rect 55865 49314 55958 49380
tri 55865 49298 55881 49314 ne
rect 55881 49298 55958 49314
rect 55698 49199 55846 49281
rect 55586 49166 55663 49182
tri 55663 49166 55679 49182 sw
rect 55586 49100 55679 49166
rect 55715 49041 55829 49199
tri 55865 49166 55881 49182 se
rect 55881 49166 55958 49182
rect 55865 49100 55958 49166
rect 55586 48965 55958 49041
rect 55586 48840 55679 48906
rect 55586 48824 55663 48840
tri 55663 48824 55679 48840 nw
rect 55715 48807 55829 48965
rect 55865 48840 55958 48906
tri 55865 48824 55881 48840 ne
rect 55881 48824 55958 48840
rect 55698 48725 55846 48807
rect 55586 48692 55663 48708
tri 55663 48692 55679 48708 sw
rect 55586 48626 55679 48692
rect 55586 48524 55679 48590
rect 55586 48508 55663 48524
tri 55663 48508 55679 48524 nw
rect 55715 48491 55829 48725
tri 55865 48692 55881 48708 se
rect 55881 48692 55958 48708
rect 55865 48626 55958 48692
rect 55865 48524 55958 48590
tri 55865 48508 55881 48524 ne
rect 55881 48508 55958 48524
rect 55698 48409 55846 48491
rect 55586 48376 55663 48392
tri 55663 48376 55679 48392 sw
rect 55586 48310 55679 48376
rect 55715 48251 55829 48409
tri 55865 48376 55881 48392 se
rect 55881 48376 55958 48392
rect 55865 48310 55958 48376
rect 55586 48175 55958 48251
rect 55586 48050 55679 48116
rect 55586 48034 55663 48050
tri 55663 48034 55679 48050 nw
rect 55715 48017 55829 48175
rect 55865 48050 55958 48116
tri 55865 48034 55881 48050 ne
rect 55881 48034 55958 48050
rect 55698 47935 55846 48017
rect 55586 47902 55663 47918
tri 55663 47902 55679 47918 sw
rect 55586 47836 55679 47902
rect 55586 47734 55679 47800
rect 55586 47718 55663 47734
tri 55663 47718 55679 47734 nw
rect 55715 47701 55829 47935
tri 55865 47902 55881 47918 se
rect 55881 47902 55958 47918
rect 55865 47836 55958 47902
rect 55865 47734 55958 47800
tri 55865 47718 55881 47734 ne
rect 55881 47718 55958 47734
rect 55698 47619 55846 47701
rect 55586 47586 55663 47602
tri 55663 47586 55679 47602 sw
rect 55586 47520 55679 47586
rect 55715 47461 55829 47619
tri 55865 47586 55881 47602 se
rect 55881 47586 55958 47602
rect 55865 47520 55958 47586
rect 55586 47385 55958 47461
rect 55586 47260 55679 47326
rect 55586 47244 55663 47260
tri 55663 47244 55679 47260 nw
rect 55715 47227 55829 47385
rect 55865 47260 55958 47326
tri 55865 47244 55881 47260 ne
rect 55881 47244 55958 47260
rect 55698 47145 55846 47227
rect 55586 47112 55663 47128
tri 55663 47112 55679 47128 sw
rect 55586 47046 55679 47112
rect 55586 46944 55679 47010
rect 55586 46928 55663 46944
tri 55663 46928 55679 46944 nw
rect 55715 46911 55829 47145
tri 55865 47112 55881 47128 se
rect 55881 47112 55958 47128
rect 55865 47046 55958 47112
rect 55865 46944 55958 47010
tri 55865 46928 55881 46944 ne
rect 55881 46928 55958 46944
rect 55698 46829 55846 46911
rect 55586 46796 55663 46812
tri 55663 46796 55679 46812 sw
rect 55586 46730 55679 46796
rect 55715 46671 55829 46829
tri 55865 46796 55881 46812 se
rect 55881 46796 55958 46812
rect 55865 46730 55958 46796
rect 55586 46595 55958 46671
rect 55586 46470 55679 46536
rect 55586 46454 55663 46470
tri 55663 46454 55679 46470 nw
rect 55715 46437 55829 46595
rect 55865 46470 55958 46536
tri 55865 46454 55881 46470 ne
rect 55881 46454 55958 46470
rect 55698 46355 55846 46437
rect 55586 46322 55663 46338
tri 55663 46322 55679 46338 sw
rect 55586 46256 55679 46322
rect 55586 46154 55679 46220
rect 55586 46138 55663 46154
tri 55663 46138 55679 46154 nw
rect 55715 46121 55829 46355
tri 55865 46322 55881 46338 se
rect 55881 46322 55958 46338
rect 55865 46256 55958 46322
rect 55865 46154 55958 46220
tri 55865 46138 55881 46154 ne
rect 55881 46138 55958 46154
rect 55698 46039 55846 46121
rect 55586 46006 55663 46022
tri 55663 46006 55679 46022 sw
rect 55586 45940 55679 46006
rect 55715 45881 55829 46039
tri 55865 46006 55881 46022 se
rect 55881 46006 55958 46022
rect 55865 45940 55958 46006
rect 55586 45805 55958 45881
rect 55586 45680 55679 45746
rect 55586 45664 55663 45680
tri 55663 45664 55679 45680 nw
rect 55715 45647 55829 45805
rect 55865 45680 55958 45746
tri 55865 45664 55881 45680 ne
rect 55881 45664 55958 45680
rect 55698 45565 55846 45647
rect 55586 45532 55663 45548
tri 55663 45532 55679 45548 sw
rect 55586 45466 55679 45532
rect 55586 45364 55679 45430
rect 55586 45348 55663 45364
tri 55663 45348 55679 45364 nw
rect 55715 45331 55829 45565
tri 55865 45532 55881 45548 se
rect 55881 45532 55958 45548
rect 55865 45466 55958 45532
rect 55865 45364 55958 45430
tri 55865 45348 55881 45364 ne
rect 55881 45348 55958 45364
rect 55698 45249 55846 45331
rect 55586 45216 55663 45232
tri 55663 45216 55679 45232 sw
rect 55586 45150 55679 45216
rect 55715 45091 55829 45249
tri 55865 45216 55881 45232 se
rect 55881 45216 55958 45232
rect 55865 45150 55958 45216
rect 55586 45015 55958 45091
rect 55586 44890 55679 44956
rect 55586 44874 55663 44890
tri 55663 44874 55679 44890 nw
rect 55715 44857 55829 45015
rect 55865 44890 55958 44956
tri 55865 44874 55881 44890 ne
rect 55881 44874 55958 44890
rect 55698 44775 55846 44857
rect 55586 44742 55663 44758
tri 55663 44742 55679 44758 sw
rect 55586 44676 55679 44742
rect 55586 44574 55679 44640
rect 55586 44558 55663 44574
tri 55663 44558 55679 44574 nw
rect 55715 44541 55829 44775
tri 55865 44742 55881 44758 se
rect 55881 44742 55958 44758
rect 55865 44676 55958 44742
rect 55865 44574 55958 44640
tri 55865 44558 55881 44574 ne
rect 55881 44558 55958 44574
rect 55698 44459 55846 44541
rect 55586 44426 55663 44442
tri 55663 44426 55679 44442 sw
rect 55586 44360 55679 44426
rect 55715 44301 55829 44459
tri 55865 44426 55881 44442 se
rect 55881 44426 55958 44442
rect 55865 44360 55958 44426
rect 55586 44225 55958 44301
rect 55586 44100 55679 44166
rect 55586 44084 55663 44100
tri 55663 44084 55679 44100 nw
rect 55715 44067 55829 44225
rect 55865 44100 55958 44166
tri 55865 44084 55881 44100 ne
rect 55881 44084 55958 44100
rect 55698 43985 55846 44067
rect 55586 43952 55663 43968
tri 55663 43952 55679 43968 sw
rect 55586 43886 55679 43952
rect 55586 43784 55679 43850
rect 55586 43768 55663 43784
tri 55663 43768 55679 43784 nw
rect 55715 43751 55829 43985
tri 55865 43952 55881 43968 se
rect 55881 43952 55958 43968
rect 55865 43886 55958 43952
rect 55865 43784 55958 43850
tri 55865 43768 55881 43784 ne
rect 55881 43768 55958 43784
rect 55698 43669 55846 43751
rect 55586 43636 55663 43652
tri 55663 43636 55679 43652 sw
rect 55586 43570 55679 43636
rect 55715 43511 55829 43669
tri 55865 43636 55881 43652 se
rect 55881 43636 55958 43652
rect 55865 43570 55958 43636
rect 55586 43435 55958 43511
rect 55586 43310 55679 43376
rect 55586 43294 55663 43310
tri 55663 43294 55679 43310 nw
rect 55715 43277 55829 43435
rect 55865 43310 55958 43376
tri 55865 43294 55881 43310 ne
rect 55881 43294 55958 43310
rect 55698 43195 55846 43277
rect 55586 43162 55663 43178
tri 55663 43162 55679 43178 sw
rect 55586 43096 55679 43162
rect 55586 42994 55679 43060
rect 55586 42978 55663 42994
tri 55663 42978 55679 42994 nw
rect 55715 42961 55829 43195
tri 55865 43162 55881 43178 se
rect 55881 43162 55958 43178
rect 55865 43096 55958 43162
rect 55865 42994 55958 43060
tri 55865 42978 55881 42994 ne
rect 55881 42978 55958 42994
rect 55698 42879 55846 42961
rect 55586 42846 55663 42862
tri 55663 42846 55679 42862 sw
rect 55586 42780 55679 42846
rect 55715 42721 55829 42879
tri 55865 42846 55881 42862 se
rect 55881 42846 55958 42862
rect 55865 42780 55958 42846
rect 55586 42645 55958 42721
rect 55586 42520 55679 42586
rect 55586 42504 55663 42520
tri 55663 42504 55679 42520 nw
rect 55715 42487 55829 42645
rect 55865 42520 55958 42586
tri 55865 42504 55881 42520 ne
rect 55881 42504 55958 42520
rect 55698 42405 55846 42487
rect 55586 42372 55663 42388
tri 55663 42372 55679 42388 sw
rect 55586 42306 55679 42372
rect 55586 42204 55679 42270
rect 55586 42188 55663 42204
tri 55663 42188 55679 42204 nw
rect 55715 42171 55829 42405
tri 55865 42372 55881 42388 se
rect 55881 42372 55958 42388
rect 55865 42306 55958 42372
rect 55865 42204 55958 42270
tri 55865 42188 55881 42204 ne
rect 55881 42188 55958 42204
rect 55698 42089 55846 42171
rect 55586 42056 55663 42072
tri 55663 42056 55679 42072 sw
rect 55586 41990 55679 42056
rect 55715 41931 55829 42089
tri 55865 42056 55881 42072 se
rect 55881 42056 55958 42072
rect 55865 41990 55958 42056
rect 55586 41855 55958 41931
rect 55586 41730 55679 41796
rect 55586 41714 55663 41730
tri 55663 41714 55679 41730 nw
rect 55715 41697 55829 41855
rect 55865 41730 55958 41796
tri 55865 41714 55881 41730 ne
rect 55881 41714 55958 41730
rect 55698 41615 55846 41697
rect 55586 41582 55663 41598
tri 55663 41582 55679 41598 sw
rect 55586 41516 55679 41582
rect 55586 41414 55679 41480
rect 55586 41398 55663 41414
tri 55663 41398 55679 41414 nw
rect 55715 41381 55829 41615
tri 55865 41582 55881 41598 se
rect 55881 41582 55958 41598
rect 55865 41516 55958 41582
rect 55865 41414 55958 41480
tri 55865 41398 55881 41414 ne
rect 55881 41398 55958 41414
rect 55698 41299 55846 41381
rect 55586 41266 55663 41282
tri 55663 41266 55679 41282 sw
rect 55586 41200 55679 41266
rect 55715 41141 55829 41299
tri 55865 41266 55881 41282 se
rect 55881 41266 55958 41282
rect 55865 41200 55958 41266
rect 55586 41065 55958 41141
rect 55586 40940 55679 41006
rect 55586 40924 55663 40940
tri 55663 40924 55679 40940 nw
rect 55715 40907 55829 41065
rect 55865 40940 55958 41006
tri 55865 40924 55881 40940 ne
rect 55881 40924 55958 40940
rect 55698 40825 55846 40907
rect 55586 40792 55663 40808
tri 55663 40792 55679 40808 sw
rect 55586 40726 55679 40792
rect 55586 40624 55679 40690
rect 55586 40608 55663 40624
tri 55663 40608 55679 40624 nw
rect 55715 40591 55829 40825
tri 55865 40792 55881 40808 se
rect 55881 40792 55958 40808
rect 55865 40726 55958 40792
rect 55865 40624 55958 40690
tri 55865 40608 55881 40624 ne
rect 55881 40608 55958 40624
rect 55698 40509 55846 40591
rect 55586 40476 55663 40492
tri 55663 40476 55679 40492 sw
rect 55586 40410 55679 40476
rect 55715 40351 55829 40509
tri 55865 40476 55881 40492 se
rect 55881 40476 55958 40492
rect 55865 40410 55958 40476
rect 55586 40275 55958 40351
rect 55586 40150 55679 40216
rect 55586 40134 55663 40150
tri 55663 40134 55679 40150 nw
rect 55715 40117 55829 40275
rect 55865 40150 55958 40216
tri 55865 40134 55881 40150 ne
rect 55881 40134 55958 40150
rect 55698 40035 55846 40117
rect 55586 40002 55663 40018
tri 55663 40002 55679 40018 sw
rect 55586 39936 55679 40002
rect 55586 39834 55679 39900
rect 55586 39818 55663 39834
tri 55663 39818 55679 39834 nw
rect 55715 39801 55829 40035
tri 55865 40002 55881 40018 se
rect 55881 40002 55958 40018
rect 55865 39936 55958 40002
rect 55865 39834 55958 39900
tri 55865 39818 55881 39834 ne
rect 55881 39818 55958 39834
rect 55698 39719 55846 39801
rect 55586 39686 55663 39702
tri 55663 39686 55679 39702 sw
rect 55586 39620 55679 39686
rect 55715 39561 55829 39719
tri 55865 39686 55881 39702 se
rect 55881 39686 55958 39702
rect 55865 39620 55958 39686
rect 55586 39485 55958 39561
rect 55586 39360 55679 39426
rect 55586 39344 55663 39360
tri 55663 39344 55679 39360 nw
rect 55715 39327 55829 39485
rect 55865 39360 55958 39426
tri 55865 39344 55881 39360 ne
rect 55881 39344 55958 39360
rect 55698 39245 55846 39327
rect 55586 39212 55663 39228
tri 55663 39212 55679 39228 sw
rect 55586 39146 55679 39212
rect 55586 39044 55679 39110
rect 55586 39028 55663 39044
tri 55663 39028 55679 39044 nw
rect 55715 39011 55829 39245
tri 55865 39212 55881 39228 se
rect 55881 39212 55958 39228
rect 55865 39146 55958 39212
rect 55865 39044 55958 39110
tri 55865 39028 55881 39044 ne
rect 55881 39028 55958 39044
rect 55698 38929 55846 39011
rect 55586 38896 55663 38912
tri 55663 38896 55679 38912 sw
rect 55586 38830 55679 38896
rect 55715 38771 55829 38929
tri 55865 38896 55881 38912 se
rect 55881 38896 55958 38912
rect 55865 38830 55958 38896
rect 55586 38695 55958 38771
rect 55586 38570 55679 38636
rect 55586 38554 55663 38570
tri 55663 38554 55679 38570 nw
rect 55715 38537 55829 38695
rect 55865 38570 55958 38636
tri 55865 38554 55881 38570 ne
rect 55881 38554 55958 38570
rect 55698 38455 55846 38537
rect 55586 38422 55663 38438
tri 55663 38422 55679 38438 sw
rect 55586 38356 55679 38422
rect 55586 38254 55679 38320
rect 55586 38238 55663 38254
tri 55663 38238 55679 38254 nw
rect 55715 38221 55829 38455
tri 55865 38422 55881 38438 se
rect 55881 38422 55958 38438
rect 55865 38356 55958 38422
rect 55865 38254 55958 38320
tri 55865 38238 55881 38254 ne
rect 55881 38238 55958 38254
rect 55698 38139 55846 38221
rect 55586 38106 55663 38122
tri 55663 38106 55679 38122 sw
rect 55586 38040 55679 38106
rect 55715 37981 55829 38139
tri 55865 38106 55881 38122 se
rect 55881 38106 55958 38122
rect 55865 38040 55958 38106
rect 55586 37905 55958 37981
rect 55586 37780 55679 37846
rect 55586 37764 55663 37780
tri 55663 37764 55679 37780 nw
rect 55715 37747 55829 37905
rect 55865 37780 55958 37846
tri 55865 37764 55881 37780 ne
rect 55881 37764 55958 37780
rect 55698 37665 55846 37747
rect 55586 37632 55663 37648
tri 55663 37632 55679 37648 sw
rect 55586 37566 55679 37632
rect 55586 37464 55679 37530
rect 55586 37448 55663 37464
tri 55663 37448 55679 37464 nw
rect 55715 37431 55829 37665
tri 55865 37632 55881 37648 se
rect 55881 37632 55958 37648
rect 55865 37566 55958 37632
rect 55865 37464 55958 37530
tri 55865 37448 55881 37464 ne
rect 55881 37448 55958 37464
rect 55698 37349 55846 37431
rect 55586 37316 55663 37332
tri 55663 37316 55679 37332 sw
rect 55586 37250 55679 37316
rect 55715 37191 55829 37349
tri 55865 37316 55881 37332 se
rect 55881 37316 55958 37332
rect 55865 37250 55958 37316
rect 55586 37115 55958 37191
rect 55586 36990 55679 37056
rect 55586 36974 55663 36990
tri 55663 36974 55679 36990 nw
rect 55715 36957 55829 37115
rect 55865 36990 55958 37056
tri 55865 36974 55881 36990 ne
rect 55881 36974 55958 36990
rect 55698 36875 55846 36957
rect 55586 36842 55663 36858
tri 55663 36842 55679 36858 sw
rect 55586 36776 55679 36842
rect 55586 36674 55679 36740
rect 55586 36658 55663 36674
tri 55663 36658 55679 36674 nw
rect 55715 36641 55829 36875
tri 55865 36842 55881 36858 se
rect 55881 36842 55958 36858
rect 55865 36776 55958 36842
rect 55865 36674 55958 36740
tri 55865 36658 55881 36674 ne
rect 55881 36658 55958 36674
rect 55698 36559 55846 36641
rect 55586 36526 55663 36542
tri 55663 36526 55679 36542 sw
rect 55586 36460 55679 36526
rect 55715 36401 55829 36559
tri 55865 36526 55881 36542 se
rect 55881 36526 55958 36542
rect 55865 36460 55958 36526
rect 55586 36325 55958 36401
rect 55586 36200 55679 36266
rect 55586 36184 55663 36200
tri 55663 36184 55679 36200 nw
rect 55715 36167 55829 36325
rect 55865 36200 55958 36266
tri 55865 36184 55881 36200 ne
rect 55881 36184 55958 36200
rect 55698 36085 55846 36167
rect 55586 36052 55663 36068
tri 55663 36052 55679 36068 sw
rect 55586 35986 55679 36052
rect 55586 35884 55679 35950
rect 55586 35868 55663 35884
tri 55663 35868 55679 35884 nw
rect 55715 35851 55829 36085
tri 55865 36052 55881 36068 se
rect 55881 36052 55958 36068
rect 55865 35986 55958 36052
rect 55865 35884 55958 35950
tri 55865 35868 55881 35884 ne
rect 55881 35868 55958 35884
rect 55698 35769 55846 35851
rect 55586 35736 55663 35752
tri 55663 35736 55679 35752 sw
rect 55586 35670 55679 35736
rect 55715 35611 55829 35769
tri 55865 35736 55881 35752 se
rect 55881 35736 55958 35752
rect 55865 35670 55958 35736
rect 55586 35535 55958 35611
rect 55586 35410 55679 35476
rect 55586 35394 55663 35410
tri 55663 35394 55679 35410 nw
rect 55715 35377 55829 35535
rect 55865 35410 55958 35476
tri 55865 35394 55881 35410 ne
rect 55881 35394 55958 35410
rect 55698 35295 55846 35377
rect 55586 35262 55663 35278
tri 55663 35262 55679 35278 sw
rect 55586 35196 55679 35262
rect 55586 35094 55679 35160
rect 55586 35078 55663 35094
tri 55663 35078 55679 35094 nw
rect 55715 35061 55829 35295
tri 55865 35262 55881 35278 se
rect 55881 35262 55958 35278
rect 55865 35196 55958 35262
rect 55865 35094 55958 35160
tri 55865 35078 55881 35094 ne
rect 55881 35078 55958 35094
rect 55698 34979 55846 35061
rect 55586 34946 55663 34962
tri 55663 34946 55679 34962 sw
rect 55586 34880 55679 34946
rect 55715 34821 55829 34979
tri 55865 34946 55881 34962 se
rect 55881 34946 55958 34962
rect 55865 34880 55958 34946
rect 55586 34745 55958 34821
rect 55586 34620 55679 34686
rect 55586 34604 55663 34620
tri 55663 34604 55679 34620 nw
rect 55715 34587 55829 34745
rect 55865 34620 55958 34686
tri 55865 34604 55881 34620 ne
rect 55881 34604 55958 34620
rect 55698 34505 55846 34587
rect 55586 34472 55663 34488
tri 55663 34472 55679 34488 sw
rect 55586 34406 55679 34472
rect 55586 34304 55679 34370
rect 55586 34288 55663 34304
tri 55663 34288 55679 34304 nw
rect 55715 34271 55829 34505
tri 55865 34472 55881 34488 se
rect 55881 34472 55958 34488
rect 55865 34406 55958 34472
rect 55865 34304 55958 34370
tri 55865 34288 55881 34304 ne
rect 55881 34288 55958 34304
rect 55698 34189 55846 34271
rect 55586 34156 55663 34172
tri 55663 34156 55679 34172 sw
rect 55586 34090 55679 34156
rect 55715 34031 55829 34189
tri 55865 34156 55881 34172 se
rect 55881 34156 55958 34172
rect 55865 34090 55958 34156
rect 55586 33955 55958 34031
rect 55586 33830 55679 33896
rect 55586 33814 55663 33830
tri 55663 33814 55679 33830 nw
rect 55715 33797 55829 33955
rect 55865 33830 55958 33896
tri 55865 33814 55881 33830 ne
rect 55881 33814 55958 33830
rect 55698 33715 55846 33797
rect 55586 33682 55663 33698
tri 55663 33682 55679 33698 sw
rect 55586 33616 55679 33682
rect 55586 33514 55679 33580
rect 55586 33498 55663 33514
tri 55663 33498 55679 33514 nw
rect 55715 33481 55829 33715
tri 55865 33682 55881 33698 se
rect 55881 33682 55958 33698
rect 55865 33616 55958 33682
rect 55865 33514 55958 33580
tri 55865 33498 55881 33514 ne
rect 55881 33498 55958 33514
rect 55698 33399 55846 33481
rect 55586 33366 55663 33382
tri 55663 33366 55679 33382 sw
rect 55586 33300 55679 33366
rect 55715 33241 55829 33399
tri 55865 33366 55881 33382 se
rect 55881 33366 55958 33382
rect 55865 33300 55958 33366
rect 55586 33165 55958 33241
rect 55586 33040 55679 33106
rect 55586 33024 55663 33040
tri 55663 33024 55679 33040 nw
rect 55715 33007 55829 33165
rect 55865 33040 55958 33106
tri 55865 33024 55881 33040 ne
rect 55881 33024 55958 33040
rect 55698 32925 55846 33007
rect 55586 32892 55663 32908
tri 55663 32892 55679 32908 sw
rect 55586 32826 55679 32892
rect 55586 32724 55679 32790
rect 55586 32708 55663 32724
tri 55663 32708 55679 32724 nw
rect 55715 32691 55829 32925
tri 55865 32892 55881 32908 se
rect 55881 32892 55958 32908
rect 55865 32826 55958 32892
rect 55865 32724 55958 32790
tri 55865 32708 55881 32724 ne
rect 55881 32708 55958 32724
rect 55698 32609 55846 32691
rect 55586 32576 55663 32592
tri 55663 32576 55679 32592 sw
rect 55586 32510 55679 32576
rect 55715 32451 55829 32609
tri 55865 32576 55881 32592 se
rect 55881 32576 55958 32592
rect 55865 32510 55958 32576
rect 55586 32375 55958 32451
rect 55586 32250 55679 32316
rect 55586 32234 55663 32250
tri 55663 32234 55679 32250 nw
rect 55715 32217 55829 32375
rect 55865 32250 55958 32316
tri 55865 32234 55881 32250 ne
rect 55881 32234 55958 32250
rect 55698 32135 55846 32217
rect 55586 32102 55663 32118
tri 55663 32102 55679 32118 sw
rect 55586 32036 55679 32102
rect 55586 31934 55679 32000
rect 55586 31918 55663 31934
tri 55663 31918 55679 31934 nw
rect 55715 31901 55829 32135
tri 55865 32102 55881 32118 se
rect 55881 32102 55958 32118
rect 55865 32036 55958 32102
rect 55865 31934 55958 32000
tri 55865 31918 55881 31934 ne
rect 55881 31918 55958 31934
rect 55698 31819 55846 31901
rect 55586 31786 55663 31802
tri 55663 31786 55679 31802 sw
rect 55586 31720 55679 31786
rect 55715 31661 55829 31819
tri 55865 31786 55881 31802 se
rect 55881 31786 55958 31802
rect 55865 31720 55958 31786
rect 55586 31585 55958 31661
rect 55586 31460 55679 31526
rect 55586 31444 55663 31460
tri 55663 31444 55679 31460 nw
rect 55715 31427 55829 31585
rect 55865 31460 55958 31526
tri 55865 31444 55881 31460 ne
rect 55881 31444 55958 31460
rect 55698 31345 55846 31427
rect 55586 31312 55663 31328
tri 55663 31312 55679 31328 sw
rect 55586 31246 55679 31312
rect 55586 31144 55679 31210
rect 55586 31128 55663 31144
tri 55663 31128 55679 31144 nw
rect 55715 31111 55829 31345
tri 55865 31312 55881 31328 se
rect 55881 31312 55958 31328
rect 55865 31246 55958 31312
rect 55865 31144 55958 31210
tri 55865 31128 55881 31144 ne
rect 55881 31128 55958 31144
rect 55698 31029 55846 31111
rect 55586 30996 55663 31012
tri 55663 30996 55679 31012 sw
rect 55586 30930 55679 30996
rect 55715 30871 55829 31029
tri 55865 30996 55881 31012 se
rect 55881 30996 55958 31012
rect 55865 30930 55958 30996
rect 55586 30795 55958 30871
rect 55586 30670 55679 30736
rect 55586 30654 55663 30670
tri 55663 30654 55679 30670 nw
rect 55715 30637 55829 30795
rect 55865 30670 55958 30736
tri 55865 30654 55881 30670 ne
rect 55881 30654 55958 30670
rect 55698 30555 55846 30637
rect 55586 30522 55663 30538
tri 55663 30522 55679 30538 sw
rect 55586 30456 55679 30522
rect 55586 30354 55679 30420
rect 55586 30338 55663 30354
tri 55663 30338 55679 30354 nw
rect 55715 30321 55829 30555
tri 55865 30522 55881 30538 se
rect 55881 30522 55958 30538
rect 55865 30456 55958 30522
rect 55865 30354 55958 30420
tri 55865 30338 55881 30354 ne
rect 55881 30338 55958 30354
rect 55698 30239 55846 30321
rect 55586 30206 55663 30222
tri 55663 30206 55679 30222 sw
rect 55586 30140 55679 30206
rect 55715 30081 55829 30239
tri 55865 30206 55881 30222 se
rect 55881 30206 55958 30222
rect 55865 30140 55958 30206
rect 55586 30005 55958 30081
rect 55586 29880 55679 29946
rect 55586 29864 55663 29880
tri 55663 29864 55679 29880 nw
rect 55715 29847 55829 30005
rect 55865 29880 55958 29946
tri 55865 29864 55881 29880 ne
rect 55881 29864 55958 29880
rect 55698 29765 55846 29847
rect 55586 29732 55663 29748
tri 55663 29732 55679 29748 sw
rect 55586 29666 55679 29732
rect 55586 29564 55679 29630
rect 55586 29548 55663 29564
tri 55663 29548 55679 29564 nw
rect 55715 29531 55829 29765
tri 55865 29732 55881 29748 se
rect 55881 29732 55958 29748
rect 55865 29666 55958 29732
rect 55865 29564 55958 29630
tri 55865 29548 55881 29564 ne
rect 55881 29548 55958 29564
rect 55698 29449 55846 29531
rect 55586 29416 55663 29432
tri 55663 29416 55679 29432 sw
rect 55586 29350 55679 29416
rect 55715 29291 55829 29449
tri 55865 29416 55881 29432 se
rect 55881 29416 55958 29432
rect 55865 29350 55958 29416
rect 55586 29215 55958 29291
rect 55586 29090 55679 29156
rect 55586 29074 55663 29090
tri 55663 29074 55679 29090 nw
rect 55715 29057 55829 29215
rect 55865 29090 55958 29156
tri 55865 29074 55881 29090 ne
rect 55881 29074 55958 29090
rect 55698 28975 55846 29057
rect 55586 28942 55663 28958
tri 55663 28942 55679 28958 sw
rect 55586 28876 55679 28942
rect 55715 28833 55829 28975
tri 55865 28942 55881 28958 se
rect 55881 28942 55958 28958
rect 55865 28876 55958 28942
rect 55994 28463 56030 80603
rect 56066 28463 56102 80603
rect 56138 80445 56174 80603
rect 56130 80303 56182 80445
rect 56138 28763 56174 80303
rect 56130 28621 56182 28763
rect 56138 28463 56174 28621
rect 56210 28463 56246 80603
rect 56282 28463 56318 80603
rect 56354 28833 56438 80233
rect 56474 28463 56510 80603
rect 56546 28463 56582 80603
rect 56618 80445 56654 80603
rect 56610 80303 56662 80445
rect 56618 28763 56654 80303
rect 56610 28621 56662 28763
rect 56618 28463 56654 28621
rect 56690 28463 56726 80603
rect 56762 28463 56798 80603
rect 56834 80124 56927 80190
rect 56834 80108 56911 80124
tri 56911 80108 56927 80124 nw
rect 56963 80091 57077 80233
rect 57113 80124 57206 80190
tri 57113 80108 57129 80124 ne
rect 57129 80108 57206 80124
rect 56946 80009 57094 80091
rect 56834 79976 56911 79992
tri 56911 79976 56927 79992 sw
rect 56834 79910 56927 79976
rect 56963 79851 57077 80009
tri 57113 79976 57129 79992 se
rect 57129 79976 57206 79992
rect 57113 79910 57206 79976
rect 56834 79775 57206 79851
rect 56834 79650 56927 79716
rect 56834 79634 56911 79650
tri 56911 79634 56927 79650 nw
rect 56963 79617 57077 79775
rect 57113 79650 57206 79716
tri 57113 79634 57129 79650 ne
rect 57129 79634 57206 79650
rect 56946 79535 57094 79617
rect 56834 79502 56911 79518
tri 56911 79502 56927 79518 sw
rect 56834 79436 56927 79502
rect 56834 79334 56927 79400
rect 56834 79318 56911 79334
tri 56911 79318 56927 79334 nw
rect 56963 79301 57077 79535
tri 57113 79502 57129 79518 se
rect 57129 79502 57206 79518
rect 57113 79436 57206 79502
rect 57113 79334 57206 79400
tri 57113 79318 57129 79334 ne
rect 57129 79318 57206 79334
rect 56946 79219 57094 79301
rect 56834 79186 56911 79202
tri 56911 79186 56927 79202 sw
rect 56834 79120 56927 79186
rect 56963 79061 57077 79219
tri 57113 79186 57129 79202 se
rect 57129 79186 57206 79202
rect 57113 79120 57206 79186
rect 56834 78985 57206 79061
rect 56834 78860 56927 78926
rect 56834 78844 56911 78860
tri 56911 78844 56927 78860 nw
rect 56963 78827 57077 78985
rect 57113 78860 57206 78926
tri 57113 78844 57129 78860 ne
rect 57129 78844 57206 78860
rect 56946 78745 57094 78827
rect 56834 78712 56911 78728
tri 56911 78712 56927 78728 sw
rect 56834 78646 56927 78712
rect 56834 78544 56927 78610
rect 56834 78528 56911 78544
tri 56911 78528 56927 78544 nw
rect 56963 78511 57077 78745
tri 57113 78712 57129 78728 se
rect 57129 78712 57206 78728
rect 57113 78646 57206 78712
rect 57113 78544 57206 78610
tri 57113 78528 57129 78544 ne
rect 57129 78528 57206 78544
rect 56946 78429 57094 78511
rect 56834 78396 56911 78412
tri 56911 78396 56927 78412 sw
rect 56834 78330 56927 78396
rect 56963 78271 57077 78429
tri 57113 78396 57129 78412 se
rect 57129 78396 57206 78412
rect 57113 78330 57206 78396
rect 56834 78195 57206 78271
rect 56834 78070 56927 78136
rect 56834 78054 56911 78070
tri 56911 78054 56927 78070 nw
rect 56963 78037 57077 78195
rect 57113 78070 57206 78136
tri 57113 78054 57129 78070 ne
rect 57129 78054 57206 78070
rect 56946 77955 57094 78037
rect 56834 77922 56911 77938
tri 56911 77922 56927 77938 sw
rect 56834 77856 56927 77922
rect 56834 77754 56927 77820
rect 56834 77738 56911 77754
tri 56911 77738 56927 77754 nw
rect 56963 77721 57077 77955
tri 57113 77922 57129 77938 se
rect 57129 77922 57206 77938
rect 57113 77856 57206 77922
rect 57113 77754 57206 77820
tri 57113 77738 57129 77754 ne
rect 57129 77738 57206 77754
rect 56946 77639 57094 77721
rect 56834 77606 56911 77622
tri 56911 77606 56927 77622 sw
rect 56834 77540 56927 77606
rect 56963 77481 57077 77639
tri 57113 77606 57129 77622 se
rect 57129 77606 57206 77622
rect 57113 77540 57206 77606
rect 56834 77405 57206 77481
rect 56834 77280 56927 77346
rect 56834 77264 56911 77280
tri 56911 77264 56927 77280 nw
rect 56963 77247 57077 77405
rect 57113 77280 57206 77346
tri 57113 77264 57129 77280 ne
rect 57129 77264 57206 77280
rect 56946 77165 57094 77247
rect 56834 77132 56911 77148
tri 56911 77132 56927 77148 sw
rect 56834 77066 56927 77132
rect 56834 76964 56927 77030
rect 56834 76948 56911 76964
tri 56911 76948 56927 76964 nw
rect 56963 76931 57077 77165
tri 57113 77132 57129 77148 se
rect 57129 77132 57206 77148
rect 57113 77066 57206 77132
rect 57113 76964 57206 77030
tri 57113 76948 57129 76964 ne
rect 57129 76948 57206 76964
rect 56946 76849 57094 76931
rect 56834 76816 56911 76832
tri 56911 76816 56927 76832 sw
rect 56834 76750 56927 76816
rect 56963 76691 57077 76849
tri 57113 76816 57129 76832 se
rect 57129 76816 57206 76832
rect 57113 76750 57206 76816
rect 56834 76615 57206 76691
rect 56834 76490 56927 76556
rect 56834 76474 56911 76490
tri 56911 76474 56927 76490 nw
rect 56963 76457 57077 76615
rect 57113 76490 57206 76556
tri 57113 76474 57129 76490 ne
rect 57129 76474 57206 76490
rect 56946 76375 57094 76457
rect 56834 76342 56911 76358
tri 56911 76342 56927 76358 sw
rect 56834 76276 56927 76342
rect 56834 76174 56927 76240
rect 56834 76158 56911 76174
tri 56911 76158 56927 76174 nw
rect 56963 76141 57077 76375
tri 57113 76342 57129 76358 se
rect 57129 76342 57206 76358
rect 57113 76276 57206 76342
rect 57113 76174 57206 76240
tri 57113 76158 57129 76174 ne
rect 57129 76158 57206 76174
rect 56946 76059 57094 76141
rect 56834 76026 56911 76042
tri 56911 76026 56927 76042 sw
rect 56834 75960 56927 76026
rect 56963 75901 57077 76059
tri 57113 76026 57129 76042 se
rect 57129 76026 57206 76042
rect 57113 75960 57206 76026
rect 56834 75825 57206 75901
rect 56834 75700 56927 75766
rect 56834 75684 56911 75700
tri 56911 75684 56927 75700 nw
rect 56963 75667 57077 75825
rect 57113 75700 57206 75766
tri 57113 75684 57129 75700 ne
rect 57129 75684 57206 75700
rect 56946 75585 57094 75667
rect 56834 75552 56911 75568
tri 56911 75552 56927 75568 sw
rect 56834 75486 56927 75552
rect 56834 75384 56927 75450
rect 56834 75368 56911 75384
tri 56911 75368 56927 75384 nw
rect 56963 75351 57077 75585
tri 57113 75552 57129 75568 se
rect 57129 75552 57206 75568
rect 57113 75486 57206 75552
rect 57113 75384 57206 75450
tri 57113 75368 57129 75384 ne
rect 57129 75368 57206 75384
rect 56946 75269 57094 75351
rect 56834 75236 56911 75252
tri 56911 75236 56927 75252 sw
rect 56834 75170 56927 75236
rect 56963 75111 57077 75269
tri 57113 75236 57129 75252 se
rect 57129 75236 57206 75252
rect 57113 75170 57206 75236
rect 56834 75035 57206 75111
rect 56834 74910 56927 74976
rect 56834 74894 56911 74910
tri 56911 74894 56927 74910 nw
rect 56963 74877 57077 75035
rect 57113 74910 57206 74976
tri 57113 74894 57129 74910 ne
rect 57129 74894 57206 74910
rect 56946 74795 57094 74877
rect 56834 74762 56911 74778
tri 56911 74762 56927 74778 sw
rect 56834 74696 56927 74762
rect 56834 74594 56927 74660
rect 56834 74578 56911 74594
tri 56911 74578 56927 74594 nw
rect 56963 74561 57077 74795
tri 57113 74762 57129 74778 se
rect 57129 74762 57206 74778
rect 57113 74696 57206 74762
rect 57113 74594 57206 74660
tri 57113 74578 57129 74594 ne
rect 57129 74578 57206 74594
rect 56946 74479 57094 74561
rect 56834 74446 56911 74462
tri 56911 74446 56927 74462 sw
rect 56834 74380 56927 74446
rect 56963 74321 57077 74479
tri 57113 74446 57129 74462 se
rect 57129 74446 57206 74462
rect 57113 74380 57206 74446
rect 56834 74245 57206 74321
rect 56834 74120 56927 74186
rect 56834 74104 56911 74120
tri 56911 74104 56927 74120 nw
rect 56963 74087 57077 74245
rect 57113 74120 57206 74186
tri 57113 74104 57129 74120 ne
rect 57129 74104 57206 74120
rect 56946 74005 57094 74087
rect 56834 73972 56911 73988
tri 56911 73972 56927 73988 sw
rect 56834 73906 56927 73972
rect 56834 73804 56927 73870
rect 56834 73788 56911 73804
tri 56911 73788 56927 73804 nw
rect 56963 73771 57077 74005
tri 57113 73972 57129 73988 se
rect 57129 73972 57206 73988
rect 57113 73906 57206 73972
rect 57113 73804 57206 73870
tri 57113 73788 57129 73804 ne
rect 57129 73788 57206 73804
rect 56946 73689 57094 73771
rect 56834 73656 56911 73672
tri 56911 73656 56927 73672 sw
rect 56834 73590 56927 73656
rect 56963 73531 57077 73689
tri 57113 73656 57129 73672 se
rect 57129 73656 57206 73672
rect 57113 73590 57206 73656
rect 56834 73455 57206 73531
rect 56834 73330 56927 73396
rect 56834 73314 56911 73330
tri 56911 73314 56927 73330 nw
rect 56963 73297 57077 73455
rect 57113 73330 57206 73396
tri 57113 73314 57129 73330 ne
rect 57129 73314 57206 73330
rect 56946 73215 57094 73297
rect 56834 73182 56911 73198
tri 56911 73182 56927 73198 sw
rect 56834 73116 56927 73182
rect 56834 73014 56927 73080
rect 56834 72998 56911 73014
tri 56911 72998 56927 73014 nw
rect 56963 72981 57077 73215
tri 57113 73182 57129 73198 se
rect 57129 73182 57206 73198
rect 57113 73116 57206 73182
rect 57113 73014 57206 73080
tri 57113 72998 57129 73014 ne
rect 57129 72998 57206 73014
rect 56946 72899 57094 72981
rect 56834 72866 56911 72882
tri 56911 72866 56927 72882 sw
rect 56834 72800 56927 72866
rect 56963 72741 57077 72899
tri 57113 72866 57129 72882 se
rect 57129 72866 57206 72882
rect 57113 72800 57206 72866
rect 56834 72665 57206 72741
rect 56834 72540 56927 72606
rect 56834 72524 56911 72540
tri 56911 72524 56927 72540 nw
rect 56963 72507 57077 72665
rect 57113 72540 57206 72606
tri 57113 72524 57129 72540 ne
rect 57129 72524 57206 72540
rect 56946 72425 57094 72507
rect 56834 72392 56911 72408
tri 56911 72392 56927 72408 sw
rect 56834 72326 56927 72392
rect 56834 72224 56927 72290
rect 56834 72208 56911 72224
tri 56911 72208 56927 72224 nw
rect 56963 72191 57077 72425
tri 57113 72392 57129 72408 se
rect 57129 72392 57206 72408
rect 57113 72326 57206 72392
rect 57113 72224 57206 72290
tri 57113 72208 57129 72224 ne
rect 57129 72208 57206 72224
rect 56946 72109 57094 72191
rect 56834 72076 56911 72092
tri 56911 72076 56927 72092 sw
rect 56834 72010 56927 72076
rect 56963 71951 57077 72109
tri 57113 72076 57129 72092 se
rect 57129 72076 57206 72092
rect 57113 72010 57206 72076
rect 56834 71875 57206 71951
rect 56834 71750 56927 71816
rect 56834 71734 56911 71750
tri 56911 71734 56927 71750 nw
rect 56963 71717 57077 71875
rect 57113 71750 57206 71816
tri 57113 71734 57129 71750 ne
rect 57129 71734 57206 71750
rect 56946 71635 57094 71717
rect 56834 71602 56911 71618
tri 56911 71602 56927 71618 sw
rect 56834 71536 56927 71602
rect 56834 71434 56927 71500
rect 56834 71418 56911 71434
tri 56911 71418 56927 71434 nw
rect 56963 71401 57077 71635
tri 57113 71602 57129 71618 se
rect 57129 71602 57206 71618
rect 57113 71536 57206 71602
rect 57113 71434 57206 71500
tri 57113 71418 57129 71434 ne
rect 57129 71418 57206 71434
rect 56946 71319 57094 71401
rect 56834 71286 56911 71302
tri 56911 71286 56927 71302 sw
rect 56834 71220 56927 71286
rect 56963 71161 57077 71319
tri 57113 71286 57129 71302 se
rect 57129 71286 57206 71302
rect 57113 71220 57206 71286
rect 56834 71085 57206 71161
rect 56834 70960 56927 71026
rect 56834 70944 56911 70960
tri 56911 70944 56927 70960 nw
rect 56963 70927 57077 71085
rect 57113 70960 57206 71026
tri 57113 70944 57129 70960 ne
rect 57129 70944 57206 70960
rect 56946 70845 57094 70927
rect 56834 70812 56911 70828
tri 56911 70812 56927 70828 sw
rect 56834 70746 56927 70812
rect 56834 70644 56927 70710
rect 56834 70628 56911 70644
tri 56911 70628 56927 70644 nw
rect 56963 70611 57077 70845
tri 57113 70812 57129 70828 se
rect 57129 70812 57206 70828
rect 57113 70746 57206 70812
rect 57113 70644 57206 70710
tri 57113 70628 57129 70644 ne
rect 57129 70628 57206 70644
rect 56946 70529 57094 70611
rect 56834 70496 56911 70512
tri 56911 70496 56927 70512 sw
rect 56834 70430 56927 70496
rect 56963 70371 57077 70529
tri 57113 70496 57129 70512 se
rect 57129 70496 57206 70512
rect 57113 70430 57206 70496
rect 56834 70295 57206 70371
rect 56834 70170 56927 70236
rect 56834 70154 56911 70170
tri 56911 70154 56927 70170 nw
rect 56963 70137 57077 70295
rect 57113 70170 57206 70236
tri 57113 70154 57129 70170 ne
rect 57129 70154 57206 70170
rect 56946 70055 57094 70137
rect 56834 70022 56911 70038
tri 56911 70022 56927 70038 sw
rect 56834 69956 56927 70022
rect 56834 69854 56927 69920
rect 56834 69838 56911 69854
tri 56911 69838 56927 69854 nw
rect 56963 69821 57077 70055
tri 57113 70022 57129 70038 se
rect 57129 70022 57206 70038
rect 57113 69956 57206 70022
rect 57113 69854 57206 69920
tri 57113 69838 57129 69854 ne
rect 57129 69838 57206 69854
rect 56946 69739 57094 69821
rect 56834 69706 56911 69722
tri 56911 69706 56927 69722 sw
rect 56834 69640 56927 69706
rect 56963 69581 57077 69739
tri 57113 69706 57129 69722 se
rect 57129 69706 57206 69722
rect 57113 69640 57206 69706
rect 56834 69505 57206 69581
rect 56834 69380 56927 69446
rect 56834 69364 56911 69380
tri 56911 69364 56927 69380 nw
rect 56963 69347 57077 69505
rect 57113 69380 57206 69446
tri 57113 69364 57129 69380 ne
rect 57129 69364 57206 69380
rect 56946 69265 57094 69347
rect 56834 69232 56911 69248
tri 56911 69232 56927 69248 sw
rect 56834 69166 56927 69232
rect 56834 69064 56927 69130
rect 56834 69048 56911 69064
tri 56911 69048 56927 69064 nw
rect 56963 69031 57077 69265
tri 57113 69232 57129 69248 se
rect 57129 69232 57206 69248
rect 57113 69166 57206 69232
rect 57113 69064 57206 69130
tri 57113 69048 57129 69064 ne
rect 57129 69048 57206 69064
rect 56946 68949 57094 69031
rect 56834 68916 56911 68932
tri 56911 68916 56927 68932 sw
rect 56834 68850 56927 68916
rect 56963 68791 57077 68949
tri 57113 68916 57129 68932 se
rect 57129 68916 57206 68932
rect 57113 68850 57206 68916
rect 56834 68715 57206 68791
rect 56834 68590 56927 68656
rect 56834 68574 56911 68590
tri 56911 68574 56927 68590 nw
rect 56963 68557 57077 68715
rect 57113 68590 57206 68656
tri 57113 68574 57129 68590 ne
rect 57129 68574 57206 68590
rect 56946 68475 57094 68557
rect 56834 68442 56911 68458
tri 56911 68442 56927 68458 sw
rect 56834 68376 56927 68442
rect 56834 68274 56927 68340
rect 56834 68258 56911 68274
tri 56911 68258 56927 68274 nw
rect 56963 68241 57077 68475
tri 57113 68442 57129 68458 se
rect 57129 68442 57206 68458
rect 57113 68376 57206 68442
rect 57113 68274 57206 68340
tri 57113 68258 57129 68274 ne
rect 57129 68258 57206 68274
rect 56946 68159 57094 68241
rect 56834 68126 56911 68142
tri 56911 68126 56927 68142 sw
rect 56834 68060 56927 68126
rect 56963 68001 57077 68159
tri 57113 68126 57129 68142 se
rect 57129 68126 57206 68142
rect 57113 68060 57206 68126
rect 56834 67925 57206 68001
rect 56834 67800 56927 67866
rect 56834 67784 56911 67800
tri 56911 67784 56927 67800 nw
rect 56963 67767 57077 67925
rect 57113 67800 57206 67866
tri 57113 67784 57129 67800 ne
rect 57129 67784 57206 67800
rect 56946 67685 57094 67767
rect 56834 67652 56911 67668
tri 56911 67652 56927 67668 sw
rect 56834 67586 56927 67652
rect 56834 67484 56927 67550
rect 56834 67468 56911 67484
tri 56911 67468 56927 67484 nw
rect 56963 67451 57077 67685
tri 57113 67652 57129 67668 se
rect 57129 67652 57206 67668
rect 57113 67586 57206 67652
rect 57113 67484 57206 67550
tri 57113 67468 57129 67484 ne
rect 57129 67468 57206 67484
rect 56946 67369 57094 67451
rect 56834 67336 56911 67352
tri 56911 67336 56927 67352 sw
rect 56834 67270 56927 67336
rect 56963 67211 57077 67369
tri 57113 67336 57129 67352 se
rect 57129 67336 57206 67352
rect 57113 67270 57206 67336
rect 56834 67135 57206 67211
rect 56834 67010 56927 67076
rect 56834 66994 56911 67010
tri 56911 66994 56927 67010 nw
rect 56963 66977 57077 67135
rect 57113 67010 57206 67076
tri 57113 66994 57129 67010 ne
rect 57129 66994 57206 67010
rect 56946 66895 57094 66977
rect 56834 66862 56911 66878
tri 56911 66862 56927 66878 sw
rect 56834 66796 56927 66862
rect 56834 66694 56927 66760
rect 56834 66678 56911 66694
tri 56911 66678 56927 66694 nw
rect 56963 66661 57077 66895
tri 57113 66862 57129 66878 se
rect 57129 66862 57206 66878
rect 57113 66796 57206 66862
rect 57113 66694 57206 66760
tri 57113 66678 57129 66694 ne
rect 57129 66678 57206 66694
rect 56946 66579 57094 66661
rect 56834 66546 56911 66562
tri 56911 66546 56927 66562 sw
rect 56834 66480 56927 66546
rect 56963 66421 57077 66579
tri 57113 66546 57129 66562 se
rect 57129 66546 57206 66562
rect 57113 66480 57206 66546
rect 56834 66345 57206 66421
rect 56834 66220 56927 66286
rect 56834 66204 56911 66220
tri 56911 66204 56927 66220 nw
rect 56963 66187 57077 66345
rect 57113 66220 57206 66286
tri 57113 66204 57129 66220 ne
rect 57129 66204 57206 66220
rect 56946 66105 57094 66187
rect 56834 66072 56911 66088
tri 56911 66072 56927 66088 sw
rect 56834 66006 56927 66072
rect 56834 65904 56927 65970
rect 56834 65888 56911 65904
tri 56911 65888 56927 65904 nw
rect 56963 65871 57077 66105
tri 57113 66072 57129 66088 se
rect 57129 66072 57206 66088
rect 57113 66006 57206 66072
rect 57113 65904 57206 65970
tri 57113 65888 57129 65904 ne
rect 57129 65888 57206 65904
rect 56946 65789 57094 65871
rect 56834 65756 56911 65772
tri 56911 65756 56927 65772 sw
rect 56834 65690 56927 65756
rect 56963 65631 57077 65789
tri 57113 65756 57129 65772 se
rect 57129 65756 57206 65772
rect 57113 65690 57206 65756
rect 56834 65555 57206 65631
rect 56834 65430 56927 65496
rect 56834 65414 56911 65430
tri 56911 65414 56927 65430 nw
rect 56963 65397 57077 65555
rect 57113 65430 57206 65496
tri 57113 65414 57129 65430 ne
rect 57129 65414 57206 65430
rect 56946 65315 57094 65397
rect 56834 65282 56911 65298
tri 56911 65282 56927 65298 sw
rect 56834 65216 56927 65282
rect 56834 65114 56927 65180
rect 56834 65098 56911 65114
tri 56911 65098 56927 65114 nw
rect 56963 65081 57077 65315
tri 57113 65282 57129 65298 se
rect 57129 65282 57206 65298
rect 57113 65216 57206 65282
rect 57113 65114 57206 65180
tri 57113 65098 57129 65114 ne
rect 57129 65098 57206 65114
rect 56946 64999 57094 65081
rect 56834 64966 56911 64982
tri 56911 64966 56927 64982 sw
rect 56834 64900 56927 64966
rect 56963 64841 57077 64999
tri 57113 64966 57129 64982 se
rect 57129 64966 57206 64982
rect 57113 64900 57206 64966
rect 56834 64765 57206 64841
rect 56834 64640 56927 64706
rect 56834 64624 56911 64640
tri 56911 64624 56927 64640 nw
rect 56963 64607 57077 64765
rect 57113 64640 57206 64706
tri 57113 64624 57129 64640 ne
rect 57129 64624 57206 64640
rect 56946 64525 57094 64607
rect 56834 64492 56911 64508
tri 56911 64492 56927 64508 sw
rect 56834 64426 56927 64492
rect 56834 64324 56927 64390
rect 56834 64308 56911 64324
tri 56911 64308 56927 64324 nw
rect 56963 64291 57077 64525
tri 57113 64492 57129 64508 se
rect 57129 64492 57206 64508
rect 57113 64426 57206 64492
rect 57113 64324 57206 64390
tri 57113 64308 57129 64324 ne
rect 57129 64308 57206 64324
rect 56946 64209 57094 64291
rect 56834 64176 56911 64192
tri 56911 64176 56927 64192 sw
rect 56834 64110 56927 64176
rect 56963 64051 57077 64209
tri 57113 64176 57129 64192 se
rect 57129 64176 57206 64192
rect 57113 64110 57206 64176
rect 56834 63975 57206 64051
rect 56834 63850 56927 63916
rect 56834 63834 56911 63850
tri 56911 63834 56927 63850 nw
rect 56963 63817 57077 63975
rect 57113 63850 57206 63916
tri 57113 63834 57129 63850 ne
rect 57129 63834 57206 63850
rect 56946 63735 57094 63817
rect 56834 63702 56911 63718
tri 56911 63702 56927 63718 sw
rect 56834 63636 56927 63702
rect 56834 63534 56927 63600
rect 56834 63518 56911 63534
tri 56911 63518 56927 63534 nw
rect 56963 63501 57077 63735
tri 57113 63702 57129 63718 se
rect 57129 63702 57206 63718
rect 57113 63636 57206 63702
rect 57113 63534 57206 63600
tri 57113 63518 57129 63534 ne
rect 57129 63518 57206 63534
rect 56946 63419 57094 63501
rect 56834 63386 56911 63402
tri 56911 63386 56927 63402 sw
rect 56834 63320 56927 63386
rect 56963 63261 57077 63419
tri 57113 63386 57129 63402 se
rect 57129 63386 57206 63402
rect 57113 63320 57206 63386
rect 56834 63185 57206 63261
rect 56834 63060 56927 63126
rect 56834 63044 56911 63060
tri 56911 63044 56927 63060 nw
rect 56963 63027 57077 63185
rect 57113 63060 57206 63126
tri 57113 63044 57129 63060 ne
rect 57129 63044 57206 63060
rect 56946 62945 57094 63027
rect 56834 62912 56911 62928
tri 56911 62912 56927 62928 sw
rect 56834 62846 56927 62912
rect 56834 62744 56927 62810
rect 56834 62728 56911 62744
tri 56911 62728 56927 62744 nw
rect 56963 62711 57077 62945
tri 57113 62912 57129 62928 se
rect 57129 62912 57206 62928
rect 57113 62846 57206 62912
rect 57113 62744 57206 62810
tri 57113 62728 57129 62744 ne
rect 57129 62728 57206 62744
rect 56946 62629 57094 62711
rect 56834 62596 56911 62612
tri 56911 62596 56927 62612 sw
rect 56834 62530 56927 62596
rect 56963 62471 57077 62629
tri 57113 62596 57129 62612 se
rect 57129 62596 57206 62612
rect 57113 62530 57206 62596
rect 56834 62395 57206 62471
rect 56834 62270 56927 62336
rect 56834 62254 56911 62270
tri 56911 62254 56927 62270 nw
rect 56963 62237 57077 62395
rect 57113 62270 57206 62336
tri 57113 62254 57129 62270 ne
rect 57129 62254 57206 62270
rect 56946 62155 57094 62237
rect 56834 62122 56911 62138
tri 56911 62122 56927 62138 sw
rect 56834 62056 56927 62122
rect 56834 61954 56927 62020
rect 56834 61938 56911 61954
tri 56911 61938 56927 61954 nw
rect 56963 61921 57077 62155
tri 57113 62122 57129 62138 se
rect 57129 62122 57206 62138
rect 57113 62056 57206 62122
rect 57113 61954 57206 62020
tri 57113 61938 57129 61954 ne
rect 57129 61938 57206 61954
rect 56946 61839 57094 61921
rect 56834 61806 56911 61822
tri 56911 61806 56927 61822 sw
rect 56834 61740 56927 61806
rect 56963 61681 57077 61839
tri 57113 61806 57129 61822 se
rect 57129 61806 57206 61822
rect 57113 61740 57206 61806
rect 56834 61605 57206 61681
rect 56834 61480 56927 61546
rect 56834 61464 56911 61480
tri 56911 61464 56927 61480 nw
rect 56963 61447 57077 61605
rect 57113 61480 57206 61546
tri 57113 61464 57129 61480 ne
rect 57129 61464 57206 61480
rect 56946 61365 57094 61447
rect 56834 61332 56911 61348
tri 56911 61332 56927 61348 sw
rect 56834 61266 56927 61332
rect 56834 61164 56927 61230
rect 56834 61148 56911 61164
tri 56911 61148 56927 61164 nw
rect 56963 61131 57077 61365
tri 57113 61332 57129 61348 se
rect 57129 61332 57206 61348
rect 57113 61266 57206 61332
rect 57113 61164 57206 61230
tri 57113 61148 57129 61164 ne
rect 57129 61148 57206 61164
rect 56946 61049 57094 61131
rect 56834 61016 56911 61032
tri 56911 61016 56927 61032 sw
rect 56834 60950 56927 61016
rect 56963 60891 57077 61049
tri 57113 61016 57129 61032 se
rect 57129 61016 57206 61032
rect 57113 60950 57206 61016
rect 56834 60815 57206 60891
rect 56834 60690 56927 60756
rect 56834 60674 56911 60690
tri 56911 60674 56927 60690 nw
rect 56963 60657 57077 60815
rect 57113 60690 57206 60756
tri 57113 60674 57129 60690 ne
rect 57129 60674 57206 60690
rect 56946 60575 57094 60657
rect 56834 60542 56911 60558
tri 56911 60542 56927 60558 sw
rect 56834 60476 56927 60542
rect 56834 60374 56927 60440
rect 56834 60358 56911 60374
tri 56911 60358 56927 60374 nw
rect 56963 60341 57077 60575
tri 57113 60542 57129 60558 se
rect 57129 60542 57206 60558
rect 57113 60476 57206 60542
rect 57113 60374 57206 60440
tri 57113 60358 57129 60374 ne
rect 57129 60358 57206 60374
rect 56946 60259 57094 60341
rect 56834 60226 56911 60242
tri 56911 60226 56927 60242 sw
rect 56834 60160 56927 60226
rect 56963 60101 57077 60259
tri 57113 60226 57129 60242 se
rect 57129 60226 57206 60242
rect 57113 60160 57206 60226
rect 56834 60025 57206 60101
rect 56834 59900 56927 59966
rect 56834 59884 56911 59900
tri 56911 59884 56927 59900 nw
rect 56963 59867 57077 60025
rect 57113 59900 57206 59966
tri 57113 59884 57129 59900 ne
rect 57129 59884 57206 59900
rect 56946 59785 57094 59867
rect 56834 59752 56911 59768
tri 56911 59752 56927 59768 sw
rect 56834 59686 56927 59752
rect 56834 59584 56927 59650
rect 56834 59568 56911 59584
tri 56911 59568 56927 59584 nw
rect 56963 59551 57077 59785
tri 57113 59752 57129 59768 se
rect 57129 59752 57206 59768
rect 57113 59686 57206 59752
rect 57113 59584 57206 59650
tri 57113 59568 57129 59584 ne
rect 57129 59568 57206 59584
rect 56946 59469 57094 59551
rect 56834 59436 56911 59452
tri 56911 59436 56927 59452 sw
rect 56834 59370 56927 59436
rect 56963 59311 57077 59469
tri 57113 59436 57129 59452 se
rect 57129 59436 57206 59452
rect 57113 59370 57206 59436
rect 56834 59235 57206 59311
rect 56834 59110 56927 59176
rect 56834 59094 56911 59110
tri 56911 59094 56927 59110 nw
rect 56963 59077 57077 59235
rect 57113 59110 57206 59176
tri 57113 59094 57129 59110 ne
rect 57129 59094 57206 59110
rect 56946 58995 57094 59077
rect 56834 58962 56911 58978
tri 56911 58962 56927 58978 sw
rect 56834 58896 56927 58962
rect 56834 58794 56927 58860
rect 56834 58778 56911 58794
tri 56911 58778 56927 58794 nw
rect 56963 58761 57077 58995
tri 57113 58962 57129 58978 se
rect 57129 58962 57206 58978
rect 57113 58896 57206 58962
rect 57113 58794 57206 58860
tri 57113 58778 57129 58794 ne
rect 57129 58778 57206 58794
rect 56946 58679 57094 58761
rect 56834 58646 56911 58662
tri 56911 58646 56927 58662 sw
rect 56834 58580 56927 58646
rect 56963 58521 57077 58679
tri 57113 58646 57129 58662 se
rect 57129 58646 57206 58662
rect 57113 58580 57206 58646
rect 56834 58445 57206 58521
rect 56834 58320 56927 58386
rect 56834 58304 56911 58320
tri 56911 58304 56927 58320 nw
rect 56963 58287 57077 58445
rect 57113 58320 57206 58386
tri 57113 58304 57129 58320 ne
rect 57129 58304 57206 58320
rect 56946 58205 57094 58287
rect 56834 58172 56911 58188
tri 56911 58172 56927 58188 sw
rect 56834 58106 56927 58172
rect 56834 58004 56927 58070
rect 56834 57988 56911 58004
tri 56911 57988 56927 58004 nw
rect 56963 57971 57077 58205
tri 57113 58172 57129 58188 se
rect 57129 58172 57206 58188
rect 57113 58106 57206 58172
rect 57113 58004 57206 58070
tri 57113 57988 57129 58004 ne
rect 57129 57988 57206 58004
rect 56946 57889 57094 57971
rect 56834 57856 56911 57872
tri 56911 57856 56927 57872 sw
rect 56834 57790 56927 57856
rect 56963 57731 57077 57889
tri 57113 57856 57129 57872 se
rect 57129 57856 57206 57872
rect 57113 57790 57206 57856
rect 56834 57655 57206 57731
rect 56834 57530 56927 57596
rect 56834 57514 56911 57530
tri 56911 57514 56927 57530 nw
rect 56963 57497 57077 57655
rect 57113 57530 57206 57596
tri 57113 57514 57129 57530 ne
rect 57129 57514 57206 57530
rect 56946 57415 57094 57497
rect 56834 57382 56911 57398
tri 56911 57382 56927 57398 sw
rect 56834 57316 56927 57382
rect 56834 57214 56927 57280
rect 56834 57198 56911 57214
tri 56911 57198 56927 57214 nw
rect 56963 57181 57077 57415
tri 57113 57382 57129 57398 se
rect 57129 57382 57206 57398
rect 57113 57316 57206 57382
rect 57113 57214 57206 57280
tri 57113 57198 57129 57214 ne
rect 57129 57198 57206 57214
rect 56946 57099 57094 57181
rect 56834 57066 56911 57082
tri 56911 57066 56927 57082 sw
rect 56834 57000 56927 57066
rect 56963 56941 57077 57099
tri 57113 57066 57129 57082 se
rect 57129 57066 57206 57082
rect 57113 57000 57206 57066
rect 56834 56865 57206 56941
rect 56834 56740 56927 56806
rect 56834 56724 56911 56740
tri 56911 56724 56927 56740 nw
rect 56963 56707 57077 56865
rect 57113 56740 57206 56806
tri 57113 56724 57129 56740 ne
rect 57129 56724 57206 56740
rect 56946 56625 57094 56707
rect 56834 56592 56911 56608
tri 56911 56592 56927 56608 sw
rect 56834 56526 56927 56592
rect 56834 56424 56927 56490
rect 56834 56408 56911 56424
tri 56911 56408 56927 56424 nw
rect 56963 56391 57077 56625
tri 57113 56592 57129 56608 se
rect 57129 56592 57206 56608
rect 57113 56526 57206 56592
rect 57113 56424 57206 56490
tri 57113 56408 57129 56424 ne
rect 57129 56408 57206 56424
rect 56946 56309 57094 56391
rect 56834 56276 56911 56292
tri 56911 56276 56927 56292 sw
rect 56834 56210 56927 56276
rect 56963 56151 57077 56309
tri 57113 56276 57129 56292 se
rect 57129 56276 57206 56292
rect 57113 56210 57206 56276
rect 56834 56075 57206 56151
rect 56834 55950 56927 56016
rect 56834 55934 56911 55950
tri 56911 55934 56927 55950 nw
rect 56963 55917 57077 56075
rect 57113 55950 57206 56016
tri 57113 55934 57129 55950 ne
rect 57129 55934 57206 55950
rect 56946 55835 57094 55917
rect 56834 55802 56911 55818
tri 56911 55802 56927 55818 sw
rect 56834 55736 56927 55802
rect 56834 55634 56927 55700
rect 56834 55618 56911 55634
tri 56911 55618 56927 55634 nw
rect 56963 55601 57077 55835
tri 57113 55802 57129 55818 se
rect 57129 55802 57206 55818
rect 57113 55736 57206 55802
rect 57113 55634 57206 55700
tri 57113 55618 57129 55634 ne
rect 57129 55618 57206 55634
rect 56946 55519 57094 55601
rect 56834 55486 56911 55502
tri 56911 55486 56927 55502 sw
rect 56834 55420 56927 55486
rect 56963 55361 57077 55519
tri 57113 55486 57129 55502 se
rect 57129 55486 57206 55502
rect 57113 55420 57206 55486
rect 56834 55285 57206 55361
rect 56834 55160 56927 55226
rect 56834 55144 56911 55160
tri 56911 55144 56927 55160 nw
rect 56963 55127 57077 55285
rect 57113 55160 57206 55226
tri 57113 55144 57129 55160 ne
rect 57129 55144 57206 55160
rect 56946 55045 57094 55127
rect 56834 55012 56911 55028
tri 56911 55012 56927 55028 sw
rect 56834 54946 56927 55012
rect 56834 54844 56927 54910
rect 56834 54828 56911 54844
tri 56911 54828 56927 54844 nw
rect 56963 54811 57077 55045
tri 57113 55012 57129 55028 se
rect 57129 55012 57206 55028
rect 57113 54946 57206 55012
rect 57113 54844 57206 54910
tri 57113 54828 57129 54844 ne
rect 57129 54828 57206 54844
rect 56946 54729 57094 54811
rect 56834 54696 56911 54712
tri 56911 54696 56927 54712 sw
rect 56834 54630 56927 54696
rect 56963 54571 57077 54729
tri 57113 54696 57129 54712 se
rect 57129 54696 57206 54712
rect 57113 54630 57206 54696
rect 56834 54495 57206 54571
rect 56834 54370 56927 54436
rect 56834 54354 56911 54370
tri 56911 54354 56927 54370 nw
rect 56963 54337 57077 54495
rect 57113 54370 57206 54436
tri 57113 54354 57129 54370 ne
rect 57129 54354 57206 54370
rect 56946 54255 57094 54337
rect 56834 54222 56911 54238
tri 56911 54222 56927 54238 sw
rect 56834 54156 56927 54222
rect 56834 54054 56927 54120
rect 56834 54038 56911 54054
tri 56911 54038 56927 54054 nw
rect 56963 54021 57077 54255
tri 57113 54222 57129 54238 se
rect 57129 54222 57206 54238
rect 57113 54156 57206 54222
rect 57113 54054 57206 54120
tri 57113 54038 57129 54054 ne
rect 57129 54038 57206 54054
rect 56946 53939 57094 54021
rect 56834 53906 56911 53922
tri 56911 53906 56927 53922 sw
rect 56834 53840 56927 53906
rect 56963 53781 57077 53939
tri 57113 53906 57129 53922 se
rect 57129 53906 57206 53922
rect 57113 53840 57206 53906
rect 56834 53705 57206 53781
rect 56834 53580 56927 53646
rect 56834 53564 56911 53580
tri 56911 53564 56927 53580 nw
rect 56963 53547 57077 53705
rect 57113 53580 57206 53646
tri 57113 53564 57129 53580 ne
rect 57129 53564 57206 53580
rect 56946 53465 57094 53547
rect 56834 53432 56911 53448
tri 56911 53432 56927 53448 sw
rect 56834 53366 56927 53432
rect 56834 53264 56927 53330
rect 56834 53248 56911 53264
tri 56911 53248 56927 53264 nw
rect 56963 53231 57077 53465
tri 57113 53432 57129 53448 se
rect 57129 53432 57206 53448
rect 57113 53366 57206 53432
rect 57113 53264 57206 53330
tri 57113 53248 57129 53264 ne
rect 57129 53248 57206 53264
rect 56946 53149 57094 53231
rect 56834 53116 56911 53132
tri 56911 53116 56927 53132 sw
rect 56834 53050 56927 53116
rect 56963 52991 57077 53149
tri 57113 53116 57129 53132 se
rect 57129 53116 57206 53132
rect 57113 53050 57206 53116
rect 56834 52915 57206 52991
rect 56834 52790 56927 52856
rect 56834 52774 56911 52790
tri 56911 52774 56927 52790 nw
rect 56963 52757 57077 52915
rect 57113 52790 57206 52856
tri 57113 52774 57129 52790 ne
rect 57129 52774 57206 52790
rect 56946 52675 57094 52757
rect 56834 52642 56911 52658
tri 56911 52642 56927 52658 sw
rect 56834 52576 56927 52642
rect 56834 52474 56927 52540
rect 56834 52458 56911 52474
tri 56911 52458 56927 52474 nw
rect 56963 52441 57077 52675
tri 57113 52642 57129 52658 se
rect 57129 52642 57206 52658
rect 57113 52576 57206 52642
rect 57113 52474 57206 52540
tri 57113 52458 57129 52474 ne
rect 57129 52458 57206 52474
rect 56946 52359 57094 52441
rect 56834 52326 56911 52342
tri 56911 52326 56927 52342 sw
rect 56834 52260 56927 52326
rect 56963 52201 57077 52359
tri 57113 52326 57129 52342 se
rect 57129 52326 57206 52342
rect 57113 52260 57206 52326
rect 56834 52125 57206 52201
rect 56834 52000 56927 52066
rect 56834 51984 56911 52000
tri 56911 51984 56927 52000 nw
rect 56963 51967 57077 52125
rect 57113 52000 57206 52066
tri 57113 51984 57129 52000 ne
rect 57129 51984 57206 52000
rect 56946 51885 57094 51967
rect 56834 51852 56911 51868
tri 56911 51852 56927 51868 sw
rect 56834 51786 56927 51852
rect 56834 51684 56927 51750
rect 56834 51668 56911 51684
tri 56911 51668 56927 51684 nw
rect 56963 51651 57077 51885
tri 57113 51852 57129 51868 se
rect 57129 51852 57206 51868
rect 57113 51786 57206 51852
rect 57113 51684 57206 51750
tri 57113 51668 57129 51684 ne
rect 57129 51668 57206 51684
rect 56946 51569 57094 51651
rect 56834 51536 56911 51552
tri 56911 51536 56927 51552 sw
rect 56834 51470 56927 51536
rect 56963 51411 57077 51569
tri 57113 51536 57129 51552 se
rect 57129 51536 57206 51552
rect 57113 51470 57206 51536
rect 56834 51335 57206 51411
rect 56834 51210 56927 51276
rect 56834 51194 56911 51210
tri 56911 51194 56927 51210 nw
rect 56963 51177 57077 51335
rect 57113 51210 57206 51276
tri 57113 51194 57129 51210 ne
rect 57129 51194 57206 51210
rect 56946 51095 57094 51177
rect 56834 51062 56911 51078
tri 56911 51062 56927 51078 sw
rect 56834 50996 56927 51062
rect 56834 50894 56927 50960
rect 56834 50878 56911 50894
tri 56911 50878 56927 50894 nw
rect 56963 50861 57077 51095
tri 57113 51062 57129 51078 se
rect 57129 51062 57206 51078
rect 57113 50996 57206 51062
rect 57113 50894 57206 50960
tri 57113 50878 57129 50894 ne
rect 57129 50878 57206 50894
rect 56946 50779 57094 50861
rect 56834 50746 56911 50762
tri 56911 50746 56927 50762 sw
rect 56834 50680 56927 50746
rect 56963 50621 57077 50779
tri 57113 50746 57129 50762 se
rect 57129 50746 57206 50762
rect 57113 50680 57206 50746
rect 56834 50545 57206 50621
rect 56834 50420 56927 50486
rect 56834 50404 56911 50420
tri 56911 50404 56927 50420 nw
rect 56963 50387 57077 50545
rect 57113 50420 57206 50486
tri 57113 50404 57129 50420 ne
rect 57129 50404 57206 50420
rect 56946 50305 57094 50387
rect 56834 50272 56911 50288
tri 56911 50272 56927 50288 sw
rect 56834 50206 56927 50272
rect 56834 50104 56927 50170
rect 56834 50088 56911 50104
tri 56911 50088 56927 50104 nw
rect 56963 50071 57077 50305
tri 57113 50272 57129 50288 se
rect 57129 50272 57206 50288
rect 57113 50206 57206 50272
rect 57113 50104 57206 50170
tri 57113 50088 57129 50104 ne
rect 57129 50088 57206 50104
rect 56946 49989 57094 50071
rect 56834 49956 56911 49972
tri 56911 49956 56927 49972 sw
rect 56834 49890 56927 49956
rect 56963 49831 57077 49989
tri 57113 49956 57129 49972 se
rect 57129 49956 57206 49972
rect 57113 49890 57206 49956
rect 56834 49755 57206 49831
rect 56834 49630 56927 49696
rect 56834 49614 56911 49630
tri 56911 49614 56927 49630 nw
rect 56963 49597 57077 49755
rect 57113 49630 57206 49696
tri 57113 49614 57129 49630 ne
rect 57129 49614 57206 49630
rect 56946 49515 57094 49597
rect 56834 49482 56911 49498
tri 56911 49482 56927 49498 sw
rect 56834 49416 56927 49482
rect 56834 49314 56927 49380
rect 56834 49298 56911 49314
tri 56911 49298 56927 49314 nw
rect 56963 49281 57077 49515
tri 57113 49482 57129 49498 se
rect 57129 49482 57206 49498
rect 57113 49416 57206 49482
rect 57113 49314 57206 49380
tri 57113 49298 57129 49314 ne
rect 57129 49298 57206 49314
rect 56946 49199 57094 49281
rect 56834 49166 56911 49182
tri 56911 49166 56927 49182 sw
rect 56834 49100 56927 49166
rect 56963 49041 57077 49199
tri 57113 49166 57129 49182 se
rect 57129 49166 57206 49182
rect 57113 49100 57206 49166
rect 56834 48965 57206 49041
rect 56834 48840 56927 48906
rect 56834 48824 56911 48840
tri 56911 48824 56927 48840 nw
rect 56963 48807 57077 48965
rect 57113 48840 57206 48906
tri 57113 48824 57129 48840 ne
rect 57129 48824 57206 48840
rect 56946 48725 57094 48807
rect 56834 48692 56911 48708
tri 56911 48692 56927 48708 sw
rect 56834 48626 56927 48692
rect 56834 48524 56927 48590
rect 56834 48508 56911 48524
tri 56911 48508 56927 48524 nw
rect 56963 48491 57077 48725
tri 57113 48692 57129 48708 se
rect 57129 48692 57206 48708
rect 57113 48626 57206 48692
rect 57113 48524 57206 48590
tri 57113 48508 57129 48524 ne
rect 57129 48508 57206 48524
rect 56946 48409 57094 48491
rect 56834 48376 56911 48392
tri 56911 48376 56927 48392 sw
rect 56834 48310 56927 48376
rect 56963 48251 57077 48409
tri 57113 48376 57129 48392 se
rect 57129 48376 57206 48392
rect 57113 48310 57206 48376
rect 56834 48175 57206 48251
rect 56834 48050 56927 48116
rect 56834 48034 56911 48050
tri 56911 48034 56927 48050 nw
rect 56963 48017 57077 48175
rect 57113 48050 57206 48116
tri 57113 48034 57129 48050 ne
rect 57129 48034 57206 48050
rect 56946 47935 57094 48017
rect 56834 47902 56911 47918
tri 56911 47902 56927 47918 sw
rect 56834 47836 56927 47902
rect 56834 47734 56927 47800
rect 56834 47718 56911 47734
tri 56911 47718 56927 47734 nw
rect 56963 47701 57077 47935
tri 57113 47902 57129 47918 se
rect 57129 47902 57206 47918
rect 57113 47836 57206 47902
rect 57113 47734 57206 47800
tri 57113 47718 57129 47734 ne
rect 57129 47718 57206 47734
rect 56946 47619 57094 47701
rect 56834 47586 56911 47602
tri 56911 47586 56927 47602 sw
rect 56834 47520 56927 47586
rect 56963 47461 57077 47619
tri 57113 47586 57129 47602 se
rect 57129 47586 57206 47602
rect 57113 47520 57206 47586
rect 56834 47385 57206 47461
rect 56834 47260 56927 47326
rect 56834 47244 56911 47260
tri 56911 47244 56927 47260 nw
rect 56963 47227 57077 47385
rect 57113 47260 57206 47326
tri 57113 47244 57129 47260 ne
rect 57129 47244 57206 47260
rect 56946 47145 57094 47227
rect 56834 47112 56911 47128
tri 56911 47112 56927 47128 sw
rect 56834 47046 56927 47112
rect 56834 46944 56927 47010
rect 56834 46928 56911 46944
tri 56911 46928 56927 46944 nw
rect 56963 46911 57077 47145
tri 57113 47112 57129 47128 se
rect 57129 47112 57206 47128
rect 57113 47046 57206 47112
rect 57113 46944 57206 47010
tri 57113 46928 57129 46944 ne
rect 57129 46928 57206 46944
rect 56946 46829 57094 46911
rect 56834 46796 56911 46812
tri 56911 46796 56927 46812 sw
rect 56834 46730 56927 46796
rect 56963 46671 57077 46829
tri 57113 46796 57129 46812 se
rect 57129 46796 57206 46812
rect 57113 46730 57206 46796
rect 56834 46595 57206 46671
rect 56834 46470 56927 46536
rect 56834 46454 56911 46470
tri 56911 46454 56927 46470 nw
rect 56963 46437 57077 46595
rect 57113 46470 57206 46536
tri 57113 46454 57129 46470 ne
rect 57129 46454 57206 46470
rect 56946 46355 57094 46437
rect 56834 46322 56911 46338
tri 56911 46322 56927 46338 sw
rect 56834 46256 56927 46322
rect 56834 46154 56927 46220
rect 56834 46138 56911 46154
tri 56911 46138 56927 46154 nw
rect 56963 46121 57077 46355
tri 57113 46322 57129 46338 se
rect 57129 46322 57206 46338
rect 57113 46256 57206 46322
rect 57113 46154 57206 46220
tri 57113 46138 57129 46154 ne
rect 57129 46138 57206 46154
rect 56946 46039 57094 46121
rect 56834 46006 56911 46022
tri 56911 46006 56927 46022 sw
rect 56834 45940 56927 46006
rect 56963 45881 57077 46039
tri 57113 46006 57129 46022 se
rect 57129 46006 57206 46022
rect 57113 45940 57206 46006
rect 56834 45805 57206 45881
rect 56834 45680 56927 45746
rect 56834 45664 56911 45680
tri 56911 45664 56927 45680 nw
rect 56963 45647 57077 45805
rect 57113 45680 57206 45746
tri 57113 45664 57129 45680 ne
rect 57129 45664 57206 45680
rect 56946 45565 57094 45647
rect 56834 45532 56911 45548
tri 56911 45532 56927 45548 sw
rect 56834 45466 56927 45532
rect 56834 45364 56927 45430
rect 56834 45348 56911 45364
tri 56911 45348 56927 45364 nw
rect 56963 45331 57077 45565
tri 57113 45532 57129 45548 se
rect 57129 45532 57206 45548
rect 57113 45466 57206 45532
rect 57113 45364 57206 45430
tri 57113 45348 57129 45364 ne
rect 57129 45348 57206 45364
rect 56946 45249 57094 45331
rect 56834 45216 56911 45232
tri 56911 45216 56927 45232 sw
rect 56834 45150 56927 45216
rect 56963 45091 57077 45249
tri 57113 45216 57129 45232 se
rect 57129 45216 57206 45232
rect 57113 45150 57206 45216
rect 56834 45015 57206 45091
rect 56834 44890 56927 44956
rect 56834 44874 56911 44890
tri 56911 44874 56927 44890 nw
rect 56963 44857 57077 45015
rect 57113 44890 57206 44956
tri 57113 44874 57129 44890 ne
rect 57129 44874 57206 44890
rect 56946 44775 57094 44857
rect 56834 44742 56911 44758
tri 56911 44742 56927 44758 sw
rect 56834 44676 56927 44742
rect 56834 44574 56927 44640
rect 56834 44558 56911 44574
tri 56911 44558 56927 44574 nw
rect 56963 44541 57077 44775
tri 57113 44742 57129 44758 se
rect 57129 44742 57206 44758
rect 57113 44676 57206 44742
rect 57113 44574 57206 44640
tri 57113 44558 57129 44574 ne
rect 57129 44558 57206 44574
rect 56946 44459 57094 44541
rect 56834 44426 56911 44442
tri 56911 44426 56927 44442 sw
rect 56834 44360 56927 44426
rect 56963 44301 57077 44459
tri 57113 44426 57129 44442 se
rect 57129 44426 57206 44442
rect 57113 44360 57206 44426
rect 56834 44225 57206 44301
rect 56834 44100 56927 44166
rect 56834 44084 56911 44100
tri 56911 44084 56927 44100 nw
rect 56963 44067 57077 44225
rect 57113 44100 57206 44166
tri 57113 44084 57129 44100 ne
rect 57129 44084 57206 44100
rect 56946 43985 57094 44067
rect 56834 43952 56911 43968
tri 56911 43952 56927 43968 sw
rect 56834 43886 56927 43952
rect 56834 43784 56927 43850
rect 56834 43768 56911 43784
tri 56911 43768 56927 43784 nw
rect 56963 43751 57077 43985
tri 57113 43952 57129 43968 se
rect 57129 43952 57206 43968
rect 57113 43886 57206 43952
rect 57113 43784 57206 43850
tri 57113 43768 57129 43784 ne
rect 57129 43768 57206 43784
rect 56946 43669 57094 43751
rect 56834 43636 56911 43652
tri 56911 43636 56927 43652 sw
rect 56834 43570 56927 43636
rect 56963 43511 57077 43669
tri 57113 43636 57129 43652 se
rect 57129 43636 57206 43652
rect 57113 43570 57206 43636
rect 56834 43435 57206 43511
rect 56834 43310 56927 43376
rect 56834 43294 56911 43310
tri 56911 43294 56927 43310 nw
rect 56963 43277 57077 43435
rect 57113 43310 57206 43376
tri 57113 43294 57129 43310 ne
rect 57129 43294 57206 43310
rect 56946 43195 57094 43277
rect 56834 43162 56911 43178
tri 56911 43162 56927 43178 sw
rect 56834 43096 56927 43162
rect 56834 42994 56927 43060
rect 56834 42978 56911 42994
tri 56911 42978 56927 42994 nw
rect 56963 42961 57077 43195
tri 57113 43162 57129 43178 se
rect 57129 43162 57206 43178
rect 57113 43096 57206 43162
rect 57113 42994 57206 43060
tri 57113 42978 57129 42994 ne
rect 57129 42978 57206 42994
rect 56946 42879 57094 42961
rect 56834 42846 56911 42862
tri 56911 42846 56927 42862 sw
rect 56834 42780 56927 42846
rect 56963 42721 57077 42879
tri 57113 42846 57129 42862 se
rect 57129 42846 57206 42862
rect 57113 42780 57206 42846
rect 56834 42645 57206 42721
rect 56834 42520 56927 42586
rect 56834 42504 56911 42520
tri 56911 42504 56927 42520 nw
rect 56963 42487 57077 42645
rect 57113 42520 57206 42586
tri 57113 42504 57129 42520 ne
rect 57129 42504 57206 42520
rect 56946 42405 57094 42487
rect 56834 42372 56911 42388
tri 56911 42372 56927 42388 sw
rect 56834 42306 56927 42372
rect 56834 42204 56927 42270
rect 56834 42188 56911 42204
tri 56911 42188 56927 42204 nw
rect 56963 42171 57077 42405
tri 57113 42372 57129 42388 se
rect 57129 42372 57206 42388
rect 57113 42306 57206 42372
rect 57113 42204 57206 42270
tri 57113 42188 57129 42204 ne
rect 57129 42188 57206 42204
rect 56946 42089 57094 42171
rect 56834 42056 56911 42072
tri 56911 42056 56927 42072 sw
rect 56834 41990 56927 42056
rect 56963 41931 57077 42089
tri 57113 42056 57129 42072 se
rect 57129 42056 57206 42072
rect 57113 41990 57206 42056
rect 56834 41855 57206 41931
rect 56834 41730 56927 41796
rect 56834 41714 56911 41730
tri 56911 41714 56927 41730 nw
rect 56963 41697 57077 41855
rect 57113 41730 57206 41796
tri 57113 41714 57129 41730 ne
rect 57129 41714 57206 41730
rect 56946 41615 57094 41697
rect 56834 41582 56911 41598
tri 56911 41582 56927 41598 sw
rect 56834 41516 56927 41582
rect 56834 41414 56927 41480
rect 56834 41398 56911 41414
tri 56911 41398 56927 41414 nw
rect 56963 41381 57077 41615
tri 57113 41582 57129 41598 se
rect 57129 41582 57206 41598
rect 57113 41516 57206 41582
rect 57113 41414 57206 41480
tri 57113 41398 57129 41414 ne
rect 57129 41398 57206 41414
rect 56946 41299 57094 41381
rect 56834 41266 56911 41282
tri 56911 41266 56927 41282 sw
rect 56834 41200 56927 41266
rect 56963 41141 57077 41299
tri 57113 41266 57129 41282 se
rect 57129 41266 57206 41282
rect 57113 41200 57206 41266
rect 56834 41065 57206 41141
rect 56834 40940 56927 41006
rect 56834 40924 56911 40940
tri 56911 40924 56927 40940 nw
rect 56963 40907 57077 41065
rect 57113 40940 57206 41006
tri 57113 40924 57129 40940 ne
rect 57129 40924 57206 40940
rect 56946 40825 57094 40907
rect 56834 40792 56911 40808
tri 56911 40792 56927 40808 sw
rect 56834 40726 56927 40792
rect 56834 40624 56927 40690
rect 56834 40608 56911 40624
tri 56911 40608 56927 40624 nw
rect 56963 40591 57077 40825
tri 57113 40792 57129 40808 se
rect 57129 40792 57206 40808
rect 57113 40726 57206 40792
rect 57113 40624 57206 40690
tri 57113 40608 57129 40624 ne
rect 57129 40608 57206 40624
rect 56946 40509 57094 40591
rect 56834 40476 56911 40492
tri 56911 40476 56927 40492 sw
rect 56834 40410 56927 40476
rect 56963 40351 57077 40509
tri 57113 40476 57129 40492 se
rect 57129 40476 57206 40492
rect 57113 40410 57206 40476
rect 56834 40275 57206 40351
rect 56834 40150 56927 40216
rect 56834 40134 56911 40150
tri 56911 40134 56927 40150 nw
rect 56963 40117 57077 40275
rect 57113 40150 57206 40216
tri 57113 40134 57129 40150 ne
rect 57129 40134 57206 40150
rect 56946 40035 57094 40117
rect 56834 40002 56911 40018
tri 56911 40002 56927 40018 sw
rect 56834 39936 56927 40002
rect 56834 39834 56927 39900
rect 56834 39818 56911 39834
tri 56911 39818 56927 39834 nw
rect 56963 39801 57077 40035
tri 57113 40002 57129 40018 se
rect 57129 40002 57206 40018
rect 57113 39936 57206 40002
rect 57113 39834 57206 39900
tri 57113 39818 57129 39834 ne
rect 57129 39818 57206 39834
rect 56946 39719 57094 39801
rect 56834 39686 56911 39702
tri 56911 39686 56927 39702 sw
rect 56834 39620 56927 39686
rect 56963 39561 57077 39719
tri 57113 39686 57129 39702 se
rect 57129 39686 57206 39702
rect 57113 39620 57206 39686
rect 56834 39485 57206 39561
rect 56834 39360 56927 39426
rect 56834 39344 56911 39360
tri 56911 39344 56927 39360 nw
rect 56963 39327 57077 39485
rect 57113 39360 57206 39426
tri 57113 39344 57129 39360 ne
rect 57129 39344 57206 39360
rect 56946 39245 57094 39327
rect 56834 39212 56911 39228
tri 56911 39212 56927 39228 sw
rect 56834 39146 56927 39212
rect 56834 39044 56927 39110
rect 56834 39028 56911 39044
tri 56911 39028 56927 39044 nw
rect 56963 39011 57077 39245
tri 57113 39212 57129 39228 se
rect 57129 39212 57206 39228
rect 57113 39146 57206 39212
rect 57113 39044 57206 39110
tri 57113 39028 57129 39044 ne
rect 57129 39028 57206 39044
rect 56946 38929 57094 39011
rect 56834 38896 56911 38912
tri 56911 38896 56927 38912 sw
rect 56834 38830 56927 38896
rect 56963 38771 57077 38929
tri 57113 38896 57129 38912 se
rect 57129 38896 57206 38912
rect 57113 38830 57206 38896
rect 56834 38695 57206 38771
rect 56834 38570 56927 38636
rect 56834 38554 56911 38570
tri 56911 38554 56927 38570 nw
rect 56963 38537 57077 38695
rect 57113 38570 57206 38636
tri 57113 38554 57129 38570 ne
rect 57129 38554 57206 38570
rect 56946 38455 57094 38537
rect 56834 38422 56911 38438
tri 56911 38422 56927 38438 sw
rect 56834 38356 56927 38422
rect 56834 38254 56927 38320
rect 56834 38238 56911 38254
tri 56911 38238 56927 38254 nw
rect 56963 38221 57077 38455
tri 57113 38422 57129 38438 se
rect 57129 38422 57206 38438
rect 57113 38356 57206 38422
rect 57113 38254 57206 38320
tri 57113 38238 57129 38254 ne
rect 57129 38238 57206 38254
rect 56946 38139 57094 38221
rect 56834 38106 56911 38122
tri 56911 38106 56927 38122 sw
rect 56834 38040 56927 38106
rect 56963 37981 57077 38139
tri 57113 38106 57129 38122 se
rect 57129 38106 57206 38122
rect 57113 38040 57206 38106
rect 56834 37905 57206 37981
rect 56834 37780 56927 37846
rect 56834 37764 56911 37780
tri 56911 37764 56927 37780 nw
rect 56963 37747 57077 37905
rect 57113 37780 57206 37846
tri 57113 37764 57129 37780 ne
rect 57129 37764 57206 37780
rect 56946 37665 57094 37747
rect 56834 37632 56911 37648
tri 56911 37632 56927 37648 sw
rect 56834 37566 56927 37632
rect 56834 37464 56927 37530
rect 56834 37448 56911 37464
tri 56911 37448 56927 37464 nw
rect 56963 37431 57077 37665
tri 57113 37632 57129 37648 se
rect 57129 37632 57206 37648
rect 57113 37566 57206 37632
rect 57113 37464 57206 37530
tri 57113 37448 57129 37464 ne
rect 57129 37448 57206 37464
rect 56946 37349 57094 37431
rect 56834 37316 56911 37332
tri 56911 37316 56927 37332 sw
rect 56834 37250 56927 37316
rect 56963 37191 57077 37349
tri 57113 37316 57129 37332 se
rect 57129 37316 57206 37332
rect 57113 37250 57206 37316
rect 56834 37115 57206 37191
rect 56834 36990 56927 37056
rect 56834 36974 56911 36990
tri 56911 36974 56927 36990 nw
rect 56963 36957 57077 37115
rect 57113 36990 57206 37056
tri 57113 36974 57129 36990 ne
rect 57129 36974 57206 36990
rect 56946 36875 57094 36957
rect 56834 36842 56911 36858
tri 56911 36842 56927 36858 sw
rect 56834 36776 56927 36842
rect 56834 36674 56927 36740
rect 56834 36658 56911 36674
tri 56911 36658 56927 36674 nw
rect 56963 36641 57077 36875
tri 57113 36842 57129 36858 se
rect 57129 36842 57206 36858
rect 57113 36776 57206 36842
rect 57113 36674 57206 36740
tri 57113 36658 57129 36674 ne
rect 57129 36658 57206 36674
rect 56946 36559 57094 36641
rect 56834 36526 56911 36542
tri 56911 36526 56927 36542 sw
rect 56834 36460 56927 36526
rect 56963 36401 57077 36559
tri 57113 36526 57129 36542 se
rect 57129 36526 57206 36542
rect 57113 36460 57206 36526
rect 56834 36325 57206 36401
rect 56834 36200 56927 36266
rect 56834 36184 56911 36200
tri 56911 36184 56927 36200 nw
rect 56963 36167 57077 36325
rect 57113 36200 57206 36266
tri 57113 36184 57129 36200 ne
rect 57129 36184 57206 36200
rect 56946 36085 57094 36167
rect 56834 36052 56911 36068
tri 56911 36052 56927 36068 sw
rect 56834 35986 56927 36052
rect 56834 35884 56927 35950
rect 56834 35868 56911 35884
tri 56911 35868 56927 35884 nw
rect 56963 35851 57077 36085
tri 57113 36052 57129 36068 se
rect 57129 36052 57206 36068
rect 57113 35986 57206 36052
rect 57113 35884 57206 35950
tri 57113 35868 57129 35884 ne
rect 57129 35868 57206 35884
rect 56946 35769 57094 35851
rect 56834 35736 56911 35752
tri 56911 35736 56927 35752 sw
rect 56834 35670 56927 35736
rect 56963 35611 57077 35769
tri 57113 35736 57129 35752 se
rect 57129 35736 57206 35752
rect 57113 35670 57206 35736
rect 56834 35535 57206 35611
rect 56834 35410 56927 35476
rect 56834 35394 56911 35410
tri 56911 35394 56927 35410 nw
rect 56963 35377 57077 35535
rect 57113 35410 57206 35476
tri 57113 35394 57129 35410 ne
rect 57129 35394 57206 35410
rect 56946 35295 57094 35377
rect 56834 35262 56911 35278
tri 56911 35262 56927 35278 sw
rect 56834 35196 56927 35262
rect 56834 35094 56927 35160
rect 56834 35078 56911 35094
tri 56911 35078 56927 35094 nw
rect 56963 35061 57077 35295
tri 57113 35262 57129 35278 se
rect 57129 35262 57206 35278
rect 57113 35196 57206 35262
rect 57113 35094 57206 35160
tri 57113 35078 57129 35094 ne
rect 57129 35078 57206 35094
rect 56946 34979 57094 35061
rect 56834 34946 56911 34962
tri 56911 34946 56927 34962 sw
rect 56834 34880 56927 34946
rect 56963 34821 57077 34979
tri 57113 34946 57129 34962 se
rect 57129 34946 57206 34962
rect 57113 34880 57206 34946
rect 56834 34745 57206 34821
rect 56834 34620 56927 34686
rect 56834 34604 56911 34620
tri 56911 34604 56927 34620 nw
rect 56963 34587 57077 34745
rect 57113 34620 57206 34686
tri 57113 34604 57129 34620 ne
rect 57129 34604 57206 34620
rect 56946 34505 57094 34587
rect 56834 34472 56911 34488
tri 56911 34472 56927 34488 sw
rect 56834 34406 56927 34472
rect 56834 34304 56927 34370
rect 56834 34288 56911 34304
tri 56911 34288 56927 34304 nw
rect 56963 34271 57077 34505
tri 57113 34472 57129 34488 se
rect 57129 34472 57206 34488
rect 57113 34406 57206 34472
rect 57113 34304 57206 34370
tri 57113 34288 57129 34304 ne
rect 57129 34288 57206 34304
rect 56946 34189 57094 34271
rect 56834 34156 56911 34172
tri 56911 34156 56927 34172 sw
rect 56834 34090 56927 34156
rect 56963 34031 57077 34189
tri 57113 34156 57129 34172 se
rect 57129 34156 57206 34172
rect 57113 34090 57206 34156
rect 56834 33955 57206 34031
rect 56834 33830 56927 33896
rect 56834 33814 56911 33830
tri 56911 33814 56927 33830 nw
rect 56963 33797 57077 33955
rect 57113 33830 57206 33896
tri 57113 33814 57129 33830 ne
rect 57129 33814 57206 33830
rect 56946 33715 57094 33797
rect 56834 33682 56911 33698
tri 56911 33682 56927 33698 sw
rect 56834 33616 56927 33682
rect 56834 33514 56927 33580
rect 56834 33498 56911 33514
tri 56911 33498 56927 33514 nw
rect 56963 33481 57077 33715
tri 57113 33682 57129 33698 se
rect 57129 33682 57206 33698
rect 57113 33616 57206 33682
rect 57113 33514 57206 33580
tri 57113 33498 57129 33514 ne
rect 57129 33498 57206 33514
rect 56946 33399 57094 33481
rect 56834 33366 56911 33382
tri 56911 33366 56927 33382 sw
rect 56834 33300 56927 33366
rect 56963 33241 57077 33399
tri 57113 33366 57129 33382 se
rect 57129 33366 57206 33382
rect 57113 33300 57206 33366
rect 56834 33165 57206 33241
rect 56834 33040 56927 33106
rect 56834 33024 56911 33040
tri 56911 33024 56927 33040 nw
rect 56963 33007 57077 33165
rect 57113 33040 57206 33106
tri 57113 33024 57129 33040 ne
rect 57129 33024 57206 33040
rect 56946 32925 57094 33007
rect 56834 32892 56911 32908
tri 56911 32892 56927 32908 sw
rect 56834 32826 56927 32892
rect 56834 32724 56927 32790
rect 56834 32708 56911 32724
tri 56911 32708 56927 32724 nw
rect 56963 32691 57077 32925
tri 57113 32892 57129 32908 se
rect 57129 32892 57206 32908
rect 57113 32826 57206 32892
rect 57113 32724 57206 32790
tri 57113 32708 57129 32724 ne
rect 57129 32708 57206 32724
rect 56946 32609 57094 32691
rect 56834 32576 56911 32592
tri 56911 32576 56927 32592 sw
rect 56834 32510 56927 32576
rect 56963 32451 57077 32609
tri 57113 32576 57129 32592 se
rect 57129 32576 57206 32592
rect 57113 32510 57206 32576
rect 56834 32375 57206 32451
rect 56834 32250 56927 32316
rect 56834 32234 56911 32250
tri 56911 32234 56927 32250 nw
rect 56963 32217 57077 32375
rect 57113 32250 57206 32316
tri 57113 32234 57129 32250 ne
rect 57129 32234 57206 32250
rect 56946 32135 57094 32217
rect 56834 32102 56911 32118
tri 56911 32102 56927 32118 sw
rect 56834 32036 56927 32102
rect 56834 31934 56927 32000
rect 56834 31918 56911 31934
tri 56911 31918 56927 31934 nw
rect 56963 31901 57077 32135
tri 57113 32102 57129 32118 se
rect 57129 32102 57206 32118
rect 57113 32036 57206 32102
rect 57113 31934 57206 32000
tri 57113 31918 57129 31934 ne
rect 57129 31918 57206 31934
rect 56946 31819 57094 31901
rect 56834 31786 56911 31802
tri 56911 31786 56927 31802 sw
rect 56834 31720 56927 31786
rect 56963 31661 57077 31819
tri 57113 31786 57129 31802 se
rect 57129 31786 57206 31802
rect 57113 31720 57206 31786
rect 56834 31585 57206 31661
rect 56834 31460 56927 31526
rect 56834 31444 56911 31460
tri 56911 31444 56927 31460 nw
rect 56963 31427 57077 31585
rect 57113 31460 57206 31526
tri 57113 31444 57129 31460 ne
rect 57129 31444 57206 31460
rect 56946 31345 57094 31427
rect 56834 31312 56911 31328
tri 56911 31312 56927 31328 sw
rect 56834 31246 56927 31312
rect 56834 31144 56927 31210
rect 56834 31128 56911 31144
tri 56911 31128 56927 31144 nw
rect 56963 31111 57077 31345
tri 57113 31312 57129 31328 se
rect 57129 31312 57206 31328
rect 57113 31246 57206 31312
rect 57113 31144 57206 31210
tri 57113 31128 57129 31144 ne
rect 57129 31128 57206 31144
rect 56946 31029 57094 31111
rect 56834 30996 56911 31012
tri 56911 30996 56927 31012 sw
rect 56834 30930 56927 30996
rect 56963 30871 57077 31029
tri 57113 30996 57129 31012 se
rect 57129 30996 57206 31012
rect 57113 30930 57206 30996
rect 56834 30795 57206 30871
rect 56834 30670 56927 30736
rect 56834 30654 56911 30670
tri 56911 30654 56927 30670 nw
rect 56963 30637 57077 30795
rect 57113 30670 57206 30736
tri 57113 30654 57129 30670 ne
rect 57129 30654 57206 30670
rect 56946 30555 57094 30637
rect 56834 30522 56911 30538
tri 56911 30522 56927 30538 sw
rect 56834 30456 56927 30522
rect 56834 30354 56927 30420
rect 56834 30338 56911 30354
tri 56911 30338 56927 30354 nw
rect 56963 30321 57077 30555
tri 57113 30522 57129 30538 se
rect 57129 30522 57206 30538
rect 57113 30456 57206 30522
rect 57113 30354 57206 30420
tri 57113 30338 57129 30354 ne
rect 57129 30338 57206 30354
rect 56946 30239 57094 30321
rect 56834 30206 56911 30222
tri 56911 30206 56927 30222 sw
rect 56834 30140 56927 30206
rect 56963 30081 57077 30239
tri 57113 30206 57129 30222 se
rect 57129 30206 57206 30222
rect 57113 30140 57206 30206
rect 56834 30005 57206 30081
rect 56834 29880 56927 29946
rect 56834 29864 56911 29880
tri 56911 29864 56927 29880 nw
rect 56963 29847 57077 30005
rect 57113 29880 57206 29946
tri 57113 29864 57129 29880 ne
rect 57129 29864 57206 29880
rect 56946 29765 57094 29847
rect 56834 29732 56911 29748
tri 56911 29732 56927 29748 sw
rect 56834 29666 56927 29732
rect 56834 29564 56927 29630
rect 56834 29548 56911 29564
tri 56911 29548 56927 29564 nw
rect 56963 29531 57077 29765
tri 57113 29732 57129 29748 se
rect 57129 29732 57206 29748
rect 57113 29666 57206 29732
rect 57113 29564 57206 29630
tri 57113 29548 57129 29564 ne
rect 57129 29548 57206 29564
rect 56946 29449 57094 29531
rect 56834 29416 56911 29432
tri 56911 29416 56927 29432 sw
rect 56834 29350 56927 29416
rect 56963 29291 57077 29449
tri 57113 29416 57129 29432 se
rect 57129 29416 57206 29432
rect 57113 29350 57206 29416
rect 56834 29215 57206 29291
rect 56834 29090 56927 29156
rect 56834 29074 56911 29090
tri 56911 29074 56927 29090 nw
rect 56963 29057 57077 29215
rect 57113 29090 57206 29156
tri 57113 29074 57129 29090 ne
rect 57129 29074 57206 29090
rect 56946 28975 57094 29057
rect 56834 28942 56911 28958
tri 56911 28942 56927 28958 sw
rect 56834 28876 56927 28942
rect 56963 28833 57077 28975
tri 57113 28942 57129 28958 se
rect 57129 28942 57206 28958
rect 57113 28876 57206 28942
rect 57242 28463 57278 80603
rect 57314 28463 57350 80603
rect 57386 80445 57422 80603
rect 57378 80303 57430 80445
rect 57386 28763 57422 80303
rect 57378 28621 57430 28763
rect 57386 28463 57422 28621
rect 57458 28463 57494 80603
rect 57530 28463 57566 80603
rect 57602 28833 57686 80233
rect 57722 28463 57758 80603
rect 57794 28463 57830 80603
rect 57866 80445 57902 80603
rect 57858 80303 57910 80445
rect 57866 28763 57902 80303
rect 57858 28621 57910 28763
rect 57866 28463 57902 28621
rect 57938 28463 57974 80603
rect 58010 28463 58046 80603
rect 58082 80124 58175 80190
rect 58082 80108 58159 80124
tri 58159 80108 58175 80124 nw
rect 58211 80091 58268 80233
rect 58194 80009 58268 80091
rect 58082 79976 58159 79992
tri 58159 79976 58175 79992 sw
rect 58082 79910 58175 79976
rect 58211 79851 58268 80009
rect 58082 79775 58268 79851
rect 58082 79650 58175 79716
rect 58082 79634 58159 79650
tri 58159 79634 58175 79650 nw
rect 58211 79617 58268 79775
rect 58194 79535 58268 79617
rect 58082 79502 58159 79518
tri 58159 79502 58175 79518 sw
rect 58082 79436 58175 79502
rect 58082 79334 58175 79400
rect 58082 79318 58159 79334
tri 58159 79318 58175 79334 nw
rect 58211 79301 58268 79535
rect 58194 79219 58268 79301
rect 58082 79186 58159 79202
tri 58159 79186 58175 79202 sw
rect 58082 79120 58175 79186
rect 58211 79061 58268 79219
rect 58082 78985 58268 79061
rect 58082 78860 58175 78926
rect 58082 78844 58159 78860
tri 58159 78844 58175 78860 nw
rect 58211 78827 58268 78985
rect 58194 78745 58268 78827
rect 58082 78712 58159 78728
tri 58159 78712 58175 78728 sw
rect 58082 78646 58175 78712
rect 58082 78544 58175 78610
rect 58082 78528 58159 78544
tri 58159 78528 58175 78544 nw
rect 58211 78511 58268 78745
rect 58194 78429 58268 78511
rect 58082 78396 58159 78412
tri 58159 78396 58175 78412 sw
rect 58082 78330 58175 78396
rect 58211 78271 58268 78429
rect 58082 78195 58268 78271
rect 58082 78070 58175 78136
rect 58082 78054 58159 78070
tri 58159 78054 58175 78070 nw
rect 58211 78037 58268 78195
rect 58194 77955 58268 78037
rect 58082 77922 58159 77938
tri 58159 77922 58175 77938 sw
rect 58082 77856 58175 77922
rect 58082 77754 58175 77820
rect 58082 77738 58159 77754
tri 58159 77738 58175 77754 nw
rect 58211 77721 58268 77955
rect 58194 77639 58268 77721
rect 58082 77606 58159 77622
tri 58159 77606 58175 77622 sw
rect 58082 77540 58175 77606
rect 58211 77481 58268 77639
rect 58082 77405 58268 77481
rect 58082 77280 58175 77346
rect 58082 77264 58159 77280
tri 58159 77264 58175 77280 nw
rect 58211 77247 58268 77405
rect 58194 77165 58268 77247
rect 58082 77132 58159 77148
tri 58159 77132 58175 77148 sw
rect 58082 77066 58175 77132
rect 58082 76964 58175 77030
rect 58082 76948 58159 76964
tri 58159 76948 58175 76964 nw
rect 58211 76931 58268 77165
rect 58194 76849 58268 76931
rect 58082 76816 58159 76832
tri 58159 76816 58175 76832 sw
rect 58082 76750 58175 76816
rect 58211 76691 58268 76849
rect 58082 76615 58268 76691
rect 58082 76490 58175 76556
rect 58082 76474 58159 76490
tri 58159 76474 58175 76490 nw
rect 58211 76457 58268 76615
rect 58194 76375 58268 76457
rect 58082 76342 58159 76358
tri 58159 76342 58175 76358 sw
rect 58082 76276 58175 76342
rect 58082 76174 58175 76240
rect 58082 76158 58159 76174
tri 58159 76158 58175 76174 nw
rect 58211 76141 58268 76375
rect 58194 76059 58268 76141
rect 58082 76026 58159 76042
tri 58159 76026 58175 76042 sw
rect 58082 75960 58175 76026
rect 58211 75901 58268 76059
rect 58082 75825 58268 75901
rect 58082 75700 58175 75766
rect 58082 75684 58159 75700
tri 58159 75684 58175 75700 nw
rect 58211 75667 58268 75825
rect 58194 75585 58268 75667
rect 58082 75552 58159 75568
tri 58159 75552 58175 75568 sw
rect 58082 75486 58175 75552
rect 58082 75384 58175 75450
rect 58082 75368 58159 75384
tri 58159 75368 58175 75384 nw
rect 58211 75351 58268 75585
rect 58194 75269 58268 75351
rect 58082 75236 58159 75252
tri 58159 75236 58175 75252 sw
rect 58082 75170 58175 75236
rect 58211 75111 58268 75269
rect 58082 75035 58268 75111
rect 58082 74910 58175 74976
rect 58082 74894 58159 74910
tri 58159 74894 58175 74910 nw
rect 58211 74877 58268 75035
rect 58194 74795 58268 74877
rect 58082 74762 58159 74778
tri 58159 74762 58175 74778 sw
rect 58082 74696 58175 74762
rect 58082 74594 58175 74660
rect 58082 74578 58159 74594
tri 58159 74578 58175 74594 nw
rect 58211 74561 58268 74795
rect 58194 74479 58268 74561
rect 58082 74446 58159 74462
tri 58159 74446 58175 74462 sw
rect 58082 74380 58175 74446
rect 58211 74321 58268 74479
rect 58082 74245 58268 74321
rect 58082 74120 58175 74186
rect 58082 74104 58159 74120
tri 58159 74104 58175 74120 nw
rect 58211 74087 58268 74245
rect 58194 74005 58268 74087
rect 58082 73972 58159 73988
tri 58159 73972 58175 73988 sw
rect 58082 73906 58175 73972
rect 58082 73804 58175 73870
rect 58082 73788 58159 73804
tri 58159 73788 58175 73804 nw
rect 58211 73771 58268 74005
rect 58194 73689 58268 73771
rect 58082 73656 58159 73672
tri 58159 73656 58175 73672 sw
rect 58082 73590 58175 73656
rect 58211 73531 58268 73689
rect 58082 73455 58268 73531
rect 58082 73330 58175 73396
rect 58082 73314 58159 73330
tri 58159 73314 58175 73330 nw
rect 58211 73297 58268 73455
rect 58194 73215 58268 73297
rect 58082 73182 58159 73198
tri 58159 73182 58175 73198 sw
rect 58082 73116 58175 73182
rect 58082 73014 58175 73080
rect 58082 72998 58159 73014
tri 58159 72998 58175 73014 nw
rect 58211 72981 58268 73215
rect 58194 72899 58268 72981
rect 58082 72866 58159 72882
tri 58159 72866 58175 72882 sw
rect 58082 72800 58175 72866
rect 58211 72741 58268 72899
rect 58082 72665 58268 72741
rect 58082 72540 58175 72606
rect 58082 72524 58159 72540
tri 58159 72524 58175 72540 nw
rect 58211 72507 58268 72665
rect 58194 72425 58268 72507
rect 58082 72392 58159 72408
tri 58159 72392 58175 72408 sw
rect 58082 72326 58175 72392
rect 58082 72224 58175 72290
rect 58082 72208 58159 72224
tri 58159 72208 58175 72224 nw
rect 58211 72191 58268 72425
rect 58194 72109 58268 72191
rect 58082 72076 58159 72092
tri 58159 72076 58175 72092 sw
rect 58082 72010 58175 72076
rect 58211 71951 58268 72109
rect 58082 71875 58268 71951
rect 58082 71750 58175 71816
rect 58082 71734 58159 71750
tri 58159 71734 58175 71750 nw
rect 58211 71717 58268 71875
rect 58194 71635 58268 71717
rect 58082 71602 58159 71618
tri 58159 71602 58175 71618 sw
rect 58082 71536 58175 71602
rect 58082 71434 58175 71500
rect 58082 71418 58159 71434
tri 58159 71418 58175 71434 nw
rect 58211 71401 58268 71635
rect 58194 71319 58268 71401
rect 58082 71286 58159 71302
tri 58159 71286 58175 71302 sw
rect 58082 71220 58175 71286
rect 58211 71161 58268 71319
rect 58082 71085 58268 71161
rect 58082 70960 58175 71026
rect 58082 70944 58159 70960
tri 58159 70944 58175 70960 nw
rect 58211 70927 58268 71085
rect 58194 70845 58268 70927
rect 58082 70812 58159 70828
tri 58159 70812 58175 70828 sw
rect 58082 70746 58175 70812
rect 58082 70644 58175 70710
rect 58082 70628 58159 70644
tri 58159 70628 58175 70644 nw
rect 58211 70611 58268 70845
rect 58194 70529 58268 70611
rect 58082 70496 58159 70512
tri 58159 70496 58175 70512 sw
rect 58082 70430 58175 70496
rect 58211 70371 58268 70529
rect 58082 70295 58268 70371
rect 58082 70170 58175 70236
rect 58082 70154 58159 70170
tri 58159 70154 58175 70170 nw
rect 58211 70137 58268 70295
rect 58194 70055 58268 70137
rect 58082 70022 58159 70038
tri 58159 70022 58175 70038 sw
rect 58082 69956 58175 70022
rect 58082 69854 58175 69920
rect 58082 69838 58159 69854
tri 58159 69838 58175 69854 nw
rect 58211 69821 58268 70055
rect 58194 69739 58268 69821
rect 58082 69706 58159 69722
tri 58159 69706 58175 69722 sw
rect 58082 69640 58175 69706
rect 58211 69581 58268 69739
rect 58082 69505 58268 69581
rect 58082 69380 58175 69446
rect 58082 69364 58159 69380
tri 58159 69364 58175 69380 nw
rect 58211 69347 58268 69505
rect 58194 69265 58268 69347
rect 58082 69232 58159 69248
tri 58159 69232 58175 69248 sw
rect 58082 69166 58175 69232
rect 58082 69064 58175 69130
rect 58082 69048 58159 69064
tri 58159 69048 58175 69064 nw
rect 58211 69031 58268 69265
rect 58194 68949 58268 69031
rect 58082 68916 58159 68932
tri 58159 68916 58175 68932 sw
rect 58082 68850 58175 68916
rect 58211 68791 58268 68949
rect 58082 68715 58268 68791
rect 58082 68590 58175 68656
rect 58082 68574 58159 68590
tri 58159 68574 58175 68590 nw
rect 58211 68557 58268 68715
rect 58194 68475 58268 68557
rect 58082 68442 58159 68458
tri 58159 68442 58175 68458 sw
rect 58082 68376 58175 68442
rect 58082 68274 58175 68340
rect 58082 68258 58159 68274
tri 58159 68258 58175 68274 nw
rect 58211 68241 58268 68475
rect 58194 68159 58268 68241
rect 58082 68126 58159 68142
tri 58159 68126 58175 68142 sw
rect 58082 68060 58175 68126
rect 58211 68001 58268 68159
rect 58082 67925 58268 68001
rect 58082 67800 58175 67866
rect 58082 67784 58159 67800
tri 58159 67784 58175 67800 nw
rect 58211 67767 58268 67925
rect 58194 67685 58268 67767
rect 58082 67652 58159 67668
tri 58159 67652 58175 67668 sw
rect 58082 67586 58175 67652
rect 58082 67484 58175 67550
rect 58082 67468 58159 67484
tri 58159 67468 58175 67484 nw
rect 58211 67451 58268 67685
rect 58194 67369 58268 67451
rect 58082 67336 58159 67352
tri 58159 67336 58175 67352 sw
rect 58082 67270 58175 67336
rect 58211 67211 58268 67369
rect 58082 67135 58268 67211
rect 58082 67010 58175 67076
rect 58082 66994 58159 67010
tri 58159 66994 58175 67010 nw
rect 58211 66977 58268 67135
rect 58194 66895 58268 66977
rect 58082 66862 58159 66878
tri 58159 66862 58175 66878 sw
rect 58082 66796 58175 66862
rect 58082 66694 58175 66760
rect 58082 66678 58159 66694
tri 58159 66678 58175 66694 nw
rect 58211 66661 58268 66895
rect 58194 66579 58268 66661
rect 58082 66546 58159 66562
tri 58159 66546 58175 66562 sw
rect 58082 66480 58175 66546
rect 58211 66421 58268 66579
rect 58082 66345 58268 66421
rect 58082 66220 58175 66286
rect 58082 66204 58159 66220
tri 58159 66204 58175 66220 nw
rect 58211 66187 58268 66345
rect 58194 66105 58268 66187
rect 58082 66072 58159 66088
tri 58159 66072 58175 66088 sw
rect 58082 66006 58175 66072
rect 58082 65904 58175 65970
rect 58082 65888 58159 65904
tri 58159 65888 58175 65904 nw
rect 58211 65871 58268 66105
rect 58194 65789 58268 65871
rect 58082 65756 58159 65772
tri 58159 65756 58175 65772 sw
rect 58082 65690 58175 65756
rect 58211 65631 58268 65789
rect 58082 65555 58268 65631
rect 58082 65430 58175 65496
rect 58082 65414 58159 65430
tri 58159 65414 58175 65430 nw
rect 58211 65397 58268 65555
rect 58194 65315 58268 65397
rect 58082 65282 58159 65298
tri 58159 65282 58175 65298 sw
rect 58082 65216 58175 65282
rect 58082 65114 58175 65180
rect 58082 65098 58159 65114
tri 58159 65098 58175 65114 nw
rect 58211 65081 58268 65315
rect 58194 64999 58268 65081
rect 58082 64966 58159 64982
tri 58159 64966 58175 64982 sw
rect 58082 64900 58175 64966
rect 58211 64841 58268 64999
rect 58082 64765 58268 64841
rect 58082 64640 58175 64706
rect 58082 64624 58159 64640
tri 58159 64624 58175 64640 nw
rect 58211 64607 58268 64765
rect 58194 64525 58268 64607
rect 58082 64492 58159 64508
tri 58159 64492 58175 64508 sw
rect 58082 64426 58175 64492
rect 58082 64324 58175 64390
rect 58082 64308 58159 64324
tri 58159 64308 58175 64324 nw
rect 58211 64291 58268 64525
rect 58194 64209 58268 64291
rect 58082 64176 58159 64192
tri 58159 64176 58175 64192 sw
rect 58082 64110 58175 64176
rect 58211 64051 58268 64209
rect 58082 63975 58268 64051
rect 58082 63850 58175 63916
rect 58082 63834 58159 63850
tri 58159 63834 58175 63850 nw
rect 58211 63817 58268 63975
rect 58194 63735 58268 63817
rect 58082 63702 58159 63718
tri 58159 63702 58175 63718 sw
rect 58082 63636 58175 63702
rect 58082 63534 58175 63600
rect 58082 63518 58159 63534
tri 58159 63518 58175 63534 nw
rect 58211 63501 58268 63735
rect 58194 63419 58268 63501
rect 58082 63386 58159 63402
tri 58159 63386 58175 63402 sw
rect 58082 63320 58175 63386
rect 58211 63261 58268 63419
rect 58082 63185 58268 63261
rect 58082 63060 58175 63126
rect 58082 63044 58159 63060
tri 58159 63044 58175 63060 nw
rect 58211 63027 58268 63185
rect 58194 62945 58268 63027
rect 58082 62912 58159 62928
tri 58159 62912 58175 62928 sw
rect 58082 62846 58175 62912
rect 58082 62744 58175 62810
rect 58082 62728 58159 62744
tri 58159 62728 58175 62744 nw
rect 58211 62711 58268 62945
rect 58194 62629 58268 62711
rect 58082 62596 58159 62612
tri 58159 62596 58175 62612 sw
rect 58082 62530 58175 62596
rect 58211 62471 58268 62629
rect 58082 62395 58268 62471
rect 58082 62270 58175 62336
rect 58082 62254 58159 62270
tri 58159 62254 58175 62270 nw
rect 58211 62237 58268 62395
rect 58194 62155 58268 62237
rect 58082 62122 58159 62138
tri 58159 62122 58175 62138 sw
rect 58082 62056 58175 62122
rect 58082 61954 58175 62020
rect 58082 61938 58159 61954
tri 58159 61938 58175 61954 nw
rect 58211 61921 58268 62155
rect 58194 61839 58268 61921
rect 58082 61806 58159 61822
tri 58159 61806 58175 61822 sw
rect 58082 61740 58175 61806
rect 58211 61681 58268 61839
rect 58082 61605 58268 61681
rect 58082 61480 58175 61546
rect 58082 61464 58159 61480
tri 58159 61464 58175 61480 nw
rect 58211 61447 58268 61605
rect 58194 61365 58268 61447
rect 58082 61332 58159 61348
tri 58159 61332 58175 61348 sw
rect 58082 61266 58175 61332
rect 58082 61164 58175 61230
rect 58082 61148 58159 61164
tri 58159 61148 58175 61164 nw
rect 58211 61131 58268 61365
rect 58194 61049 58268 61131
rect 58082 61016 58159 61032
tri 58159 61016 58175 61032 sw
rect 58082 60950 58175 61016
rect 58211 60891 58268 61049
rect 58082 60815 58268 60891
rect 58082 60690 58175 60756
rect 58082 60674 58159 60690
tri 58159 60674 58175 60690 nw
rect 58211 60657 58268 60815
rect 58194 60575 58268 60657
rect 58082 60542 58159 60558
tri 58159 60542 58175 60558 sw
rect 58082 60476 58175 60542
rect 58082 60374 58175 60440
rect 58082 60358 58159 60374
tri 58159 60358 58175 60374 nw
rect 58211 60341 58268 60575
rect 58194 60259 58268 60341
rect 58082 60226 58159 60242
tri 58159 60226 58175 60242 sw
rect 58082 60160 58175 60226
rect 58211 60101 58268 60259
rect 58082 60025 58268 60101
rect 58082 59900 58175 59966
rect 58082 59884 58159 59900
tri 58159 59884 58175 59900 nw
rect 58211 59867 58268 60025
rect 58194 59785 58268 59867
rect 58082 59752 58159 59768
tri 58159 59752 58175 59768 sw
rect 58082 59686 58175 59752
rect 58082 59584 58175 59650
rect 58082 59568 58159 59584
tri 58159 59568 58175 59584 nw
rect 58211 59551 58268 59785
rect 58194 59469 58268 59551
rect 58082 59436 58159 59452
tri 58159 59436 58175 59452 sw
rect 58082 59370 58175 59436
rect 58211 59311 58268 59469
rect 58082 59235 58268 59311
rect 58082 59110 58175 59176
rect 58082 59094 58159 59110
tri 58159 59094 58175 59110 nw
rect 58211 59077 58268 59235
rect 58194 58995 58268 59077
rect 58082 58962 58159 58978
tri 58159 58962 58175 58978 sw
rect 58082 58896 58175 58962
rect 58082 58794 58175 58860
rect 58082 58778 58159 58794
tri 58159 58778 58175 58794 nw
rect 58211 58761 58268 58995
rect 58194 58679 58268 58761
rect 58082 58646 58159 58662
tri 58159 58646 58175 58662 sw
rect 58082 58580 58175 58646
rect 58211 58521 58268 58679
rect 58082 58445 58268 58521
rect 58082 58320 58175 58386
rect 58082 58304 58159 58320
tri 58159 58304 58175 58320 nw
rect 58211 58287 58268 58445
rect 58194 58205 58268 58287
rect 58082 58172 58159 58188
tri 58159 58172 58175 58188 sw
rect 58082 58106 58175 58172
rect 58082 58004 58175 58070
rect 58082 57988 58159 58004
tri 58159 57988 58175 58004 nw
rect 58211 57971 58268 58205
rect 58194 57889 58268 57971
rect 58082 57856 58159 57872
tri 58159 57856 58175 57872 sw
rect 58082 57790 58175 57856
rect 58211 57731 58268 57889
rect 58082 57655 58268 57731
rect 58082 57530 58175 57596
rect 58082 57514 58159 57530
tri 58159 57514 58175 57530 nw
rect 58211 57497 58268 57655
rect 58194 57415 58268 57497
rect 58082 57382 58159 57398
tri 58159 57382 58175 57398 sw
rect 58082 57316 58175 57382
rect 58082 57214 58175 57280
rect 58082 57198 58159 57214
tri 58159 57198 58175 57214 nw
rect 58211 57181 58268 57415
rect 58194 57099 58268 57181
rect 58082 57066 58159 57082
tri 58159 57066 58175 57082 sw
rect 58082 57000 58175 57066
rect 58211 56941 58268 57099
rect 58082 56865 58268 56941
rect 58082 56740 58175 56806
rect 58082 56724 58159 56740
tri 58159 56724 58175 56740 nw
rect 58211 56707 58268 56865
rect 58194 56625 58268 56707
rect 58082 56592 58159 56608
tri 58159 56592 58175 56608 sw
rect 58082 56526 58175 56592
rect 58082 56424 58175 56490
rect 58082 56408 58159 56424
tri 58159 56408 58175 56424 nw
rect 58211 56391 58268 56625
rect 58194 56309 58268 56391
rect 58082 56276 58159 56292
tri 58159 56276 58175 56292 sw
rect 58082 56210 58175 56276
rect 58211 56151 58268 56309
rect 58082 56075 58268 56151
rect 58082 55950 58175 56016
rect 58082 55934 58159 55950
tri 58159 55934 58175 55950 nw
rect 58211 55917 58268 56075
rect 58194 55835 58268 55917
rect 58082 55802 58159 55818
tri 58159 55802 58175 55818 sw
rect 58082 55736 58175 55802
rect 58082 55634 58175 55700
rect 58082 55618 58159 55634
tri 58159 55618 58175 55634 nw
rect 58211 55601 58268 55835
rect 58194 55519 58268 55601
rect 58082 55486 58159 55502
tri 58159 55486 58175 55502 sw
rect 58082 55420 58175 55486
rect 58211 55361 58268 55519
rect 58082 55285 58268 55361
rect 58082 55160 58175 55226
rect 58082 55144 58159 55160
tri 58159 55144 58175 55160 nw
rect 58211 55127 58268 55285
rect 58194 55045 58268 55127
rect 58082 55012 58159 55028
tri 58159 55012 58175 55028 sw
rect 58082 54946 58175 55012
rect 58082 54844 58175 54910
rect 58082 54828 58159 54844
tri 58159 54828 58175 54844 nw
rect 58211 54811 58268 55045
rect 58194 54729 58268 54811
rect 58082 54696 58159 54712
tri 58159 54696 58175 54712 sw
rect 58082 54630 58175 54696
rect 58211 54571 58268 54729
rect 58082 54495 58268 54571
rect 58082 54370 58175 54436
rect 58082 54354 58159 54370
tri 58159 54354 58175 54370 nw
rect 58211 54337 58268 54495
rect 58194 54255 58268 54337
rect 58082 54222 58159 54238
tri 58159 54222 58175 54238 sw
rect 58082 54156 58175 54222
rect 58082 54054 58175 54120
rect 58082 54038 58159 54054
tri 58159 54038 58175 54054 nw
rect 58211 54021 58268 54255
rect 58194 53939 58268 54021
rect 58082 53906 58159 53922
tri 58159 53906 58175 53922 sw
rect 58082 53840 58175 53906
rect 58211 53781 58268 53939
rect 58082 53705 58268 53781
rect 58082 53580 58175 53646
rect 58082 53564 58159 53580
tri 58159 53564 58175 53580 nw
rect 58211 53547 58268 53705
rect 58194 53465 58268 53547
rect 58082 53432 58159 53448
tri 58159 53432 58175 53448 sw
rect 58082 53366 58175 53432
rect 58082 53264 58175 53330
rect 58082 53248 58159 53264
tri 58159 53248 58175 53264 nw
rect 58211 53231 58268 53465
rect 58194 53149 58268 53231
rect 58082 53116 58159 53132
tri 58159 53116 58175 53132 sw
rect 58082 53050 58175 53116
rect 58211 52991 58268 53149
rect 58082 52915 58268 52991
rect 58082 52790 58175 52856
rect 58082 52774 58159 52790
tri 58159 52774 58175 52790 nw
rect 58211 52757 58268 52915
rect 58194 52675 58268 52757
rect 58082 52642 58159 52658
tri 58159 52642 58175 52658 sw
rect 58082 52576 58175 52642
rect 58082 52474 58175 52540
rect 58082 52458 58159 52474
tri 58159 52458 58175 52474 nw
rect 58211 52441 58268 52675
rect 58194 52359 58268 52441
rect 58082 52326 58159 52342
tri 58159 52326 58175 52342 sw
rect 58082 52260 58175 52326
rect 58211 52201 58268 52359
rect 58082 52125 58268 52201
rect 58082 52000 58175 52066
rect 58082 51984 58159 52000
tri 58159 51984 58175 52000 nw
rect 58211 51967 58268 52125
rect 58194 51885 58268 51967
rect 58082 51852 58159 51868
tri 58159 51852 58175 51868 sw
rect 58082 51786 58175 51852
rect 58082 51684 58175 51750
rect 58082 51668 58159 51684
tri 58159 51668 58175 51684 nw
rect 58211 51651 58268 51885
rect 58194 51569 58268 51651
rect 58082 51536 58159 51552
tri 58159 51536 58175 51552 sw
rect 58082 51470 58175 51536
rect 58211 51411 58268 51569
rect 58082 51335 58268 51411
rect 58082 51210 58175 51276
rect 58082 51194 58159 51210
tri 58159 51194 58175 51210 nw
rect 58211 51177 58268 51335
rect 58194 51095 58268 51177
rect 58082 51062 58159 51078
tri 58159 51062 58175 51078 sw
rect 58082 50996 58175 51062
rect 58082 50894 58175 50960
rect 58082 50878 58159 50894
tri 58159 50878 58175 50894 nw
rect 58211 50861 58268 51095
rect 58194 50779 58268 50861
rect 58082 50746 58159 50762
tri 58159 50746 58175 50762 sw
rect 58082 50680 58175 50746
rect 58211 50621 58268 50779
rect 58082 50545 58268 50621
rect 58082 50420 58175 50486
rect 58082 50404 58159 50420
tri 58159 50404 58175 50420 nw
rect 58211 50387 58268 50545
rect 58194 50305 58268 50387
rect 58082 50272 58159 50288
tri 58159 50272 58175 50288 sw
rect 58082 50206 58175 50272
rect 58082 50104 58175 50170
rect 58082 50088 58159 50104
tri 58159 50088 58175 50104 nw
rect 58211 50071 58268 50305
rect 58194 49989 58268 50071
rect 58082 49956 58159 49972
tri 58159 49956 58175 49972 sw
rect 58082 49890 58175 49956
rect 58211 49831 58268 49989
rect 58082 49755 58268 49831
rect 58082 49630 58175 49696
rect 58082 49614 58159 49630
tri 58159 49614 58175 49630 nw
rect 58211 49597 58268 49755
rect 58194 49515 58268 49597
rect 58082 49482 58159 49498
tri 58159 49482 58175 49498 sw
rect 58082 49416 58175 49482
rect 58082 49314 58175 49380
rect 58082 49298 58159 49314
tri 58159 49298 58175 49314 nw
rect 58211 49281 58268 49515
rect 58194 49199 58268 49281
rect 58082 49166 58159 49182
tri 58159 49166 58175 49182 sw
rect 58082 49100 58175 49166
rect 58211 49041 58268 49199
rect 58082 48965 58268 49041
rect 58082 48840 58175 48906
rect 58082 48824 58159 48840
tri 58159 48824 58175 48840 nw
rect 58211 48807 58268 48965
rect 58194 48725 58268 48807
rect 58082 48692 58159 48708
tri 58159 48692 58175 48708 sw
rect 58082 48626 58175 48692
rect 58082 48524 58175 48590
rect 58082 48508 58159 48524
tri 58159 48508 58175 48524 nw
rect 58211 48491 58268 48725
rect 58194 48409 58268 48491
rect 58082 48376 58159 48392
tri 58159 48376 58175 48392 sw
rect 58082 48310 58175 48376
rect 58211 48251 58268 48409
rect 58082 48175 58268 48251
rect 58082 48050 58175 48116
rect 58082 48034 58159 48050
tri 58159 48034 58175 48050 nw
rect 58211 48017 58268 48175
rect 58194 47935 58268 48017
rect 58082 47902 58159 47918
tri 58159 47902 58175 47918 sw
rect 58082 47836 58175 47902
rect 58082 47734 58175 47800
rect 58082 47718 58159 47734
tri 58159 47718 58175 47734 nw
rect 58211 47701 58268 47935
rect 58194 47619 58268 47701
rect 58082 47586 58159 47602
tri 58159 47586 58175 47602 sw
rect 58082 47520 58175 47586
rect 58211 47461 58268 47619
rect 58082 47385 58268 47461
rect 58082 47260 58175 47326
rect 58082 47244 58159 47260
tri 58159 47244 58175 47260 nw
rect 58211 47227 58268 47385
rect 58194 47145 58268 47227
rect 58082 47112 58159 47128
tri 58159 47112 58175 47128 sw
rect 58082 47046 58175 47112
rect 58082 46944 58175 47010
rect 58082 46928 58159 46944
tri 58159 46928 58175 46944 nw
rect 58211 46911 58268 47145
rect 58194 46829 58268 46911
rect 58082 46796 58159 46812
tri 58159 46796 58175 46812 sw
rect 58082 46730 58175 46796
rect 58211 46671 58268 46829
rect 58082 46595 58268 46671
rect 58082 46470 58175 46536
rect 58082 46454 58159 46470
tri 58159 46454 58175 46470 nw
rect 58211 46437 58268 46595
rect 58194 46355 58268 46437
rect 58082 46322 58159 46338
tri 58159 46322 58175 46338 sw
rect 58082 46256 58175 46322
rect 58082 46154 58175 46220
rect 58082 46138 58159 46154
tri 58159 46138 58175 46154 nw
rect 58211 46121 58268 46355
rect 58194 46039 58268 46121
rect 58082 46006 58159 46022
tri 58159 46006 58175 46022 sw
rect 58082 45940 58175 46006
rect 58211 45881 58268 46039
rect 58082 45805 58268 45881
rect 58082 45680 58175 45746
rect 58082 45664 58159 45680
tri 58159 45664 58175 45680 nw
rect 58211 45647 58268 45805
rect 58194 45565 58268 45647
rect 58082 45532 58159 45548
tri 58159 45532 58175 45548 sw
rect 58082 45466 58175 45532
rect 58082 45364 58175 45430
rect 58082 45348 58159 45364
tri 58159 45348 58175 45364 nw
rect 58211 45331 58268 45565
rect 58194 45249 58268 45331
rect 58082 45216 58159 45232
tri 58159 45216 58175 45232 sw
rect 58082 45150 58175 45216
rect 58211 45091 58268 45249
rect 58082 45015 58268 45091
rect 58082 44890 58175 44956
rect 58082 44874 58159 44890
tri 58159 44874 58175 44890 nw
rect 58211 44857 58268 45015
rect 58194 44775 58268 44857
rect 58082 44742 58159 44758
tri 58159 44742 58175 44758 sw
rect 58082 44676 58175 44742
rect 58082 44574 58175 44640
rect 58082 44558 58159 44574
tri 58159 44558 58175 44574 nw
rect 58211 44541 58268 44775
rect 58194 44459 58268 44541
rect 58082 44426 58159 44442
tri 58159 44426 58175 44442 sw
rect 58082 44360 58175 44426
rect 58211 44301 58268 44459
rect 58082 44225 58268 44301
rect 58082 44100 58175 44166
rect 58082 44084 58159 44100
tri 58159 44084 58175 44100 nw
rect 58211 44067 58268 44225
rect 58194 43985 58268 44067
rect 58082 43952 58159 43968
tri 58159 43952 58175 43968 sw
rect 58082 43886 58175 43952
rect 58082 43784 58175 43850
rect 58082 43768 58159 43784
tri 58159 43768 58175 43784 nw
rect 58211 43751 58268 43985
rect 58194 43669 58268 43751
rect 58082 43636 58159 43652
tri 58159 43636 58175 43652 sw
rect 58082 43570 58175 43636
rect 58211 43511 58268 43669
rect 58082 43435 58268 43511
rect 58082 43310 58175 43376
rect 58082 43294 58159 43310
tri 58159 43294 58175 43310 nw
rect 58211 43277 58268 43435
rect 58194 43195 58268 43277
rect 58082 43162 58159 43178
tri 58159 43162 58175 43178 sw
rect 58082 43096 58175 43162
rect 58082 42994 58175 43060
rect 58082 42978 58159 42994
tri 58159 42978 58175 42994 nw
rect 58211 42961 58268 43195
rect 58194 42879 58268 42961
rect 58082 42846 58159 42862
tri 58159 42846 58175 42862 sw
rect 58082 42780 58175 42846
rect 58211 42721 58268 42879
rect 58082 42645 58268 42721
rect 58082 42520 58175 42586
rect 58082 42504 58159 42520
tri 58159 42504 58175 42520 nw
rect 58211 42487 58268 42645
rect 58194 42405 58268 42487
rect 58082 42372 58159 42388
tri 58159 42372 58175 42388 sw
rect 58082 42306 58175 42372
rect 58082 42204 58175 42270
rect 58082 42188 58159 42204
tri 58159 42188 58175 42204 nw
rect 58211 42171 58268 42405
rect 58194 42089 58268 42171
rect 58082 42056 58159 42072
tri 58159 42056 58175 42072 sw
rect 58082 41990 58175 42056
rect 58211 41931 58268 42089
rect 58082 41855 58268 41931
rect 58082 41730 58175 41796
rect 58082 41714 58159 41730
tri 58159 41714 58175 41730 nw
rect 58211 41697 58268 41855
rect 58194 41615 58268 41697
rect 58082 41582 58159 41598
tri 58159 41582 58175 41598 sw
rect 58082 41516 58175 41582
rect 58082 41414 58175 41480
rect 58082 41398 58159 41414
tri 58159 41398 58175 41414 nw
rect 58211 41381 58268 41615
rect 58194 41299 58268 41381
rect 58082 41266 58159 41282
tri 58159 41266 58175 41282 sw
rect 58082 41200 58175 41266
rect 58211 41141 58268 41299
rect 58082 41065 58268 41141
rect 58082 40940 58175 41006
rect 58082 40924 58159 40940
tri 58159 40924 58175 40940 nw
rect 58211 40907 58268 41065
rect 58194 40825 58268 40907
rect 58082 40792 58159 40808
tri 58159 40792 58175 40808 sw
rect 58082 40726 58175 40792
rect 58082 40624 58175 40690
rect 58082 40608 58159 40624
tri 58159 40608 58175 40624 nw
rect 58211 40591 58268 40825
rect 58194 40509 58268 40591
rect 58082 40476 58159 40492
tri 58159 40476 58175 40492 sw
rect 58082 40410 58175 40476
rect 58211 40351 58268 40509
rect 58082 40275 58268 40351
rect 58082 40150 58175 40216
rect 58082 40134 58159 40150
tri 58159 40134 58175 40150 nw
rect 58211 40117 58268 40275
rect 58194 40035 58268 40117
rect 58082 40002 58159 40018
tri 58159 40002 58175 40018 sw
rect 58082 39936 58175 40002
rect 58082 39834 58175 39900
rect 58082 39818 58159 39834
tri 58159 39818 58175 39834 nw
rect 58211 39801 58268 40035
rect 58194 39719 58268 39801
rect 58082 39686 58159 39702
tri 58159 39686 58175 39702 sw
rect 58082 39620 58175 39686
rect 58211 39561 58268 39719
rect 58082 39485 58268 39561
rect 58082 39360 58175 39426
rect 58082 39344 58159 39360
tri 58159 39344 58175 39360 nw
rect 58211 39327 58268 39485
rect 58194 39245 58268 39327
rect 58082 39212 58159 39228
tri 58159 39212 58175 39228 sw
rect 58082 39146 58175 39212
rect 58082 39044 58175 39110
rect 58082 39028 58159 39044
tri 58159 39028 58175 39044 nw
rect 58211 39011 58268 39245
rect 58194 38929 58268 39011
rect 58082 38896 58159 38912
tri 58159 38896 58175 38912 sw
rect 58082 38830 58175 38896
rect 58211 38771 58268 38929
rect 58082 38695 58268 38771
rect 58082 38570 58175 38636
rect 58082 38554 58159 38570
tri 58159 38554 58175 38570 nw
rect 58211 38537 58268 38695
rect 58194 38455 58268 38537
rect 58082 38422 58159 38438
tri 58159 38422 58175 38438 sw
rect 58082 38356 58175 38422
rect 58082 38254 58175 38320
rect 58082 38238 58159 38254
tri 58159 38238 58175 38254 nw
rect 58211 38221 58268 38455
rect 58194 38139 58268 38221
rect 58082 38106 58159 38122
tri 58159 38106 58175 38122 sw
rect 58082 38040 58175 38106
rect 58211 37981 58268 38139
rect 58082 37905 58268 37981
rect 58082 37780 58175 37846
rect 58082 37764 58159 37780
tri 58159 37764 58175 37780 nw
rect 58211 37747 58268 37905
rect 58194 37665 58268 37747
rect 58082 37632 58159 37648
tri 58159 37632 58175 37648 sw
rect 58082 37566 58175 37632
rect 58082 37464 58175 37530
rect 58082 37448 58159 37464
tri 58159 37448 58175 37464 nw
rect 58211 37431 58268 37665
rect 58194 37349 58268 37431
rect 58082 37316 58159 37332
tri 58159 37316 58175 37332 sw
rect 58082 37250 58175 37316
rect 58211 37191 58268 37349
rect 58082 37115 58268 37191
rect 58082 36990 58175 37056
rect 58082 36974 58159 36990
tri 58159 36974 58175 36990 nw
rect 58211 36957 58268 37115
rect 58194 36875 58268 36957
rect 58082 36842 58159 36858
tri 58159 36842 58175 36858 sw
rect 58082 36776 58175 36842
rect 58082 36674 58175 36740
rect 58082 36658 58159 36674
tri 58159 36658 58175 36674 nw
rect 58211 36641 58268 36875
rect 58194 36559 58268 36641
rect 58082 36526 58159 36542
tri 58159 36526 58175 36542 sw
rect 58082 36460 58175 36526
rect 58211 36401 58268 36559
rect 58082 36325 58268 36401
rect 58082 36200 58175 36266
rect 58082 36184 58159 36200
tri 58159 36184 58175 36200 nw
rect 58211 36167 58268 36325
rect 58194 36085 58268 36167
rect 58082 36052 58159 36068
tri 58159 36052 58175 36068 sw
rect 58082 35986 58175 36052
rect 58082 35884 58175 35950
rect 58082 35868 58159 35884
tri 58159 35868 58175 35884 nw
rect 58211 35851 58268 36085
rect 58194 35769 58268 35851
rect 58082 35736 58159 35752
tri 58159 35736 58175 35752 sw
rect 58082 35670 58175 35736
rect 58211 35611 58268 35769
rect 58082 35535 58268 35611
rect 58082 35410 58175 35476
rect 58082 35394 58159 35410
tri 58159 35394 58175 35410 nw
rect 58211 35377 58268 35535
rect 58194 35295 58268 35377
rect 58082 35262 58159 35278
tri 58159 35262 58175 35278 sw
rect 58082 35196 58175 35262
rect 58082 35094 58175 35160
rect 58082 35078 58159 35094
tri 58159 35078 58175 35094 nw
rect 58211 35061 58268 35295
rect 58194 34979 58268 35061
rect 58082 34946 58159 34962
tri 58159 34946 58175 34962 sw
rect 58082 34880 58175 34946
rect 58211 34821 58268 34979
rect 58082 34745 58268 34821
rect 58082 34620 58175 34686
rect 58082 34604 58159 34620
tri 58159 34604 58175 34620 nw
rect 58211 34587 58268 34745
rect 58194 34505 58268 34587
rect 58082 34472 58159 34488
tri 58159 34472 58175 34488 sw
rect 58082 34406 58175 34472
rect 58082 34304 58175 34370
rect 58082 34288 58159 34304
tri 58159 34288 58175 34304 nw
rect 58211 34271 58268 34505
rect 58194 34189 58268 34271
rect 58082 34156 58159 34172
tri 58159 34156 58175 34172 sw
rect 58082 34090 58175 34156
rect 58211 34031 58268 34189
rect 58082 33955 58268 34031
rect 58082 33830 58175 33896
rect 58082 33814 58159 33830
tri 58159 33814 58175 33830 nw
rect 58211 33797 58268 33955
rect 58194 33715 58268 33797
rect 58082 33682 58159 33698
tri 58159 33682 58175 33698 sw
rect 58082 33616 58175 33682
rect 58082 33514 58175 33580
rect 58082 33498 58159 33514
tri 58159 33498 58175 33514 nw
rect 58211 33481 58268 33715
rect 58194 33399 58268 33481
rect 58082 33366 58159 33382
tri 58159 33366 58175 33382 sw
rect 58082 33300 58175 33366
rect 58211 33241 58268 33399
rect 58082 33165 58268 33241
rect 58082 33040 58175 33106
rect 58082 33024 58159 33040
tri 58159 33024 58175 33040 nw
rect 58211 33007 58268 33165
rect 58194 32925 58268 33007
rect 58082 32892 58159 32908
tri 58159 32892 58175 32908 sw
rect 58082 32826 58175 32892
rect 58082 32724 58175 32790
rect 58082 32708 58159 32724
tri 58159 32708 58175 32724 nw
rect 58211 32691 58268 32925
rect 58194 32609 58268 32691
rect 58082 32576 58159 32592
tri 58159 32576 58175 32592 sw
rect 58082 32510 58175 32576
rect 58211 32451 58268 32609
rect 58082 32375 58268 32451
rect 58082 32250 58175 32316
rect 58082 32234 58159 32250
tri 58159 32234 58175 32250 nw
rect 58211 32217 58268 32375
rect 58194 32135 58268 32217
rect 58082 32102 58159 32118
tri 58159 32102 58175 32118 sw
rect 58082 32036 58175 32102
rect 58082 31934 58175 32000
rect 58082 31918 58159 31934
tri 58159 31918 58175 31934 nw
rect 58211 31901 58268 32135
rect 58194 31819 58268 31901
rect 58082 31786 58159 31802
tri 58159 31786 58175 31802 sw
rect 58082 31720 58175 31786
rect 58211 31661 58268 31819
rect 58082 31585 58268 31661
rect 58082 31460 58175 31526
rect 58082 31444 58159 31460
tri 58159 31444 58175 31460 nw
rect 58211 31427 58268 31585
rect 58194 31345 58268 31427
rect 58082 31312 58159 31328
tri 58159 31312 58175 31328 sw
rect 58082 31246 58175 31312
rect 58082 31144 58175 31210
rect 58082 31128 58159 31144
tri 58159 31128 58175 31144 nw
rect 58211 31111 58268 31345
rect 58194 31029 58268 31111
rect 58082 30996 58159 31012
tri 58159 30996 58175 31012 sw
rect 58082 30930 58175 30996
rect 58211 30871 58268 31029
rect 58082 30795 58268 30871
rect 58082 30670 58175 30736
rect 58082 30654 58159 30670
tri 58159 30654 58175 30670 nw
rect 58211 30637 58268 30795
rect 58194 30555 58268 30637
rect 58082 30522 58159 30538
tri 58159 30522 58175 30538 sw
rect 58082 30456 58175 30522
rect 58082 30354 58175 30420
rect 58082 30338 58159 30354
tri 58159 30338 58175 30354 nw
rect 58211 30321 58268 30555
rect 58194 30239 58268 30321
rect 58082 30206 58159 30222
tri 58159 30206 58175 30222 sw
rect 58082 30140 58175 30206
rect 58211 30081 58268 30239
rect 58082 30005 58268 30081
rect 58082 29880 58175 29946
rect 58082 29864 58159 29880
tri 58159 29864 58175 29880 nw
rect 58211 29847 58268 30005
rect 58194 29765 58268 29847
rect 58082 29732 58159 29748
tri 58159 29732 58175 29748 sw
rect 58082 29666 58175 29732
rect 58082 29564 58175 29630
rect 58082 29548 58159 29564
tri 58159 29548 58175 29564 nw
rect 58211 29531 58268 29765
rect 58194 29449 58268 29531
rect 58082 29416 58159 29432
tri 58159 29416 58175 29432 sw
rect 58082 29350 58175 29416
rect 58211 29291 58268 29449
rect 58082 29215 58268 29291
rect 59902 29253 59930 79813
rect 61426 29253 61454 79813
rect 62458 29221 62508 79845
rect 62884 29223 62932 79843
rect 63340 29282 63368 79842
rect 63612 29282 63640 79842
rect 63984 79066 64032 79828
rect 64416 79066 64464 79828
rect 63984 78276 64032 79038
rect 64416 78276 64464 79038
rect 63984 77486 64032 78248
rect 64416 77486 64464 78248
rect 63984 76696 64032 77458
rect 64416 76696 64464 77458
rect 63984 75906 64032 76668
rect 64416 75906 64464 76668
rect 63984 75116 64032 75878
rect 64416 75116 64464 75878
rect 63984 74326 64032 75088
rect 64416 74326 64464 75088
rect 63984 73536 64032 74298
rect 64416 73536 64464 74298
rect 63984 72746 64032 73508
rect 64416 72746 64464 73508
rect 63984 71956 64032 72718
rect 64416 71956 64464 72718
rect 63984 71166 64032 71928
rect 64416 71166 64464 71928
rect 63984 70376 64032 71138
rect 64416 70376 64464 71138
rect 63984 69586 64032 70348
rect 64416 69586 64464 70348
rect 63984 68796 64032 69558
rect 64416 68796 64464 69558
rect 63984 68006 64032 68768
rect 64416 68006 64464 68768
rect 63984 67216 64032 67978
rect 64416 67216 64464 67978
rect 63984 66426 64032 67188
rect 64416 66426 64464 67188
rect 63984 65636 64032 66398
rect 64416 65636 64464 66398
rect 63984 64846 64032 65608
rect 64416 64846 64464 65608
rect 63984 64056 64032 64818
rect 64416 64056 64464 64818
rect 63984 63266 64032 64028
rect 64416 63266 64464 64028
rect 63984 62476 64032 63238
rect 64416 62476 64464 63238
rect 63984 61686 64032 62448
rect 64416 61686 64464 62448
rect 63984 60896 64032 61658
rect 64416 60896 64464 61658
rect 63984 60106 64032 60868
rect 64416 60106 64464 60868
rect 63984 59316 64032 60078
rect 64416 59316 64464 60078
rect 63984 58526 64032 59288
rect 64416 58526 64464 59288
rect 63984 57736 64032 58498
rect 64416 57736 64464 58498
rect 63984 56946 64032 57708
rect 64416 56946 64464 57708
rect 63984 56156 64032 56918
rect 64416 56156 64464 56918
rect 63984 55366 64032 56128
rect 64416 55366 64464 56128
rect 63984 54576 64032 55338
rect 64416 54576 64464 55338
rect 63984 53786 64032 54548
rect 64416 53786 64464 54548
rect 63984 52996 64032 53758
rect 64416 52996 64464 53758
rect 63984 52206 64032 52968
rect 64416 52206 64464 52968
rect 63984 51416 64032 52178
rect 64416 51416 64464 52178
rect 63984 50626 64032 51388
rect 64416 50626 64464 51388
rect 63984 49836 64032 50598
rect 64416 49836 64464 50598
rect 63984 49046 64032 49808
rect 64416 49046 64464 49808
rect 63984 48256 64032 49018
rect 64416 48256 64464 49018
rect 63984 47466 64032 48228
rect 64416 47466 64464 48228
rect 63984 46676 64032 47438
rect 64416 46676 64464 47438
rect 63984 45886 64032 46648
rect 64416 45886 64464 46648
rect 63984 45096 64032 45858
rect 64416 45096 64464 45858
rect 63984 44306 64032 45068
rect 64416 44306 64464 45068
rect 63984 43516 64032 44278
rect 64416 43516 64464 44278
rect 63984 42726 64032 43488
rect 64416 42726 64464 43488
rect 63984 41936 64032 42698
rect 64416 41936 64464 42698
rect 63984 41146 64032 41908
rect 64416 41146 64464 41908
rect 63984 40356 64032 41118
rect 64416 40356 64464 41118
rect 63984 39566 64032 40328
rect 64416 39566 64464 40328
rect 63984 38776 64032 39538
rect 64416 38776 64464 39538
rect 63984 37986 64032 38748
rect 64416 37986 64464 38748
rect 63984 37196 64032 37958
rect 64416 37196 64464 37958
rect 63984 36406 64032 37168
rect 64416 36406 64464 37168
rect 63984 35616 64032 36378
rect 64416 35616 64464 36378
rect 63984 34826 64032 35588
rect 64416 34826 64464 35588
rect 63984 34036 64032 34798
rect 64416 34036 64464 34798
rect 63984 33246 64032 34008
rect 64416 33246 64464 34008
rect 63984 32456 64032 33218
rect 64416 32456 64464 33218
rect 63984 31666 64032 32428
rect 64416 31666 64464 32428
rect 63984 30876 64032 31638
rect 64416 30876 64464 31638
rect 63984 30086 64032 30848
rect 64416 30086 64464 30848
rect 63984 29296 64032 30058
rect 64416 29296 64464 30058
rect 64842 29238 64888 79886
rect 66630 34022 66658 37182
rect 66902 34022 66930 37182
rect 67274 36406 67322 37168
rect 67706 36406 67754 37168
rect 67274 35616 67322 36378
rect 67706 35616 67754 36378
rect 67274 34826 67322 35588
rect 67706 34826 67754 35588
rect 67274 34036 67322 34798
rect 67706 34036 67754 34798
rect 68132 33978 68178 37226
rect 69200 34022 69228 35207
rect 69472 34022 69500 35207
rect 69804 34977 69856 35041
rect 69884 34583 69936 34647
rect 69964 34187 70016 34251
rect 66630 31652 66658 33232
rect 66902 31652 66930 33232
rect 67270 31620 67320 33264
rect 67696 31622 67744 33262
rect 68604 31652 68632 32442
rect 68876 31652 68904 32442
rect 69208 32213 69260 32277
rect 69288 31817 69340 31881
rect 66630 29282 66658 30862
rect 66902 29282 66930 30862
rect 67270 29250 67320 30894
rect 67696 29252 67744 30892
rect 68604 29282 68632 30072
rect 68876 29282 68904 30072
rect 69208 29843 69260 29907
rect 69288 29447 69340 29511
rect 70164 29282 70192 37182
rect 70244 29282 70272 37182
rect 70324 29282 70352 37182
rect 70404 29282 70432 37182
rect 70484 29282 70512 37182
rect 70564 29282 70592 37182
rect 70644 29282 70672 37182
rect 58082 29090 58175 29156
rect 58082 29074 58159 29090
tri 58159 29074 58175 29090 nw
rect 58211 29057 58268 29215
rect 58194 28975 58268 29057
rect 58082 28942 58159 28958
tri 58159 28942 58175 28958 sw
rect 58082 28876 58175 28942
rect 58211 28833 58268 28975
rect 70966 28709 71024 28755
rect 71156 28709 71214 28755
rect 71417 28709 71475 28755
rect 71767 28709 71825 28755
rect 72028 28709 72086 28755
rect 70978 28367 71012 28709
rect 71040 28466 71106 28518
rect 71168 28515 71202 28709
rect 71156 28469 71214 28515
rect 70962 28315 71028 28367
rect 17150 27457 17178 28211
rect 17614 27457 17642 28211
rect 17774 27457 17802 28211
rect 18238 27457 18266 28211
rect 18398 27457 18426 28211
rect 18862 27457 18890 28211
rect 19022 27457 19050 28211
rect 19486 27457 19514 28211
rect 19646 27457 19674 28211
rect 20110 27457 20138 28211
rect 20270 27457 20298 28211
rect 20734 27457 20762 28211
rect 20894 27457 20922 28211
rect 21358 27457 21386 28211
rect 21518 27457 21546 28211
rect 21982 27457 22010 28211
rect 22142 27457 22170 28211
rect 22606 27457 22634 28211
rect 22766 27457 22794 28211
rect 23230 27457 23258 28211
rect 23390 27457 23418 28211
rect 23854 27457 23882 28211
rect 24014 27457 24042 28211
rect 24478 27457 24506 28211
rect 24638 27457 24666 28211
rect 25102 27457 25130 28211
rect 25262 27457 25290 28211
rect 25726 27457 25754 28211
rect 25886 27457 25914 28211
rect 26350 27457 26378 28211
rect 26510 27457 26538 28211
rect 26974 27457 27002 28211
rect 27134 27457 27162 28211
rect 27598 27457 27626 28211
rect 27758 27457 27786 28211
rect 28222 27457 28250 28211
rect 28382 27457 28410 28211
rect 28846 27457 28874 28211
rect 29006 27457 29034 28211
rect 29470 27457 29498 28211
rect 29630 27457 29658 28211
rect 30094 27457 30122 28211
rect 30254 27457 30282 28211
rect 30718 27457 30746 28211
rect 30878 27457 30906 28211
rect 31342 27457 31370 28211
rect 31502 27457 31530 28211
rect 31966 27457 31994 28211
rect 32126 27457 32154 28211
rect 32590 27457 32618 28211
rect 32750 27457 32778 28211
rect 33214 27457 33242 28211
rect 33374 27457 33402 28211
rect 33838 27457 33866 28211
rect 33998 27457 34026 28211
rect 34462 27457 34490 28211
rect 34622 27457 34650 28211
rect 35086 27457 35114 28211
rect 35246 27457 35274 28211
rect 35710 27457 35738 28211
rect 35870 27457 35898 28211
rect 36334 27457 36362 28211
rect 36494 27457 36522 28211
rect 36958 27457 36986 28211
rect 37118 27457 37146 28211
rect 37582 27457 37610 28211
rect 37742 27457 37770 28211
rect 38206 27457 38234 28211
rect 38366 27457 38394 28211
rect 38830 27457 38858 28211
rect 38990 27457 39018 28211
rect 39454 27457 39482 28211
rect 39614 27457 39642 28211
rect 40078 27457 40106 28211
rect 40238 27457 40266 28211
rect 40702 27457 40730 28211
rect 40862 27457 40890 28211
rect 41326 27457 41354 28211
rect 41486 27457 41514 28211
rect 41950 27457 41978 28211
rect 42110 27457 42138 28211
rect 42574 27457 42602 28211
rect 42734 27457 42762 28211
rect 43198 27457 43226 28211
rect 43358 27457 43386 28211
rect 43822 27457 43850 28211
rect 43982 27457 44010 28211
rect 44446 27457 44474 28211
rect 44606 27457 44634 28211
rect 45070 27457 45098 28211
rect 45230 27457 45258 28211
rect 45694 27457 45722 28211
rect 45854 27457 45882 28211
rect 46318 27457 46346 28211
rect 46478 27457 46506 28211
rect 46942 27457 46970 28211
rect 47102 27457 47130 28211
rect 47566 27457 47594 28211
rect 47726 27457 47754 28211
rect 48190 27457 48218 28211
rect 48350 27457 48378 28211
rect 48814 27457 48842 28211
rect 48974 27457 49002 28211
rect 49438 27457 49466 28211
rect 49598 27457 49626 28211
rect 50062 27457 50090 28211
rect 50222 27457 50250 28211
rect 50686 27457 50714 28211
rect 50846 27457 50874 28211
rect 51310 27457 51338 28211
rect 51470 27457 51498 28211
rect 51934 27457 51962 28211
rect 52094 27457 52122 28211
rect 52558 27457 52586 28211
rect 52718 27457 52746 28211
rect 53182 27457 53210 28211
rect 53342 27457 53370 28211
rect 53806 27457 53834 28211
rect 53966 27457 53994 28211
rect 54430 27457 54458 28211
rect 54590 27457 54618 28211
rect 55054 27457 55082 28211
rect 55214 27457 55242 28211
rect 55678 27457 55706 28211
rect 55838 27457 55866 28211
rect 56302 27457 56330 28211
rect 56462 27457 56490 28211
rect 56926 27457 56954 28211
rect 57086 27457 57114 28211
rect 57550 27457 57578 28211
rect 70978 28195 71012 28315
rect 71168 28195 71202 28469
rect 71429 28195 71463 28709
rect 71687 28595 71741 28604
rect 71685 28549 71743 28595
rect 71687 28540 71741 28549
rect 71697 28284 71731 28540
rect 71779 28349 71813 28709
rect 72040 28515 72074 28709
rect 72028 28469 72086 28515
rect 71907 28386 71973 28438
rect 71951 28349 72009 28355
rect 71779 28315 72009 28349
rect 71687 28275 71741 28284
rect 71685 28229 71743 28275
rect 71687 28220 71741 28229
rect 71779 28195 71813 28315
rect 71951 28309 72009 28315
rect 72040 28195 72074 28469
rect 70966 28149 71024 28195
rect 71156 28149 71214 28195
rect 71417 28149 71475 28195
rect 71767 28149 71825 28195
rect 72028 28149 72086 28195
rect 17788 27149 17816 27205
rect 18252 27149 18280 27205
rect 18384 27149 18412 27205
rect 18848 27149 18876 27205
rect 19036 27149 19064 27205
rect 19500 27149 19528 27205
rect 19632 27149 19660 27205
rect 20096 27149 20124 27205
rect 20284 27149 20312 27205
rect 20748 27149 20776 27205
rect 20880 27149 20908 27205
rect 21344 27149 21372 27205
rect 21532 27149 21560 27205
rect 21996 27149 22024 27205
rect 22128 27149 22156 27205
rect 22592 27149 22620 27205
rect 22780 27149 22808 27205
rect 23244 27149 23272 27205
rect 23376 27149 23404 27205
rect 23840 27149 23868 27205
rect 24028 27149 24056 27205
rect 24492 27149 24520 27205
rect 24624 27149 24652 27205
rect 25088 27149 25116 27205
rect 25276 27149 25304 27205
rect 25740 27149 25768 27205
rect 25872 27149 25900 27205
rect 26336 27149 26364 27205
rect 26524 27149 26552 27205
rect 26988 27149 27016 27205
rect 27120 27149 27148 27205
rect 27584 27149 27612 27205
rect 27772 27149 27800 27205
rect 28236 27149 28264 27205
rect 28368 27149 28396 27205
rect 28832 27149 28860 27205
rect 29020 27149 29048 27205
rect 29484 27149 29512 27205
rect 29616 27149 29644 27205
rect 30080 27149 30108 27205
rect 30268 27149 30296 27205
rect 30732 27149 30760 27205
rect 30864 27149 30892 27205
rect 31328 27149 31356 27205
rect 31516 27149 31544 27205
rect 31980 27149 32008 27205
rect 32112 27149 32140 27205
rect 32576 27149 32604 27205
rect 32764 27149 32792 27205
rect 33228 27149 33256 27205
rect 33360 27149 33388 27205
rect 33824 27149 33852 27205
rect 34012 27149 34040 27205
rect 34476 27149 34504 27205
rect 34608 27149 34636 27205
rect 35072 27149 35100 27205
rect 35260 27149 35288 27205
rect 35724 27149 35752 27205
rect 35856 27149 35884 27205
rect 36320 27149 36348 27205
rect 36508 27149 36536 27205
rect 36972 27149 37000 27205
rect 37104 27149 37132 27205
rect 37568 27149 37596 27205
rect 37756 27149 37784 27205
rect 38220 27149 38248 27205
rect 38352 27149 38380 27205
rect 38816 27149 38844 27205
rect 39004 27149 39032 27205
rect 39468 27149 39496 27205
rect 39600 27149 39628 27205
rect 40064 27149 40092 27205
rect 40252 27149 40280 27205
rect 40716 27149 40744 27205
rect 40848 27149 40876 27205
rect 41312 27149 41340 27205
rect 41500 27149 41528 27205
rect 41964 27149 41992 27205
rect 42096 27149 42124 27205
rect 42560 27149 42588 27205
rect 42748 27149 42776 27205
rect 43212 27149 43240 27205
rect 43344 27149 43372 27205
rect 43808 27149 43836 27205
rect 43996 27149 44024 27205
rect 44460 27149 44488 27205
rect 44592 27149 44620 27205
rect 45056 27149 45084 27205
rect 45244 27149 45272 27205
rect 45708 27149 45736 27205
rect 45840 27149 45868 27205
rect 46304 27149 46332 27205
rect 46492 27149 46520 27205
rect 46956 27149 46984 27205
rect 47088 27149 47116 27205
rect 47552 27149 47580 27205
rect 47740 27149 47768 27205
rect 48204 27149 48232 27205
rect 48336 27149 48364 27205
rect 48800 27149 48828 27205
rect 48988 27149 49016 27205
rect 49452 27149 49480 27205
rect 49584 27149 49612 27205
rect 50048 27149 50076 27205
rect 50236 27149 50264 27205
rect 50700 27149 50728 27205
rect 50832 27149 50860 27205
rect 51296 27149 51324 27205
rect 51484 27149 51512 27205
rect 51948 27149 51976 27205
rect 52080 27149 52108 27205
rect 52544 27149 52572 27205
rect 52732 27149 52760 27205
rect 53196 27149 53224 27205
rect 53328 27149 53356 27205
rect 53792 27149 53820 27205
rect 53980 27149 54008 27205
rect 54444 27149 54472 27205
rect 54576 27149 54604 27205
rect 55040 27149 55068 27205
rect 55228 27149 55256 27205
rect 55692 27149 55720 27205
rect 55824 27149 55852 27205
rect 56288 27149 56316 27205
rect 56476 27149 56504 27205
rect 56940 27149 56968 27205
rect 57072 27149 57100 27205
rect 57536 27149 57564 27205
rect 70966 26929 71024 26975
rect 71156 26929 71214 26975
rect 71417 26929 71475 26975
rect 71767 26929 71825 26975
rect 72028 26929 72086 26975
rect 70978 26809 71012 26929
rect 70962 26757 71028 26809
rect 70978 26415 71012 26757
rect 71040 26606 71106 26658
rect 71168 26655 71202 26929
rect 71156 26609 71214 26655
rect 71168 26415 71202 26609
rect 71429 26415 71463 26929
rect 71687 26895 71741 26904
rect 71685 26849 71743 26895
rect 71687 26840 71741 26849
rect 71697 26584 71731 26840
rect 71779 26809 71813 26929
rect 71951 26809 72009 26815
rect 71779 26775 72009 26809
rect 71687 26575 71741 26584
rect 71685 26529 71743 26575
rect 71687 26520 71741 26529
rect 71779 26415 71813 26775
rect 71951 26769 72009 26775
rect 71907 26686 71973 26738
rect 72040 26655 72074 26929
rect 72028 26609 72086 26655
rect 72040 26415 72074 26609
rect 70966 26369 71024 26415
rect 71156 26369 71214 26415
rect 71417 26369 71475 26415
rect 71767 26369 71825 26415
rect 72028 26369 72086 26415
rect 17788 25469 17816 25897
rect 18252 25345 18280 25897
rect 18384 25841 18412 25897
rect 18848 25841 18876 25897
rect 19036 25469 19064 25897
rect 19500 25345 19528 25897
rect 19632 25841 19660 25897
rect 20096 25841 20124 25897
rect 20284 25469 20312 25897
rect 20748 25345 20776 25897
rect 20880 25841 20908 25897
rect 21344 25841 21372 25897
rect 21532 25469 21560 25897
rect 21996 25345 22024 25897
rect 22128 25841 22156 25897
rect 22592 25841 22620 25897
rect 22780 25469 22808 25897
rect 23244 25345 23272 25897
rect 23376 25841 23404 25897
rect 23840 25841 23868 25897
rect 24028 25469 24056 25897
rect 24492 25345 24520 25897
rect 24624 25841 24652 25897
rect 25088 25841 25116 25897
rect 25276 25469 25304 25897
rect 25740 25345 25768 25897
rect 25872 25841 25900 25897
rect 26336 25841 26364 25897
rect 26524 25469 26552 25897
rect 26988 25345 27016 25897
rect 27120 25841 27148 25897
rect 27584 25841 27612 25897
rect 27772 25469 27800 25897
rect 28236 25345 28264 25897
rect 28368 25841 28396 25897
rect 28832 25841 28860 25897
rect 29020 25469 29048 25897
rect 29484 25345 29512 25897
rect 29616 25841 29644 25897
rect 30080 25841 30108 25897
rect 30268 25469 30296 25897
rect 30732 25345 30760 25897
rect 30864 25841 30892 25897
rect 31328 25841 31356 25897
rect 31516 25469 31544 25897
rect 31980 25345 32008 25897
rect 32112 25841 32140 25897
rect 32576 25841 32604 25897
rect 32764 25469 32792 25897
rect 33228 25345 33256 25897
rect 33360 25841 33388 25897
rect 33824 25841 33852 25897
rect 34012 25469 34040 25897
rect 34476 25345 34504 25897
rect 34608 25841 34636 25897
rect 35072 25841 35100 25897
rect 35260 25469 35288 25897
rect 35724 25345 35752 25897
rect 35856 25841 35884 25897
rect 36320 25841 36348 25897
rect 36508 25469 36536 25897
rect 36972 25345 37000 25897
rect 37104 25841 37132 25897
rect 37568 25841 37596 25897
rect 37756 25469 37784 25897
rect 38220 25345 38248 25897
rect 38352 25841 38380 25897
rect 38816 25841 38844 25897
rect 39004 25469 39032 25897
rect 39468 25345 39496 25897
rect 39600 25841 39628 25897
rect 40064 25841 40092 25897
rect 40252 25469 40280 25897
rect 40716 25345 40744 25897
rect 40848 25841 40876 25897
rect 41312 25841 41340 25897
rect 41500 25469 41528 25897
rect 41964 25345 41992 25897
rect 42096 25841 42124 25897
rect 42560 25841 42588 25897
rect 42748 25469 42776 25897
rect 43212 25345 43240 25897
rect 43344 25841 43372 25897
rect 43808 25841 43836 25897
rect 43996 25469 44024 25897
rect 44460 25345 44488 25897
rect 44592 25841 44620 25897
rect 45056 25841 45084 25897
rect 45244 25469 45272 25897
rect 45708 25345 45736 25897
rect 45840 25841 45868 25897
rect 46304 25841 46332 25897
rect 46492 25469 46520 25897
rect 46956 25345 46984 25897
rect 47088 25841 47116 25897
rect 47552 25841 47580 25897
rect 47740 25469 47768 25897
rect 48204 25345 48232 25897
rect 48336 25841 48364 25897
rect 48800 25841 48828 25897
rect 48988 25469 49016 25897
rect 49452 25345 49480 25897
rect 49584 25841 49612 25897
rect 50048 25841 50076 25897
rect 50236 25469 50264 25897
rect 50700 25345 50728 25897
rect 50832 25841 50860 25897
rect 51296 25841 51324 25897
rect 51484 25469 51512 25897
rect 51948 25345 51976 25897
rect 52080 25841 52108 25897
rect 52544 25841 52572 25897
rect 52732 25469 52760 25897
rect 53196 25345 53224 25897
rect 53328 25841 53356 25897
rect 53792 25841 53820 25897
rect 53980 25469 54008 25897
rect 54444 25345 54472 25897
rect 54576 25841 54604 25897
rect 55040 25841 55068 25897
rect 55228 25469 55256 25897
rect 55692 25345 55720 25897
rect 55824 25841 55852 25897
rect 56288 25841 56316 25897
rect 56476 25469 56504 25897
rect 56940 25345 56968 25897
rect 57072 25841 57100 25897
rect 57536 25841 57564 25897
rect 70966 25881 71024 25927
rect 71156 25881 71214 25927
rect 71417 25881 71475 25927
rect 71767 25881 71825 25927
rect 72028 25881 72086 25927
rect 70978 25539 71012 25881
rect 71040 25638 71106 25690
rect 71168 25687 71202 25881
rect 71156 25641 71214 25687
rect 70962 25487 71028 25539
rect 70978 25367 71012 25487
rect 71168 25367 71202 25641
rect 71429 25367 71463 25881
rect 71687 25767 71741 25776
rect 71685 25721 71743 25767
rect 71687 25712 71741 25721
rect 71697 25456 71731 25712
rect 71779 25521 71813 25881
rect 72040 25687 72074 25881
rect 72028 25641 72086 25687
rect 71907 25558 71973 25610
rect 71951 25521 72009 25527
rect 71779 25487 72009 25521
rect 71687 25447 71741 25456
rect 71685 25401 71743 25447
rect 71687 25392 71741 25401
rect 71779 25367 71813 25487
rect 71951 25481 72009 25487
rect 72040 25367 72074 25641
rect 70966 25321 71024 25367
rect 71156 25321 71214 25367
rect 71417 25321 71475 25367
rect 71767 25321 71825 25367
rect 72028 25321 72086 25367
rect 17802 24877 17860 24937
rect 17904 23843 17938 24969
rect 17980 23855 18008 24969
rect 19050 24877 19108 24937
rect 18136 24718 18182 24792
rect 18046 23947 18108 24015
rect 17892 23797 17950 23843
rect 17980 23797 18048 23855
rect 19152 23843 19186 24969
rect 19228 23855 19256 24969
rect 20298 24877 20356 24937
rect 19384 24718 19430 24792
rect 19294 23947 19356 24015
rect 19140 23797 19198 23843
rect 19228 23797 19296 23855
rect 20400 23843 20434 24969
rect 20476 23855 20504 24969
rect 21546 24877 21604 24937
rect 20632 24718 20678 24792
rect 20542 23947 20604 24015
rect 20388 23797 20446 23843
rect 20476 23797 20544 23855
rect 21648 23843 21682 24969
rect 21724 23855 21752 24969
rect 22794 24877 22852 24937
rect 21880 24718 21926 24792
rect 21790 23947 21852 24015
rect 21636 23797 21694 23843
rect 21724 23797 21792 23855
rect 22896 23843 22930 24969
rect 22972 23855 23000 24969
rect 24042 24877 24100 24937
rect 23128 24718 23174 24792
rect 23038 23947 23100 24015
rect 22884 23797 22942 23843
rect 22972 23797 23040 23855
rect 24144 23843 24178 24969
rect 24220 23855 24248 24969
rect 25290 24877 25348 24937
rect 24376 24718 24422 24792
rect 24286 23947 24348 24015
rect 24132 23797 24190 23843
rect 24220 23797 24288 23855
rect 25392 23843 25426 24969
rect 25468 23855 25496 24969
rect 26538 24877 26596 24937
rect 25624 24718 25670 24792
rect 25534 23947 25596 24015
rect 25380 23797 25438 23843
rect 25468 23797 25536 23855
rect 26640 23843 26674 24969
rect 26716 23855 26744 24969
rect 27786 24877 27844 24937
rect 26872 24718 26918 24792
rect 26782 23947 26844 24015
rect 26628 23797 26686 23843
rect 26716 23797 26784 23855
rect 27888 23843 27922 24969
rect 27964 23855 27992 24969
rect 29034 24877 29092 24937
rect 28120 24718 28166 24792
rect 28030 23947 28092 24015
rect 27876 23797 27934 23843
rect 27964 23797 28032 23855
rect 29136 23843 29170 24969
rect 29212 23855 29240 24969
rect 30282 24877 30340 24937
rect 29368 24718 29414 24792
rect 29278 23947 29340 24015
rect 29124 23797 29182 23843
rect 29212 23797 29280 23855
rect 30384 23843 30418 24969
rect 30460 23855 30488 24969
rect 31530 24877 31588 24937
rect 30616 24718 30662 24792
rect 30526 23947 30588 24015
rect 30372 23797 30430 23843
rect 30460 23797 30528 23855
rect 31632 23843 31666 24969
rect 31708 23855 31736 24969
rect 32778 24877 32836 24937
rect 31864 24718 31910 24792
rect 31774 23947 31836 24015
rect 31620 23797 31678 23843
rect 31708 23797 31776 23855
rect 32880 23843 32914 24969
rect 32956 23855 32984 24969
rect 34026 24877 34084 24937
rect 33112 24718 33158 24792
rect 33022 23947 33084 24015
rect 32868 23797 32926 23843
rect 32956 23797 33024 23855
rect 34128 23843 34162 24969
rect 34204 23855 34232 24969
rect 35274 24877 35332 24937
rect 34360 24718 34406 24792
rect 34270 23947 34332 24015
rect 34116 23797 34174 23843
rect 34204 23797 34272 23855
rect 35376 23843 35410 24969
rect 35452 23855 35480 24969
rect 36522 24877 36580 24937
rect 35608 24718 35654 24792
rect 35518 23947 35580 24015
rect 35364 23797 35422 23843
rect 35452 23797 35520 23855
rect 36624 23843 36658 24969
rect 36700 23855 36728 24969
rect 37770 24877 37828 24937
rect 36856 24718 36902 24792
rect 36766 23947 36828 24015
rect 36612 23797 36670 23843
rect 36700 23797 36768 23855
rect 37872 23843 37906 24969
rect 37948 23855 37976 24969
rect 39018 24877 39076 24937
rect 38104 24718 38150 24792
rect 38014 23947 38076 24015
rect 37860 23797 37918 23843
rect 37948 23797 38016 23855
rect 39120 23843 39154 24969
rect 39196 23855 39224 24969
rect 40266 24877 40324 24937
rect 39352 24718 39398 24792
rect 39262 23947 39324 24015
rect 39108 23797 39166 23843
rect 39196 23797 39264 23855
rect 40368 23843 40402 24969
rect 40444 23855 40472 24969
rect 41514 24877 41572 24937
rect 40600 24718 40646 24792
rect 40510 23947 40572 24015
rect 40356 23797 40414 23843
rect 40444 23797 40512 23855
rect 41616 23843 41650 24969
rect 41692 23855 41720 24969
rect 42762 24877 42820 24937
rect 41848 24718 41894 24792
rect 41758 23947 41820 24015
rect 41604 23797 41662 23843
rect 41692 23797 41760 23855
rect 42864 23843 42898 24969
rect 42940 23855 42968 24969
rect 44010 24877 44068 24937
rect 43096 24718 43142 24792
rect 43006 23947 43068 24015
rect 42852 23797 42910 23843
rect 42940 23797 43008 23855
rect 44112 23843 44146 24969
rect 44188 23855 44216 24969
rect 45258 24877 45316 24937
rect 44344 24718 44390 24792
rect 44254 23947 44316 24015
rect 44100 23797 44158 23843
rect 44188 23797 44256 23855
rect 45360 23843 45394 24969
rect 45436 23855 45464 24969
rect 46506 24877 46564 24937
rect 45592 24718 45638 24792
rect 45502 23947 45564 24015
rect 45348 23797 45406 23843
rect 45436 23797 45504 23855
rect 46608 23843 46642 24969
rect 46684 23855 46712 24969
rect 47754 24877 47812 24937
rect 46840 24718 46886 24792
rect 46750 23947 46812 24015
rect 46596 23797 46654 23843
rect 46684 23797 46752 23855
rect 47856 23843 47890 24969
rect 47932 23855 47960 24969
rect 49002 24877 49060 24937
rect 48088 24718 48134 24792
rect 47998 23947 48060 24015
rect 47844 23797 47902 23843
rect 47932 23797 48000 23855
rect 49104 23843 49138 24969
rect 49180 23855 49208 24969
rect 50250 24877 50308 24937
rect 49336 24718 49382 24792
rect 49246 23947 49308 24015
rect 49092 23797 49150 23843
rect 49180 23797 49248 23855
rect 50352 23843 50386 24969
rect 50428 23855 50456 24969
rect 51498 24877 51556 24937
rect 50584 24718 50630 24792
rect 50494 23947 50556 24015
rect 50340 23797 50398 23843
rect 50428 23797 50496 23855
rect 51600 23843 51634 24969
rect 51676 23855 51704 24969
rect 52746 24877 52804 24937
rect 51832 24718 51878 24792
rect 51742 23947 51804 24015
rect 51588 23797 51646 23843
rect 51676 23797 51744 23855
rect 52848 23843 52882 24969
rect 52924 23855 52952 24969
rect 53994 24877 54052 24937
rect 53080 24718 53126 24792
rect 52990 23947 53052 24015
rect 52836 23797 52894 23843
rect 52924 23797 52992 23855
rect 54096 23843 54130 24969
rect 54172 23855 54200 24969
rect 55242 24877 55300 24937
rect 54328 24718 54374 24792
rect 54238 23947 54300 24015
rect 54084 23797 54142 23843
rect 54172 23797 54240 23855
rect 55344 23843 55378 24969
rect 55420 23855 55448 24969
rect 56490 24877 56548 24937
rect 55576 24718 55622 24792
rect 55486 23947 55548 24015
rect 55332 23797 55390 23843
rect 55420 23797 55488 23855
rect 56592 23843 56626 24969
rect 56668 23855 56696 24969
rect 56824 24718 56870 24792
rect 70966 24101 71024 24147
rect 71156 24101 71214 24147
rect 71417 24101 71475 24147
rect 71767 24101 71825 24147
rect 72028 24101 72086 24147
rect 56734 23947 56796 24015
rect 70978 23981 71012 24101
rect 70962 23929 71028 23981
rect 56580 23797 56638 23843
rect 56668 23797 56736 23855
rect 17812 22713 17858 22967
rect 17904 22713 17938 23797
rect 17980 22713 18008 23797
rect 18066 23105 18112 23181
rect 18066 22784 18112 22858
rect 19060 22713 19106 22967
rect 19152 22713 19186 23797
rect 19228 22713 19256 23797
rect 19314 23105 19360 23181
rect 19314 22784 19360 22858
rect 20308 22713 20354 22967
rect 20400 22713 20434 23797
rect 20476 22713 20504 23797
rect 20562 23105 20608 23181
rect 20562 22784 20608 22858
rect 21556 22713 21602 22967
rect 21648 22713 21682 23797
rect 21724 22713 21752 23797
rect 21810 23105 21856 23181
rect 21810 22784 21856 22858
rect 22804 22713 22850 22967
rect 22896 22713 22930 23797
rect 22972 22713 23000 23797
rect 23058 23105 23104 23181
rect 23058 22784 23104 22858
rect 24052 22713 24098 22967
rect 24144 22713 24178 23797
rect 24220 22713 24248 23797
rect 24306 23105 24352 23181
rect 24306 22784 24352 22858
rect 25300 22713 25346 22967
rect 25392 22713 25426 23797
rect 25468 22713 25496 23797
rect 25554 23105 25600 23181
rect 25554 22784 25600 22858
rect 26548 22713 26594 22967
rect 26640 22713 26674 23797
rect 26716 22713 26744 23797
rect 26802 23105 26848 23181
rect 26802 22784 26848 22858
rect 27796 22713 27842 22967
rect 27888 22713 27922 23797
rect 27964 22713 27992 23797
rect 28050 23105 28096 23181
rect 28050 22784 28096 22858
rect 29044 22713 29090 22967
rect 29136 22713 29170 23797
rect 29212 22713 29240 23797
rect 29298 23105 29344 23181
rect 29298 22784 29344 22858
rect 30292 22713 30338 22967
rect 30384 22713 30418 23797
rect 30460 22713 30488 23797
rect 30546 23105 30592 23181
rect 30546 22784 30592 22858
rect 31540 22713 31586 22967
rect 31632 22713 31666 23797
rect 31708 22713 31736 23797
rect 31794 23105 31840 23181
rect 31794 22784 31840 22858
rect 32788 22713 32834 22967
rect 32880 22713 32914 23797
rect 32956 22713 32984 23797
rect 33042 23105 33088 23181
rect 33042 22784 33088 22858
rect 34036 22713 34082 22967
rect 34128 22713 34162 23797
rect 34204 22713 34232 23797
rect 34290 23105 34336 23181
rect 34290 22784 34336 22858
rect 35284 22713 35330 22967
rect 35376 22713 35410 23797
rect 35452 22713 35480 23797
rect 35538 23105 35584 23181
rect 35538 22784 35584 22858
rect 36532 22713 36578 22967
rect 36624 22713 36658 23797
rect 36700 22713 36728 23797
rect 36786 23105 36832 23181
rect 36786 22784 36832 22858
rect 37780 22713 37826 22967
rect 37872 22713 37906 23797
rect 37948 22713 37976 23797
rect 38034 23105 38080 23181
rect 38034 22784 38080 22858
rect 39028 22713 39074 22967
rect 39120 22713 39154 23797
rect 39196 22713 39224 23797
rect 39282 23105 39328 23181
rect 39282 22784 39328 22858
rect 40276 22713 40322 22967
rect 40368 22713 40402 23797
rect 40444 22713 40472 23797
rect 40530 23105 40576 23181
rect 40530 22784 40576 22858
rect 41524 22713 41570 22967
rect 41616 22713 41650 23797
rect 41692 22713 41720 23797
rect 41778 23105 41824 23181
rect 41778 22784 41824 22858
rect 42772 22713 42818 22967
rect 42864 22713 42898 23797
rect 42940 22713 42968 23797
rect 43026 23105 43072 23181
rect 43026 22784 43072 22858
rect 44020 22713 44066 22967
rect 44112 22713 44146 23797
rect 44188 22713 44216 23797
rect 44274 23105 44320 23181
rect 44274 22784 44320 22858
rect 45268 22713 45314 22967
rect 45360 22713 45394 23797
rect 45436 22713 45464 23797
rect 45522 23105 45568 23181
rect 45522 22784 45568 22858
rect 46516 22713 46562 22967
rect 46608 22713 46642 23797
rect 46684 22713 46712 23797
rect 46770 23105 46816 23181
rect 46770 22784 46816 22858
rect 47764 22713 47810 22967
rect 47856 22713 47890 23797
rect 47932 22713 47960 23797
rect 48018 23105 48064 23181
rect 48018 22784 48064 22858
rect 49012 22713 49058 22967
rect 49104 22713 49138 23797
rect 49180 22713 49208 23797
rect 49266 23105 49312 23181
rect 49266 22784 49312 22858
rect 50260 22713 50306 22967
rect 50352 22713 50386 23797
rect 50428 22713 50456 23797
rect 50514 23105 50560 23181
rect 50514 22784 50560 22858
rect 51508 22713 51554 22967
rect 51600 22713 51634 23797
rect 51676 22713 51704 23797
rect 51762 23105 51808 23181
rect 51762 22784 51808 22858
rect 52756 22713 52802 22967
rect 52848 22713 52882 23797
rect 52924 22713 52952 23797
rect 53010 23105 53056 23181
rect 53010 22784 53056 22858
rect 54004 22713 54050 22967
rect 54096 22713 54130 23797
rect 54172 22713 54200 23797
rect 54258 23105 54304 23181
rect 54258 22784 54304 22858
rect 55252 22713 55298 22967
rect 55344 22713 55378 23797
rect 55420 22713 55448 23797
rect 55506 23105 55552 23181
rect 55506 22784 55552 22858
rect 56500 22713 56546 22967
rect 56592 22713 56626 23797
rect 56668 22713 56696 23797
rect 70978 23587 71012 23929
rect 71040 23778 71106 23830
rect 71168 23827 71202 24101
rect 71156 23781 71214 23827
rect 71168 23587 71202 23781
rect 71429 23587 71463 24101
rect 71687 24067 71741 24076
rect 71685 24021 71743 24067
rect 71687 24012 71741 24021
rect 71697 23756 71731 24012
rect 71779 23981 71813 24101
rect 71951 23981 72009 23987
rect 71779 23947 72009 23981
rect 71687 23747 71741 23756
rect 71685 23701 71743 23747
rect 71687 23692 71741 23701
rect 71779 23587 71813 23947
rect 71951 23941 72009 23947
rect 71907 23858 71973 23910
rect 72040 23827 72074 24101
rect 72028 23781 72086 23827
rect 72040 23587 72074 23781
rect 70966 23541 71024 23587
rect 71156 23541 71214 23587
rect 71417 23541 71475 23587
rect 71767 23541 71825 23587
rect 72028 23541 72086 23587
rect 56754 23105 56800 23181
rect 70966 23053 71024 23099
rect 71156 23053 71214 23099
rect 71417 23053 71475 23099
rect 71767 23053 71825 23099
rect 72028 23053 72086 23099
rect 56754 22784 56800 22858
rect 70978 22711 71012 23053
rect 71040 22810 71106 22862
rect 71168 22859 71202 23053
rect 71156 22813 71214 22859
rect 70962 22659 71028 22711
rect 70978 22539 71012 22659
rect 71168 22539 71202 22813
rect 71429 22539 71463 23053
rect 71687 22939 71741 22948
rect 71685 22893 71743 22939
rect 71687 22884 71741 22893
rect 71697 22628 71731 22884
rect 71779 22693 71813 23053
rect 72040 22859 72074 23053
rect 72028 22813 72086 22859
rect 71907 22730 71973 22782
rect 71951 22693 72009 22699
rect 71779 22659 72009 22693
rect 71687 22619 71741 22628
rect 71685 22573 71743 22619
rect 71687 22564 71741 22573
rect 71779 22539 71813 22659
rect 71951 22653 72009 22659
rect 72040 22539 72074 22813
rect 70966 22493 71024 22539
rect 71156 22493 71214 22539
rect 71417 22493 71475 22539
rect 71767 22493 71825 22539
rect 72028 22493 72086 22539
rect 17834 22409 17864 22461
rect 18036 22409 18066 22461
rect 19082 22409 19112 22461
rect 19284 22409 19314 22461
rect 20330 22409 20360 22461
rect 20532 22409 20562 22461
rect 21578 22409 21608 22461
rect 21780 22409 21810 22461
rect 22826 22409 22856 22461
rect 23028 22409 23058 22461
rect 24074 22409 24104 22461
rect 24276 22409 24306 22461
rect 25322 22409 25352 22461
rect 25524 22409 25554 22461
rect 26570 22409 26600 22461
rect 26772 22409 26802 22461
rect 27818 22409 27848 22461
rect 28020 22409 28050 22461
rect 29066 22409 29096 22461
rect 29268 22409 29298 22461
rect 30314 22409 30344 22461
rect 30516 22409 30546 22461
rect 31562 22409 31592 22461
rect 31764 22409 31794 22461
rect 32810 22409 32840 22461
rect 33012 22409 33042 22461
rect 34058 22409 34088 22461
rect 34260 22409 34290 22461
rect 35306 22409 35336 22461
rect 35508 22409 35538 22461
rect 36554 22409 36584 22461
rect 36756 22409 36786 22461
rect 37802 22409 37832 22461
rect 38004 22409 38034 22461
rect 39050 22409 39080 22461
rect 39252 22409 39282 22461
rect 40298 22409 40328 22461
rect 40500 22409 40530 22461
rect 41546 22409 41576 22461
rect 41748 22409 41778 22461
rect 42794 22409 42824 22461
rect 42996 22409 43026 22461
rect 44042 22409 44072 22461
rect 44244 22409 44274 22461
rect 45290 22409 45320 22461
rect 45492 22409 45522 22461
rect 46538 22409 46568 22461
rect 46740 22409 46770 22461
rect 47786 22409 47816 22461
rect 47988 22409 48018 22461
rect 49034 22409 49064 22461
rect 49236 22409 49266 22461
rect 50282 22409 50312 22461
rect 50484 22409 50514 22461
rect 51530 22409 51560 22461
rect 51732 22409 51762 22461
rect 52778 22409 52808 22461
rect 52980 22409 53010 22461
rect 54026 22409 54056 22461
rect 54228 22409 54258 22461
rect 55274 22409 55304 22461
rect 55476 22409 55506 22461
rect 56522 22409 56552 22461
rect 56724 22409 56754 22461
rect 17833 22351 17890 22409
rect 18010 22351 18067 22409
rect 19081 22351 19138 22409
rect 19258 22351 19315 22409
rect 20329 22351 20386 22409
rect 20506 22351 20563 22409
rect 21577 22351 21634 22409
rect 21754 22351 21811 22409
rect 22825 22351 22882 22409
rect 23002 22351 23059 22409
rect 24073 22351 24130 22409
rect 24250 22351 24307 22409
rect 25321 22351 25378 22409
rect 25498 22351 25555 22409
rect 26569 22351 26626 22409
rect 26746 22351 26803 22409
rect 27817 22351 27874 22409
rect 27994 22351 28051 22409
rect 29065 22351 29122 22409
rect 29242 22351 29299 22409
rect 30313 22351 30370 22409
rect 30490 22351 30547 22409
rect 31561 22351 31618 22409
rect 31738 22351 31795 22409
rect 32809 22351 32866 22409
rect 32986 22351 33043 22409
rect 34057 22351 34114 22409
rect 34234 22351 34291 22409
rect 35305 22351 35362 22409
rect 35482 22351 35539 22409
rect 36553 22351 36610 22409
rect 36730 22351 36787 22409
rect 37801 22351 37858 22409
rect 37978 22351 38035 22409
rect 39049 22351 39106 22409
rect 39226 22351 39283 22409
rect 40297 22351 40354 22409
rect 40474 22351 40531 22409
rect 41545 22351 41602 22409
rect 41722 22351 41779 22409
rect 42793 22351 42850 22409
rect 42970 22351 43027 22409
rect 44041 22351 44098 22409
rect 44218 22351 44275 22409
rect 45289 22351 45346 22409
rect 45466 22351 45523 22409
rect 46537 22351 46594 22409
rect 46714 22351 46771 22409
rect 47785 22351 47842 22409
rect 47962 22351 48019 22409
rect 49033 22351 49090 22409
rect 49210 22351 49267 22409
rect 50281 22351 50338 22409
rect 50458 22351 50515 22409
rect 51529 22351 51586 22409
rect 51706 22351 51763 22409
rect 52777 22351 52834 22409
rect 52954 22351 53011 22409
rect 54025 22351 54082 22409
rect 54202 22351 54259 22409
rect 55273 22351 55330 22409
rect 55450 22351 55507 22409
rect 56521 22351 56578 22409
rect 56698 22351 56755 22409
rect 17921 22045 18007 22051
rect 19169 22045 19255 22051
rect 20417 22045 20503 22051
rect 21665 22045 21751 22051
rect 22913 22045 22999 22051
rect 24161 22045 24247 22051
rect 25409 22045 25495 22051
rect 26657 22045 26743 22051
rect 27905 22045 27991 22051
rect 29153 22045 29239 22051
rect 30401 22045 30487 22051
rect 31649 22045 31735 22051
rect 32897 22045 32983 22051
rect 34145 22045 34231 22051
rect 35393 22045 35479 22051
rect 36641 22045 36727 22051
rect 37889 22045 37975 22051
rect 39137 22045 39223 22051
rect 40385 22045 40471 22051
rect 41633 22045 41719 22051
rect 42881 22045 42967 22051
rect 44129 22045 44215 22051
rect 45377 22045 45463 22051
rect 46625 22045 46711 22051
rect 47873 22045 47959 22051
rect 49121 22045 49207 22051
rect 50369 22045 50455 22051
rect 51617 22045 51703 22051
rect 52865 22045 52951 22051
rect 54113 22045 54199 22051
rect 55361 22045 55447 22051
rect 56609 22045 56695 22051
rect 17921 22011 18029 22045
rect 19169 22011 19277 22045
rect 20417 22011 20525 22045
rect 21665 22011 21773 22045
rect 22913 22011 23021 22045
rect 24161 22011 24269 22045
rect 25409 22011 25517 22045
rect 26657 22011 26765 22045
rect 27905 22011 28013 22045
rect 29153 22011 29261 22045
rect 30401 22011 30509 22045
rect 31649 22011 31757 22045
rect 32897 22011 33005 22045
rect 34145 22011 34253 22045
rect 35393 22011 35501 22045
rect 36641 22011 36749 22045
rect 37889 22011 37997 22045
rect 39137 22011 39245 22045
rect 40385 22011 40493 22045
rect 41633 22011 41741 22045
rect 42881 22011 42989 22045
rect 44129 22011 44237 22045
rect 45377 22011 45485 22045
rect 46625 22011 46733 22045
rect 47873 22011 47981 22045
rect 49121 22011 49229 22045
rect 50369 22011 50477 22045
rect 51617 22011 51725 22045
rect 52865 22011 52973 22045
rect 54113 22011 54221 22045
rect 55361 22011 55469 22045
rect 56609 22011 56717 22045
rect 17921 22005 18007 22011
rect 19169 22005 19255 22011
rect 20417 22005 20503 22011
rect 21665 22005 21751 22011
rect 22913 22005 22999 22011
rect 24161 22005 24247 22011
rect 25409 22005 25495 22011
rect 26657 22005 26743 22011
rect 27905 22005 27991 22011
rect 29153 22005 29239 22011
rect 30401 22005 30487 22011
rect 31649 22005 31735 22011
rect 32897 22005 32983 22011
rect 34145 22005 34231 22011
rect 35393 22005 35479 22011
rect 36641 22005 36727 22011
rect 37889 22005 37975 22011
rect 39137 22005 39223 22011
rect 40385 22005 40471 22011
rect 41633 22005 41719 22011
rect 42881 22005 42967 22011
rect 44129 22005 44215 22011
rect 45377 22005 45463 22011
rect 46625 22005 46711 22011
rect 47873 22005 47959 22011
rect 49121 22005 49207 22011
rect 50369 22005 50455 22011
rect 51617 22005 51703 22011
rect 52865 22005 52951 22011
rect 54113 22005 54199 22011
rect 55361 22005 55447 22011
rect 56609 22005 56695 22011
rect 17921 21568 18007 21614
rect 19169 21568 19255 21614
rect 20417 21568 20503 21614
rect 21665 21568 21751 21614
rect 22913 21568 22999 21614
rect 24161 21568 24247 21614
rect 25409 21568 25495 21614
rect 26657 21568 26743 21614
rect 27905 21568 27991 21614
rect 29153 21568 29239 21614
rect 30401 21568 30487 21614
rect 31649 21568 31735 21614
rect 32897 21568 32983 21614
rect 34145 21568 34231 21614
rect 35393 21568 35479 21614
rect 36641 21568 36727 21614
rect 37889 21568 37975 21614
rect 39137 21568 39223 21614
rect 40385 21568 40471 21614
rect 41633 21568 41719 21614
rect 42881 21568 42967 21614
rect 44129 21568 44215 21614
rect 45377 21568 45463 21614
rect 46625 21568 46711 21614
rect 47873 21568 47959 21614
rect 49121 21568 49207 21614
rect 50369 21568 50455 21614
rect 51617 21568 51703 21614
rect 52865 21568 52951 21614
rect 54113 21568 54199 21614
rect 55361 21568 55447 21614
rect 56609 21568 56695 21614
rect 18042 21239 18128 21280
rect 19290 21239 19376 21280
rect 20538 21239 20624 21280
rect 21786 21239 21872 21280
rect 23034 21239 23120 21280
rect 24282 21239 24368 21280
rect 25530 21239 25616 21280
rect 26778 21239 26864 21280
rect 28026 21239 28112 21280
rect 29274 21239 29360 21280
rect 30522 21239 30608 21280
rect 31770 21239 31856 21280
rect 33018 21239 33104 21280
rect 34266 21239 34352 21280
rect 35514 21239 35600 21280
rect 36762 21239 36848 21280
rect 38010 21239 38096 21280
rect 39258 21239 39344 21280
rect 40506 21239 40592 21280
rect 41754 21239 41840 21280
rect 43002 21239 43088 21280
rect 44250 21239 44336 21280
rect 45498 21239 45584 21280
rect 46746 21239 46832 21280
rect 47994 21239 48080 21280
rect 49242 21239 49328 21280
rect 50490 21239 50576 21280
rect 51738 21239 51824 21280
rect 52986 21239 53072 21280
rect 54234 21239 54320 21280
rect 55482 21239 55568 21280
rect 56730 21239 56816 21280
rect 70966 21273 71024 21319
rect 71156 21273 71214 21319
rect 71417 21273 71475 21319
rect 71767 21273 71825 21319
rect 72028 21273 72086 21319
rect 18055 21234 18128 21239
rect 19303 21234 19376 21239
rect 20551 21234 20624 21239
rect 21799 21234 21872 21239
rect 23047 21234 23120 21239
rect 24295 21234 24368 21239
rect 25543 21234 25616 21239
rect 26791 21234 26864 21239
rect 28039 21234 28112 21239
rect 29287 21234 29360 21239
rect 30535 21234 30608 21239
rect 31783 21234 31856 21239
rect 33031 21234 33104 21239
rect 34279 21234 34352 21239
rect 35527 21234 35600 21239
rect 36775 21234 36848 21239
rect 38023 21234 38096 21239
rect 39271 21234 39344 21239
rect 40519 21234 40592 21239
rect 41767 21234 41840 21239
rect 43015 21234 43088 21239
rect 44263 21234 44336 21239
rect 45511 21234 45584 21239
rect 46759 21234 46832 21239
rect 48007 21234 48080 21239
rect 49255 21234 49328 21239
rect 50503 21234 50576 21239
rect 51751 21234 51824 21239
rect 52999 21234 53072 21239
rect 54247 21234 54320 21239
rect 55495 21234 55568 21239
rect 56743 21234 56816 21239
rect 70978 21153 71012 21273
rect 70962 21101 71028 21153
rect 17927 21034 18013 21080
rect 19175 21034 19261 21080
rect 20423 21034 20509 21080
rect 21671 21034 21757 21080
rect 22919 21034 23005 21080
rect 24167 21034 24253 21080
rect 25415 21034 25501 21080
rect 26663 21034 26749 21080
rect 27911 21034 27997 21080
rect 29159 21034 29245 21080
rect 30407 21034 30493 21080
rect 31655 21034 31741 21080
rect 32903 21034 32989 21080
rect 34151 21034 34237 21080
rect 35399 21034 35485 21080
rect 36647 21034 36733 21080
rect 37895 21034 37981 21080
rect 39143 21034 39229 21080
rect 40391 21034 40477 21080
rect 41639 21034 41725 21080
rect 42887 21034 42973 21080
rect 44135 21034 44221 21080
rect 45383 21034 45469 21080
rect 46631 21034 46717 21080
rect 47879 21034 47965 21080
rect 49127 21034 49213 21080
rect 50375 21034 50461 21080
rect 51623 21034 51709 21080
rect 52871 21034 52957 21080
rect 54119 21034 54205 21080
rect 55367 21034 55453 21080
rect 56615 21034 56701 21080
rect 70978 20759 71012 21101
rect 71040 20950 71106 21002
rect 71168 20999 71202 21273
rect 71156 20953 71214 20999
rect 71168 20759 71202 20953
rect 71429 20759 71463 21273
rect 71687 21239 71741 21248
rect 71685 21193 71743 21239
rect 71687 21184 71741 21193
rect 71697 20928 71731 21184
rect 71779 21153 71813 21273
rect 71951 21153 72009 21159
rect 71779 21119 72009 21153
rect 71687 20919 71741 20928
rect 71685 20873 71743 20919
rect 71687 20864 71741 20873
rect 71779 20759 71813 21119
rect 71951 21113 72009 21119
rect 71907 21030 71973 21082
rect 72040 20999 72074 21273
rect 72028 20953 72086 20999
rect 72040 20759 72074 20953
rect 70966 20713 71024 20759
rect 71156 20713 71214 20759
rect 71417 20713 71475 20759
rect 71767 20713 71825 20759
rect 72028 20713 72086 20759
rect 17941 20618 18027 20664
rect 19189 20618 19275 20664
rect 20437 20618 20523 20664
rect 21685 20618 21771 20664
rect 22933 20618 23019 20664
rect 24181 20618 24267 20664
rect 25429 20618 25515 20664
rect 26677 20618 26763 20664
rect 27925 20618 28011 20664
rect 29173 20618 29259 20664
rect 30421 20618 30507 20664
rect 31669 20618 31755 20664
rect 32917 20618 33003 20664
rect 34165 20618 34251 20664
rect 35413 20618 35499 20664
rect 36661 20618 36747 20664
rect 37909 20618 37995 20664
rect 39157 20618 39243 20664
rect 40405 20618 40491 20664
rect 41653 20618 41739 20664
rect 42901 20618 42987 20664
rect 44149 20618 44235 20664
rect 45397 20618 45483 20664
rect 46645 20618 46731 20664
rect 47893 20618 47979 20664
rect 49141 20618 49227 20664
rect 50389 20618 50475 20664
rect 51637 20618 51723 20664
rect 52885 20618 52971 20664
rect 54133 20618 54219 20664
rect 55381 20618 55467 20664
rect 56629 20618 56715 20664
rect 17807 20578 17865 20606
rect 19055 20578 19113 20606
rect 20303 20578 20361 20606
rect 21551 20578 21609 20606
rect 22799 20578 22857 20606
rect 24047 20578 24105 20606
rect 25295 20578 25353 20606
rect 26543 20578 26601 20606
rect 27791 20578 27849 20606
rect 29039 20578 29097 20606
rect 30287 20578 30345 20606
rect 31535 20578 31593 20606
rect 32783 20578 32841 20606
rect 34031 20578 34089 20606
rect 35279 20578 35337 20606
rect 36527 20578 36585 20606
rect 37775 20578 37833 20606
rect 39023 20578 39081 20606
rect 40271 20578 40329 20606
rect 41519 20578 41577 20606
rect 42767 20578 42825 20606
rect 44015 20578 44073 20606
rect 45263 20578 45321 20606
rect 46511 20578 46569 20606
rect 47759 20578 47817 20606
rect 49007 20578 49065 20606
rect 50255 20578 50313 20606
rect 51503 20578 51561 20606
rect 52751 20578 52809 20606
rect 53999 20578 54057 20606
rect 55247 20578 55305 20606
rect 56495 20578 56553 20606
rect 17807 20544 27167 20578
rect 27791 20544 37151 20578
rect 37775 20544 47135 20578
rect 47759 20544 57119 20578
rect 17963 20454 18023 20510
rect 19211 20454 19271 20510
rect 20459 20454 20519 20510
rect 21707 20454 21767 20510
rect 22955 20454 23015 20510
rect 24203 20454 24263 20510
rect 25451 20454 25511 20510
rect 26699 20454 26759 20510
rect 27947 20454 28007 20510
rect 29195 20454 29255 20510
rect 30443 20454 30503 20510
rect 31691 20454 31751 20510
rect 32939 20454 32999 20510
rect 34187 20454 34247 20510
rect 35435 20454 35495 20510
rect 36683 20454 36743 20510
rect 37931 20454 37991 20510
rect 39179 20454 39239 20510
rect 40427 20454 40487 20510
rect 41675 20454 41735 20510
rect 42923 20454 42983 20510
rect 44171 20454 44231 20510
rect 45419 20454 45479 20510
rect 46667 20454 46727 20510
rect 47915 20454 47975 20510
rect 49163 20454 49223 20510
rect 50411 20454 50471 20510
rect 51659 20454 51719 20510
rect 52907 20454 52967 20510
rect 54155 20454 54215 20510
rect 55403 20454 55463 20510
rect 56651 20454 56711 20510
rect 70966 20225 71024 20271
rect 71156 20225 71214 20271
rect 71417 20225 71475 20271
rect 71767 20225 71825 20271
rect 72028 20225 72086 20271
rect 70978 19883 71012 20225
rect 71040 19982 71106 20034
rect 71168 20031 71202 20225
rect 71156 19985 71214 20031
rect 70962 19831 71028 19883
rect 70978 19711 71012 19831
rect 71168 19711 71202 19985
rect 71429 19711 71463 20225
rect 71687 20111 71741 20120
rect 71685 20065 71743 20111
rect 71687 20056 71741 20065
rect 71697 19800 71731 20056
rect 71779 19865 71813 20225
rect 72040 20031 72074 20225
rect 72028 19985 72086 20031
rect 71907 19902 71973 19954
rect 71951 19865 72009 19871
rect 71779 19831 72009 19865
rect 71687 19791 71741 19800
rect 71685 19745 71743 19791
rect 71687 19736 71741 19745
rect 71779 19711 71813 19831
rect 71951 19825 72009 19831
rect 72040 19711 72074 19985
rect 70966 19665 71024 19711
rect 71156 19665 71214 19711
rect 71417 19665 71475 19711
rect 71767 19665 71825 19711
rect 72028 19665 72086 19711
rect 80 19552 138 19598
rect 341 19552 399 19598
rect 691 19552 749 19598
rect 952 19552 1010 19598
rect 1142 19552 1200 19598
rect 92 19358 126 19552
rect 80 19312 138 19358
rect 92 19038 126 19312
rect 193 19229 259 19281
rect 157 19192 215 19198
rect 353 19192 387 19552
rect 425 19438 479 19447
rect 423 19392 481 19438
rect 425 19383 479 19392
rect 157 19158 387 19192
rect 157 19152 215 19158
rect 353 19038 387 19158
rect 435 19127 469 19383
rect 425 19118 479 19127
rect 423 19072 481 19118
rect 425 19063 479 19072
rect 703 19038 737 19552
rect 964 19358 998 19552
rect 952 19312 1010 19358
rect 964 19038 998 19312
rect 1060 19309 1126 19361
rect 1154 19210 1188 19552
rect 1138 19158 1204 19210
rect 1154 19038 1188 19158
rect 80 18992 138 19038
rect 341 18992 399 19038
rect 691 18992 749 19038
rect 952 18992 1010 19038
rect 1142 18992 1200 19038
rect 80 17772 138 17818
rect 341 17772 399 17818
rect 691 17772 749 17818
rect 952 17772 1010 17818
rect 1142 17772 1200 17818
rect 92 17498 126 17772
rect 157 17652 215 17658
rect 353 17652 387 17772
rect 425 17738 479 17747
rect 423 17692 481 17738
rect 425 17683 479 17692
rect 157 17618 387 17652
rect 157 17612 215 17618
rect 193 17529 259 17581
rect 80 17452 138 17498
rect 92 17258 126 17452
rect 353 17258 387 17618
rect 435 17427 469 17683
rect 425 17418 479 17427
rect 423 17372 481 17418
rect 425 17363 479 17372
rect 703 17258 737 17772
rect 964 17498 998 17772
rect 1154 17652 1188 17772
rect 1138 17600 1204 17652
rect 952 17452 1010 17498
rect 964 17258 998 17452
rect 1060 17449 1126 17501
rect 1154 17258 1188 17600
rect 80 17212 138 17258
rect 341 17212 399 17258
rect 691 17212 749 17258
rect 952 17212 1010 17258
rect 1142 17212 1200 17258
rect 5686 877 5744 923
rect 5947 877 6005 923
rect 6297 877 6355 923
rect 6558 877 6616 923
rect 6748 877 6806 923
rect 6854 877 6912 923
rect 7115 877 7173 923
rect 7465 877 7523 923
rect 7726 877 7784 923
rect 7916 877 7974 923
rect 8022 877 8080 923
rect 8283 877 8341 923
rect 8633 877 8691 923
rect 8894 877 8952 923
rect 9084 877 9142 923
rect 9190 877 9248 923
rect 9451 877 9509 923
rect 9801 877 9859 923
rect 10062 877 10120 923
rect 10252 877 10310 923
rect 10358 877 10416 923
rect 10619 877 10677 923
rect 10969 877 11027 923
rect 11230 877 11288 923
rect 11420 877 11478 923
rect 11526 877 11584 923
rect 11787 877 11845 923
rect 12137 877 12195 923
rect 12398 877 12456 923
rect 12588 877 12646 923
rect 12694 877 12752 923
rect 12955 877 13013 923
rect 13305 877 13363 923
rect 13566 877 13624 923
rect 13756 877 13814 923
rect 13862 877 13920 923
rect 14123 877 14181 923
rect 14473 877 14531 923
rect 14734 877 14792 923
rect 14924 877 14982 923
rect 15030 877 15088 923
rect 15291 877 15349 923
rect 15641 877 15699 923
rect 15902 877 15960 923
rect 16092 877 16150 923
rect 16198 877 16256 923
rect 16459 877 16517 923
rect 16809 877 16867 923
rect 17070 877 17128 923
rect 17260 877 17318 923
rect 17366 877 17424 923
rect 17627 877 17685 923
rect 17977 877 18035 923
rect 18238 877 18296 923
rect 18428 877 18486 923
rect 18534 877 18592 923
rect 18795 877 18853 923
rect 19145 877 19203 923
rect 19406 877 19464 923
rect 19596 877 19654 923
rect 19702 877 19760 923
rect 19963 877 20021 923
rect 20313 877 20371 923
rect 20574 877 20632 923
rect 20764 877 20822 923
rect 20870 877 20928 923
rect 21131 877 21189 923
rect 21481 877 21539 923
rect 21742 877 21800 923
rect 21932 877 21990 923
rect 22038 877 22096 923
rect 22299 877 22357 923
rect 22649 877 22707 923
rect 22910 877 22968 923
rect 23100 877 23158 923
rect 23206 877 23264 923
rect 23467 877 23525 923
rect 23817 877 23875 923
rect 24078 877 24136 923
rect 24268 877 24326 923
rect 24374 877 24432 923
rect 24635 877 24693 923
rect 24985 877 25043 923
rect 25246 877 25304 923
rect 25436 877 25494 923
rect 25542 877 25600 923
rect 25803 877 25861 923
rect 26153 877 26211 923
rect 26414 877 26472 923
rect 26604 877 26662 923
rect 26710 877 26768 923
rect 26971 877 27029 923
rect 27321 877 27379 923
rect 27582 877 27640 923
rect 27772 877 27830 923
rect 27878 877 27936 923
rect 28139 877 28197 923
rect 28489 877 28547 923
rect 28750 877 28808 923
rect 28940 877 28998 923
rect 29046 877 29104 923
rect 29307 877 29365 923
rect 29657 877 29715 923
rect 29918 877 29976 923
rect 30108 877 30166 923
rect 30214 877 30272 923
rect 30475 877 30533 923
rect 30825 877 30883 923
rect 31086 877 31144 923
rect 31276 877 31334 923
rect 31382 877 31440 923
rect 31643 877 31701 923
rect 31993 877 32051 923
rect 32254 877 32312 923
rect 32444 877 32502 923
rect 32550 877 32608 923
rect 32811 877 32869 923
rect 33161 877 33219 923
rect 33422 877 33480 923
rect 33612 877 33670 923
rect 33718 877 33776 923
rect 33979 877 34037 923
rect 34329 877 34387 923
rect 34590 877 34648 923
rect 34780 877 34838 923
rect 34886 877 34944 923
rect 35147 877 35205 923
rect 35497 877 35555 923
rect 35758 877 35816 923
rect 35948 877 36006 923
rect 36054 877 36112 923
rect 36315 877 36373 923
rect 36665 877 36723 923
rect 36926 877 36984 923
rect 37116 877 37174 923
rect 37222 877 37280 923
rect 37483 877 37541 923
rect 37833 877 37891 923
rect 38094 877 38152 923
rect 38284 877 38342 923
rect 38390 877 38448 923
rect 38651 877 38709 923
rect 39001 877 39059 923
rect 39262 877 39320 923
rect 39452 877 39510 923
rect 39558 877 39616 923
rect 39819 877 39877 923
rect 40169 877 40227 923
rect 40430 877 40488 923
rect 40620 877 40678 923
rect 40726 877 40784 923
rect 40987 877 41045 923
rect 41337 877 41395 923
rect 41598 877 41656 923
rect 41788 877 41846 923
rect 41894 877 41952 923
rect 42155 877 42213 923
rect 42505 877 42563 923
rect 42766 877 42824 923
rect 42956 877 43014 923
rect 43062 877 43120 923
rect 43323 877 43381 923
rect 43673 877 43731 923
rect 43934 877 43992 923
rect 44124 877 44182 923
rect 44230 877 44288 923
rect 44491 877 44549 923
rect 44841 877 44899 923
rect 45102 877 45160 923
rect 45292 877 45350 923
rect 45398 877 45456 923
rect 45659 877 45717 923
rect 46009 877 46067 923
rect 46270 877 46328 923
rect 46460 877 46518 923
rect 46566 877 46624 923
rect 46827 877 46885 923
rect 47177 877 47235 923
rect 47438 877 47496 923
rect 47628 877 47686 923
rect 47734 877 47792 923
rect 47995 877 48053 923
rect 48345 877 48403 923
rect 48606 877 48664 923
rect 48796 877 48854 923
rect 5698 603 5732 877
rect 5763 757 5821 763
rect 5959 757 5993 877
rect 6031 843 6085 852
rect 6029 797 6087 843
rect 6031 788 6085 797
rect 5763 723 5993 757
rect 5763 717 5821 723
rect 5799 634 5865 686
rect 5686 557 5744 603
rect 5698 363 5732 557
rect 5959 363 5993 723
rect 6041 532 6075 788
rect 6031 523 6085 532
rect 6029 477 6087 523
rect 6031 468 6085 477
rect 6309 363 6343 877
rect 6570 603 6604 877
rect 6760 757 6794 877
rect 6744 705 6810 757
rect 6558 557 6616 603
rect 6570 363 6604 557
rect 6666 554 6732 606
rect 6760 363 6794 705
rect 6866 603 6900 877
rect 6931 757 6989 763
rect 7127 757 7161 877
rect 7199 843 7253 852
rect 7197 797 7255 843
rect 7199 788 7253 797
rect 6931 723 7161 757
rect 6931 717 6989 723
rect 6967 634 7033 686
rect 6854 557 6912 603
rect 6866 363 6900 557
rect 7127 363 7161 723
rect 7209 532 7243 788
rect 7199 523 7253 532
rect 7197 477 7255 523
rect 7199 468 7253 477
rect 7477 363 7511 877
rect 7738 603 7772 877
rect 7928 757 7962 877
rect 7912 705 7978 757
rect 7726 557 7784 603
rect 7738 363 7772 557
rect 7834 554 7900 606
rect 7928 363 7962 705
rect 8034 603 8068 877
rect 8099 757 8157 763
rect 8295 757 8329 877
rect 8367 843 8421 852
rect 8365 797 8423 843
rect 8367 788 8421 797
rect 8099 723 8329 757
rect 8099 717 8157 723
rect 8135 634 8201 686
rect 8022 557 8080 603
rect 8034 363 8068 557
rect 8295 363 8329 723
rect 8377 532 8411 788
rect 8367 523 8421 532
rect 8365 477 8423 523
rect 8367 468 8421 477
rect 8645 363 8679 877
rect 8906 603 8940 877
rect 9096 757 9130 877
rect 9080 705 9146 757
rect 8894 557 8952 603
rect 8906 363 8940 557
rect 9002 554 9068 606
rect 9096 363 9130 705
rect 9202 603 9236 877
rect 9267 757 9325 763
rect 9463 757 9497 877
rect 9535 843 9589 852
rect 9533 797 9591 843
rect 9535 788 9589 797
rect 9267 723 9497 757
rect 9267 717 9325 723
rect 9303 634 9369 686
rect 9190 557 9248 603
rect 9202 363 9236 557
rect 9463 363 9497 723
rect 9545 532 9579 788
rect 9535 523 9589 532
rect 9533 477 9591 523
rect 9535 468 9589 477
rect 9813 363 9847 877
rect 10074 603 10108 877
rect 10264 757 10298 877
rect 10248 705 10314 757
rect 10062 557 10120 603
rect 10074 363 10108 557
rect 10170 554 10236 606
rect 10264 363 10298 705
rect 10370 603 10404 877
rect 10435 757 10493 763
rect 10631 757 10665 877
rect 10703 843 10757 852
rect 10701 797 10759 843
rect 10703 788 10757 797
rect 10435 723 10665 757
rect 10435 717 10493 723
rect 10471 634 10537 686
rect 10358 557 10416 603
rect 10370 363 10404 557
rect 10631 363 10665 723
rect 10713 532 10747 788
rect 10703 523 10757 532
rect 10701 477 10759 523
rect 10703 468 10757 477
rect 10981 363 11015 877
rect 11242 603 11276 877
rect 11432 757 11466 877
rect 11416 705 11482 757
rect 11230 557 11288 603
rect 11242 363 11276 557
rect 11338 554 11404 606
rect 11432 363 11466 705
rect 11538 603 11572 877
rect 11603 757 11661 763
rect 11799 757 11833 877
rect 11871 843 11925 852
rect 11869 797 11927 843
rect 11871 788 11925 797
rect 11603 723 11833 757
rect 11603 717 11661 723
rect 11639 634 11705 686
rect 11526 557 11584 603
rect 11538 363 11572 557
rect 11799 363 11833 723
rect 11881 532 11915 788
rect 11871 523 11925 532
rect 11869 477 11927 523
rect 11871 468 11925 477
rect 12149 363 12183 877
rect 12410 603 12444 877
rect 12600 757 12634 877
rect 12584 705 12650 757
rect 12398 557 12456 603
rect 12410 363 12444 557
rect 12506 554 12572 606
rect 12600 363 12634 705
rect 12706 603 12740 877
rect 12771 757 12829 763
rect 12967 757 13001 877
rect 13039 843 13093 852
rect 13037 797 13095 843
rect 13039 788 13093 797
rect 12771 723 13001 757
rect 12771 717 12829 723
rect 12807 634 12873 686
rect 12694 557 12752 603
rect 12706 363 12740 557
rect 12967 363 13001 723
rect 13049 532 13083 788
rect 13039 523 13093 532
rect 13037 477 13095 523
rect 13039 468 13093 477
rect 13317 363 13351 877
rect 13578 603 13612 877
rect 13768 757 13802 877
rect 13752 705 13818 757
rect 13566 557 13624 603
rect 13578 363 13612 557
rect 13674 554 13740 606
rect 13768 363 13802 705
rect 13874 603 13908 877
rect 13939 757 13997 763
rect 14135 757 14169 877
rect 14207 843 14261 852
rect 14205 797 14263 843
rect 14207 788 14261 797
rect 13939 723 14169 757
rect 13939 717 13997 723
rect 13975 634 14041 686
rect 13862 557 13920 603
rect 13874 363 13908 557
rect 14135 363 14169 723
rect 14217 532 14251 788
rect 14207 523 14261 532
rect 14205 477 14263 523
rect 14207 468 14261 477
rect 14485 363 14519 877
rect 14746 603 14780 877
rect 14936 757 14970 877
rect 14920 705 14986 757
rect 14734 557 14792 603
rect 14746 363 14780 557
rect 14842 554 14908 606
rect 14936 363 14970 705
rect 15042 603 15076 877
rect 15107 757 15165 763
rect 15303 757 15337 877
rect 15375 843 15429 852
rect 15373 797 15431 843
rect 15375 788 15429 797
rect 15107 723 15337 757
rect 15107 717 15165 723
rect 15143 634 15209 686
rect 15030 557 15088 603
rect 15042 363 15076 557
rect 15303 363 15337 723
rect 15385 532 15419 788
rect 15375 523 15429 532
rect 15373 477 15431 523
rect 15375 468 15429 477
rect 15653 363 15687 877
rect 15914 603 15948 877
rect 16104 757 16138 877
rect 16088 705 16154 757
rect 15902 557 15960 603
rect 15914 363 15948 557
rect 16010 554 16076 606
rect 16104 363 16138 705
rect 16210 603 16244 877
rect 16275 757 16333 763
rect 16471 757 16505 877
rect 16543 843 16597 852
rect 16541 797 16599 843
rect 16543 788 16597 797
rect 16275 723 16505 757
rect 16275 717 16333 723
rect 16311 634 16377 686
rect 16198 557 16256 603
rect 16210 363 16244 557
rect 16471 363 16505 723
rect 16553 532 16587 788
rect 16543 523 16597 532
rect 16541 477 16599 523
rect 16543 468 16597 477
rect 16821 363 16855 877
rect 17082 603 17116 877
rect 17272 757 17306 877
rect 17256 705 17322 757
rect 17070 557 17128 603
rect 17082 363 17116 557
rect 17178 554 17244 606
rect 17272 363 17306 705
rect 17378 603 17412 877
rect 17443 757 17501 763
rect 17639 757 17673 877
rect 17711 843 17765 852
rect 17709 797 17767 843
rect 17711 788 17765 797
rect 17443 723 17673 757
rect 17443 717 17501 723
rect 17479 634 17545 686
rect 17366 557 17424 603
rect 17378 363 17412 557
rect 17639 363 17673 723
rect 17721 532 17755 788
rect 17711 523 17765 532
rect 17709 477 17767 523
rect 17711 468 17765 477
rect 17989 363 18023 877
rect 18250 603 18284 877
rect 18440 757 18474 877
rect 18424 705 18490 757
rect 18238 557 18296 603
rect 18250 363 18284 557
rect 18346 554 18412 606
rect 18440 363 18474 705
rect 18546 603 18580 877
rect 18611 757 18669 763
rect 18807 757 18841 877
rect 18879 843 18933 852
rect 18877 797 18935 843
rect 18879 788 18933 797
rect 18611 723 18841 757
rect 18611 717 18669 723
rect 18647 634 18713 686
rect 18534 557 18592 603
rect 18546 363 18580 557
rect 18807 363 18841 723
rect 18889 532 18923 788
rect 18879 523 18933 532
rect 18877 477 18935 523
rect 18879 468 18933 477
rect 19157 363 19191 877
rect 19418 603 19452 877
rect 19608 757 19642 877
rect 19592 705 19658 757
rect 19406 557 19464 603
rect 19418 363 19452 557
rect 19514 554 19580 606
rect 19608 363 19642 705
rect 19714 603 19748 877
rect 19779 757 19837 763
rect 19975 757 20009 877
rect 20047 843 20101 852
rect 20045 797 20103 843
rect 20047 788 20101 797
rect 19779 723 20009 757
rect 19779 717 19837 723
rect 19815 634 19881 686
rect 19702 557 19760 603
rect 19714 363 19748 557
rect 19975 363 20009 723
rect 20057 532 20091 788
rect 20047 523 20101 532
rect 20045 477 20103 523
rect 20047 468 20101 477
rect 20325 363 20359 877
rect 20586 603 20620 877
rect 20776 757 20810 877
rect 20760 705 20826 757
rect 20574 557 20632 603
rect 20586 363 20620 557
rect 20682 554 20748 606
rect 20776 363 20810 705
rect 20882 603 20916 877
rect 20947 757 21005 763
rect 21143 757 21177 877
rect 21215 843 21269 852
rect 21213 797 21271 843
rect 21215 788 21269 797
rect 20947 723 21177 757
rect 20947 717 21005 723
rect 20983 634 21049 686
rect 20870 557 20928 603
rect 20882 363 20916 557
rect 21143 363 21177 723
rect 21225 532 21259 788
rect 21215 523 21269 532
rect 21213 477 21271 523
rect 21215 468 21269 477
rect 21493 363 21527 877
rect 21754 603 21788 877
rect 21944 757 21978 877
rect 21928 705 21994 757
rect 21742 557 21800 603
rect 21754 363 21788 557
rect 21850 554 21916 606
rect 21944 363 21978 705
rect 22050 603 22084 877
rect 22115 757 22173 763
rect 22311 757 22345 877
rect 22383 843 22437 852
rect 22381 797 22439 843
rect 22383 788 22437 797
rect 22115 723 22345 757
rect 22115 717 22173 723
rect 22151 634 22217 686
rect 22038 557 22096 603
rect 22050 363 22084 557
rect 22311 363 22345 723
rect 22393 532 22427 788
rect 22383 523 22437 532
rect 22381 477 22439 523
rect 22383 468 22437 477
rect 22661 363 22695 877
rect 22922 603 22956 877
rect 23112 757 23146 877
rect 23096 705 23162 757
rect 22910 557 22968 603
rect 22922 363 22956 557
rect 23018 554 23084 606
rect 23112 363 23146 705
rect 23218 603 23252 877
rect 23283 757 23341 763
rect 23479 757 23513 877
rect 23551 843 23605 852
rect 23549 797 23607 843
rect 23551 788 23605 797
rect 23283 723 23513 757
rect 23283 717 23341 723
rect 23319 634 23385 686
rect 23206 557 23264 603
rect 23218 363 23252 557
rect 23479 363 23513 723
rect 23561 532 23595 788
rect 23551 523 23605 532
rect 23549 477 23607 523
rect 23551 468 23605 477
rect 23829 363 23863 877
rect 24090 603 24124 877
rect 24280 757 24314 877
rect 24264 705 24330 757
rect 24078 557 24136 603
rect 24090 363 24124 557
rect 24186 554 24252 606
rect 24280 363 24314 705
rect 24386 603 24420 877
rect 24451 757 24509 763
rect 24647 757 24681 877
rect 24719 843 24773 852
rect 24717 797 24775 843
rect 24719 788 24773 797
rect 24451 723 24681 757
rect 24451 717 24509 723
rect 24487 634 24553 686
rect 24374 557 24432 603
rect 24386 363 24420 557
rect 24647 363 24681 723
rect 24729 532 24763 788
rect 24719 523 24773 532
rect 24717 477 24775 523
rect 24719 468 24773 477
rect 24997 363 25031 877
rect 25258 603 25292 877
rect 25448 757 25482 877
rect 25432 705 25498 757
rect 25246 557 25304 603
rect 25258 363 25292 557
rect 25354 554 25420 606
rect 25448 363 25482 705
rect 25554 603 25588 877
rect 25619 757 25677 763
rect 25815 757 25849 877
rect 25887 843 25941 852
rect 25885 797 25943 843
rect 25887 788 25941 797
rect 25619 723 25849 757
rect 25619 717 25677 723
rect 25655 634 25721 686
rect 25542 557 25600 603
rect 25554 363 25588 557
rect 25815 363 25849 723
rect 25897 532 25931 788
rect 25887 523 25941 532
rect 25885 477 25943 523
rect 25887 468 25941 477
rect 26165 363 26199 877
rect 26426 603 26460 877
rect 26616 757 26650 877
rect 26600 705 26666 757
rect 26414 557 26472 603
rect 26426 363 26460 557
rect 26522 554 26588 606
rect 26616 363 26650 705
rect 26722 603 26756 877
rect 26787 757 26845 763
rect 26983 757 27017 877
rect 27055 843 27109 852
rect 27053 797 27111 843
rect 27055 788 27109 797
rect 26787 723 27017 757
rect 26787 717 26845 723
rect 26823 634 26889 686
rect 26710 557 26768 603
rect 26722 363 26756 557
rect 26983 363 27017 723
rect 27065 532 27099 788
rect 27055 523 27109 532
rect 27053 477 27111 523
rect 27055 468 27109 477
rect 27333 363 27367 877
rect 27594 603 27628 877
rect 27784 757 27818 877
rect 27768 705 27834 757
rect 27582 557 27640 603
rect 27594 363 27628 557
rect 27690 554 27756 606
rect 27784 363 27818 705
rect 27890 603 27924 877
rect 27955 757 28013 763
rect 28151 757 28185 877
rect 28223 843 28277 852
rect 28221 797 28279 843
rect 28223 788 28277 797
rect 27955 723 28185 757
rect 27955 717 28013 723
rect 27991 634 28057 686
rect 27878 557 27936 603
rect 27890 363 27924 557
rect 28151 363 28185 723
rect 28233 532 28267 788
rect 28223 523 28277 532
rect 28221 477 28279 523
rect 28223 468 28277 477
rect 28501 363 28535 877
rect 28762 603 28796 877
rect 28952 757 28986 877
rect 28936 705 29002 757
rect 28750 557 28808 603
rect 28762 363 28796 557
rect 28858 554 28924 606
rect 28952 363 28986 705
rect 29058 603 29092 877
rect 29123 757 29181 763
rect 29319 757 29353 877
rect 29391 843 29445 852
rect 29389 797 29447 843
rect 29391 788 29445 797
rect 29123 723 29353 757
rect 29123 717 29181 723
rect 29159 634 29225 686
rect 29046 557 29104 603
rect 29058 363 29092 557
rect 29319 363 29353 723
rect 29401 532 29435 788
rect 29391 523 29445 532
rect 29389 477 29447 523
rect 29391 468 29445 477
rect 29669 363 29703 877
rect 29930 603 29964 877
rect 30120 757 30154 877
rect 30104 705 30170 757
rect 29918 557 29976 603
rect 29930 363 29964 557
rect 30026 554 30092 606
rect 30120 363 30154 705
rect 30226 603 30260 877
rect 30291 757 30349 763
rect 30487 757 30521 877
rect 30559 843 30613 852
rect 30557 797 30615 843
rect 30559 788 30613 797
rect 30291 723 30521 757
rect 30291 717 30349 723
rect 30327 634 30393 686
rect 30214 557 30272 603
rect 30226 363 30260 557
rect 30487 363 30521 723
rect 30569 532 30603 788
rect 30559 523 30613 532
rect 30557 477 30615 523
rect 30559 468 30613 477
rect 30837 363 30871 877
rect 31098 603 31132 877
rect 31288 757 31322 877
rect 31272 705 31338 757
rect 31086 557 31144 603
rect 31098 363 31132 557
rect 31194 554 31260 606
rect 31288 363 31322 705
rect 31394 603 31428 877
rect 31459 757 31517 763
rect 31655 757 31689 877
rect 31727 843 31781 852
rect 31725 797 31783 843
rect 31727 788 31781 797
rect 31459 723 31689 757
rect 31459 717 31517 723
rect 31495 634 31561 686
rect 31382 557 31440 603
rect 31394 363 31428 557
rect 31655 363 31689 723
rect 31737 532 31771 788
rect 31727 523 31781 532
rect 31725 477 31783 523
rect 31727 468 31781 477
rect 32005 363 32039 877
rect 32266 603 32300 877
rect 32456 757 32490 877
rect 32440 705 32506 757
rect 32254 557 32312 603
rect 32266 363 32300 557
rect 32362 554 32428 606
rect 32456 363 32490 705
rect 32562 603 32596 877
rect 32627 757 32685 763
rect 32823 757 32857 877
rect 32895 843 32949 852
rect 32893 797 32951 843
rect 32895 788 32949 797
rect 32627 723 32857 757
rect 32627 717 32685 723
rect 32663 634 32729 686
rect 32550 557 32608 603
rect 32562 363 32596 557
rect 32823 363 32857 723
rect 32905 532 32939 788
rect 32895 523 32949 532
rect 32893 477 32951 523
rect 32895 468 32949 477
rect 33173 363 33207 877
rect 33434 603 33468 877
rect 33624 757 33658 877
rect 33608 705 33674 757
rect 33422 557 33480 603
rect 33434 363 33468 557
rect 33530 554 33596 606
rect 33624 363 33658 705
rect 33730 603 33764 877
rect 33795 757 33853 763
rect 33991 757 34025 877
rect 34063 843 34117 852
rect 34061 797 34119 843
rect 34063 788 34117 797
rect 33795 723 34025 757
rect 33795 717 33853 723
rect 33831 634 33897 686
rect 33718 557 33776 603
rect 33730 363 33764 557
rect 33991 363 34025 723
rect 34073 532 34107 788
rect 34063 523 34117 532
rect 34061 477 34119 523
rect 34063 468 34117 477
rect 34341 363 34375 877
rect 34602 603 34636 877
rect 34792 757 34826 877
rect 34776 705 34842 757
rect 34590 557 34648 603
rect 34602 363 34636 557
rect 34698 554 34764 606
rect 34792 363 34826 705
rect 34898 603 34932 877
rect 34963 757 35021 763
rect 35159 757 35193 877
rect 35231 843 35285 852
rect 35229 797 35287 843
rect 35231 788 35285 797
rect 34963 723 35193 757
rect 34963 717 35021 723
rect 34999 634 35065 686
rect 34886 557 34944 603
rect 34898 363 34932 557
rect 35159 363 35193 723
rect 35241 532 35275 788
rect 35231 523 35285 532
rect 35229 477 35287 523
rect 35231 468 35285 477
rect 35509 363 35543 877
rect 35770 603 35804 877
rect 35960 757 35994 877
rect 35944 705 36010 757
rect 35758 557 35816 603
rect 35770 363 35804 557
rect 35866 554 35932 606
rect 35960 363 35994 705
rect 36066 603 36100 877
rect 36131 757 36189 763
rect 36327 757 36361 877
rect 36399 843 36453 852
rect 36397 797 36455 843
rect 36399 788 36453 797
rect 36131 723 36361 757
rect 36131 717 36189 723
rect 36167 634 36233 686
rect 36054 557 36112 603
rect 36066 363 36100 557
rect 36327 363 36361 723
rect 36409 532 36443 788
rect 36399 523 36453 532
rect 36397 477 36455 523
rect 36399 468 36453 477
rect 36677 363 36711 877
rect 36938 603 36972 877
rect 37128 757 37162 877
rect 37112 705 37178 757
rect 36926 557 36984 603
rect 36938 363 36972 557
rect 37034 554 37100 606
rect 37128 363 37162 705
rect 37234 603 37268 877
rect 37299 757 37357 763
rect 37495 757 37529 877
rect 37567 843 37621 852
rect 37565 797 37623 843
rect 37567 788 37621 797
rect 37299 723 37529 757
rect 37299 717 37357 723
rect 37335 634 37401 686
rect 37222 557 37280 603
rect 37234 363 37268 557
rect 37495 363 37529 723
rect 37577 532 37611 788
rect 37567 523 37621 532
rect 37565 477 37623 523
rect 37567 468 37621 477
rect 37845 363 37879 877
rect 38106 603 38140 877
rect 38296 757 38330 877
rect 38280 705 38346 757
rect 38094 557 38152 603
rect 38106 363 38140 557
rect 38202 554 38268 606
rect 38296 363 38330 705
rect 38402 603 38436 877
rect 38467 757 38525 763
rect 38663 757 38697 877
rect 38735 843 38789 852
rect 38733 797 38791 843
rect 38735 788 38789 797
rect 38467 723 38697 757
rect 38467 717 38525 723
rect 38503 634 38569 686
rect 38390 557 38448 603
rect 38402 363 38436 557
rect 38663 363 38697 723
rect 38745 532 38779 788
rect 38735 523 38789 532
rect 38733 477 38791 523
rect 38735 468 38789 477
rect 39013 363 39047 877
rect 39274 603 39308 877
rect 39464 757 39498 877
rect 39448 705 39514 757
rect 39262 557 39320 603
rect 39274 363 39308 557
rect 39370 554 39436 606
rect 39464 363 39498 705
rect 39570 603 39604 877
rect 39635 757 39693 763
rect 39831 757 39865 877
rect 39903 843 39957 852
rect 39901 797 39959 843
rect 39903 788 39957 797
rect 39635 723 39865 757
rect 39635 717 39693 723
rect 39671 634 39737 686
rect 39558 557 39616 603
rect 39570 363 39604 557
rect 39831 363 39865 723
rect 39913 532 39947 788
rect 39903 523 39957 532
rect 39901 477 39959 523
rect 39903 468 39957 477
rect 40181 363 40215 877
rect 40442 603 40476 877
rect 40632 757 40666 877
rect 40616 705 40682 757
rect 40430 557 40488 603
rect 40442 363 40476 557
rect 40538 554 40604 606
rect 40632 363 40666 705
rect 40738 603 40772 877
rect 40803 757 40861 763
rect 40999 757 41033 877
rect 41071 843 41125 852
rect 41069 797 41127 843
rect 41071 788 41125 797
rect 40803 723 41033 757
rect 40803 717 40861 723
rect 40839 634 40905 686
rect 40726 557 40784 603
rect 40738 363 40772 557
rect 40999 363 41033 723
rect 41081 532 41115 788
rect 41071 523 41125 532
rect 41069 477 41127 523
rect 41071 468 41125 477
rect 41349 363 41383 877
rect 41610 603 41644 877
rect 41800 757 41834 877
rect 41784 705 41850 757
rect 41598 557 41656 603
rect 41610 363 41644 557
rect 41706 554 41772 606
rect 41800 363 41834 705
rect 41906 603 41940 877
rect 41971 757 42029 763
rect 42167 757 42201 877
rect 42239 843 42293 852
rect 42237 797 42295 843
rect 42239 788 42293 797
rect 41971 723 42201 757
rect 41971 717 42029 723
rect 42007 634 42073 686
rect 41894 557 41952 603
rect 41906 363 41940 557
rect 42167 363 42201 723
rect 42249 532 42283 788
rect 42239 523 42293 532
rect 42237 477 42295 523
rect 42239 468 42293 477
rect 42517 363 42551 877
rect 42778 603 42812 877
rect 42968 757 43002 877
rect 42952 705 43018 757
rect 42766 557 42824 603
rect 42778 363 42812 557
rect 42874 554 42940 606
rect 42968 363 43002 705
rect 43074 603 43108 877
rect 43139 757 43197 763
rect 43335 757 43369 877
rect 43407 843 43461 852
rect 43405 797 43463 843
rect 43407 788 43461 797
rect 43139 723 43369 757
rect 43139 717 43197 723
rect 43175 634 43241 686
rect 43062 557 43120 603
rect 43074 363 43108 557
rect 43335 363 43369 723
rect 43417 532 43451 788
rect 43407 523 43461 532
rect 43405 477 43463 523
rect 43407 468 43461 477
rect 43685 363 43719 877
rect 43946 603 43980 877
rect 44136 757 44170 877
rect 44120 705 44186 757
rect 43934 557 43992 603
rect 43946 363 43980 557
rect 44042 554 44108 606
rect 44136 363 44170 705
rect 44242 603 44276 877
rect 44307 757 44365 763
rect 44503 757 44537 877
rect 44575 843 44629 852
rect 44573 797 44631 843
rect 44575 788 44629 797
rect 44307 723 44537 757
rect 44307 717 44365 723
rect 44343 634 44409 686
rect 44230 557 44288 603
rect 44242 363 44276 557
rect 44503 363 44537 723
rect 44585 532 44619 788
rect 44575 523 44629 532
rect 44573 477 44631 523
rect 44575 468 44629 477
rect 44853 363 44887 877
rect 45114 603 45148 877
rect 45304 757 45338 877
rect 45288 705 45354 757
rect 45102 557 45160 603
rect 45114 363 45148 557
rect 45210 554 45276 606
rect 45304 363 45338 705
rect 45410 603 45444 877
rect 45475 757 45533 763
rect 45671 757 45705 877
rect 45743 843 45797 852
rect 45741 797 45799 843
rect 45743 788 45797 797
rect 45475 723 45705 757
rect 45475 717 45533 723
rect 45511 634 45577 686
rect 45398 557 45456 603
rect 45410 363 45444 557
rect 45671 363 45705 723
rect 45753 532 45787 788
rect 45743 523 45797 532
rect 45741 477 45799 523
rect 45743 468 45797 477
rect 46021 363 46055 877
rect 46282 603 46316 877
rect 46472 757 46506 877
rect 46456 705 46522 757
rect 46270 557 46328 603
rect 46282 363 46316 557
rect 46378 554 46444 606
rect 46472 363 46506 705
rect 46578 603 46612 877
rect 46643 757 46701 763
rect 46839 757 46873 877
rect 46911 843 46965 852
rect 46909 797 46967 843
rect 46911 788 46965 797
rect 46643 723 46873 757
rect 46643 717 46701 723
rect 46679 634 46745 686
rect 46566 557 46624 603
rect 46578 363 46612 557
rect 46839 363 46873 723
rect 46921 532 46955 788
rect 46911 523 46965 532
rect 46909 477 46967 523
rect 46911 468 46965 477
rect 47189 363 47223 877
rect 47450 603 47484 877
rect 47640 757 47674 877
rect 47624 705 47690 757
rect 47438 557 47496 603
rect 47450 363 47484 557
rect 47546 554 47612 606
rect 47640 363 47674 705
rect 47746 603 47780 877
rect 47811 757 47869 763
rect 48007 757 48041 877
rect 48079 843 48133 852
rect 48077 797 48135 843
rect 48079 788 48133 797
rect 47811 723 48041 757
rect 47811 717 47869 723
rect 47847 634 47913 686
rect 47734 557 47792 603
rect 47746 363 47780 557
rect 48007 363 48041 723
rect 48089 532 48123 788
rect 48079 523 48133 532
rect 48077 477 48135 523
rect 48079 468 48133 477
rect 48357 363 48391 877
rect 48618 603 48652 877
rect 48808 757 48842 877
rect 48792 705 48858 757
rect 48606 557 48664 603
rect 48618 363 48652 557
rect 48714 554 48780 606
rect 48808 363 48842 705
rect 5686 317 5744 363
rect 5947 317 6005 363
rect 6297 317 6355 363
rect 6558 317 6616 363
rect 6748 317 6806 363
rect 6854 317 6912 363
rect 7115 317 7173 363
rect 7465 317 7523 363
rect 7726 317 7784 363
rect 7916 317 7974 363
rect 8022 317 8080 363
rect 8283 317 8341 363
rect 8633 317 8691 363
rect 8894 317 8952 363
rect 9084 317 9142 363
rect 9190 317 9248 363
rect 9451 317 9509 363
rect 9801 317 9859 363
rect 10062 317 10120 363
rect 10252 317 10310 363
rect 10358 317 10416 363
rect 10619 317 10677 363
rect 10969 317 11027 363
rect 11230 317 11288 363
rect 11420 317 11478 363
rect 11526 317 11584 363
rect 11787 317 11845 363
rect 12137 317 12195 363
rect 12398 317 12456 363
rect 12588 317 12646 363
rect 12694 317 12752 363
rect 12955 317 13013 363
rect 13305 317 13363 363
rect 13566 317 13624 363
rect 13756 317 13814 363
rect 13862 317 13920 363
rect 14123 317 14181 363
rect 14473 317 14531 363
rect 14734 317 14792 363
rect 14924 317 14982 363
rect 15030 317 15088 363
rect 15291 317 15349 363
rect 15641 317 15699 363
rect 15902 317 15960 363
rect 16092 317 16150 363
rect 16198 317 16256 363
rect 16459 317 16517 363
rect 16809 317 16867 363
rect 17070 317 17128 363
rect 17260 317 17318 363
rect 17366 317 17424 363
rect 17627 317 17685 363
rect 17977 317 18035 363
rect 18238 317 18296 363
rect 18428 317 18486 363
rect 18534 317 18592 363
rect 18795 317 18853 363
rect 19145 317 19203 363
rect 19406 317 19464 363
rect 19596 317 19654 363
rect 19702 317 19760 363
rect 19963 317 20021 363
rect 20313 317 20371 363
rect 20574 317 20632 363
rect 20764 317 20822 363
rect 20870 317 20928 363
rect 21131 317 21189 363
rect 21481 317 21539 363
rect 21742 317 21800 363
rect 21932 317 21990 363
rect 22038 317 22096 363
rect 22299 317 22357 363
rect 22649 317 22707 363
rect 22910 317 22968 363
rect 23100 317 23158 363
rect 23206 317 23264 363
rect 23467 317 23525 363
rect 23817 317 23875 363
rect 24078 317 24136 363
rect 24268 317 24326 363
rect 24374 317 24432 363
rect 24635 317 24693 363
rect 24985 317 25043 363
rect 25246 317 25304 363
rect 25436 317 25494 363
rect 25542 317 25600 363
rect 25803 317 25861 363
rect 26153 317 26211 363
rect 26414 317 26472 363
rect 26604 317 26662 363
rect 26710 317 26768 363
rect 26971 317 27029 363
rect 27321 317 27379 363
rect 27582 317 27640 363
rect 27772 317 27830 363
rect 27878 317 27936 363
rect 28139 317 28197 363
rect 28489 317 28547 363
rect 28750 317 28808 363
rect 28940 317 28998 363
rect 29046 317 29104 363
rect 29307 317 29365 363
rect 29657 317 29715 363
rect 29918 317 29976 363
rect 30108 317 30166 363
rect 30214 317 30272 363
rect 30475 317 30533 363
rect 30825 317 30883 363
rect 31086 317 31144 363
rect 31276 317 31334 363
rect 31382 317 31440 363
rect 31643 317 31701 363
rect 31993 317 32051 363
rect 32254 317 32312 363
rect 32444 317 32502 363
rect 32550 317 32608 363
rect 32811 317 32869 363
rect 33161 317 33219 363
rect 33422 317 33480 363
rect 33612 317 33670 363
rect 33718 317 33776 363
rect 33979 317 34037 363
rect 34329 317 34387 363
rect 34590 317 34648 363
rect 34780 317 34838 363
rect 34886 317 34944 363
rect 35147 317 35205 363
rect 35497 317 35555 363
rect 35758 317 35816 363
rect 35948 317 36006 363
rect 36054 317 36112 363
rect 36315 317 36373 363
rect 36665 317 36723 363
rect 36926 317 36984 363
rect 37116 317 37174 363
rect 37222 317 37280 363
rect 37483 317 37541 363
rect 37833 317 37891 363
rect 38094 317 38152 363
rect 38284 317 38342 363
rect 38390 317 38448 363
rect 38651 317 38709 363
rect 39001 317 39059 363
rect 39262 317 39320 363
rect 39452 317 39510 363
rect 39558 317 39616 363
rect 39819 317 39877 363
rect 40169 317 40227 363
rect 40430 317 40488 363
rect 40620 317 40678 363
rect 40726 317 40784 363
rect 40987 317 41045 363
rect 41337 317 41395 363
rect 41598 317 41656 363
rect 41788 317 41846 363
rect 41894 317 41952 363
rect 42155 317 42213 363
rect 42505 317 42563 363
rect 42766 317 42824 363
rect 42956 317 43014 363
rect 43062 317 43120 363
rect 43323 317 43381 363
rect 43673 317 43731 363
rect 43934 317 43992 363
rect 44124 317 44182 363
rect 44230 317 44288 363
rect 44491 317 44549 363
rect 44841 317 44899 363
rect 45102 317 45160 363
rect 45292 317 45350 363
rect 45398 317 45456 363
rect 45659 317 45717 363
rect 46009 317 46067 363
rect 46270 317 46328 363
rect 46460 317 46518 363
rect 46566 317 46624 363
rect 46827 317 46885 363
rect 47177 317 47235 363
rect 47438 317 47496 363
rect 47628 317 47686 363
rect 47734 317 47792 363
rect 47995 317 48053 363
rect 48345 317 48403 363
rect 48606 317 48664 363
rect 48796 317 48854 363
<< obsm2 >>
rect 73412 88728 73440 88756
rect 74226 88737 74292 88789
rect 72589 88564 72617 88592
rect 74148 88586 74214 88638
rect 74899 88555 74927 89247
rect 75093 88657 75159 88709
rect 70942 88526 71088 88554
rect 74873 88491 74927 88555
rect 68442 88317 68508 88369
rect 73756 88341 73784 88369
rect 67575 88237 67641 88289
rect 68520 88166 68586 88218
rect 67807 88071 67861 88135
rect 74899 87833 74927 88491
rect 3695 85715 3749 85779
rect 4408 85632 4474 85684
rect 3463 85561 3529 85613
rect 4330 85481 4396 85533
rect 4330 84513 4396 84565
rect 3463 84433 3529 84485
rect 4408 84362 4474 84414
rect 3695 84267 3749 84331
rect 3695 82887 3749 82951
rect 4408 82804 4474 82856
rect 3463 82733 3529 82785
rect 4330 82653 4396 82705
rect 4330 81685 4396 81737
rect 3463 81605 3529 81657
rect 4408 81534 4474 81586
rect 17708 81570 58268 81598
rect 3695 81439 3749 81503
rect 17084 80319 58268 80429
rect 16418 80136 58934 80184
rect 3695 80059 3749 80123
rect 16898 80122 16980 80136
rect 17188 80122 17270 80136
rect 18146 80122 18228 80136
rect 18436 80122 18518 80136
rect 19394 80122 19476 80136
rect 19684 80122 19766 80136
rect 20642 80122 20724 80136
rect 20932 80122 21014 80136
rect 21890 80122 21972 80136
rect 22180 80122 22262 80136
rect 23138 80122 23220 80136
rect 23428 80122 23510 80136
rect 24386 80122 24468 80136
rect 24676 80122 24758 80136
rect 25634 80122 25716 80136
rect 25924 80122 26006 80136
rect 26882 80122 26964 80136
rect 27172 80122 27254 80136
rect 28130 80122 28212 80136
rect 28420 80122 28502 80136
rect 29378 80122 29460 80136
rect 29668 80122 29750 80136
rect 30626 80122 30708 80136
rect 30916 80122 30998 80136
rect 31874 80122 31956 80136
rect 32164 80122 32246 80136
rect 33122 80122 33204 80136
rect 33412 80122 33494 80136
rect 34370 80122 34452 80136
rect 34660 80122 34742 80136
rect 35618 80122 35700 80136
rect 35908 80122 35990 80136
rect 36866 80122 36948 80136
rect 37156 80122 37238 80136
rect 38114 80122 38196 80136
rect 38404 80122 38486 80136
rect 39362 80122 39444 80136
rect 39652 80122 39734 80136
rect 40610 80122 40692 80136
rect 40900 80122 40982 80136
rect 41858 80122 41940 80136
rect 42148 80122 42230 80136
rect 43106 80122 43188 80136
rect 43396 80122 43478 80136
rect 44354 80122 44436 80136
rect 44644 80122 44726 80136
rect 45602 80122 45684 80136
rect 45892 80122 45974 80136
rect 46850 80122 46932 80136
rect 47140 80122 47222 80136
rect 48098 80122 48180 80136
rect 48388 80122 48470 80136
rect 49346 80122 49428 80136
rect 49636 80122 49718 80136
rect 50594 80122 50676 80136
rect 50884 80122 50966 80136
rect 51842 80122 51924 80136
rect 52132 80122 52214 80136
rect 53090 80122 53172 80136
rect 53380 80122 53462 80136
rect 54338 80122 54420 80136
rect 54628 80122 54710 80136
rect 55586 80122 55668 80136
rect 55876 80122 55958 80136
rect 56834 80122 56916 80136
rect 57124 80122 57206 80136
rect 58082 80122 58164 80136
rect 58372 80122 58454 80136
rect 16418 80074 16864 80088
rect 17014 80074 17154 80088
rect 17304 80074 18112 80088
rect 18262 80074 18402 80088
rect 18552 80074 19360 80088
rect 19510 80074 19650 80088
rect 19800 80074 20608 80088
rect 20758 80074 20898 80088
rect 21048 80074 21856 80088
rect 22006 80074 22146 80088
rect 22296 80074 23104 80088
rect 23254 80074 23394 80088
rect 23544 80074 24352 80088
rect 24502 80074 24642 80088
rect 24792 80074 25600 80088
rect 25750 80074 25890 80088
rect 26040 80074 26848 80088
rect 26998 80074 27138 80088
rect 27288 80074 28096 80088
rect 28246 80074 28386 80088
rect 28536 80074 29344 80088
rect 29494 80074 29634 80088
rect 29784 80074 30592 80088
rect 30742 80074 30882 80088
rect 31032 80074 31840 80088
rect 31990 80074 32130 80088
rect 32280 80074 33088 80088
rect 33238 80074 33378 80088
rect 33528 80074 34336 80088
rect 34486 80074 34626 80088
rect 34776 80074 35584 80088
rect 35734 80074 35874 80088
rect 36024 80074 36832 80088
rect 36982 80074 37122 80088
rect 37272 80074 38080 80088
rect 38230 80074 38370 80088
rect 38520 80074 39328 80088
rect 39478 80074 39618 80088
rect 39768 80074 40576 80088
rect 40726 80074 40866 80088
rect 41016 80074 41824 80088
rect 41974 80074 42114 80088
rect 42264 80074 43072 80088
rect 43222 80074 43362 80088
rect 43512 80074 44320 80088
rect 44470 80074 44610 80088
rect 44760 80074 45568 80088
rect 45718 80074 45858 80088
rect 46008 80074 46816 80088
rect 46966 80074 47106 80088
rect 47256 80074 48064 80088
rect 48214 80074 48354 80088
rect 48504 80074 49312 80088
rect 49462 80074 49602 80088
rect 49752 80074 50560 80088
rect 50710 80074 50850 80088
rect 51000 80074 51808 80088
rect 51958 80074 52098 80088
rect 52248 80074 53056 80088
rect 53206 80074 53346 80088
rect 53496 80074 54304 80088
rect 54454 80074 54594 80088
rect 54744 80074 55552 80088
rect 55702 80074 55842 80088
rect 55992 80074 56800 80088
rect 56950 80074 57090 80088
rect 57240 80074 58048 80088
rect 58198 80074 58338 80088
rect 58488 80074 58934 80088
rect 4408 79976 4474 80028
rect 16418 80026 58934 80074
rect 16418 80012 16864 80026
rect 17014 80012 17154 80026
rect 17304 80012 18112 80026
rect 18262 80012 18402 80026
rect 18552 80012 19360 80026
rect 19510 80012 19650 80026
rect 19800 80012 20608 80026
rect 20758 80012 20898 80026
rect 21048 80012 21856 80026
rect 22006 80012 22146 80026
rect 22296 80012 23104 80026
rect 23254 80012 23394 80026
rect 23544 80012 24352 80026
rect 24502 80012 24642 80026
rect 24792 80012 25600 80026
rect 25750 80012 25890 80026
rect 26040 80012 26848 80026
rect 26998 80012 27138 80026
rect 27288 80012 28096 80026
rect 28246 80012 28386 80026
rect 28536 80012 29344 80026
rect 29494 80012 29634 80026
rect 29784 80012 30592 80026
rect 30742 80012 30882 80026
rect 31032 80012 31840 80026
rect 31990 80012 32130 80026
rect 32280 80012 33088 80026
rect 33238 80012 33378 80026
rect 33528 80012 34336 80026
rect 34486 80012 34626 80026
rect 34776 80012 35584 80026
rect 35734 80012 35874 80026
rect 36024 80012 36832 80026
rect 36982 80012 37122 80026
rect 37272 80012 38080 80026
rect 38230 80012 38370 80026
rect 38520 80012 39328 80026
rect 39478 80012 39618 80026
rect 39768 80012 40576 80026
rect 40726 80012 40866 80026
rect 41016 80012 41824 80026
rect 41974 80012 42114 80026
rect 42264 80012 43072 80026
rect 43222 80012 43362 80026
rect 43512 80012 44320 80026
rect 44470 80012 44610 80026
rect 44760 80012 45568 80026
rect 45718 80012 45858 80026
rect 46008 80012 46816 80026
rect 46966 80012 47106 80026
rect 47256 80012 48064 80026
rect 48214 80012 48354 80026
rect 48504 80012 49312 80026
rect 49462 80012 49602 80026
rect 49752 80012 50560 80026
rect 50710 80012 50850 80026
rect 51000 80012 51808 80026
rect 51958 80012 52098 80026
rect 52248 80012 53056 80026
rect 53206 80012 53346 80026
rect 53496 80012 54304 80026
rect 54454 80012 54594 80026
rect 54744 80012 55552 80026
rect 55702 80012 55842 80026
rect 55992 80012 56800 80026
rect 56950 80012 57090 80026
rect 57240 80012 58048 80026
rect 58198 80012 58338 80026
rect 58488 80012 58934 80026
rect 16898 79964 16980 79978
rect 17188 79964 17270 79978
rect 18146 79964 18228 79978
rect 18436 79964 18518 79978
rect 19394 79964 19476 79978
rect 19684 79964 19766 79978
rect 20642 79964 20724 79978
rect 20932 79964 21014 79978
rect 21890 79964 21972 79978
rect 22180 79964 22262 79978
rect 23138 79964 23220 79978
rect 23428 79964 23510 79978
rect 24386 79964 24468 79978
rect 24676 79964 24758 79978
rect 25634 79964 25716 79978
rect 25924 79964 26006 79978
rect 26882 79964 26964 79978
rect 27172 79964 27254 79978
rect 28130 79964 28212 79978
rect 28420 79964 28502 79978
rect 29378 79964 29460 79978
rect 29668 79964 29750 79978
rect 30626 79964 30708 79978
rect 30916 79964 30998 79978
rect 31874 79964 31956 79978
rect 32164 79964 32246 79978
rect 33122 79964 33204 79978
rect 33412 79964 33494 79978
rect 34370 79964 34452 79978
rect 34660 79964 34742 79978
rect 35618 79964 35700 79978
rect 35908 79964 35990 79978
rect 36866 79964 36948 79978
rect 37156 79964 37238 79978
rect 38114 79964 38196 79978
rect 38404 79964 38486 79978
rect 39362 79964 39444 79978
rect 39652 79964 39734 79978
rect 40610 79964 40692 79978
rect 40900 79964 40982 79978
rect 41858 79964 41940 79978
rect 42148 79964 42230 79978
rect 43106 79964 43188 79978
rect 43396 79964 43478 79978
rect 44354 79964 44436 79978
rect 44644 79964 44726 79978
rect 45602 79964 45684 79978
rect 45892 79964 45974 79978
rect 46850 79964 46932 79978
rect 47140 79964 47222 79978
rect 48098 79964 48180 79978
rect 48388 79964 48470 79978
rect 49346 79964 49428 79978
rect 49636 79964 49718 79978
rect 50594 79964 50676 79978
rect 50884 79964 50966 79978
rect 51842 79964 51924 79978
rect 52132 79964 52214 79978
rect 53090 79964 53172 79978
rect 53380 79964 53462 79978
rect 54338 79964 54420 79978
rect 54628 79964 54710 79978
rect 55586 79964 55668 79978
rect 55876 79964 55958 79978
rect 56834 79964 56916 79978
rect 57124 79964 57206 79978
rect 58082 79964 58164 79978
rect 58372 79964 58454 79978
rect 59016 79973 59044 86437
rect 59140 79973 59168 86437
rect 59264 79973 59292 86437
rect 70942 84284 71088 84312
rect 70942 82870 71136 82898
rect 70942 81456 72010 81484
rect 73520 80081 73548 80603
rect 3463 79905 3529 79957
rect 16418 79916 58934 79964
rect 4330 79825 4396 79877
rect 4330 78857 4396 78909
rect 3463 78777 3529 78829
rect 4408 78706 4474 78758
rect 3695 78611 3749 78675
rect 3695 77231 3749 77295
rect 4408 77148 4474 77200
rect 3463 77077 3529 77129
rect 4330 76997 4396 77049
rect 245 28463 273 37945
rect 12244 29253 12272 79813
rect 16418 79758 58934 79868
rect 16418 79662 58934 79710
rect 16898 79648 16980 79662
rect 17188 79648 17270 79662
rect 18146 79648 18228 79662
rect 18436 79648 18518 79662
rect 19394 79648 19476 79662
rect 19684 79648 19766 79662
rect 20642 79648 20724 79662
rect 20932 79648 21014 79662
rect 21890 79648 21972 79662
rect 22180 79648 22262 79662
rect 23138 79648 23220 79662
rect 23428 79648 23510 79662
rect 24386 79648 24468 79662
rect 24676 79648 24758 79662
rect 25634 79648 25716 79662
rect 25924 79648 26006 79662
rect 26882 79648 26964 79662
rect 27172 79648 27254 79662
rect 28130 79648 28212 79662
rect 28420 79648 28502 79662
rect 29378 79648 29460 79662
rect 29668 79648 29750 79662
rect 30626 79648 30708 79662
rect 30916 79648 30998 79662
rect 31874 79648 31956 79662
rect 32164 79648 32246 79662
rect 33122 79648 33204 79662
rect 33412 79648 33494 79662
rect 34370 79648 34452 79662
rect 34660 79648 34742 79662
rect 35618 79648 35700 79662
rect 35908 79648 35990 79662
rect 36866 79648 36948 79662
rect 37156 79648 37238 79662
rect 38114 79648 38196 79662
rect 38404 79648 38486 79662
rect 39362 79648 39444 79662
rect 39652 79648 39734 79662
rect 40610 79648 40692 79662
rect 40900 79648 40982 79662
rect 41858 79648 41940 79662
rect 42148 79648 42230 79662
rect 43106 79648 43188 79662
rect 43396 79648 43478 79662
rect 44354 79648 44436 79662
rect 44644 79648 44726 79662
rect 45602 79648 45684 79662
rect 45892 79648 45974 79662
rect 46850 79648 46932 79662
rect 47140 79648 47222 79662
rect 48098 79648 48180 79662
rect 48388 79648 48470 79662
rect 49346 79648 49428 79662
rect 49636 79648 49718 79662
rect 50594 79648 50676 79662
rect 50884 79648 50966 79662
rect 51842 79648 51924 79662
rect 52132 79648 52214 79662
rect 53090 79648 53172 79662
rect 53380 79648 53462 79662
rect 54338 79648 54420 79662
rect 54628 79648 54710 79662
rect 55586 79648 55668 79662
rect 55876 79648 55958 79662
rect 56834 79648 56916 79662
rect 57124 79648 57206 79662
rect 58082 79648 58164 79662
rect 58372 79648 58454 79662
rect 16418 79600 16864 79614
rect 17014 79600 17154 79614
rect 17304 79600 18112 79614
rect 18262 79600 18402 79614
rect 18552 79600 19360 79614
rect 19510 79600 19650 79614
rect 19800 79600 20608 79614
rect 20758 79600 20898 79614
rect 21048 79600 21856 79614
rect 22006 79600 22146 79614
rect 22296 79600 23104 79614
rect 23254 79600 23394 79614
rect 23544 79600 24352 79614
rect 24502 79600 24642 79614
rect 24792 79600 25600 79614
rect 25750 79600 25890 79614
rect 26040 79600 26848 79614
rect 26998 79600 27138 79614
rect 27288 79600 28096 79614
rect 28246 79600 28386 79614
rect 28536 79600 29344 79614
rect 29494 79600 29634 79614
rect 29784 79600 30592 79614
rect 30742 79600 30882 79614
rect 31032 79600 31840 79614
rect 31990 79600 32130 79614
rect 32280 79600 33088 79614
rect 33238 79600 33378 79614
rect 33528 79600 34336 79614
rect 34486 79600 34626 79614
rect 34776 79600 35584 79614
rect 35734 79600 35874 79614
rect 36024 79600 36832 79614
rect 36982 79600 37122 79614
rect 37272 79600 38080 79614
rect 38230 79600 38370 79614
rect 38520 79600 39328 79614
rect 39478 79600 39618 79614
rect 39768 79600 40576 79614
rect 40726 79600 40866 79614
rect 41016 79600 41824 79614
rect 41974 79600 42114 79614
rect 42264 79600 43072 79614
rect 43222 79600 43362 79614
rect 43512 79600 44320 79614
rect 44470 79600 44610 79614
rect 44760 79600 45568 79614
rect 45718 79600 45858 79614
rect 46008 79600 46816 79614
rect 46966 79600 47106 79614
rect 47256 79600 48064 79614
rect 48214 79600 48354 79614
rect 48504 79600 49312 79614
rect 49462 79600 49602 79614
rect 49752 79600 50560 79614
rect 50710 79600 50850 79614
rect 51000 79600 51808 79614
rect 51958 79600 52098 79614
rect 52248 79600 53056 79614
rect 53206 79600 53346 79614
rect 53496 79600 54304 79614
rect 54454 79600 54594 79614
rect 54744 79600 55552 79614
rect 55702 79600 55842 79614
rect 55992 79600 56800 79614
rect 56950 79600 57090 79614
rect 57240 79600 58048 79614
rect 58198 79600 58338 79614
rect 58488 79600 58934 79614
rect 16418 79552 58934 79600
rect 16418 79538 16864 79552
rect 17014 79538 17154 79552
rect 17304 79538 18112 79552
rect 18262 79538 18402 79552
rect 18552 79538 19360 79552
rect 19510 79538 19650 79552
rect 19800 79538 20608 79552
rect 20758 79538 20898 79552
rect 21048 79538 21856 79552
rect 22006 79538 22146 79552
rect 22296 79538 23104 79552
rect 23254 79538 23394 79552
rect 23544 79538 24352 79552
rect 24502 79538 24642 79552
rect 24792 79538 25600 79552
rect 25750 79538 25890 79552
rect 26040 79538 26848 79552
rect 26998 79538 27138 79552
rect 27288 79538 28096 79552
rect 28246 79538 28386 79552
rect 28536 79538 29344 79552
rect 29494 79538 29634 79552
rect 29784 79538 30592 79552
rect 30742 79538 30882 79552
rect 31032 79538 31840 79552
rect 31990 79538 32130 79552
rect 32280 79538 33088 79552
rect 33238 79538 33378 79552
rect 33528 79538 34336 79552
rect 34486 79538 34626 79552
rect 34776 79538 35584 79552
rect 35734 79538 35874 79552
rect 36024 79538 36832 79552
rect 36982 79538 37122 79552
rect 37272 79538 38080 79552
rect 38230 79538 38370 79552
rect 38520 79538 39328 79552
rect 39478 79538 39618 79552
rect 39768 79538 40576 79552
rect 40726 79538 40866 79552
rect 41016 79538 41824 79552
rect 41974 79538 42114 79552
rect 42264 79538 43072 79552
rect 43222 79538 43362 79552
rect 43512 79538 44320 79552
rect 44470 79538 44610 79552
rect 44760 79538 45568 79552
rect 45718 79538 45858 79552
rect 46008 79538 46816 79552
rect 46966 79538 47106 79552
rect 47256 79538 48064 79552
rect 48214 79538 48354 79552
rect 48504 79538 49312 79552
rect 49462 79538 49602 79552
rect 49752 79538 50560 79552
rect 50710 79538 50850 79552
rect 51000 79538 51808 79552
rect 51958 79538 52098 79552
rect 52248 79538 53056 79552
rect 53206 79538 53346 79552
rect 53496 79538 54304 79552
rect 54454 79538 54594 79552
rect 54744 79538 55552 79552
rect 55702 79538 55842 79552
rect 55992 79538 56800 79552
rect 56950 79538 57090 79552
rect 57240 79538 58048 79552
rect 58198 79538 58338 79552
rect 58488 79538 58934 79552
rect 16898 79490 16980 79504
rect 17188 79490 17270 79504
rect 18146 79490 18228 79504
rect 18436 79490 18518 79504
rect 19394 79490 19476 79504
rect 19684 79490 19766 79504
rect 20642 79490 20724 79504
rect 20932 79490 21014 79504
rect 21890 79490 21972 79504
rect 22180 79490 22262 79504
rect 23138 79490 23220 79504
rect 23428 79490 23510 79504
rect 24386 79490 24468 79504
rect 24676 79490 24758 79504
rect 25634 79490 25716 79504
rect 25924 79490 26006 79504
rect 26882 79490 26964 79504
rect 27172 79490 27254 79504
rect 28130 79490 28212 79504
rect 28420 79490 28502 79504
rect 29378 79490 29460 79504
rect 29668 79490 29750 79504
rect 30626 79490 30708 79504
rect 30916 79490 30998 79504
rect 31874 79490 31956 79504
rect 32164 79490 32246 79504
rect 33122 79490 33204 79504
rect 33412 79490 33494 79504
rect 34370 79490 34452 79504
rect 34660 79490 34742 79504
rect 35618 79490 35700 79504
rect 35908 79490 35990 79504
rect 36866 79490 36948 79504
rect 37156 79490 37238 79504
rect 38114 79490 38196 79504
rect 38404 79490 38486 79504
rect 39362 79490 39444 79504
rect 39652 79490 39734 79504
rect 40610 79490 40692 79504
rect 40900 79490 40982 79504
rect 41858 79490 41940 79504
rect 42148 79490 42230 79504
rect 43106 79490 43188 79504
rect 43396 79490 43478 79504
rect 44354 79490 44436 79504
rect 44644 79490 44726 79504
rect 45602 79490 45684 79504
rect 45892 79490 45974 79504
rect 46850 79490 46932 79504
rect 47140 79490 47222 79504
rect 48098 79490 48180 79504
rect 48388 79490 48470 79504
rect 49346 79490 49428 79504
rect 49636 79490 49718 79504
rect 50594 79490 50676 79504
rect 50884 79490 50966 79504
rect 51842 79490 51924 79504
rect 52132 79490 52214 79504
rect 53090 79490 53172 79504
rect 53380 79490 53462 79504
rect 54338 79490 54420 79504
rect 54628 79490 54710 79504
rect 55586 79490 55668 79504
rect 55876 79490 55958 79504
rect 56834 79490 56916 79504
rect 57124 79490 57206 79504
rect 58082 79490 58164 79504
rect 58372 79490 58454 79504
rect 16418 79442 58934 79490
rect 16418 79346 58934 79394
rect 16898 79332 16980 79346
rect 17188 79332 17270 79346
rect 18146 79332 18228 79346
rect 18436 79332 18518 79346
rect 19394 79332 19476 79346
rect 19684 79332 19766 79346
rect 20642 79332 20724 79346
rect 20932 79332 21014 79346
rect 21890 79332 21972 79346
rect 22180 79332 22262 79346
rect 23138 79332 23220 79346
rect 23428 79332 23510 79346
rect 24386 79332 24468 79346
rect 24676 79332 24758 79346
rect 25634 79332 25716 79346
rect 25924 79332 26006 79346
rect 26882 79332 26964 79346
rect 27172 79332 27254 79346
rect 28130 79332 28212 79346
rect 28420 79332 28502 79346
rect 29378 79332 29460 79346
rect 29668 79332 29750 79346
rect 30626 79332 30708 79346
rect 30916 79332 30998 79346
rect 31874 79332 31956 79346
rect 32164 79332 32246 79346
rect 33122 79332 33204 79346
rect 33412 79332 33494 79346
rect 34370 79332 34452 79346
rect 34660 79332 34742 79346
rect 35618 79332 35700 79346
rect 35908 79332 35990 79346
rect 36866 79332 36948 79346
rect 37156 79332 37238 79346
rect 38114 79332 38196 79346
rect 38404 79332 38486 79346
rect 39362 79332 39444 79346
rect 39652 79332 39734 79346
rect 40610 79332 40692 79346
rect 40900 79332 40982 79346
rect 41858 79332 41940 79346
rect 42148 79332 42230 79346
rect 43106 79332 43188 79346
rect 43396 79332 43478 79346
rect 44354 79332 44436 79346
rect 44644 79332 44726 79346
rect 45602 79332 45684 79346
rect 45892 79332 45974 79346
rect 46850 79332 46932 79346
rect 47140 79332 47222 79346
rect 48098 79332 48180 79346
rect 48388 79332 48470 79346
rect 49346 79332 49428 79346
rect 49636 79332 49718 79346
rect 50594 79332 50676 79346
rect 50884 79332 50966 79346
rect 51842 79332 51924 79346
rect 52132 79332 52214 79346
rect 53090 79332 53172 79346
rect 53380 79332 53462 79346
rect 54338 79332 54420 79346
rect 54628 79332 54710 79346
rect 55586 79332 55668 79346
rect 55876 79332 55958 79346
rect 56834 79332 56916 79346
rect 57124 79332 57206 79346
rect 58082 79332 58164 79346
rect 58372 79332 58454 79346
rect 16418 79284 16864 79298
rect 17014 79284 17154 79298
rect 17304 79284 18112 79298
rect 18262 79284 18402 79298
rect 18552 79284 19360 79298
rect 19510 79284 19650 79298
rect 19800 79284 20608 79298
rect 20758 79284 20898 79298
rect 21048 79284 21856 79298
rect 22006 79284 22146 79298
rect 22296 79284 23104 79298
rect 23254 79284 23394 79298
rect 23544 79284 24352 79298
rect 24502 79284 24642 79298
rect 24792 79284 25600 79298
rect 25750 79284 25890 79298
rect 26040 79284 26848 79298
rect 26998 79284 27138 79298
rect 27288 79284 28096 79298
rect 28246 79284 28386 79298
rect 28536 79284 29344 79298
rect 29494 79284 29634 79298
rect 29784 79284 30592 79298
rect 30742 79284 30882 79298
rect 31032 79284 31840 79298
rect 31990 79284 32130 79298
rect 32280 79284 33088 79298
rect 33238 79284 33378 79298
rect 33528 79284 34336 79298
rect 34486 79284 34626 79298
rect 34776 79284 35584 79298
rect 35734 79284 35874 79298
rect 36024 79284 36832 79298
rect 36982 79284 37122 79298
rect 37272 79284 38080 79298
rect 38230 79284 38370 79298
rect 38520 79284 39328 79298
rect 39478 79284 39618 79298
rect 39768 79284 40576 79298
rect 40726 79284 40866 79298
rect 41016 79284 41824 79298
rect 41974 79284 42114 79298
rect 42264 79284 43072 79298
rect 43222 79284 43362 79298
rect 43512 79284 44320 79298
rect 44470 79284 44610 79298
rect 44760 79284 45568 79298
rect 45718 79284 45858 79298
rect 46008 79284 46816 79298
rect 46966 79284 47106 79298
rect 47256 79284 48064 79298
rect 48214 79284 48354 79298
rect 48504 79284 49312 79298
rect 49462 79284 49602 79298
rect 49752 79284 50560 79298
rect 50710 79284 50850 79298
rect 51000 79284 51808 79298
rect 51958 79284 52098 79298
rect 52248 79284 53056 79298
rect 53206 79284 53346 79298
rect 53496 79284 54304 79298
rect 54454 79284 54594 79298
rect 54744 79284 55552 79298
rect 55702 79284 55842 79298
rect 55992 79284 56800 79298
rect 56950 79284 57090 79298
rect 57240 79284 58048 79298
rect 58198 79284 58338 79298
rect 58488 79284 58934 79298
rect 16418 79236 58934 79284
rect 16418 79222 16864 79236
rect 17014 79222 17154 79236
rect 17304 79222 18112 79236
rect 18262 79222 18402 79236
rect 18552 79222 19360 79236
rect 19510 79222 19650 79236
rect 19800 79222 20608 79236
rect 20758 79222 20898 79236
rect 21048 79222 21856 79236
rect 22006 79222 22146 79236
rect 22296 79222 23104 79236
rect 23254 79222 23394 79236
rect 23544 79222 24352 79236
rect 24502 79222 24642 79236
rect 24792 79222 25600 79236
rect 25750 79222 25890 79236
rect 26040 79222 26848 79236
rect 26998 79222 27138 79236
rect 27288 79222 28096 79236
rect 28246 79222 28386 79236
rect 28536 79222 29344 79236
rect 29494 79222 29634 79236
rect 29784 79222 30592 79236
rect 30742 79222 30882 79236
rect 31032 79222 31840 79236
rect 31990 79222 32130 79236
rect 32280 79222 33088 79236
rect 33238 79222 33378 79236
rect 33528 79222 34336 79236
rect 34486 79222 34626 79236
rect 34776 79222 35584 79236
rect 35734 79222 35874 79236
rect 36024 79222 36832 79236
rect 36982 79222 37122 79236
rect 37272 79222 38080 79236
rect 38230 79222 38370 79236
rect 38520 79222 39328 79236
rect 39478 79222 39618 79236
rect 39768 79222 40576 79236
rect 40726 79222 40866 79236
rect 41016 79222 41824 79236
rect 41974 79222 42114 79236
rect 42264 79222 43072 79236
rect 43222 79222 43362 79236
rect 43512 79222 44320 79236
rect 44470 79222 44610 79236
rect 44760 79222 45568 79236
rect 45718 79222 45858 79236
rect 46008 79222 46816 79236
rect 46966 79222 47106 79236
rect 47256 79222 48064 79236
rect 48214 79222 48354 79236
rect 48504 79222 49312 79236
rect 49462 79222 49602 79236
rect 49752 79222 50560 79236
rect 50710 79222 50850 79236
rect 51000 79222 51808 79236
rect 51958 79222 52098 79236
rect 52248 79222 53056 79236
rect 53206 79222 53346 79236
rect 53496 79222 54304 79236
rect 54454 79222 54594 79236
rect 54744 79222 55552 79236
rect 55702 79222 55842 79236
rect 55992 79222 56800 79236
rect 56950 79222 57090 79236
rect 57240 79222 58048 79236
rect 58198 79222 58338 79236
rect 58488 79222 58934 79236
rect 16898 79174 16980 79188
rect 17188 79174 17270 79188
rect 18146 79174 18228 79188
rect 18436 79174 18518 79188
rect 19394 79174 19476 79188
rect 19684 79174 19766 79188
rect 20642 79174 20724 79188
rect 20932 79174 21014 79188
rect 21890 79174 21972 79188
rect 22180 79174 22262 79188
rect 23138 79174 23220 79188
rect 23428 79174 23510 79188
rect 24386 79174 24468 79188
rect 24676 79174 24758 79188
rect 25634 79174 25716 79188
rect 25924 79174 26006 79188
rect 26882 79174 26964 79188
rect 27172 79174 27254 79188
rect 28130 79174 28212 79188
rect 28420 79174 28502 79188
rect 29378 79174 29460 79188
rect 29668 79174 29750 79188
rect 30626 79174 30708 79188
rect 30916 79174 30998 79188
rect 31874 79174 31956 79188
rect 32164 79174 32246 79188
rect 33122 79174 33204 79188
rect 33412 79174 33494 79188
rect 34370 79174 34452 79188
rect 34660 79174 34742 79188
rect 35618 79174 35700 79188
rect 35908 79174 35990 79188
rect 36866 79174 36948 79188
rect 37156 79174 37238 79188
rect 38114 79174 38196 79188
rect 38404 79174 38486 79188
rect 39362 79174 39444 79188
rect 39652 79174 39734 79188
rect 40610 79174 40692 79188
rect 40900 79174 40982 79188
rect 41858 79174 41940 79188
rect 42148 79174 42230 79188
rect 43106 79174 43188 79188
rect 43396 79174 43478 79188
rect 44354 79174 44436 79188
rect 44644 79174 44726 79188
rect 45602 79174 45684 79188
rect 45892 79174 45974 79188
rect 46850 79174 46932 79188
rect 47140 79174 47222 79188
rect 48098 79174 48180 79188
rect 48388 79174 48470 79188
rect 49346 79174 49428 79188
rect 49636 79174 49718 79188
rect 50594 79174 50676 79188
rect 50884 79174 50966 79188
rect 51842 79174 51924 79188
rect 52132 79174 52214 79188
rect 53090 79174 53172 79188
rect 53380 79174 53462 79188
rect 54338 79174 54420 79188
rect 54628 79174 54710 79188
rect 55586 79174 55668 79188
rect 55876 79174 55958 79188
rect 56834 79174 56916 79188
rect 57124 79174 57206 79188
rect 58082 79174 58164 79188
rect 58372 79174 58454 79188
rect 16418 79126 58934 79174
rect 16418 78968 58934 79078
rect 16418 78872 58934 78920
rect 16898 78858 16980 78872
rect 17188 78858 17270 78872
rect 18146 78858 18228 78872
rect 18436 78858 18518 78872
rect 19394 78858 19476 78872
rect 19684 78858 19766 78872
rect 20642 78858 20724 78872
rect 20932 78858 21014 78872
rect 21890 78858 21972 78872
rect 22180 78858 22262 78872
rect 23138 78858 23220 78872
rect 23428 78858 23510 78872
rect 24386 78858 24468 78872
rect 24676 78858 24758 78872
rect 25634 78858 25716 78872
rect 25924 78858 26006 78872
rect 26882 78858 26964 78872
rect 27172 78858 27254 78872
rect 28130 78858 28212 78872
rect 28420 78858 28502 78872
rect 29378 78858 29460 78872
rect 29668 78858 29750 78872
rect 30626 78858 30708 78872
rect 30916 78858 30998 78872
rect 31874 78858 31956 78872
rect 32164 78858 32246 78872
rect 33122 78858 33204 78872
rect 33412 78858 33494 78872
rect 34370 78858 34452 78872
rect 34660 78858 34742 78872
rect 35618 78858 35700 78872
rect 35908 78858 35990 78872
rect 36866 78858 36948 78872
rect 37156 78858 37238 78872
rect 38114 78858 38196 78872
rect 38404 78858 38486 78872
rect 39362 78858 39444 78872
rect 39652 78858 39734 78872
rect 40610 78858 40692 78872
rect 40900 78858 40982 78872
rect 41858 78858 41940 78872
rect 42148 78858 42230 78872
rect 43106 78858 43188 78872
rect 43396 78858 43478 78872
rect 44354 78858 44436 78872
rect 44644 78858 44726 78872
rect 45602 78858 45684 78872
rect 45892 78858 45974 78872
rect 46850 78858 46932 78872
rect 47140 78858 47222 78872
rect 48098 78858 48180 78872
rect 48388 78858 48470 78872
rect 49346 78858 49428 78872
rect 49636 78858 49718 78872
rect 50594 78858 50676 78872
rect 50884 78858 50966 78872
rect 51842 78858 51924 78872
rect 52132 78858 52214 78872
rect 53090 78858 53172 78872
rect 53380 78858 53462 78872
rect 54338 78858 54420 78872
rect 54628 78858 54710 78872
rect 55586 78858 55668 78872
rect 55876 78858 55958 78872
rect 56834 78858 56916 78872
rect 57124 78858 57206 78872
rect 58082 78858 58164 78872
rect 58372 78858 58454 78872
rect 16418 78810 16864 78824
rect 17014 78810 17154 78824
rect 17304 78810 18112 78824
rect 18262 78810 18402 78824
rect 18552 78810 19360 78824
rect 19510 78810 19650 78824
rect 19800 78810 20608 78824
rect 20758 78810 20898 78824
rect 21048 78810 21856 78824
rect 22006 78810 22146 78824
rect 22296 78810 23104 78824
rect 23254 78810 23394 78824
rect 23544 78810 24352 78824
rect 24502 78810 24642 78824
rect 24792 78810 25600 78824
rect 25750 78810 25890 78824
rect 26040 78810 26848 78824
rect 26998 78810 27138 78824
rect 27288 78810 28096 78824
rect 28246 78810 28386 78824
rect 28536 78810 29344 78824
rect 29494 78810 29634 78824
rect 29784 78810 30592 78824
rect 30742 78810 30882 78824
rect 31032 78810 31840 78824
rect 31990 78810 32130 78824
rect 32280 78810 33088 78824
rect 33238 78810 33378 78824
rect 33528 78810 34336 78824
rect 34486 78810 34626 78824
rect 34776 78810 35584 78824
rect 35734 78810 35874 78824
rect 36024 78810 36832 78824
rect 36982 78810 37122 78824
rect 37272 78810 38080 78824
rect 38230 78810 38370 78824
rect 38520 78810 39328 78824
rect 39478 78810 39618 78824
rect 39768 78810 40576 78824
rect 40726 78810 40866 78824
rect 41016 78810 41824 78824
rect 41974 78810 42114 78824
rect 42264 78810 43072 78824
rect 43222 78810 43362 78824
rect 43512 78810 44320 78824
rect 44470 78810 44610 78824
rect 44760 78810 45568 78824
rect 45718 78810 45858 78824
rect 46008 78810 46816 78824
rect 46966 78810 47106 78824
rect 47256 78810 48064 78824
rect 48214 78810 48354 78824
rect 48504 78810 49312 78824
rect 49462 78810 49602 78824
rect 49752 78810 50560 78824
rect 50710 78810 50850 78824
rect 51000 78810 51808 78824
rect 51958 78810 52098 78824
rect 52248 78810 53056 78824
rect 53206 78810 53346 78824
rect 53496 78810 54304 78824
rect 54454 78810 54594 78824
rect 54744 78810 55552 78824
rect 55702 78810 55842 78824
rect 55992 78810 56800 78824
rect 56950 78810 57090 78824
rect 57240 78810 58048 78824
rect 58198 78810 58338 78824
rect 58488 78810 58934 78824
rect 16418 78762 58934 78810
rect 16418 78748 16864 78762
rect 17014 78748 17154 78762
rect 17304 78748 18112 78762
rect 18262 78748 18402 78762
rect 18552 78748 19360 78762
rect 19510 78748 19650 78762
rect 19800 78748 20608 78762
rect 20758 78748 20898 78762
rect 21048 78748 21856 78762
rect 22006 78748 22146 78762
rect 22296 78748 23104 78762
rect 23254 78748 23394 78762
rect 23544 78748 24352 78762
rect 24502 78748 24642 78762
rect 24792 78748 25600 78762
rect 25750 78748 25890 78762
rect 26040 78748 26848 78762
rect 26998 78748 27138 78762
rect 27288 78748 28096 78762
rect 28246 78748 28386 78762
rect 28536 78748 29344 78762
rect 29494 78748 29634 78762
rect 29784 78748 30592 78762
rect 30742 78748 30882 78762
rect 31032 78748 31840 78762
rect 31990 78748 32130 78762
rect 32280 78748 33088 78762
rect 33238 78748 33378 78762
rect 33528 78748 34336 78762
rect 34486 78748 34626 78762
rect 34776 78748 35584 78762
rect 35734 78748 35874 78762
rect 36024 78748 36832 78762
rect 36982 78748 37122 78762
rect 37272 78748 38080 78762
rect 38230 78748 38370 78762
rect 38520 78748 39328 78762
rect 39478 78748 39618 78762
rect 39768 78748 40576 78762
rect 40726 78748 40866 78762
rect 41016 78748 41824 78762
rect 41974 78748 42114 78762
rect 42264 78748 43072 78762
rect 43222 78748 43362 78762
rect 43512 78748 44320 78762
rect 44470 78748 44610 78762
rect 44760 78748 45568 78762
rect 45718 78748 45858 78762
rect 46008 78748 46816 78762
rect 46966 78748 47106 78762
rect 47256 78748 48064 78762
rect 48214 78748 48354 78762
rect 48504 78748 49312 78762
rect 49462 78748 49602 78762
rect 49752 78748 50560 78762
rect 50710 78748 50850 78762
rect 51000 78748 51808 78762
rect 51958 78748 52098 78762
rect 52248 78748 53056 78762
rect 53206 78748 53346 78762
rect 53496 78748 54304 78762
rect 54454 78748 54594 78762
rect 54744 78748 55552 78762
rect 55702 78748 55842 78762
rect 55992 78748 56800 78762
rect 56950 78748 57090 78762
rect 57240 78748 58048 78762
rect 58198 78748 58338 78762
rect 58488 78748 58934 78762
rect 16898 78700 16980 78714
rect 17188 78700 17270 78714
rect 18146 78700 18228 78714
rect 18436 78700 18518 78714
rect 19394 78700 19476 78714
rect 19684 78700 19766 78714
rect 20642 78700 20724 78714
rect 20932 78700 21014 78714
rect 21890 78700 21972 78714
rect 22180 78700 22262 78714
rect 23138 78700 23220 78714
rect 23428 78700 23510 78714
rect 24386 78700 24468 78714
rect 24676 78700 24758 78714
rect 25634 78700 25716 78714
rect 25924 78700 26006 78714
rect 26882 78700 26964 78714
rect 27172 78700 27254 78714
rect 28130 78700 28212 78714
rect 28420 78700 28502 78714
rect 29378 78700 29460 78714
rect 29668 78700 29750 78714
rect 30626 78700 30708 78714
rect 30916 78700 30998 78714
rect 31874 78700 31956 78714
rect 32164 78700 32246 78714
rect 33122 78700 33204 78714
rect 33412 78700 33494 78714
rect 34370 78700 34452 78714
rect 34660 78700 34742 78714
rect 35618 78700 35700 78714
rect 35908 78700 35990 78714
rect 36866 78700 36948 78714
rect 37156 78700 37238 78714
rect 38114 78700 38196 78714
rect 38404 78700 38486 78714
rect 39362 78700 39444 78714
rect 39652 78700 39734 78714
rect 40610 78700 40692 78714
rect 40900 78700 40982 78714
rect 41858 78700 41940 78714
rect 42148 78700 42230 78714
rect 43106 78700 43188 78714
rect 43396 78700 43478 78714
rect 44354 78700 44436 78714
rect 44644 78700 44726 78714
rect 45602 78700 45684 78714
rect 45892 78700 45974 78714
rect 46850 78700 46932 78714
rect 47140 78700 47222 78714
rect 48098 78700 48180 78714
rect 48388 78700 48470 78714
rect 49346 78700 49428 78714
rect 49636 78700 49718 78714
rect 50594 78700 50676 78714
rect 50884 78700 50966 78714
rect 51842 78700 51924 78714
rect 52132 78700 52214 78714
rect 53090 78700 53172 78714
rect 53380 78700 53462 78714
rect 54338 78700 54420 78714
rect 54628 78700 54710 78714
rect 55586 78700 55668 78714
rect 55876 78700 55958 78714
rect 56834 78700 56916 78714
rect 57124 78700 57206 78714
rect 58082 78700 58164 78714
rect 58372 78700 58454 78714
rect 16418 78652 58934 78700
rect 16418 78556 58934 78604
rect 16898 78542 16980 78556
rect 17188 78542 17270 78556
rect 18146 78542 18228 78556
rect 18436 78542 18518 78556
rect 19394 78542 19476 78556
rect 19684 78542 19766 78556
rect 20642 78542 20724 78556
rect 20932 78542 21014 78556
rect 21890 78542 21972 78556
rect 22180 78542 22262 78556
rect 23138 78542 23220 78556
rect 23428 78542 23510 78556
rect 24386 78542 24468 78556
rect 24676 78542 24758 78556
rect 25634 78542 25716 78556
rect 25924 78542 26006 78556
rect 26882 78542 26964 78556
rect 27172 78542 27254 78556
rect 28130 78542 28212 78556
rect 28420 78542 28502 78556
rect 29378 78542 29460 78556
rect 29668 78542 29750 78556
rect 30626 78542 30708 78556
rect 30916 78542 30998 78556
rect 31874 78542 31956 78556
rect 32164 78542 32246 78556
rect 33122 78542 33204 78556
rect 33412 78542 33494 78556
rect 34370 78542 34452 78556
rect 34660 78542 34742 78556
rect 35618 78542 35700 78556
rect 35908 78542 35990 78556
rect 36866 78542 36948 78556
rect 37156 78542 37238 78556
rect 38114 78542 38196 78556
rect 38404 78542 38486 78556
rect 39362 78542 39444 78556
rect 39652 78542 39734 78556
rect 40610 78542 40692 78556
rect 40900 78542 40982 78556
rect 41858 78542 41940 78556
rect 42148 78542 42230 78556
rect 43106 78542 43188 78556
rect 43396 78542 43478 78556
rect 44354 78542 44436 78556
rect 44644 78542 44726 78556
rect 45602 78542 45684 78556
rect 45892 78542 45974 78556
rect 46850 78542 46932 78556
rect 47140 78542 47222 78556
rect 48098 78542 48180 78556
rect 48388 78542 48470 78556
rect 49346 78542 49428 78556
rect 49636 78542 49718 78556
rect 50594 78542 50676 78556
rect 50884 78542 50966 78556
rect 51842 78542 51924 78556
rect 52132 78542 52214 78556
rect 53090 78542 53172 78556
rect 53380 78542 53462 78556
rect 54338 78542 54420 78556
rect 54628 78542 54710 78556
rect 55586 78542 55668 78556
rect 55876 78542 55958 78556
rect 56834 78542 56916 78556
rect 57124 78542 57206 78556
rect 58082 78542 58164 78556
rect 58372 78542 58454 78556
rect 16418 78494 16864 78508
rect 17014 78494 17154 78508
rect 17304 78494 18112 78508
rect 18262 78494 18402 78508
rect 18552 78494 19360 78508
rect 19510 78494 19650 78508
rect 19800 78494 20608 78508
rect 20758 78494 20898 78508
rect 21048 78494 21856 78508
rect 22006 78494 22146 78508
rect 22296 78494 23104 78508
rect 23254 78494 23394 78508
rect 23544 78494 24352 78508
rect 24502 78494 24642 78508
rect 24792 78494 25600 78508
rect 25750 78494 25890 78508
rect 26040 78494 26848 78508
rect 26998 78494 27138 78508
rect 27288 78494 28096 78508
rect 28246 78494 28386 78508
rect 28536 78494 29344 78508
rect 29494 78494 29634 78508
rect 29784 78494 30592 78508
rect 30742 78494 30882 78508
rect 31032 78494 31840 78508
rect 31990 78494 32130 78508
rect 32280 78494 33088 78508
rect 33238 78494 33378 78508
rect 33528 78494 34336 78508
rect 34486 78494 34626 78508
rect 34776 78494 35584 78508
rect 35734 78494 35874 78508
rect 36024 78494 36832 78508
rect 36982 78494 37122 78508
rect 37272 78494 38080 78508
rect 38230 78494 38370 78508
rect 38520 78494 39328 78508
rect 39478 78494 39618 78508
rect 39768 78494 40576 78508
rect 40726 78494 40866 78508
rect 41016 78494 41824 78508
rect 41974 78494 42114 78508
rect 42264 78494 43072 78508
rect 43222 78494 43362 78508
rect 43512 78494 44320 78508
rect 44470 78494 44610 78508
rect 44760 78494 45568 78508
rect 45718 78494 45858 78508
rect 46008 78494 46816 78508
rect 46966 78494 47106 78508
rect 47256 78494 48064 78508
rect 48214 78494 48354 78508
rect 48504 78494 49312 78508
rect 49462 78494 49602 78508
rect 49752 78494 50560 78508
rect 50710 78494 50850 78508
rect 51000 78494 51808 78508
rect 51958 78494 52098 78508
rect 52248 78494 53056 78508
rect 53206 78494 53346 78508
rect 53496 78494 54304 78508
rect 54454 78494 54594 78508
rect 54744 78494 55552 78508
rect 55702 78494 55842 78508
rect 55992 78494 56800 78508
rect 56950 78494 57090 78508
rect 57240 78494 58048 78508
rect 58198 78494 58338 78508
rect 58488 78494 58934 78508
rect 16418 78446 58934 78494
rect 16418 78432 16864 78446
rect 17014 78432 17154 78446
rect 17304 78432 18112 78446
rect 18262 78432 18402 78446
rect 18552 78432 19360 78446
rect 19510 78432 19650 78446
rect 19800 78432 20608 78446
rect 20758 78432 20898 78446
rect 21048 78432 21856 78446
rect 22006 78432 22146 78446
rect 22296 78432 23104 78446
rect 23254 78432 23394 78446
rect 23544 78432 24352 78446
rect 24502 78432 24642 78446
rect 24792 78432 25600 78446
rect 25750 78432 25890 78446
rect 26040 78432 26848 78446
rect 26998 78432 27138 78446
rect 27288 78432 28096 78446
rect 28246 78432 28386 78446
rect 28536 78432 29344 78446
rect 29494 78432 29634 78446
rect 29784 78432 30592 78446
rect 30742 78432 30882 78446
rect 31032 78432 31840 78446
rect 31990 78432 32130 78446
rect 32280 78432 33088 78446
rect 33238 78432 33378 78446
rect 33528 78432 34336 78446
rect 34486 78432 34626 78446
rect 34776 78432 35584 78446
rect 35734 78432 35874 78446
rect 36024 78432 36832 78446
rect 36982 78432 37122 78446
rect 37272 78432 38080 78446
rect 38230 78432 38370 78446
rect 38520 78432 39328 78446
rect 39478 78432 39618 78446
rect 39768 78432 40576 78446
rect 40726 78432 40866 78446
rect 41016 78432 41824 78446
rect 41974 78432 42114 78446
rect 42264 78432 43072 78446
rect 43222 78432 43362 78446
rect 43512 78432 44320 78446
rect 44470 78432 44610 78446
rect 44760 78432 45568 78446
rect 45718 78432 45858 78446
rect 46008 78432 46816 78446
rect 46966 78432 47106 78446
rect 47256 78432 48064 78446
rect 48214 78432 48354 78446
rect 48504 78432 49312 78446
rect 49462 78432 49602 78446
rect 49752 78432 50560 78446
rect 50710 78432 50850 78446
rect 51000 78432 51808 78446
rect 51958 78432 52098 78446
rect 52248 78432 53056 78446
rect 53206 78432 53346 78446
rect 53496 78432 54304 78446
rect 54454 78432 54594 78446
rect 54744 78432 55552 78446
rect 55702 78432 55842 78446
rect 55992 78432 56800 78446
rect 56950 78432 57090 78446
rect 57240 78432 58048 78446
rect 58198 78432 58338 78446
rect 58488 78432 58934 78446
rect 16898 78384 16980 78398
rect 17188 78384 17270 78398
rect 18146 78384 18228 78398
rect 18436 78384 18518 78398
rect 19394 78384 19476 78398
rect 19684 78384 19766 78398
rect 20642 78384 20724 78398
rect 20932 78384 21014 78398
rect 21890 78384 21972 78398
rect 22180 78384 22262 78398
rect 23138 78384 23220 78398
rect 23428 78384 23510 78398
rect 24386 78384 24468 78398
rect 24676 78384 24758 78398
rect 25634 78384 25716 78398
rect 25924 78384 26006 78398
rect 26882 78384 26964 78398
rect 27172 78384 27254 78398
rect 28130 78384 28212 78398
rect 28420 78384 28502 78398
rect 29378 78384 29460 78398
rect 29668 78384 29750 78398
rect 30626 78384 30708 78398
rect 30916 78384 30998 78398
rect 31874 78384 31956 78398
rect 32164 78384 32246 78398
rect 33122 78384 33204 78398
rect 33412 78384 33494 78398
rect 34370 78384 34452 78398
rect 34660 78384 34742 78398
rect 35618 78384 35700 78398
rect 35908 78384 35990 78398
rect 36866 78384 36948 78398
rect 37156 78384 37238 78398
rect 38114 78384 38196 78398
rect 38404 78384 38486 78398
rect 39362 78384 39444 78398
rect 39652 78384 39734 78398
rect 40610 78384 40692 78398
rect 40900 78384 40982 78398
rect 41858 78384 41940 78398
rect 42148 78384 42230 78398
rect 43106 78384 43188 78398
rect 43396 78384 43478 78398
rect 44354 78384 44436 78398
rect 44644 78384 44726 78398
rect 45602 78384 45684 78398
rect 45892 78384 45974 78398
rect 46850 78384 46932 78398
rect 47140 78384 47222 78398
rect 48098 78384 48180 78398
rect 48388 78384 48470 78398
rect 49346 78384 49428 78398
rect 49636 78384 49718 78398
rect 50594 78384 50676 78398
rect 50884 78384 50966 78398
rect 51842 78384 51924 78398
rect 52132 78384 52214 78398
rect 53090 78384 53172 78398
rect 53380 78384 53462 78398
rect 54338 78384 54420 78398
rect 54628 78384 54710 78398
rect 55586 78384 55668 78398
rect 55876 78384 55958 78398
rect 56834 78384 56916 78398
rect 57124 78384 57206 78398
rect 58082 78384 58164 78398
rect 58372 78384 58454 78398
rect 16418 78336 58934 78384
rect 16418 78178 58934 78288
rect 16418 78082 58934 78130
rect 16898 78068 16980 78082
rect 17188 78068 17270 78082
rect 18146 78068 18228 78082
rect 18436 78068 18518 78082
rect 19394 78068 19476 78082
rect 19684 78068 19766 78082
rect 20642 78068 20724 78082
rect 20932 78068 21014 78082
rect 21890 78068 21972 78082
rect 22180 78068 22262 78082
rect 23138 78068 23220 78082
rect 23428 78068 23510 78082
rect 24386 78068 24468 78082
rect 24676 78068 24758 78082
rect 25634 78068 25716 78082
rect 25924 78068 26006 78082
rect 26882 78068 26964 78082
rect 27172 78068 27254 78082
rect 28130 78068 28212 78082
rect 28420 78068 28502 78082
rect 29378 78068 29460 78082
rect 29668 78068 29750 78082
rect 30626 78068 30708 78082
rect 30916 78068 30998 78082
rect 31874 78068 31956 78082
rect 32164 78068 32246 78082
rect 33122 78068 33204 78082
rect 33412 78068 33494 78082
rect 34370 78068 34452 78082
rect 34660 78068 34742 78082
rect 35618 78068 35700 78082
rect 35908 78068 35990 78082
rect 36866 78068 36948 78082
rect 37156 78068 37238 78082
rect 38114 78068 38196 78082
rect 38404 78068 38486 78082
rect 39362 78068 39444 78082
rect 39652 78068 39734 78082
rect 40610 78068 40692 78082
rect 40900 78068 40982 78082
rect 41858 78068 41940 78082
rect 42148 78068 42230 78082
rect 43106 78068 43188 78082
rect 43396 78068 43478 78082
rect 44354 78068 44436 78082
rect 44644 78068 44726 78082
rect 45602 78068 45684 78082
rect 45892 78068 45974 78082
rect 46850 78068 46932 78082
rect 47140 78068 47222 78082
rect 48098 78068 48180 78082
rect 48388 78068 48470 78082
rect 49346 78068 49428 78082
rect 49636 78068 49718 78082
rect 50594 78068 50676 78082
rect 50884 78068 50966 78082
rect 51842 78068 51924 78082
rect 52132 78068 52214 78082
rect 53090 78068 53172 78082
rect 53380 78068 53462 78082
rect 54338 78068 54420 78082
rect 54628 78068 54710 78082
rect 55586 78068 55668 78082
rect 55876 78068 55958 78082
rect 56834 78068 56916 78082
rect 57124 78068 57206 78082
rect 58082 78068 58164 78082
rect 58372 78068 58454 78082
rect 16418 78020 16864 78034
rect 17014 78020 17154 78034
rect 17304 78020 18112 78034
rect 18262 78020 18402 78034
rect 18552 78020 19360 78034
rect 19510 78020 19650 78034
rect 19800 78020 20608 78034
rect 20758 78020 20898 78034
rect 21048 78020 21856 78034
rect 22006 78020 22146 78034
rect 22296 78020 23104 78034
rect 23254 78020 23394 78034
rect 23544 78020 24352 78034
rect 24502 78020 24642 78034
rect 24792 78020 25600 78034
rect 25750 78020 25890 78034
rect 26040 78020 26848 78034
rect 26998 78020 27138 78034
rect 27288 78020 28096 78034
rect 28246 78020 28386 78034
rect 28536 78020 29344 78034
rect 29494 78020 29634 78034
rect 29784 78020 30592 78034
rect 30742 78020 30882 78034
rect 31032 78020 31840 78034
rect 31990 78020 32130 78034
rect 32280 78020 33088 78034
rect 33238 78020 33378 78034
rect 33528 78020 34336 78034
rect 34486 78020 34626 78034
rect 34776 78020 35584 78034
rect 35734 78020 35874 78034
rect 36024 78020 36832 78034
rect 36982 78020 37122 78034
rect 37272 78020 38080 78034
rect 38230 78020 38370 78034
rect 38520 78020 39328 78034
rect 39478 78020 39618 78034
rect 39768 78020 40576 78034
rect 40726 78020 40866 78034
rect 41016 78020 41824 78034
rect 41974 78020 42114 78034
rect 42264 78020 43072 78034
rect 43222 78020 43362 78034
rect 43512 78020 44320 78034
rect 44470 78020 44610 78034
rect 44760 78020 45568 78034
rect 45718 78020 45858 78034
rect 46008 78020 46816 78034
rect 46966 78020 47106 78034
rect 47256 78020 48064 78034
rect 48214 78020 48354 78034
rect 48504 78020 49312 78034
rect 49462 78020 49602 78034
rect 49752 78020 50560 78034
rect 50710 78020 50850 78034
rect 51000 78020 51808 78034
rect 51958 78020 52098 78034
rect 52248 78020 53056 78034
rect 53206 78020 53346 78034
rect 53496 78020 54304 78034
rect 54454 78020 54594 78034
rect 54744 78020 55552 78034
rect 55702 78020 55842 78034
rect 55992 78020 56800 78034
rect 56950 78020 57090 78034
rect 57240 78020 58048 78034
rect 58198 78020 58338 78034
rect 58488 78020 58934 78034
rect 16418 77972 58934 78020
rect 16418 77958 16864 77972
rect 17014 77958 17154 77972
rect 17304 77958 18112 77972
rect 18262 77958 18402 77972
rect 18552 77958 19360 77972
rect 19510 77958 19650 77972
rect 19800 77958 20608 77972
rect 20758 77958 20898 77972
rect 21048 77958 21856 77972
rect 22006 77958 22146 77972
rect 22296 77958 23104 77972
rect 23254 77958 23394 77972
rect 23544 77958 24352 77972
rect 24502 77958 24642 77972
rect 24792 77958 25600 77972
rect 25750 77958 25890 77972
rect 26040 77958 26848 77972
rect 26998 77958 27138 77972
rect 27288 77958 28096 77972
rect 28246 77958 28386 77972
rect 28536 77958 29344 77972
rect 29494 77958 29634 77972
rect 29784 77958 30592 77972
rect 30742 77958 30882 77972
rect 31032 77958 31840 77972
rect 31990 77958 32130 77972
rect 32280 77958 33088 77972
rect 33238 77958 33378 77972
rect 33528 77958 34336 77972
rect 34486 77958 34626 77972
rect 34776 77958 35584 77972
rect 35734 77958 35874 77972
rect 36024 77958 36832 77972
rect 36982 77958 37122 77972
rect 37272 77958 38080 77972
rect 38230 77958 38370 77972
rect 38520 77958 39328 77972
rect 39478 77958 39618 77972
rect 39768 77958 40576 77972
rect 40726 77958 40866 77972
rect 41016 77958 41824 77972
rect 41974 77958 42114 77972
rect 42264 77958 43072 77972
rect 43222 77958 43362 77972
rect 43512 77958 44320 77972
rect 44470 77958 44610 77972
rect 44760 77958 45568 77972
rect 45718 77958 45858 77972
rect 46008 77958 46816 77972
rect 46966 77958 47106 77972
rect 47256 77958 48064 77972
rect 48214 77958 48354 77972
rect 48504 77958 49312 77972
rect 49462 77958 49602 77972
rect 49752 77958 50560 77972
rect 50710 77958 50850 77972
rect 51000 77958 51808 77972
rect 51958 77958 52098 77972
rect 52248 77958 53056 77972
rect 53206 77958 53346 77972
rect 53496 77958 54304 77972
rect 54454 77958 54594 77972
rect 54744 77958 55552 77972
rect 55702 77958 55842 77972
rect 55992 77958 56800 77972
rect 56950 77958 57090 77972
rect 57240 77958 58048 77972
rect 58198 77958 58338 77972
rect 58488 77958 58934 77972
rect 16898 77910 16980 77924
rect 17188 77910 17270 77924
rect 18146 77910 18228 77924
rect 18436 77910 18518 77924
rect 19394 77910 19476 77924
rect 19684 77910 19766 77924
rect 20642 77910 20724 77924
rect 20932 77910 21014 77924
rect 21890 77910 21972 77924
rect 22180 77910 22262 77924
rect 23138 77910 23220 77924
rect 23428 77910 23510 77924
rect 24386 77910 24468 77924
rect 24676 77910 24758 77924
rect 25634 77910 25716 77924
rect 25924 77910 26006 77924
rect 26882 77910 26964 77924
rect 27172 77910 27254 77924
rect 28130 77910 28212 77924
rect 28420 77910 28502 77924
rect 29378 77910 29460 77924
rect 29668 77910 29750 77924
rect 30626 77910 30708 77924
rect 30916 77910 30998 77924
rect 31874 77910 31956 77924
rect 32164 77910 32246 77924
rect 33122 77910 33204 77924
rect 33412 77910 33494 77924
rect 34370 77910 34452 77924
rect 34660 77910 34742 77924
rect 35618 77910 35700 77924
rect 35908 77910 35990 77924
rect 36866 77910 36948 77924
rect 37156 77910 37238 77924
rect 38114 77910 38196 77924
rect 38404 77910 38486 77924
rect 39362 77910 39444 77924
rect 39652 77910 39734 77924
rect 40610 77910 40692 77924
rect 40900 77910 40982 77924
rect 41858 77910 41940 77924
rect 42148 77910 42230 77924
rect 43106 77910 43188 77924
rect 43396 77910 43478 77924
rect 44354 77910 44436 77924
rect 44644 77910 44726 77924
rect 45602 77910 45684 77924
rect 45892 77910 45974 77924
rect 46850 77910 46932 77924
rect 47140 77910 47222 77924
rect 48098 77910 48180 77924
rect 48388 77910 48470 77924
rect 49346 77910 49428 77924
rect 49636 77910 49718 77924
rect 50594 77910 50676 77924
rect 50884 77910 50966 77924
rect 51842 77910 51924 77924
rect 52132 77910 52214 77924
rect 53090 77910 53172 77924
rect 53380 77910 53462 77924
rect 54338 77910 54420 77924
rect 54628 77910 54710 77924
rect 55586 77910 55668 77924
rect 55876 77910 55958 77924
rect 56834 77910 56916 77924
rect 57124 77910 57206 77924
rect 58082 77910 58164 77924
rect 58372 77910 58454 77924
rect 16418 77862 58934 77910
rect 16418 77766 58934 77814
rect 16898 77752 16980 77766
rect 17188 77752 17270 77766
rect 18146 77752 18228 77766
rect 18436 77752 18518 77766
rect 19394 77752 19476 77766
rect 19684 77752 19766 77766
rect 20642 77752 20724 77766
rect 20932 77752 21014 77766
rect 21890 77752 21972 77766
rect 22180 77752 22262 77766
rect 23138 77752 23220 77766
rect 23428 77752 23510 77766
rect 24386 77752 24468 77766
rect 24676 77752 24758 77766
rect 25634 77752 25716 77766
rect 25924 77752 26006 77766
rect 26882 77752 26964 77766
rect 27172 77752 27254 77766
rect 28130 77752 28212 77766
rect 28420 77752 28502 77766
rect 29378 77752 29460 77766
rect 29668 77752 29750 77766
rect 30626 77752 30708 77766
rect 30916 77752 30998 77766
rect 31874 77752 31956 77766
rect 32164 77752 32246 77766
rect 33122 77752 33204 77766
rect 33412 77752 33494 77766
rect 34370 77752 34452 77766
rect 34660 77752 34742 77766
rect 35618 77752 35700 77766
rect 35908 77752 35990 77766
rect 36866 77752 36948 77766
rect 37156 77752 37238 77766
rect 38114 77752 38196 77766
rect 38404 77752 38486 77766
rect 39362 77752 39444 77766
rect 39652 77752 39734 77766
rect 40610 77752 40692 77766
rect 40900 77752 40982 77766
rect 41858 77752 41940 77766
rect 42148 77752 42230 77766
rect 43106 77752 43188 77766
rect 43396 77752 43478 77766
rect 44354 77752 44436 77766
rect 44644 77752 44726 77766
rect 45602 77752 45684 77766
rect 45892 77752 45974 77766
rect 46850 77752 46932 77766
rect 47140 77752 47222 77766
rect 48098 77752 48180 77766
rect 48388 77752 48470 77766
rect 49346 77752 49428 77766
rect 49636 77752 49718 77766
rect 50594 77752 50676 77766
rect 50884 77752 50966 77766
rect 51842 77752 51924 77766
rect 52132 77752 52214 77766
rect 53090 77752 53172 77766
rect 53380 77752 53462 77766
rect 54338 77752 54420 77766
rect 54628 77752 54710 77766
rect 55586 77752 55668 77766
rect 55876 77752 55958 77766
rect 56834 77752 56916 77766
rect 57124 77752 57206 77766
rect 58082 77752 58164 77766
rect 58372 77752 58454 77766
rect 16418 77704 16864 77718
rect 17014 77704 17154 77718
rect 17304 77704 18112 77718
rect 18262 77704 18402 77718
rect 18552 77704 19360 77718
rect 19510 77704 19650 77718
rect 19800 77704 20608 77718
rect 20758 77704 20898 77718
rect 21048 77704 21856 77718
rect 22006 77704 22146 77718
rect 22296 77704 23104 77718
rect 23254 77704 23394 77718
rect 23544 77704 24352 77718
rect 24502 77704 24642 77718
rect 24792 77704 25600 77718
rect 25750 77704 25890 77718
rect 26040 77704 26848 77718
rect 26998 77704 27138 77718
rect 27288 77704 28096 77718
rect 28246 77704 28386 77718
rect 28536 77704 29344 77718
rect 29494 77704 29634 77718
rect 29784 77704 30592 77718
rect 30742 77704 30882 77718
rect 31032 77704 31840 77718
rect 31990 77704 32130 77718
rect 32280 77704 33088 77718
rect 33238 77704 33378 77718
rect 33528 77704 34336 77718
rect 34486 77704 34626 77718
rect 34776 77704 35584 77718
rect 35734 77704 35874 77718
rect 36024 77704 36832 77718
rect 36982 77704 37122 77718
rect 37272 77704 38080 77718
rect 38230 77704 38370 77718
rect 38520 77704 39328 77718
rect 39478 77704 39618 77718
rect 39768 77704 40576 77718
rect 40726 77704 40866 77718
rect 41016 77704 41824 77718
rect 41974 77704 42114 77718
rect 42264 77704 43072 77718
rect 43222 77704 43362 77718
rect 43512 77704 44320 77718
rect 44470 77704 44610 77718
rect 44760 77704 45568 77718
rect 45718 77704 45858 77718
rect 46008 77704 46816 77718
rect 46966 77704 47106 77718
rect 47256 77704 48064 77718
rect 48214 77704 48354 77718
rect 48504 77704 49312 77718
rect 49462 77704 49602 77718
rect 49752 77704 50560 77718
rect 50710 77704 50850 77718
rect 51000 77704 51808 77718
rect 51958 77704 52098 77718
rect 52248 77704 53056 77718
rect 53206 77704 53346 77718
rect 53496 77704 54304 77718
rect 54454 77704 54594 77718
rect 54744 77704 55552 77718
rect 55702 77704 55842 77718
rect 55992 77704 56800 77718
rect 56950 77704 57090 77718
rect 57240 77704 58048 77718
rect 58198 77704 58338 77718
rect 58488 77704 58934 77718
rect 16418 77656 58934 77704
rect 16418 77642 16864 77656
rect 17014 77642 17154 77656
rect 17304 77642 18112 77656
rect 18262 77642 18402 77656
rect 18552 77642 19360 77656
rect 19510 77642 19650 77656
rect 19800 77642 20608 77656
rect 20758 77642 20898 77656
rect 21048 77642 21856 77656
rect 22006 77642 22146 77656
rect 22296 77642 23104 77656
rect 23254 77642 23394 77656
rect 23544 77642 24352 77656
rect 24502 77642 24642 77656
rect 24792 77642 25600 77656
rect 25750 77642 25890 77656
rect 26040 77642 26848 77656
rect 26998 77642 27138 77656
rect 27288 77642 28096 77656
rect 28246 77642 28386 77656
rect 28536 77642 29344 77656
rect 29494 77642 29634 77656
rect 29784 77642 30592 77656
rect 30742 77642 30882 77656
rect 31032 77642 31840 77656
rect 31990 77642 32130 77656
rect 32280 77642 33088 77656
rect 33238 77642 33378 77656
rect 33528 77642 34336 77656
rect 34486 77642 34626 77656
rect 34776 77642 35584 77656
rect 35734 77642 35874 77656
rect 36024 77642 36832 77656
rect 36982 77642 37122 77656
rect 37272 77642 38080 77656
rect 38230 77642 38370 77656
rect 38520 77642 39328 77656
rect 39478 77642 39618 77656
rect 39768 77642 40576 77656
rect 40726 77642 40866 77656
rect 41016 77642 41824 77656
rect 41974 77642 42114 77656
rect 42264 77642 43072 77656
rect 43222 77642 43362 77656
rect 43512 77642 44320 77656
rect 44470 77642 44610 77656
rect 44760 77642 45568 77656
rect 45718 77642 45858 77656
rect 46008 77642 46816 77656
rect 46966 77642 47106 77656
rect 47256 77642 48064 77656
rect 48214 77642 48354 77656
rect 48504 77642 49312 77656
rect 49462 77642 49602 77656
rect 49752 77642 50560 77656
rect 50710 77642 50850 77656
rect 51000 77642 51808 77656
rect 51958 77642 52098 77656
rect 52248 77642 53056 77656
rect 53206 77642 53346 77656
rect 53496 77642 54304 77656
rect 54454 77642 54594 77656
rect 54744 77642 55552 77656
rect 55702 77642 55842 77656
rect 55992 77642 56800 77656
rect 56950 77642 57090 77656
rect 57240 77642 58048 77656
rect 58198 77642 58338 77656
rect 58488 77642 58934 77656
rect 16898 77594 16980 77608
rect 17188 77594 17270 77608
rect 18146 77594 18228 77608
rect 18436 77594 18518 77608
rect 19394 77594 19476 77608
rect 19684 77594 19766 77608
rect 20642 77594 20724 77608
rect 20932 77594 21014 77608
rect 21890 77594 21972 77608
rect 22180 77594 22262 77608
rect 23138 77594 23220 77608
rect 23428 77594 23510 77608
rect 24386 77594 24468 77608
rect 24676 77594 24758 77608
rect 25634 77594 25716 77608
rect 25924 77594 26006 77608
rect 26882 77594 26964 77608
rect 27172 77594 27254 77608
rect 28130 77594 28212 77608
rect 28420 77594 28502 77608
rect 29378 77594 29460 77608
rect 29668 77594 29750 77608
rect 30626 77594 30708 77608
rect 30916 77594 30998 77608
rect 31874 77594 31956 77608
rect 32164 77594 32246 77608
rect 33122 77594 33204 77608
rect 33412 77594 33494 77608
rect 34370 77594 34452 77608
rect 34660 77594 34742 77608
rect 35618 77594 35700 77608
rect 35908 77594 35990 77608
rect 36866 77594 36948 77608
rect 37156 77594 37238 77608
rect 38114 77594 38196 77608
rect 38404 77594 38486 77608
rect 39362 77594 39444 77608
rect 39652 77594 39734 77608
rect 40610 77594 40692 77608
rect 40900 77594 40982 77608
rect 41858 77594 41940 77608
rect 42148 77594 42230 77608
rect 43106 77594 43188 77608
rect 43396 77594 43478 77608
rect 44354 77594 44436 77608
rect 44644 77594 44726 77608
rect 45602 77594 45684 77608
rect 45892 77594 45974 77608
rect 46850 77594 46932 77608
rect 47140 77594 47222 77608
rect 48098 77594 48180 77608
rect 48388 77594 48470 77608
rect 49346 77594 49428 77608
rect 49636 77594 49718 77608
rect 50594 77594 50676 77608
rect 50884 77594 50966 77608
rect 51842 77594 51924 77608
rect 52132 77594 52214 77608
rect 53090 77594 53172 77608
rect 53380 77594 53462 77608
rect 54338 77594 54420 77608
rect 54628 77594 54710 77608
rect 55586 77594 55668 77608
rect 55876 77594 55958 77608
rect 56834 77594 56916 77608
rect 57124 77594 57206 77608
rect 58082 77594 58164 77608
rect 58372 77594 58454 77608
rect 16418 77546 58934 77594
rect 16418 77388 58934 77498
rect 16418 77292 58934 77340
rect 16898 77278 16980 77292
rect 17188 77278 17270 77292
rect 18146 77278 18228 77292
rect 18436 77278 18518 77292
rect 19394 77278 19476 77292
rect 19684 77278 19766 77292
rect 20642 77278 20724 77292
rect 20932 77278 21014 77292
rect 21890 77278 21972 77292
rect 22180 77278 22262 77292
rect 23138 77278 23220 77292
rect 23428 77278 23510 77292
rect 24386 77278 24468 77292
rect 24676 77278 24758 77292
rect 25634 77278 25716 77292
rect 25924 77278 26006 77292
rect 26882 77278 26964 77292
rect 27172 77278 27254 77292
rect 28130 77278 28212 77292
rect 28420 77278 28502 77292
rect 29378 77278 29460 77292
rect 29668 77278 29750 77292
rect 30626 77278 30708 77292
rect 30916 77278 30998 77292
rect 31874 77278 31956 77292
rect 32164 77278 32246 77292
rect 33122 77278 33204 77292
rect 33412 77278 33494 77292
rect 34370 77278 34452 77292
rect 34660 77278 34742 77292
rect 35618 77278 35700 77292
rect 35908 77278 35990 77292
rect 36866 77278 36948 77292
rect 37156 77278 37238 77292
rect 38114 77278 38196 77292
rect 38404 77278 38486 77292
rect 39362 77278 39444 77292
rect 39652 77278 39734 77292
rect 40610 77278 40692 77292
rect 40900 77278 40982 77292
rect 41858 77278 41940 77292
rect 42148 77278 42230 77292
rect 43106 77278 43188 77292
rect 43396 77278 43478 77292
rect 44354 77278 44436 77292
rect 44644 77278 44726 77292
rect 45602 77278 45684 77292
rect 45892 77278 45974 77292
rect 46850 77278 46932 77292
rect 47140 77278 47222 77292
rect 48098 77278 48180 77292
rect 48388 77278 48470 77292
rect 49346 77278 49428 77292
rect 49636 77278 49718 77292
rect 50594 77278 50676 77292
rect 50884 77278 50966 77292
rect 51842 77278 51924 77292
rect 52132 77278 52214 77292
rect 53090 77278 53172 77292
rect 53380 77278 53462 77292
rect 54338 77278 54420 77292
rect 54628 77278 54710 77292
rect 55586 77278 55668 77292
rect 55876 77278 55958 77292
rect 56834 77278 56916 77292
rect 57124 77278 57206 77292
rect 58082 77278 58164 77292
rect 58372 77278 58454 77292
rect 16418 77230 16864 77244
rect 17014 77230 17154 77244
rect 17304 77230 18112 77244
rect 18262 77230 18402 77244
rect 18552 77230 19360 77244
rect 19510 77230 19650 77244
rect 19800 77230 20608 77244
rect 20758 77230 20898 77244
rect 21048 77230 21856 77244
rect 22006 77230 22146 77244
rect 22296 77230 23104 77244
rect 23254 77230 23394 77244
rect 23544 77230 24352 77244
rect 24502 77230 24642 77244
rect 24792 77230 25600 77244
rect 25750 77230 25890 77244
rect 26040 77230 26848 77244
rect 26998 77230 27138 77244
rect 27288 77230 28096 77244
rect 28246 77230 28386 77244
rect 28536 77230 29344 77244
rect 29494 77230 29634 77244
rect 29784 77230 30592 77244
rect 30742 77230 30882 77244
rect 31032 77230 31840 77244
rect 31990 77230 32130 77244
rect 32280 77230 33088 77244
rect 33238 77230 33378 77244
rect 33528 77230 34336 77244
rect 34486 77230 34626 77244
rect 34776 77230 35584 77244
rect 35734 77230 35874 77244
rect 36024 77230 36832 77244
rect 36982 77230 37122 77244
rect 37272 77230 38080 77244
rect 38230 77230 38370 77244
rect 38520 77230 39328 77244
rect 39478 77230 39618 77244
rect 39768 77230 40576 77244
rect 40726 77230 40866 77244
rect 41016 77230 41824 77244
rect 41974 77230 42114 77244
rect 42264 77230 43072 77244
rect 43222 77230 43362 77244
rect 43512 77230 44320 77244
rect 44470 77230 44610 77244
rect 44760 77230 45568 77244
rect 45718 77230 45858 77244
rect 46008 77230 46816 77244
rect 46966 77230 47106 77244
rect 47256 77230 48064 77244
rect 48214 77230 48354 77244
rect 48504 77230 49312 77244
rect 49462 77230 49602 77244
rect 49752 77230 50560 77244
rect 50710 77230 50850 77244
rect 51000 77230 51808 77244
rect 51958 77230 52098 77244
rect 52248 77230 53056 77244
rect 53206 77230 53346 77244
rect 53496 77230 54304 77244
rect 54454 77230 54594 77244
rect 54744 77230 55552 77244
rect 55702 77230 55842 77244
rect 55992 77230 56800 77244
rect 56950 77230 57090 77244
rect 57240 77230 58048 77244
rect 58198 77230 58338 77244
rect 58488 77230 58934 77244
rect 16418 77182 58934 77230
rect 16418 77168 16864 77182
rect 17014 77168 17154 77182
rect 17304 77168 18112 77182
rect 18262 77168 18402 77182
rect 18552 77168 19360 77182
rect 19510 77168 19650 77182
rect 19800 77168 20608 77182
rect 20758 77168 20898 77182
rect 21048 77168 21856 77182
rect 22006 77168 22146 77182
rect 22296 77168 23104 77182
rect 23254 77168 23394 77182
rect 23544 77168 24352 77182
rect 24502 77168 24642 77182
rect 24792 77168 25600 77182
rect 25750 77168 25890 77182
rect 26040 77168 26848 77182
rect 26998 77168 27138 77182
rect 27288 77168 28096 77182
rect 28246 77168 28386 77182
rect 28536 77168 29344 77182
rect 29494 77168 29634 77182
rect 29784 77168 30592 77182
rect 30742 77168 30882 77182
rect 31032 77168 31840 77182
rect 31990 77168 32130 77182
rect 32280 77168 33088 77182
rect 33238 77168 33378 77182
rect 33528 77168 34336 77182
rect 34486 77168 34626 77182
rect 34776 77168 35584 77182
rect 35734 77168 35874 77182
rect 36024 77168 36832 77182
rect 36982 77168 37122 77182
rect 37272 77168 38080 77182
rect 38230 77168 38370 77182
rect 38520 77168 39328 77182
rect 39478 77168 39618 77182
rect 39768 77168 40576 77182
rect 40726 77168 40866 77182
rect 41016 77168 41824 77182
rect 41974 77168 42114 77182
rect 42264 77168 43072 77182
rect 43222 77168 43362 77182
rect 43512 77168 44320 77182
rect 44470 77168 44610 77182
rect 44760 77168 45568 77182
rect 45718 77168 45858 77182
rect 46008 77168 46816 77182
rect 46966 77168 47106 77182
rect 47256 77168 48064 77182
rect 48214 77168 48354 77182
rect 48504 77168 49312 77182
rect 49462 77168 49602 77182
rect 49752 77168 50560 77182
rect 50710 77168 50850 77182
rect 51000 77168 51808 77182
rect 51958 77168 52098 77182
rect 52248 77168 53056 77182
rect 53206 77168 53346 77182
rect 53496 77168 54304 77182
rect 54454 77168 54594 77182
rect 54744 77168 55552 77182
rect 55702 77168 55842 77182
rect 55992 77168 56800 77182
rect 56950 77168 57090 77182
rect 57240 77168 58048 77182
rect 58198 77168 58338 77182
rect 58488 77168 58934 77182
rect 16898 77120 16980 77134
rect 17188 77120 17270 77134
rect 18146 77120 18228 77134
rect 18436 77120 18518 77134
rect 19394 77120 19476 77134
rect 19684 77120 19766 77134
rect 20642 77120 20724 77134
rect 20932 77120 21014 77134
rect 21890 77120 21972 77134
rect 22180 77120 22262 77134
rect 23138 77120 23220 77134
rect 23428 77120 23510 77134
rect 24386 77120 24468 77134
rect 24676 77120 24758 77134
rect 25634 77120 25716 77134
rect 25924 77120 26006 77134
rect 26882 77120 26964 77134
rect 27172 77120 27254 77134
rect 28130 77120 28212 77134
rect 28420 77120 28502 77134
rect 29378 77120 29460 77134
rect 29668 77120 29750 77134
rect 30626 77120 30708 77134
rect 30916 77120 30998 77134
rect 31874 77120 31956 77134
rect 32164 77120 32246 77134
rect 33122 77120 33204 77134
rect 33412 77120 33494 77134
rect 34370 77120 34452 77134
rect 34660 77120 34742 77134
rect 35618 77120 35700 77134
rect 35908 77120 35990 77134
rect 36866 77120 36948 77134
rect 37156 77120 37238 77134
rect 38114 77120 38196 77134
rect 38404 77120 38486 77134
rect 39362 77120 39444 77134
rect 39652 77120 39734 77134
rect 40610 77120 40692 77134
rect 40900 77120 40982 77134
rect 41858 77120 41940 77134
rect 42148 77120 42230 77134
rect 43106 77120 43188 77134
rect 43396 77120 43478 77134
rect 44354 77120 44436 77134
rect 44644 77120 44726 77134
rect 45602 77120 45684 77134
rect 45892 77120 45974 77134
rect 46850 77120 46932 77134
rect 47140 77120 47222 77134
rect 48098 77120 48180 77134
rect 48388 77120 48470 77134
rect 49346 77120 49428 77134
rect 49636 77120 49718 77134
rect 50594 77120 50676 77134
rect 50884 77120 50966 77134
rect 51842 77120 51924 77134
rect 52132 77120 52214 77134
rect 53090 77120 53172 77134
rect 53380 77120 53462 77134
rect 54338 77120 54420 77134
rect 54628 77120 54710 77134
rect 55586 77120 55668 77134
rect 55876 77120 55958 77134
rect 56834 77120 56916 77134
rect 57124 77120 57206 77134
rect 58082 77120 58164 77134
rect 58372 77120 58454 77134
rect 16418 77072 58934 77120
rect 16418 76976 58934 77024
rect 16898 76962 16980 76976
rect 17188 76962 17270 76976
rect 18146 76962 18228 76976
rect 18436 76962 18518 76976
rect 19394 76962 19476 76976
rect 19684 76962 19766 76976
rect 20642 76962 20724 76976
rect 20932 76962 21014 76976
rect 21890 76962 21972 76976
rect 22180 76962 22262 76976
rect 23138 76962 23220 76976
rect 23428 76962 23510 76976
rect 24386 76962 24468 76976
rect 24676 76962 24758 76976
rect 25634 76962 25716 76976
rect 25924 76962 26006 76976
rect 26882 76962 26964 76976
rect 27172 76962 27254 76976
rect 28130 76962 28212 76976
rect 28420 76962 28502 76976
rect 29378 76962 29460 76976
rect 29668 76962 29750 76976
rect 30626 76962 30708 76976
rect 30916 76962 30998 76976
rect 31874 76962 31956 76976
rect 32164 76962 32246 76976
rect 33122 76962 33204 76976
rect 33412 76962 33494 76976
rect 34370 76962 34452 76976
rect 34660 76962 34742 76976
rect 35618 76962 35700 76976
rect 35908 76962 35990 76976
rect 36866 76962 36948 76976
rect 37156 76962 37238 76976
rect 38114 76962 38196 76976
rect 38404 76962 38486 76976
rect 39362 76962 39444 76976
rect 39652 76962 39734 76976
rect 40610 76962 40692 76976
rect 40900 76962 40982 76976
rect 41858 76962 41940 76976
rect 42148 76962 42230 76976
rect 43106 76962 43188 76976
rect 43396 76962 43478 76976
rect 44354 76962 44436 76976
rect 44644 76962 44726 76976
rect 45602 76962 45684 76976
rect 45892 76962 45974 76976
rect 46850 76962 46932 76976
rect 47140 76962 47222 76976
rect 48098 76962 48180 76976
rect 48388 76962 48470 76976
rect 49346 76962 49428 76976
rect 49636 76962 49718 76976
rect 50594 76962 50676 76976
rect 50884 76962 50966 76976
rect 51842 76962 51924 76976
rect 52132 76962 52214 76976
rect 53090 76962 53172 76976
rect 53380 76962 53462 76976
rect 54338 76962 54420 76976
rect 54628 76962 54710 76976
rect 55586 76962 55668 76976
rect 55876 76962 55958 76976
rect 56834 76962 56916 76976
rect 57124 76962 57206 76976
rect 58082 76962 58164 76976
rect 58372 76962 58454 76976
rect 16418 76914 16864 76928
rect 17014 76914 17154 76928
rect 17304 76914 18112 76928
rect 18262 76914 18402 76928
rect 18552 76914 19360 76928
rect 19510 76914 19650 76928
rect 19800 76914 20608 76928
rect 20758 76914 20898 76928
rect 21048 76914 21856 76928
rect 22006 76914 22146 76928
rect 22296 76914 23104 76928
rect 23254 76914 23394 76928
rect 23544 76914 24352 76928
rect 24502 76914 24642 76928
rect 24792 76914 25600 76928
rect 25750 76914 25890 76928
rect 26040 76914 26848 76928
rect 26998 76914 27138 76928
rect 27288 76914 28096 76928
rect 28246 76914 28386 76928
rect 28536 76914 29344 76928
rect 29494 76914 29634 76928
rect 29784 76914 30592 76928
rect 30742 76914 30882 76928
rect 31032 76914 31840 76928
rect 31990 76914 32130 76928
rect 32280 76914 33088 76928
rect 33238 76914 33378 76928
rect 33528 76914 34336 76928
rect 34486 76914 34626 76928
rect 34776 76914 35584 76928
rect 35734 76914 35874 76928
rect 36024 76914 36832 76928
rect 36982 76914 37122 76928
rect 37272 76914 38080 76928
rect 38230 76914 38370 76928
rect 38520 76914 39328 76928
rect 39478 76914 39618 76928
rect 39768 76914 40576 76928
rect 40726 76914 40866 76928
rect 41016 76914 41824 76928
rect 41974 76914 42114 76928
rect 42264 76914 43072 76928
rect 43222 76914 43362 76928
rect 43512 76914 44320 76928
rect 44470 76914 44610 76928
rect 44760 76914 45568 76928
rect 45718 76914 45858 76928
rect 46008 76914 46816 76928
rect 46966 76914 47106 76928
rect 47256 76914 48064 76928
rect 48214 76914 48354 76928
rect 48504 76914 49312 76928
rect 49462 76914 49602 76928
rect 49752 76914 50560 76928
rect 50710 76914 50850 76928
rect 51000 76914 51808 76928
rect 51958 76914 52098 76928
rect 52248 76914 53056 76928
rect 53206 76914 53346 76928
rect 53496 76914 54304 76928
rect 54454 76914 54594 76928
rect 54744 76914 55552 76928
rect 55702 76914 55842 76928
rect 55992 76914 56800 76928
rect 56950 76914 57090 76928
rect 57240 76914 58048 76928
rect 58198 76914 58338 76928
rect 58488 76914 58934 76928
rect 16418 76866 58934 76914
rect 16418 76852 16864 76866
rect 17014 76852 17154 76866
rect 17304 76852 18112 76866
rect 18262 76852 18402 76866
rect 18552 76852 19360 76866
rect 19510 76852 19650 76866
rect 19800 76852 20608 76866
rect 20758 76852 20898 76866
rect 21048 76852 21856 76866
rect 22006 76852 22146 76866
rect 22296 76852 23104 76866
rect 23254 76852 23394 76866
rect 23544 76852 24352 76866
rect 24502 76852 24642 76866
rect 24792 76852 25600 76866
rect 25750 76852 25890 76866
rect 26040 76852 26848 76866
rect 26998 76852 27138 76866
rect 27288 76852 28096 76866
rect 28246 76852 28386 76866
rect 28536 76852 29344 76866
rect 29494 76852 29634 76866
rect 29784 76852 30592 76866
rect 30742 76852 30882 76866
rect 31032 76852 31840 76866
rect 31990 76852 32130 76866
rect 32280 76852 33088 76866
rect 33238 76852 33378 76866
rect 33528 76852 34336 76866
rect 34486 76852 34626 76866
rect 34776 76852 35584 76866
rect 35734 76852 35874 76866
rect 36024 76852 36832 76866
rect 36982 76852 37122 76866
rect 37272 76852 38080 76866
rect 38230 76852 38370 76866
rect 38520 76852 39328 76866
rect 39478 76852 39618 76866
rect 39768 76852 40576 76866
rect 40726 76852 40866 76866
rect 41016 76852 41824 76866
rect 41974 76852 42114 76866
rect 42264 76852 43072 76866
rect 43222 76852 43362 76866
rect 43512 76852 44320 76866
rect 44470 76852 44610 76866
rect 44760 76852 45568 76866
rect 45718 76852 45858 76866
rect 46008 76852 46816 76866
rect 46966 76852 47106 76866
rect 47256 76852 48064 76866
rect 48214 76852 48354 76866
rect 48504 76852 49312 76866
rect 49462 76852 49602 76866
rect 49752 76852 50560 76866
rect 50710 76852 50850 76866
rect 51000 76852 51808 76866
rect 51958 76852 52098 76866
rect 52248 76852 53056 76866
rect 53206 76852 53346 76866
rect 53496 76852 54304 76866
rect 54454 76852 54594 76866
rect 54744 76852 55552 76866
rect 55702 76852 55842 76866
rect 55992 76852 56800 76866
rect 56950 76852 57090 76866
rect 57240 76852 58048 76866
rect 58198 76852 58338 76866
rect 58488 76852 58934 76866
rect 16898 76804 16980 76818
rect 17188 76804 17270 76818
rect 18146 76804 18228 76818
rect 18436 76804 18518 76818
rect 19394 76804 19476 76818
rect 19684 76804 19766 76818
rect 20642 76804 20724 76818
rect 20932 76804 21014 76818
rect 21890 76804 21972 76818
rect 22180 76804 22262 76818
rect 23138 76804 23220 76818
rect 23428 76804 23510 76818
rect 24386 76804 24468 76818
rect 24676 76804 24758 76818
rect 25634 76804 25716 76818
rect 25924 76804 26006 76818
rect 26882 76804 26964 76818
rect 27172 76804 27254 76818
rect 28130 76804 28212 76818
rect 28420 76804 28502 76818
rect 29378 76804 29460 76818
rect 29668 76804 29750 76818
rect 30626 76804 30708 76818
rect 30916 76804 30998 76818
rect 31874 76804 31956 76818
rect 32164 76804 32246 76818
rect 33122 76804 33204 76818
rect 33412 76804 33494 76818
rect 34370 76804 34452 76818
rect 34660 76804 34742 76818
rect 35618 76804 35700 76818
rect 35908 76804 35990 76818
rect 36866 76804 36948 76818
rect 37156 76804 37238 76818
rect 38114 76804 38196 76818
rect 38404 76804 38486 76818
rect 39362 76804 39444 76818
rect 39652 76804 39734 76818
rect 40610 76804 40692 76818
rect 40900 76804 40982 76818
rect 41858 76804 41940 76818
rect 42148 76804 42230 76818
rect 43106 76804 43188 76818
rect 43396 76804 43478 76818
rect 44354 76804 44436 76818
rect 44644 76804 44726 76818
rect 45602 76804 45684 76818
rect 45892 76804 45974 76818
rect 46850 76804 46932 76818
rect 47140 76804 47222 76818
rect 48098 76804 48180 76818
rect 48388 76804 48470 76818
rect 49346 76804 49428 76818
rect 49636 76804 49718 76818
rect 50594 76804 50676 76818
rect 50884 76804 50966 76818
rect 51842 76804 51924 76818
rect 52132 76804 52214 76818
rect 53090 76804 53172 76818
rect 53380 76804 53462 76818
rect 54338 76804 54420 76818
rect 54628 76804 54710 76818
rect 55586 76804 55668 76818
rect 55876 76804 55958 76818
rect 56834 76804 56916 76818
rect 57124 76804 57206 76818
rect 58082 76804 58164 76818
rect 58372 76804 58454 76818
rect 16418 76756 58934 76804
rect 16418 76598 58934 76708
rect 16418 76502 58934 76550
rect 16898 76488 16980 76502
rect 17188 76488 17270 76502
rect 18146 76488 18228 76502
rect 18436 76488 18518 76502
rect 19394 76488 19476 76502
rect 19684 76488 19766 76502
rect 20642 76488 20724 76502
rect 20932 76488 21014 76502
rect 21890 76488 21972 76502
rect 22180 76488 22262 76502
rect 23138 76488 23220 76502
rect 23428 76488 23510 76502
rect 24386 76488 24468 76502
rect 24676 76488 24758 76502
rect 25634 76488 25716 76502
rect 25924 76488 26006 76502
rect 26882 76488 26964 76502
rect 27172 76488 27254 76502
rect 28130 76488 28212 76502
rect 28420 76488 28502 76502
rect 29378 76488 29460 76502
rect 29668 76488 29750 76502
rect 30626 76488 30708 76502
rect 30916 76488 30998 76502
rect 31874 76488 31956 76502
rect 32164 76488 32246 76502
rect 33122 76488 33204 76502
rect 33412 76488 33494 76502
rect 34370 76488 34452 76502
rect 34660 76488 34742 76502
rect 35618 76488 35700 76502
rect 35908 76488 35990 76502
rect 36866 76488 36948 76502
rect 37156 76488 37238 76502
rect 38114 76488 38196 76502
rect 38404 76488 38486 76502
rect 39362 76488 39444 76502
rect 39652 76488 39734 76502
rect 40610 76488 40692 76502
rect 40900 76488 40982 76502
rect 41858 76488 41940 76502
rect 42148 76488 42230 76502
rect 43106 76488 43188 76502
rect 43396 76488 43478 76502
rect 44354 76488 44436 76502
rect 44644 76488 44726 76502
rect 45602 76488 45684 76502
rect 45892 76488 45974 76502
rect 46850 76488 46932 76502
rect 47140 76488 47222 76502
rect 48098 76488 48180 76502
rect 48388 76488 48470 76502
rect 49346 76488 49428 76502
rect 49636 76488 49718 76502
rect 50594 76488 50676 76502
rect 50884 76488 50966 76502
rect 51842 76488 51924 76502
rect 52132 76488 52214 76502
rect 53090 76488 53172 76502
rect 53380 76488 53462 76502
rect 54338 76488 54420 76502
rect 54628 76488 54710 76502
rect 55586 76488 55668 76502
rect 55876 76488 55958 76502
rect 56834 76488 56916 76502
rect 57124 76488 57206 76502
rect 58082 76488 58164 76502
rect 58372 76488 58454 76502
rect 16418 76440 16864 76454
rect 17014 76440 17154 76454
rect 17304 76440 18112 76454
rect 18262 76440 18402 76454
rect 18552 76440 19360 76454
rect 19510 76440 19650 76454
rect 19800 76440 20608 76454
rect 20758 76440 20898 76454
rect 21048 76440 21856 76454
rect 22006 76440 22146 76454
rect 22296 76440 23104 76454
rect 23254 76440 23394 76454
rect 23544 76440 24352 76454
rect 24502 76440 24642 76454
rect 24792 76440 25600 76454
rect 25750 76440 25890 76454
rect 26040 76440 26848 76454
rect 26998 76440 27138 76454
rect 27288 76440 28096 76454
rect 28246 76440 28386 76454
rect 28536 76440 29344 76454
rect 29494 76440 29634 76454
rect 29784 76440 30592 76454
rect 30742 76440 30882 76454
rect 31032 76440 31840 76454
rect 31990 76440 32130 76454
rect 32280 76440 33088 76454
rect 33238 76440 33378 76454
rect 33528 76440 34336 76454
rect 34486 76440 34626 76454
rect 34776 76440 35584 76454
rect 35734 76440 35874 76454
rect 36024 76440 36832 76454
rect 36982 76440 37122 76454
rect 37272 76440 38080 76454
rect 38230 76440 38370 76454
rect 38520 76440 39328 76454
rect 39478 76440 39618 76454
rect 39768 76440 40576 76454
rect 40726 76440 40866 76454
rect 41016 76440 41824 76454
rect 41974 76440 42114 76454
rect 42264 76440 43072 76454
rect 43222 76440 43362 76454
rect 43512 76440 44320 76454
rect 44470 76440 44610 76454
rect 44760 76440 45568 76454
rect 45718 76440 45858 76454
rect 46008 76440 46816 76454
rect 46966 76440 47106 76454
rect 47256 76440 48064 76454
rect 48214 76440 48354 76454
rect 48504 76440 49312 76454
rect 49462 76440 49602 76454
rect 49752 76440 50560 76454
rect 50710 76440 50850 76454
rect 51000 76440 51808 76454
rect 51958 76440 52098 76454
rect 52248 76440 53056 76454
rect 53206 76440 53346 76454
rect 53496 76440 54304 76454
rect 54454 76440 54594 76454
rect 54744 76440 55552 76454
rect 55702 76440 55842 76454
rect 55992 76440 56800 76454
rect 56950 76440 57090 76454
rect 57240 76440 58048 76454
rect 58198 76440 58338 76454
rect 58488 76440 58934 76454
rect 16418 76392 58934 76440
rect 16418 76378 16864 76392
rect 17014 76378 17154 76392
rect 17304 76378 18112 76392
rect 18262 76378 18402 76392
rect 18552 76378 19360 76392
rect 19510 76378 19650 76392
rect 19800 76378 20608 76392
rect 20758 76378 20898 76392
rect 21048 76378 21856 76392
rect 22006 76378 22146 76392
rect 22296 76378 23104 76392
rect 23254 76378 23394 76392
rect 23544 76378 24352 76392
rect 24502 76378 24642 76392
rect 24792 76378 25600 76392
rect 25750 76378 25890 76392
rect 26040 76378 26848 76392
rect 26998 76378 27138 76392
rect 27288 76378 28096 76392
rect 28246 76378 28386 76392
rect 28536 76378 29344 76392
rect 29494 76378 29634 76392
rect 29784 76378 30592 76392
rect 30742 76378 30882 76392
rect 31032 76378 31840 76392
rect 31990 76378 32130 76392
rect 32280 76378 33088 76392
rect 33238 76378 33378 76392
rect 33528 76378 34336 76392
rect 34486 76378 34626 76392
rect 34776 76378 35584 76392
rect 35734 76378 35874 76392
rect 36024 76378 36832 76392
rect 36982 76378 37122 76392
rect 37272 76378 38080 76392
rect 38230 76378 38370 76392
rect 38520 76378 39328 76392
rect 39478 76378 39618 76392
rect 39768 76378 40576 76392
rect 40726 76378 40866 76392
rect 41016 76378 41824 76392
rect 41974 76378 42114 76392
rect 42264 76378 43072 76392
rect 43222 76378 43362 76392
rect 43512 76378 44320 76392
rect 44470 76378 44610 76392
rect 44760 76378 45568 76392
rect 45718 76378 45858 76392
rect 46008 76378 46816 76392
rect 46966 76378 47106 76392
rect 47256 76378 48064 76392
rect 48214 76378 48354 76392
rect 48504 76378 49312 76392
rect 49462 76378 49602 76392
rect 49752 76378 50560 76392
rect 50710 76378 50850 76392
rect 51000 76378 51808 76392
rect 51958 76378 52098 76392
rect 52248 76378 53056 76392
rect 53206 76378 53346 76392
rect 53496 76378 54304 76392
rect 54454 76378 54594 76392
rect 54744 76378 55552 76392
rect 55702 76378 55842 76392
rect 55992 76378 56800 76392
rect 56950 76378 57090 76392
rect 57240 76378 58048 76392
rect 58198 76378 58338 76392
rect 58488 76378 58934 76392
rect 16898 76330 16980 76344
rect 17188 76330 17270 76344
rect 18146 76330 18228 76344
rect 18436 76330 18518 76344
rect 19394 76330 19476 76344
rect 19684 76330 19766 76344
rect 20642 76330 20724 76344
rect 20932 76330 21014 76344
rect 21890 76330 21972 76344
rect 22180 76330 22262 76344
rect 23138 76330 23220 76344
rect 23428 76330 23510 76344
rect 24386 76330 24468 76344
rect 24676 76330 24758 76344
rect 25634 76330 25716 76344
rect 25924 76330 26006 76344
rect 26882 76330 26964 76344
rect 27172 76330 27254 76344
rect 28130 76330 28212 76344
rect 28420 76330 28502 76344
rect 29378 76330 29460 76344
rect 29668 76330 29750 76344
rect 30626 76330 30708 76344
rect 30916 76330 30998 76344
rect 31874 76330 31956 76344
rect 32164 76330 32246 76344
rect 33122 76330 33204 76344
rect 33412 76330 33494 76344
rect 34370 76330 34452 76344
rect 34660 76330 34742 76344
rect 35618 76330 35700 76344
rect 35908 76330 35990 76344
rect 36866 76330 36948 76344
rect 37156 76330 37238 76344
rect 38114 76330 38196 76344
rect 38404 76330 38486 76344
rect 39362 76330 39444 76344
rect 39652 76330 39734 76344
rect 40610 76330 40692 76344
rect 40900 76330 40982 76344
rect 41858 76330 41940 76344
rect 42148 76330 42230 76344
rect 43106 76330 43188 76344
rect 43396 76330 43478 76344
rect 44354 76330 44436 76344
rect 44644 76330 44726 76344
rect 45602 76330 45684 76344
rect 45892 76330 45974 76344
rect 46850 76330 46932 76344
rect 47140 76330 47222 76344
rect 48098 76330 48180 76344
rect 48388 76330 48470 76344
rect 49346 76330 49428 76344
rect 49636 76330 49718 76344
rect 50594 76330 50676 76344
rect 50884 76330 50966 76344
rect 51842 76330 51924 76344
rect 52132 76330 52214 76344
rect 53090 76330 53172 76344
rect 53380 76330 53462 76344
rect 54338 76330 54420 76344
rect 54628 76330 54710 76344
rect 55586 76330 55668 76344
rect 55876 76330 55958 76344
rect 56834 76330 56916 76344
rect 57124 76330 57206 76344
rect 58082 76330 58164 76344
rect 58372 76330 58454 76344
rect 16418 76282 58934 76330
rect 16418 76186 58934 76234
rect 16898 76172 16980 76186
rect 17188 76172 17270 76186
rect 18146 76172 18228 76186
rect 18436 76172 18518 76186
rect 19394 76172 19476 76186
rect 19684 76172 19766 76186
rect 20642 76172 20724 76186
rect 20932 76172 21014 76186
rect 21890 76172 21972 76186
rect 22180 76172 22262 76186
rect 23138 76172 23220 76186
rect 23428 76172 23510 76186
rect 24386 76172 24468 76186
rect 24676 76172 24758 76186
rect 25634 76172 25716 76186
rect 25924 76172 26006 76186
rect 26882 76172 26964 76186
rect 27172 76172 27254 76186
rect 28130 76172 28212 76186
rect 28420 76172 28502 76186
rect 29378 76172 29460 76186
rect 29668 76172 29750 76186
rect 30626 76172 30708 76186
rect 30916 76172 30998 76186
rect 31874 76172 31956 76186
rect 32164 76172 32246 76186
rect 33122 76172 33204 76186
rect 33412 76172 33494 76186
rect 34370 76172 34452 76186
rect 34660 76172 34742 76186
rect 35618 76172 35700 76186
rect 35908 76172 35990 76186
rect 36866 76172 36948 76186
rect 37156 76172 37238 76186
rect 38114 76172 38196 76186
rect 38404 76172 38486 76186
rect 39362 76172 39444 76186
rect 39652 76172 39734 76186
rect 40610 76172 40692 76186
rect 40900 76172 40982 76186
rect 41858 76172 41940 76186
rect 42148 76172 42230 76186
rect 43106 76172 43188 76186
rect 43396 76172 43478 76186
rect 44354 76172 44436 76186
rect 44644 76172 44726 76186
rect 45602 76172 45684 76186
rect 45892 76172 45974 76186
rect 46850 76172 46932 76186
rect 47140 76172 47222 76186
rect 48098 76172 48180 76186
rect 48388 76172 48470 76186
rect 49346 76172 49428 76186
rect 49636 76172 49718 76186
rect 50594 76172 50676 76186
rect 50884 76172 50966 76186
rect 51842 76172 51924 76186
rect 52132 76172 52214 76186
rect 53090 76172 53172 76186
rect 53380 76172 53462 76186
rect 54338 76172 54420 76186
rect 54628 76172 54710 76186
rect 55586 76172 55668 76186
rect 55876 76172 55958 76186
rect 56834 76172 56916 76186
rect 57124 76172 57206 76186
rect 58082 76172 58164 76186
rect 58372 76172 58454 76186
rect 16418 76124 16864 76138
rect 17014 76124 17154 76138
rect 17304 76124 18112 76138
rect 18262 76124 18402 76138
rect 18552 76124 19360 76138
rect 19510 76124 19650 76138
rect 19800 76124 20608 76138
rect 20758 76124 20898 76138
rect 21048 76124 21856 76138
rect 22006 76124 22146 76138
rect 22296 76124 23104 76138
rect 23254 76124 23394 76138
rect 23544 76124 24352 76138
rect 24502 76124 24642 76138
rect 24792 76124 25600 76138
rect 25750 76124 25890 76138
rect 26040 76124 26848 76138
rect 26998 76124 27138 76138
rect 27288 76124 28096 76138
rect 28246 76124 28386 76138
rect 28536 76124 29344 76138
rect 29494 76124 29634 76138
rect 29784 76124 30592 76138
rect 30742 76124 30882 76138
rect 31032 76124 31840 76138
rect 31990 76124 32130 76138
rect 32280 76124 33088 76138
rect 33238 76124 33378 76138
rect 33528 76124 34336 76138
rect 34486 76124 34626 76138
rect 34776 76124 35584 76138
rect 35734 76124 35874 76138
rect 36024 76124 36832 76138
rect 36982 76124 37122 76138
rect 37272 76124 38080 76138
rect 38230 76124 38370 76138
rect 38520 76124 39328 76138
rect 39478 76124 39618 76138
rect 39768 76124 40576 76138
rect 40726 76124 40866 76138
rect 41016 76124 41824 76138
rect 41974 76124 42114 76138
rect 42264 76124 43072 76138
rect 43222 76124 43362 76138
rect 43512 76124 44320 76138
rect 44470 76124 44610 76138
rect 44760 76124 45568 76138
rect 45718 76124 45858 76138
rect 46008 76124 46816 76138
rect 46966 76124 47106 76138
rect 47256 76124 48064 76138
rect 48214 76124 48354 76138
rect 48504 76124 49312 76138
rect 49462 76124 49602 76138
rect 49752 76124 50560 76138
rect 50710 76124 50850 76138
rect 51000 76124 51808 76138
rect 51958 76124 52098 76138
rect 52248 76124 53056 76138
rect 53206 76124 53346 76138
rect 53496 76124 54304 76138
rect 54454 76124 54594 76138
rect 54744 76124 55552 76138
rect 55702 76124 55842 76138
rect 55992 76124 56800 76138
rect 56950 76124 57090 76138
rect 57240 76124 58048 76138
rect 58198 76124 58338 76138
rect 58488 76124 58934 76138
rect 16418 76076 58934 76124
rect 16418 76062 16864 76076
rect 17014 76062 17154 76076
rect 17304 76062 18112 76076
rect 18262 76062 18402 76076
rect 18552 76062 19360 76076
rect 19510 76062 19650 76076
rect 19800 76062 20608 76076
rect 20758 76062 20898 76076
rect 21048 76062 21856 76076
rect 22006 76062 22146 76076
rect 22296 76062 23104 76076
rect 23254 76062 23394 76076
rect 23544 76062 24352 76076
rect 24502 76062 24642 76076
rect 24792 76062 25600 76076
rect 25750 76062 25890 76076
rect 26040 76062 26848 76076
rect 26998 76062 27138 76076
rect 27288 76062 28096 76076
rect 28246 76062 28386 76076
rect 28536 76062 29344 76076
rect 29494 76062 29634 76076
rect 29784 76062 30592 76076
rect 30742 76062 30882 76076
rect 31032 76062 31840 76076
rect 31990 76062 32130 76076
rect 32280 76062 33088 76076
rect 33238 76062 33378 76076
rect 33528 76062 34336 76076
rect 34486 76062 34626 76076
rect 34776 76062 35584 76076
rect 35734 76062 35874 76076
rect 36024 76062 36832 76076
rect 36982 76062 37122 76076
rect 37272 76062 38080 76076
rect 38230 76062 38370 76076
rect 38520 76062 39328 76076
rect 39478 76062 39618 76076
rect 39768 76062 40576 76076
rect 40726 76062 40866 76076
rect 41016 76062 41824 76076
rect 41974 76062 42114 76076
rect 42264 76062 43072 76076
rect 43222 76062 43362 76076
rect 43512 76062 44320 76076
rect 44470 76062 44610 76076
rect 44760 76062 45568 76076
rect 45718 76062 45858 76076
rect 46008 76062 46816 76076
rect 46966 76062 47106 76076
rect 47256 76062 48064 76076
rect 48214 76062 48354 76076
rect 48504 76062 49312 76076
rect 49462 76062 49602 76076
rect 49752 76062 50560 76076
rect 50710 76062 50850 76076
rect 51000 76062 51808 76076
rect 51958 76062 52098 76076
rect 52248 76062 53056 76076
rect 53206 76062 53346 76076
rect 53496 76062 54304 76076
rect 54454 76062 54594 76076
rect 54744 76062 55552 76076
rect 55702 76062 55842 76076
rect 55992 76062 56800 76076
rect 56950 76062 57090 76076
rect 57240 76062 58048 76076
rect 58198 76062 58338 76076
rect 58488 76062 58934 76076
rect 16898 76014 16980 76028
rect 17188 76014 17270 76028
rect 18146 76014 18228 76028
rect 18436 76014 18518 76028
rect 19394 76014 19476 76028
rect 19684 76014 19766 76028
rect 20642 76014 20724 76028
rect 20932 76014 21014 76028
rect 21890 76014 21972 76028
rect 22180 76014 22262 76028
rect 23138 76014 23220 76028
rect 23428 76014 23510 76028
rect 24386 76014 24468 76028
rect 24676 76014 24758 76028
rect 25634 76014 25716 76028
rect 25924 76014 26006 76028
rect 26882 76014 26964 76028
rect 27172 76014 27254 76028
rect 28130 76014 28212 76028
rect 28420 76014 28502 76028
rect 29378 76014 29460 76028
rect 29668 76014 29750 76028
rect 30626 76014 30708 76028
rect 30916 76014 30998 76028
rect 31874 76014 31956 76028
rect 32164 76014 32246 76028
rect 33122 76014 33204 76028
rect 33412 76014 33494 76028
rect 34370 76014 34452 76028
rect 34660 76014 34742 76028
rect 35618 76014 35700 76028
rect 35908 76014 35990 76028
rect 36866 76014 36948 76028
rect 37156 76014 37238 76028
rect 38114 76014 38196 76028
rect 38404 76014 38486 76028
rect 39362 76014 39444 76028
rect 39652 76014 39734 76028
rect 40610 76014 40692 76028
rect 40900 76014 40982 76028
rect 41858 76014 41940 76028
rect 42148 76014 42230 76028
rect 43106 76014 43188 76028
rect 43396 76014 43478 76028
rect 44354 76014 44436 76028
rect 44644 76014 44726 76028
rect 45602 76014 45684 76028
rect 45892 76014 45974 76028
rect 46850 76014 46932 76028
rect 47140 76014 47222 76028
rect 48098 76014 48180 76028
rect 48388 76014 48470 76028
rect 49346 76014 49428 76028
rect 49636 76014 49718 76028
rect 50594 76014 50676 76028
rect 50884 76014 50966 76028
rect 51842 76014 51924 76028
rect 52132 76014 52214 76028
rect 53090 76014 53172 76028
rect 53380 76014 53462 76028
rect 54338 76014 54420 76028
rect 54628 76014 54710 76028
rect 55586 76014 55668 76028
rect 55876 76014 55958 76028
rect 56834 76014 56916 76028
rect 57124 76014 57206 76028
rect 58082 76014 58164 76028
rect 58372 76014 58454 76028
rect 16418 75966 58934 76014
rect 16418 75808 58934 75918
rect 16418 75712 58934 75760
rect 16898 75698 16980 75712
rect 17188 75698 17270 75712
rect 18146 75698 18228 75712
rect 18436 75698 18518 75712
rect 19394 75698 19476 75712
rect 19684 75698 19766 75712
rect 20642 75698 20724 75712
rect 20932 75698 21014 75712
rect 21890 75698 21972 75712
rect 22180 75698 22262 75712
rect 23138 75698 23220 75712
rect 23428 75698 23510 75712
rect 24386 75698 24468 75712
rect 24676 75698 24758 75712
rect 25634 75698 25716 75712
rect 25924 75698 26006 75712
rect 26882 75698 26964 75712
rect 27172 75698 27254 75712
rect 28130 75698 28212 75712
rect 28420 75698 28502 75712
rect 29378 75698 29460 75712
rect 29668 75698 29750 75712
rect 30626 75698 30708 75712
rect 30916 75698 30998 75712
rect 31874 75698 31956 75712
rect 32164 75698 32246 75712
rect 33122 75698 33204 75712
rect 33412 75698 33494 75712
rect 34370 75698 34452 75712
rect 34660 75698 34742 75712
rect 35618 75698 35700 75712
rect 35908 75698 35990 75712
rect 36866 75698 36948 75712
rect 37156 75698 37238 75712
rect 38114 75698 38196 75712
rect 38404 75698 38486 75712
rect 39362 75698 39444 75712
rect 39652 75698 39734 75712
rect 40610 75698 40692 75712
rect 40900 75698 40982 75712
rect 41858 75698 41940 75712
rect 42148 75698 42230 75712
rect 43106 75698 43188 75712
rect 43396 75698 43478 75712
rect 44354 75698 44436 75712
rect 44644 75698 44726 75712
rect 45602 75698 45684 75712
rect 45892 75698 45974 75712
rect 46850 75698 46932 75712
rect 47140 75698 47222 75712
rect 48098 75698 48180 75712
rect 48388 75698 48470 75712
rect 49346 75698 49428 75712
rect 49636 75698 49718 75712
rect 50594 75698 50676 75712
rect 50884 75698 50966 75712
rect 51842 75698 51924 75712
rect 52132 75698 52214 75712
rect 53090 75698 53172 75712
rect 53380 75698 53462 75712
rect 54338 75698 54420 75712
rect 54628 75698 54710 75712
rect 55586 75698 55668 75712
rect 55876 75698 55958 75712
rect 56834 75698 56916 75712
rect 57124 75698 57206 75712
rect 58082 75698 58164 75712
rect 58372 75698 58454 75712
rect 16418 75650 16864 75664
rect 17014 75650 17154 75664
rect 17304 75650 18112 75664
rect 18262 75650 18402 75664
rect 18552 75650 19360 75664
rect 19510 75650 19650 75664
rect 19800 75650 20608 75664
rect 20758 75650 20898 75664
rect 21048 75650 21856 75664
rect 22006 75650 22146 75664
rect 22296 75650 23104 75664
rect 23254 75650 23394 75664
rect 23544 75650 24352 75664
rect 24502 75650 24642 75664
rect 24792 75650 25600 75664
rect 25750 75650 25890 75664
rect 26040 75650 26848 75664
rect 26998 75650 27138 75664
rect 27288 75650 28096 75664
rect 28246 75650 28386 75664
rect 28536 75650 29344 75664
rect 29494 75650 29634 75664
rect 29784 75650 30592 75664
rect 30742 75650 30882 75664
rect 31032 75650 31840 75664
rect 31990 75650 32130 75664
rect 32280 75650 33088 75664
rect 33238 75650 33378 75664
rect 33528 75650 34336 75664
rect 34486 75650 34626 75664
rect 34776 75650 35584 75664
rect 35734 75650 35874 75664
rect 36024 75650 36832 75664
rect 36982 75650 37122 75664
rect 37272 75650 38080 75664
rect 38230 75650 38370 75664
rect 38520 75650 39328 75664
rect 39478 75650 39618 75664
rect 39768 75650 40576 75664
rect 40726 75650 40866 75664
rect 41016 75650 41824 75664
rect 41974 75650 42114 75664
rect 42264 75650 43072 75664
rect 43222 75650 43362 75664
rect 43512 75650 44320 75664
rect 44470 75650 44610 75664
rect 44760 75650 45568 75664
rect 45718 75650 45858 75664
rect 46008 75650 46816 75664
rect 46966 75650 47106 75664
rect 47256 75650 48064 75664
rect 48214 75650 48354 75664
rect 48504 75650 49312 75664
rect 49462 75650 49602 75664
rect 49752 75650 50560 75664
rect 50710 75650 50850 75664
rect 51000 75650 51808 75664
rect 51958 75650 52098 75664
rect 52248 75650 53056 75664
rect 53206 75650 53346 75664
rect 53496 75650 54304 75664
rect 54454 75650 54594 75664
rect 54744 75650 55552 75664
rect 55702 75650 55842 75664
rect 55992 75650 56800 75664
rect 56950 75650 57090 75664
rect 57240 75650 58048 75664
rect 58198 75650 58338 75664
rect 58488 75650 58934 75664
rect 16418 75602 58934 75650
rect 16418 75588 16864 75602
rect 17014 75588 17154 75602
rect 17304 75588 18112 75602
rect 18262 75588 18402 75602
rect 18552 75588 19360 75602
rect 19510 75588 19650 75602
rect 19800 75588 20608 75602
rect 20758 75588 20898 75602
rect 21048 75588 21856 75602
rect 22006 75588 22146 75602
rect 22296 75588 23104 75602
rect 23254 75588 23394 75602
rect 23544 75588 24352 75602
rect 24502 75588 24642 75602
rect 24792 75588 25600 75602
rect 25750 75588 25890 75602
rect 26040 75588 26848 75602
rect 26998 75588 27138 75602
rect 27288 75588 28096 75602
rect 28246 75588 28386 75602
rect 28536 75588 29344 75602
rect 29494 75588 29634 75602
rect 29784 75588 30592 75602
rect 30742 75588 30882 75602
rect 31032 75588 31840 75602
rect 31990 75588 32130 75602
rect 32280 75588 33088 75602
rect 33238 75588 33378 75602
rect 33528 75588 34336 75602
rect 34486 75588 34626 75602
rect 34776 75588 35584 75602
rect 35734 75588 35874 75602
rect 36024 75588 36832 75602
rect 36982 75588 37122 75602
rect 37272 75588 38080 75602
rect 38230 75588 38370 75602
rect 38520 75588 39328 75602
rect 39478 75588 39618 75602
rect 39768 75588 40576 75602
rect 40726 75588 40866 75602
rect 41016 75588 41824 75602
rect 41974 75588 42114 75602
rect 42264 75588 43072 75602
rect 43222 75588 43362 75602
rect 43512 75588 44320 75602
rect 44470 75588 44610 75602
rect 44760 75588 45568 75602
rect 45718 75588 45858 75602
rect 46008 75588 46816 75602
rect 46966 75588 47106 75602
rect 47256 75588 48064 75602
rect 48214 75588 48354 75602
rect 48504 75588 49312 75602
rect 49462 75588 49602 75602
rect 49752 75588 50560 75602
rect 50710 75588 50850 75602
rect 51000 75588 51808 75602
rect 51958 75588 52098 75602
rect 52248 75588 53056 75602
rect 53206 75588 53346 75602
rect 53496 75588 54304 75602
rect 54454 75588 54594 75602
rect 54744 75588 55552 75602
rect 55702 75588 55842 75602
rect 55992 75588 56800 75602
rect 56950 75588 57090 75602
rect 57240 75588 58048 75602
rect 58198 75588 58338 75602
rect 58488 75588 58934 75602
rect 16898 75540 16980 75554
rect 17188 75540 17270 75554
rect 18146 75540 18228 75554
rect 18436 75540 18518 75554
rect 19394 75540 19476 75554
rect 19684 75540 19766 75554
rect 20642 75540 20724 75554
rect 20932 75540 21014 75554
rect 21890 75540 21972 75554
rect 22180 75540 22262 75554
rect 23138 75540 23220 75554
rect 23428 75540 23510 75554
rect 24386 75540 24468 75554
rect 24676 75540 24758 75554
rect 25634 75540 25716 75554
rect 25924 75540 26006 75554
rect 26882 75540 26964 75554
rect 27172 75540 27254 75554
rect 28130 75540 28212 75554
rect 28420 75540 28502 75554
rect 29378 75540 29460 75554
rect 29668 75540 29750 75554
rect 30626 75540 30708 75554
rect 30916 75540 30998 75554
rect 31874 75540 31956 75554
rect 32164 75540 32246 75554
rect 33122 75540 33204 75554
rect 33412 75540 33494 75554
rect 34370 75540 34452 75554
rect 34660 75540 34742 75554
rect 35618 75540 35700 75554
rect 35908 75540 35990 75554
rect 36866 75540 36948 75554
rect 37156 75540 37238 75554
rect 38114 75540 38196 75554
rect 38404 75540 38486 75554
rect 39362 75540 39444 75554
rect 39652 75540 39734 75554
rect 40610 75540 40692 75554
rect 40900 75540 40982 75554
rect 41858 75540 41940 75554
rect 42148 75540 42230 75554
rect 43106 75540 43188 75554
rect 43396 75540 43478 75554
rect 44354 75540 44436 75554
rect 44644 75540 44726 75554
rect 45602 75540 45684 75554
rect 45892 75540 45974 75554
rect 46850 75540 46932 75554
rect 47140 75540 47222 75554
rect 48098 75540 48180 75554
rect 48388 75540 48470 75554
rect 49346 75540 49428 75554
rect 49636 75540 49718 75554
rect 50594 75540 50676 75554
rect 50884 75540 50966 75554
rect 51842 75540 51924 75554
rect 52132 75540 52214 75554
rect 53090 75540 53172 75554
rect 53380 75540 53462 75554
rect 54338 75540 54420 75554
rect 54628 75540 54710 75554
rect 55586 75540 55668 75554
rect 55876 75540 55958 75554
rect 56834 75540 56916 75554
rect 57124 75540 57206 75554
rect 58082 75540 58164 75554
rect 58372 75540 58454 75554
rect 16418 75492 58934 75540
rect 16418 75396 58934 75444
rect 16898 75382 16980 75396
rect 17188 75382 17270 75396
rect 18146 75382 18228 75396
rect 18436 75382 18518 75396
rect 19394 75382 19476 75396
rect 19684 75382 19766 75396
rect 20642 75382 20724 75396
rect 20932 75382 21014 75396
rect 21890 75382 21972 75396
rect 22180 75382 22262 75396
rect 23138 75382 23220 75396
rect 23428 75382 23510 75396
rect 24386 75382 24468 75396
rect 24676 75382 24758 75396
rect 25634 75382 25716 75396
rect 25924 75382 26006 75396
rect 26882 75382 26964 75396
rect 27172 75382 27254 75396
rect 28130 75382 28212 75396
rect 28420 75382 28502 75396
rect 29378 75382 29460 75396
rect 29668 75382 29750 75396
rect 30626 75382 30708 75396
rect 30916 75382 30998 75396
rect 31874 75382 31956 75396
rect 32164 75382 32246 75396
rect 33122 75382 33204 75396
rect 33412 75382 33494 75396
rect 34370 75382 34452 75396
rect 34660 75382 34742 75396
rect 35618 75382 35700 75396
rect 35908 75382 35990 75396
rect 36866 75382 36948 75396
rect 37156 75382 37238 75396
rect 38114 75382 38196 75396
rect 38404 75382 38486 75396
rect 39362 75382 39444 75396
rect 39652 75382 39734 75396
rect 40610 75382 40692 75396
rect 40900 75382 40982 75396
rect 41858 75382 41940 75396
rect 42148 75382 42230 75396
rect 43106 75382 43188 75396
rect 43396 75382 43478 75396
rect 44354 75382 44436 75396
rect 44644 75382 44726 75396
rect 45602 75382 45684 75396
rect 45892 75382 45974 75396
rect 46850 75382 46932 75396
rect 47140 75382 47222 75396
rect 48098 75382 48180 75396
rect 48388 75382 48470 75396
rect 49346 75382 49428 75396
rect 49636 75382 49718 75396
rect 50594 75382 50676 75396
rect 50884 75382 50966 75396
rect 51842 75382 51924 75396
rect 52132 75382 52214 75396
rect 53090 75382 53172 75396
rect 53380 75382 53462 75396
rect 54338 75382 54420 75396
rect 54628 75382 54710 75396
rect 55586 75382 55668 75396
rect 55876 75382 55958 75396
rect 56834 75382 56916 75396
rect 57124 75382 57206 75396
rect 58082 75382 58164 75396
rect 58372 75382 58454 75396
rect 16418 75334 16864 75348
rect 17014 75334 17154 75348
rect 17304 75334 18112 75348
rect 18262 75334 18402 75348
rect 18552 75334 19360 75348
rect 19510 75334 19650 75348
rect 19800 75334 20608 75348
rect 20758 75334 20898 75348
rect 21048 75334 21856 75348
rect 22006 75334 22146 75348
rect 22296 75334 23104 75348
rect 23254 75334 23394 75348
rect 23544 75334 24352 75348
rect 24502 75334 24642 75348
rect 24792 75334 25600 75348
rect 25750 75334 25890 75348
rect 26040 75334 26848 75348
rect 26998 75334 27138 75348
rect 27288 75334 28096 75348
rect 28246 75334 28386 75348
rect 28536 75334 29344 75348
rect 29494 75334 29634 75348
rect 29784 75334 30592 75348
rect 30742 75334 30882 75348
rect 31032 75334 31840 75348
rect 31990 75334 32130 75348
rect 32280 75334 33088 75348
rect 33238 75334 33378 75348
rect 33528 75334 34336 75348
rect 34486 75334 34626 75348
rect 34776 75334 35584 75348
rect 35734 75334 35874 75348
rect 36024 75334 36832 75348
rect 36982 75334 37122 75348
rect 37272 75334 38080 75348
rect 38230 75334 38370 75348
rect 38520 75334 39328 75348
rect 39478 75334 39618 75348
rect 39768 75334 40576 75348
rect 40726 75334 40866 75348
rect 41016 75334 41824 75348
rect 41974 75334 42114 75348
rect 42264 75334 43072 75348
rect 43222 75334 43362 75348
rect 43512 75334 44320 75348
rect 44470 75334 44610 75348
rect 44760 75334 45568 75348
rect 45718 75334 45858 75348
rect 46008 75334 46816 75348
rect 46966 75334 47106 75348
rect 47256 75334 48064 75348
rect 48214 75334 48354 75348
rect 48504 75334 49312 75348
rect 49462 75334 49602 75348
rect 49752 75334 50560 75348
rect 50710 75334 50850 75348
rect 51000 75334 51808 75348
rect 51958 75334 52098 75348
rect 52248 75334 53056 75348
rect 53206 75334 53346 75348
rect 53496 75334 54304 75348
rect 54454 75334 54594 75348
rect 54744 75334 55552 75348
rect 55702 75334 55842 75348
rect 55992 75334 56800 75348
rect 56950 75334 57090 75348
rect 57240 75334 58048 75348
rect 58198 75334 58338 75348
rect 58488 75334 58934 75348
rect 16418 75286 58934 75334
rect 16418 75272 16864 75286
rect 17014 75272 17154 75286
rect 17304 75272 18112 75286
rect 18262 75272 18402 75286
rect 18552 75272 19360 75286
rect 19510 75272 19650 75286
rect 19800 75272 20608 75286
rect 20758 75272 20898 75286
rect 21048 75272 21856 75286
rect 22006 75272 22146 75286
rect 22296 75272 23104 75286
rect 23254 75272 23394 75286
rect 23544 75272 24352 75286
rect 24502 75272 24642 75286
rect 24792 75272 25600 75286
rect 25750 75272 25890 75286
rect 26040 75272 26848 75286
rect 26998 75272 27138 75286
rect 27288 75272 28096 75286
rect 28246 75272 28386 75286
rect 28536 75272 29344 75286
rect 29494 75272 29634 75286
rect 29784 75272 30592 75286
rect 30742 75272 30882 75286
rect 31032 75272 31840 75286
rect 31990 75272 32130 75286
rect 32280 75272 33088 75286
rect 33238 75272 33378 75286
rect 33528 75272 34336 75286
rect 34486 75272 34626 75286
rect 34776 75272 35584 75286
rect 35734 75272 35874 75286
rect 36024 75272 36832 75286
rect 36982 75272 37122 75286
rect 37272 75272 38080 75286
rect 38230 75272 38370 75286
rect 38520 75272 39328 75286
rect 39478 75272 39618 75286
rect 39768 75272 40576 75286
rect 40726 75272 40866 75286
rect 41016 75272 41824 75286
rect 41974 75272 42114 75286
rect 42264 75272 43072 75286
rect 43222 75272 43362 75286
rect 43512 75272 44320 75286
rect 44470 75272 44610 75286
rect 44760 75272 45568 75286
rect 45718 75272 45858 75286
rect 46008 75272 46816 75286
rect 46966 75272 47106 75286
rect 47256 75272 48064 75286
rect 48214 75272 48354 75286
rect 48504 75272 49312 75286
rect 49462 75272 49602 75286
rect 49752 75272 50560 75286
rect 50710 75272 50850 75286
rect 51000 75272 51808 75286
rect 51958 75272 52098 75286
rect 52248 75272 53056 75286
rect 53206 75272 53346 75286
rect 53496 75272 54304 75286
rect 54454 75272 54594 75286
rect 54744 75272 55552 75286
rect 55702 75272 55842 75286
rect 55992 75272 56800 75286
rect 56950 75272 57090 75286
rect 57240 75272 58048 75286
rect 58198 75272 58338 75286
rect 58488 75272 58934 75286
rect 16898 75224 16980 75238
rect 17188 75224 17270 75238
rect 18146 75224 18228 75238
rect 18436 75224 18518 75238
rect 19394 75224 19476 75238
rect 19684 75224 19766 75238
rect 20642 75224 20724 75238
rect 20932 75224 21014 75238
rect 21890 75224 21972 75238
rect 22180 75224 22262 75238
rect 23138 75224 23220 75238
rect 23428 75224 23510 75238
rect 24386 75224 24468 75238
rect 24676 75224 24758 75238
rect 25634 75224 25716 75238
rect 25924 75224 26006 75238
rect 26882 75224 26964 75238
rect 27172 75224 27254 75238
rect 28130 75224 28212 75238
rect 28420 75224 28502 75238
rect 29378 75224 29460 75238
rect 29668 75224 29750 75238
rect 30626 75224 30708 75238
rect 30916 75224 30998 75238
rect 31874 75224 31956 75238
rect 32164 75224 32246 75238
rect 33122 75224 33204 75238
rect 33412 75224 33494 75238
rect 34370 75224 34452 75238
rect 34660 75224 34742 75238
rect 35618 75224 35700 75238
rect 35908 75224 35990 75238
rect 36866 75224 36948 75238
rect 37156 75224 37238 75238
rect 38114 75224 38196 75238
rect 38404 75224 38486 75238
rect 39362 75224 39444 75238
rect 39652 75224 39734 75238
rect 40610 75224 40692 75238
rect 40900 75224 40982 75238
rect 41858 75224 41940 75238
rect 42148 75224 42230 75238
rect 43106 75224 43188 75238
rect 43396 75224 43478 75238
rect 44354 75224 44436 75238
rect 44644 75224 44726 75238
rect 45602 75224 45684 75238
rect 45892 75224 45974 75238
rect 46850 75224 46932 75238
rect 47140 75224 47222 75238
rect 48098 75224 48180 75238
rect 48388 75224 48470 75238
rect 49346 75224 49428 75238
rect 49636 75224 49718 75238
rect 50594 75224 50676 75238
rect 50884 75224 50966 75238
rect 51842 75224 51924 75238
rect 52132 75224 52214 75238
rect 53090 75224 53172 75238
rect 53380 75224 53462 75238
rect 54338 75224 54420 75238
rect 54628 75224 54710 75238
rect 55586 75224 55668 75238
rect 55876 75224 55958 75238
rect 56834 75224 56916 75238
rect 57124 75224 57206 75238
rect 58082 75224 58164 75238
rect 58372 75224 58454 75238
rect 16418 75176 58934 75224
rect 16418 75018 58934 75128
rect 16418 74922 58934 74970
rect 16898 74908 16980 74922
rect 17188 74908 17270 74922
rect 18146 74908 18228 74922
rect 18436 74908 18518 74922
rect 19394 74908 19476 74922
rect 19684 74908 19766 74922
rect 20642 74908 20724 74922
rect 20932 74908 21014 74922
rect 21890 74908 21972 74922
rect 22180 74908 22262 74922
rect 23138 74908 23220 74922
rect 23428 74908 23510 74922
rect 24386 74908 24468 74922
rect 24676 74908 24758 74922
rect 25634 74908 25716 74922
rect 25924 74908 26006 74922
rect 26882 74908 26964 74922
rect 27172 74908 27254 74922
rect 28130 74908 28212 74922
rect 28420 74908 28502 74922
rect 29378 74908 29460 74922
rect 29668 74908 29750 74922
rect 30626 74908 30708 74922
rect 30916 74908 30998 74922
rect 31874 74908 31956 74922
rect 32164 74908 32246 74922
rect 33122 74908 33204 74922
rect 33412 74908 33494 74922
rect 34370 74908 34452 74922
rect 34660 74908 34742 74922
rect 35618 74908 35700 74922
rect 35908 74908 35990 74922
rect 36866 74908 36948 74922
rect 37156 74908 37238 74922
rect 38114 74908 38196 74922
rect 38404 74908 38486 74922
rect 39362 74908 39444 74922
rect 39652 74908 39734 74922
rect 40610 74908 40692 74922
rect 40900 74908 40982 74922
rect 41858 74908 41940 74922
rect 42148 74908 42230 74922
rect 43106 74908 43188 74922
rect 43396 74908 43478 74922
rect 44354 74908 44436 74922
rect 44644 74908 44726 74922
rect 45602 74908 45684 74922
rect 45892 74908 45974 74922
rect 46850 74908 46932 74922
rect 47140 74908 47222 74922
rect 48098 74908 48180 74922
rect 48388 74908 48470 74922
rect 49346 74908 49428 74922
rect 49636 74908 49718 74922
rect 50594 74908 50676 74922
rect 50884 74908 50966 74922
rect 51842 74908 51924 74922
rect 52132 74908 52214 74922
rect 53090 74908 53172 74922
rect 53380 74908 53462 74922
rect 54338 74908 54420 74922
rect 54628 74908 54710 74922
rect 55586 74908 55668 74922
rect 55876 74908 55958 74922
rect 56834 74908 56916 74922
rect 57124 74908 57206 74922
rect 58082 74908 58164 74922
rect 58372 74908 58454 74922
rect 16418 74860 16864 74874
rect 17014 74860 17154 74874
rect 17304 74860 18112 74874
rect 18262 74860 18402 74874
rect 18552 74860 19360 74874
rect 19510 74860 19650 74874
rect 19800 74860 20608 74874
rect 20758 74860 20898 74874
rect 21048 74860 21856 74874
rect 22006 74860 22146 74874
rect 22296 74860 23104 74874
rect 23254 74860 23394 74874
rect 23544 74860 24352 74874
rect 24502 74860 24642 74874
rect 24792 74860 25600 74874
rect 25750 74860 25890 74874
rect 26040 74860 26848 74874
rect 26998 74860 27138 74874
rect 27288 74860 28096 74874
rect 28246 74860 28386 74874
rect 28536 74860 29344 74874
rect 29494 74860 29634 74874
rect 29784 74860 30592 74874
rect 30742 74860 30882 74874
rect 31032 74860 31840 74874
rect 31990 74860 32130 74874
rect 32280 74860 33088 74874
rect 33238 74860 33378 74874
rect 33528 74860 34336 74874
rect 34486 74860 34626 74874
rect 34776 74860 35584 74874
rect 35734 74860 35874 74874
rect 36024 74860 36832 74874
rect 36982 74860 37122 74874
rect 37272 74860 38080 74874
rect 38230 74860 38370 74874
rect 38520 74860 39328 74874
rect 39478 74860 39618 74874
rect 39768 74860 40576 74874
rect 40726 74860 40866 74874
rect 41016 74860 41824 74874
rect 41974 74860 42114 74874
rect 42264 74860 43072 74874
rect 43222 74860 43362 74874
rect 43512 74860 44320 74874
rect 44470 74860 44610 74874
rect 44760 74860 45568 74874
rect 45718 74860 45858 74874
rect 46008 74860 46816 74874
rect 46966 74860 47106 74874
rect 47256 74860 48064 74874
rect 48214 74860 48354 74874
rect 48504 74860 49312 74874
rect 49462 74860 49602 74874
rect 49752 74860 50560 74874
rect 50710 74860 50850 74874
rect 51000 74860 51808 74874
rect 51958 74860 52098 74874
rect 52248 74860 53056 74874
rect 53206 74860 53346 74874
rect 53496 74860 54304 74874
rect 54454 74860 54594 74874
rect 54744 74860 55552 74874
rect 55702 74860 55842 74874
rect 55992 74860 56800 74874
rect 56950 74860 57090 74874
rect 57240 74860 58048 74874
rect 58198 74860 58338 74874
rect 58488 74860 58934 74874
rect 16418 74812 58934 74860
rect 16418 74798 16864 74812
rect 17014 74798 17154 74812
rect 17304 74798 18112 74812
rect 18262 74798 18402 74812
rect 18552 74798 19360 74812
rect 19510 74798 19650 74812
rect 19800 74798 20608 74812
rect 20758 74798 20898 74812
rect 21048 74798 21856 74812
rect 22006 74798 22146 74812
rect 22296 74798 23104 74812
rect 23254 74798 23394 74812
rect 23544 74798 24352 74812
rect 24502 74798 24642 74812
rect 24792 74798 25600 74812
rect 25750 74798 25890 74812
rect 26040 74798 26848 74812
rect 26998 74798 27138 74812
rect 27288 74798 28096 74812
rect 28246 74798 28386 74812
rect 28536 74798 29344 74812
rect 29494 74798 29634 74812
rect 29784 74798 30592 74812
rect 30742 74798 30882 74812
rect 31032 74798 31840 74812
rect 31990 74798 32130 74812
rect 32280 74798 33088 74812
rect 33238 74798 33378 74812
rect 33528 74798 34336 74812
rect 34486 74798 34626 74812
rect 34776 74798 35584 74812
rect 35734 74798 35874 74812
rect 36024 74798 36832 74812
rect 36982 74798 37122 74812
rect 37272 74798 38080 74812
rect 38230 74798 38370 74812
rect 38520 74798 39328 74812
rect 39478 74798 39618 74812
rect 39768 74798 40576 74812
rect 40726 74798 40866 74812
rect 41016 74798 41824 74812
rect 41974 74798 42114 74812
rect 42264 74798 43072 74812
rect 43222 74798 43362 74812
rect 43512 74798 44320 74812
rect 44470 74798 44610 74812
rect 44760 74798 45568 74812
rect 45718 74798 45858 74812
rect 46008 74798 46816 74812
rect 46966 74798 47106 74812
rect 47256 74798 48064 74812
rect 48214 74798 48354 74812
rect 48504 74798 49312 74812
rect 49462 74798 49602 74812
rect 49752 74798 50560 74812
rect 50710 74798 50850 74812
rect 51000 74798 51808 74812
rect 51958 74798 52098 74812
rect 52248 74798 53056 74812
rect 53206 74798 53346 74812
rect 53496 74798 54304 74812
rect 54454 74798 54594 74812
rect 54744 74798 55552 74812
rect 55702 74798 55842 74812
rect 55992 74798 56800 74812
rect 56950 74798 57090 74812
rect 57240 74798 58048 74812
rect 58198 74798 58338 74812
rect 58488 74798 58934 74812
rect 16898 74750 16980 74764
rect 17188 74750 17270 74764
rect 18146 74750 18228 74764
rect 18436 74750 18518 74764
rect 19394 74750 19476 74764
rect 19684 74750 19766 74764
rect 20642 74750 20724 74764
rect 20932 74750 21014 74764
rect 21890 74750 21972 74764
rect 22180 74750 22262 74764
rect 23138 74750 23220 74764
rect 23428 74750 23510 74764
rect 24386 74750 24468 74764
rect 24676 74750 24758 74764
rect 25634 74750 25716 74764
rect 25924 74750 26006 74764
rect 26882 74750 26964 74764
rect 27172 74750 27254 74764
rect 28130 74750 28212 74764
rect 28420 74750 28502 74764
rect 29378 74750 29460 74764
rect 29668 74750 29750 74764
rect 30626 74750 30708 74764
rect 30916 74750 30998 74764
rect 31874 74750 31956 74764
rect 32164 74750 32246 74764
rect 33122 74750 33204 74764
rect 33412 74750 33494 74764
rect 34370 74750 34452 74764
rect 34660 74750 34742 74764
rect 35618 74750 35700 74764
rect 35908 74750 35990 74764
rect 36866 74750 36948 74764
rect 37156 74750 37238 74764
rect 38114 74750 38196 74764
rect 38404 74750 38486 74764
rect 39362 74750 39444 74764
rect 39652 74750 39734 74764
rect 40610 74750 40692 74764
rect 40900 74750 40982 74764
rect 41858 74750 41940 74764
rect 42148 74750 42230 74764
rect 43106 74750 43188 74764
rect 43396 74750 43478 74764
rect 44354 74750 44436 74764
rect 44644 74750 44726 74764
rect 45602 74750 45684 74764
rect 45892 74750 45974 74764
rect 46850 74750 46932 74764
rect 47140 74750 47222 74764
rect 48098 74750 48180 74764
rect 48388 74750 48470 74764
rect 49346 74750 49428 74764
rect 49636 74750 49718 74764
rect 50594 74750 50676 74764
rect 50884 74750 50966 74764
rect 51842 74750 51924 74764
rect 52132 74750 52214 74764
rect 53090 74750 53172 74764
rect 53380 74750 53462 74764
rect 54338 74750 54420 74764
rect 54628 74750 54710 74764
rect 55586 74750 55668 74764
rect 55876 74750 55958 74764
rect 56834 74750 56916 74764
rect 57124 74750 57206 74764
rect 58082 74750 58164 74764
rect 58372 74750 58454 74764
rect 16418 74702 58934 74750
rect 16418 74606 58934 74654
rect 16898 74592 16980 74606
rect 17188 74592 17270 74606
rect 18146 74592 18228 74606
rect 18436 74592 18518 74606
rect 19394 74592 19476 74606
rect 19684 74592 19766 74606
rect 20642 74592 20724 74606
rect 20932 74592 21014 74606
rect 21890 74592 21972 74606
rect 22180 74592 22262 74606
rect 23138 74592 23220 74606
rect 23428 74592 23510 74606
rect 24386 74592 24468 74606
rect 24676 74592 24758 74606
rect 25634 74592 25716 74606
rect 25924 74592 26006 74606
rect 26882 74592 26964 74606
rect 27172 74592 27254 74606
rect 28130 74592 28212 74606
rect 28420 74592 28502 74606
rect 29378 74592 29460 74606
rect 29668 74592 29750 74606
rect 30626 74592 30708 74606
rect 30916 74592 30998 74606
rect 31874 74592 31956 74606
rect 32164 74592 32246 74606
rect 33122 74592 33204 74606
rect 33412 74592 33494 74606
rect 34370 74592 34452 74606
rect 34660 74592 34742 74606
rect 35618 74592 35700 74606
rect 35908 74592 35990 74606
rect 36866 74592 36948 74606
rect 37156 74592 37238 74606
rect 38114 74592 38196 74606
rect 38404 74592 38486 74606
rect 39362 74592 39444 74606
rect 39652 74592 39734 74606
rect 40610 74592 40692 74606
rect 40900 74592 40982 74606
rect 41858 74592 41940 74606
rect 42148 74592 42230 74606
rect 43106 74592 43188 74606
rect 43396 74592 43478 74606
rect 44354 74592 44436 74606
rect 44644 74592 44726 74606
rect 45602 74592 45684 74606
rect 45892 74592 45974 74606
rect 46850 74592 46932 74606
rect 47140 74592 47222 74606
rect 48098 74592 48180 74606
rect 48388 74592 48470 74606
rect 49346 74592 49428 74606
rect 49636 74592 49718 74606
rect 50594 74592 50676 74606
rect 50884 74592 50966 74606
rect 51842 74592 51924 74606
rect 52132 74592 52214 74606
rect 53090 74592 53172 74606
rect 53380 74592 53462 74606
rect 54338 74592 54420 74606
rect 54628 74592 54710 74606
rect 55586 74592 55668 74606
rect 55876 74592 55958 74606
rect 56834 74592 56916 74606
rect 57124 74592 57206 74606
rect 58082 74592 58164 74606
rect 58372 74592 58454 74606
rect 16418 74544 16864 74558
rect 17014 74544 17154 74558
rect 17304 74544 18112 74558
rect 18262 74544 18402 74558
rect 18552 74544 19360 74558
rect 19510 74544 19650 74558
rect 19800 74544 20608 74558
rect 20758 74544 20898 74558
rect 21048 74544 21856 74558
rect 22006 74544 22146 74558
rect 22296 74544 23104 74558
rect 23254 74544 23394 74558
rect 23544 74544 24352 74558
rect 24502 74544 24642 74558
rect 24792 74544 25600 74558
rect 25750 74544 25890 74558
rect 26040 74544 26848 74558
rect 26998 74544 27138 74558
rect 27288 74544 28096 74558
rect 28246 74544 28386 74558
rect 28536 74544 29344 74558
rect 29494 74544 29634 74558
rect 29784 74544 30592 74558
rect 30742 74544 30882 74558
rect 31032 74544 31840 74558
rect 31990 74544 32130 74558
rect 32280 74544 33088 74558
rect 33238 74544 33378 74558
rect 33528 74544 34336 74558
rect 34486 74544 34626 74558
rect 34776 74544 35584 74558
rect 35734 74544 35874 74558
rect 36024 74544 36832 74558
rect 36982 74544 37122 74558
rect 37272 74544 38080 74558
rect 38230 74544 38370 74558
rect 38520 74544 39328 74558
rect 39478 74544 39618 74558
rect 39768 74544 40576 74558
rect 40726 74544 40866 74558
rect 41016 74544 41824 74558
rect 41974 74544 42114 74558
rect 42264 74544 43072 74558
rect 43222 74544 43362 74558
rect 43512 74544 44320 74558
rect 44470 74544 44610 74558
rect 44760 74544 45568 74558
rect 45718 74544 45858 74558
rect 46008 74544 46816 74558
rect 46966 74544 47106 74558
rect 47256 74544 48064 74558
rect 48214 74544 48354 74558
rect 48504 74544 49312 74558
rect 49462 74544 49602 74558
rect 49752 74544 50560 74558
rect 50710 74544 50850 74558
rect 51000 74544 51808 74558
rect 51958 74544 52098 74558
rect 52248 74544 53056 74558
rect 53206 74544 53346 74558
rect 53496 74544 54304 74558
rect 54454 74544 54594 74558
rect 54744 74544 55552 74558
rect 55702 74544 55842 74558
rect 55992 74544 56800 74558
rect 56950 74544 57090 74558
rect 57240 74544 58048 74558
rect 58198 74544 58338 74558
rect 58488 74544 58934 74558
rect 16418 74496 58934 74544
rect 16418 74482 16864 74496
rect 17014 74482 17154 74496
rect 17304 74482 18112 74496
rect 18262 74482 18402 74496
rect 18552 74482 19360 74496
rect 19510 74482 19650 74496
rect 19800 74482 20608 74496
rect 20758 74482 20898 74496
rect 21048 74482 21856 74496
rect 22006 74482 22146 74496
rect 22296 74482 23104 74496
rect 23254 74482 23394 74496
rect 23544 74482 24352 74496
rect 24502 74482 24642 74496
rect 24792 74482 25600 74496
rect 25750 74482 25890 74496
rect 26040 74482 26848 74496
rect 26998 74482 27138 74496
rect 27288 74482 28096 74496
rect 28246 74482 28386 74496
rect 28536 74482 29344 74496
rect 29494 74482 29634 74496
rect 29784 74482 30592 74496
rect 30742 74482 30882 74496
rect 31032 74482 31840 74496
rect 31990 74482 32130 74496
rect 32280 74482 33088 74496
rect 33238 74482 33378 74496
rect 33528 74482 34336 74496
rect 34486 74482 34626 74496
rect 34776 74482 35584 74496
rect 35734 74482 35874 74496
rect 36024 74482 36832 74496
rect 36982 74482 37122 74496
rect 37272 74482 38080 74496
rect 38230 74482 38370 74496
rect 38520 74482 39328 74496
rect 39478 74482 39618 74496
rect 39768 74482 40576 74496
rect 40726 74482 40866 74496
rect 41016 74482 41824 74496
rect 41974 74482 42114 74496
rect 42264 74482 43072 74496
rect 43222 74482 43362 74496
rect 43512 74482 44320 74496
rect 44470 74482 44610 74496
rect 44760 74482 45568 74496
rect 45718 74482 45858 74496
rect 46008 74482 46816 74496
rect 46966 74482 47106 74496
rect 47256 74482 48064 74496
rect 48214 74482 48354 74496
rect 48504 74482 49312 74496
rect 49462 74482 49602 74496
rect 49752 74482 50560 74496
rect 50710 74482 50850 74496
rect 51000 74482 51808 74496
rect 51958 74482 52098 74496
rect 52248 74482 53056 74496
rect 53206 74482 53346 74496
rect 53496 74482 54304 74496
rect 54454 74482 54594 74496
rect 54744 74482 55552 74496
rect 55702 74482 55842 74496
rect 55992 74482 56800 74496
rect 56950 74482 57090 74496
rect 57240 74482 58048 74496
rect 58198 74482 58338 74496
rect 58488 74482 58934 74496
rect 16898 74434 16980 74448
rect 17188 74434 17270 74448
rect 18146 74434 18228 74448
rect 18436 74434 18518 74448
rect 19394 74434 19476 74448
rect 19684 74434 19766 74448
rect 20642 74434 20724 74448
rect 20932 74434 21014 74448
rect 21890 74434 21972 74448
rect 22180 74434 22262 74448
rect 23138 74434 23220 74448
rect 23428 74434 23510 74448
rect 24386 74434 24468 74448
rect 24676 74434 24758 74448
rect 25634 74434 25716 74448
rect 25924 74434 26006 74448
rect 26882 74434 26964 74448
rect 27172 74434 27254 74448
rect 28130 74434 28212 74448
rect 28420 74434 28502 74448
rect 29378 74434 29460 74448
rect 29668 74434 29750 74448
rect 30626 74434 30708 74448
rect 30916 74434 30998 74448
rect 31874 74434 31956 74448
rect 32164 74434 32246 74448
rect 33122 74434 33204 74448
rect 33412 74434 33494 74448
rect 34370 74434 34452 74448
rect 34660 74434 34742 74448
rect 35618 74434 35700 74448
rect 35908 74434 35990 74448
rect 36866 74434 36948 74448
rect 37156 74434 37238 74448
rect 38114 74434 38196 74448
rect 38404 74434 38486 74448
rect 39362 74434 39444 74448
rect 39652 74434 39734 74448
rect 40610 74434 40692 74448
rect 40900 74434 40982 74448
rect 41858 74434 41940 74448
rect 42148 74434 42230 74448
rect 43106 74434 43188 74448
rect 43396 74434 43478 74448
rect 44354 74434 44436 74448
rect 44644 74434 44726 74448
rect 45602 74434 45684 74448
rect 45892 74434 45974 74448
rect 46850 74434 46932 74448
rect 47140 74434 47222 74448
rect 48098 74434 48180 74448
rect 48388 74434 48470 74448
rect 49346 74434 49428 74448
rect 49636 74434 49718 74448
rect 50594 74434 50676 74448
rect 50884 74434 50966 74448
rect 51842 74434 51924 74448
rect 52132 74434 52214 74448
rect 53090 74434 53172 74448
rect 53380 74434 53462 74448
rect 54338 74434 54420 74448
rect 54628 74434 54710 74448
rect 55586 74434 55668 74448
rect 55876 74434 55958 74448
rect 56834 74434 56916 74448
rect 57124 74434 57206 74448
rect 58082 74434 58164 74448
rect 58372 74434 58454 74448
rect 16418 74386 58934 74434
rect 16418 74228 58934 74338
rect 16418 74132 58934 74180
rect 16898 74118 16980 74132
rect 17188 74118 17270 74132
rect 18146 74118 18228 74132
rect 18436 74118 18518 74132
rect 19394 74118 19476 74132
rect 19684 74118 19766 74132
rect 20642 74118 20724 74132
rect 20932 74118 21014 74132
rect 21890 74118 21972 74132
rect 22180 74118 22262 74132
rect 23138 74118 23220 74132
rect 23428 74118 23510 74132
rect 24386 74118 24468 74132
rect 24676 74118 24758 74132
rect 25634 74118 25716 74132
rect 25924 74118 26006 74132
rect 26882 74118 26964 74132
rect 27172 74118 27254 74132
rect 28130 74118 28212 74132
rect 28420 74118 28502 74132
rect 29378 74118 29460 74132
rect 29668 74118 29750 74132
rect 30626 74118 30708 74132
rect 30916 74118 30998 74132
rect 31874 74118 31956 74132
rect 32164 74118 32246 74132
rect 33122 74118 33204 74132
rect 33412 74118 33494 74132
rect 34370 74118 34452 74132
rect 34660 74118 34742 74132
rect 35618 74118 35700 74132
rect 35908 74118 35990 74132
rect 36866 74118 36948 74132
rect 37156 74118 37238 74132
rect 38114 74118 38196 74132
rect 38404 74118 38486 74132
rect 39362 74118 39444 74132
rect 39652 74118 39734 74132
rect 40610 74118 40692 74132
rect 40900 74118 40982 74132
rect 41858 74118 41940 74132
rect 42148 74118 42230 74132
rect 43106 74118 43188 74132
rect 43396 74118 43478 74132
rect 44354 74118 44436 74132
rect 44644 74118 44726 74132
rect 45602 74118 45684 74132
rect 45892 74118 45974 74132
rect 46850 74118 46932 74132
rect 47140 74118 47222 74132
rect 48098 74118 48180 74132
rect 48388 74118 48470 74132
rect 49346 74118 49428 74132
rect 49636 74118 49718 74132
rect 50594 74118 50676 74132
rect 50884 74118 50966 74132
rect 51842 74118 51924 74132
rect 52132 74118 52214 74132
rect 53090 74118 53172 74132
rect 53380 74118 53462 74132
rect 54338 74118 54420 74132
rect 54628 74118 54710 74132
rect 55586 74118 55668 74132
rect 55876 74118 55958 74132
rect 56834 74118 56916 74132
rect 57124 74118 57206 74132
rect 58082 74118 58164 74132
rect 58372 74118 58454 74132
rect 16418 74070 16864 74084
rect 17014 74070 17154 74084
rect 17304 74070 18112 74084
rect 18262 74070 18402 74084
rect 18552 74070 19360 74084
rect 19510 74070 19650 74084
rect 19800 74070 20608 74084
rect 20758 74070 20898 74084
rect 21048 74070 21856 74084
rect 22006 74070 22146 74084
rect 22296 74070 23104 74084
rect 23254 74070 23394 74084
rect 23544 74070 24352 74084
rect 24502 74070 24642 74084
rect 24792 74070 25600 74084
rect 25750 74070 25890 74084
rect 26040 74070 26848 74084
rect 26998 74070 27138 74084
rect 27288 74070 28096 74084
rect 28246 74070 28386 74084
rect 28536 74070 29344 74084
rect 29494 74070 29634 74084
rect 29784 74070 30592 74084
rect 30742 74070 30882 74084
rect 31032 74070 31840 74084
rect 31990 74070 32130 74084
rect 32280 74070 33088 74084
rect 33238 74070 33378 74084
rect 33528 74070 34336 74084
rect 34486 74070 34626 74084
rect 34776 74070 35584 74084
rect 35734 74070 35874 74084
rect 36024 74070 36832 74084
rect 36982 74070 37122 74084
rect 37272 74070 38080 74084
rect 38230 74070 38370 74084
rect 38520 74070 39328 74084
rect 39478 74070 39618 74084
rect 39768 74070 40576 74084
rect 40726 74070 40866 74084
rect 41016 74070 41824 74084
rect 41974 74070 42114 74084
rect 42264 74070 43072 74084
rect 43222 74070 43362 74084
rect 43512 74070 44320 74084
rect 44470 74070 44610 74084
rect 44760 74070 45568 74084
rect 45718 74070 45858 74084
rect 46008 74070 46816 74084
rect 46966 74070 47106 74084
rect 47256 74070 48064 74084
rect 48214 74070 48354 74084
rect 48504 74070 49312 74084
rect 49462 74070 49602 74084
rect 49752 74070 50560 74084
rect 50710 74070 50850 74084
rect 51000 74070 51808 74084
rect 51958 74070 52098 74084
rect 52248 74070 53056 74084
rect 53206 74070 53346 74084
rect 53496 74070 54304 74084
rect 54454 74070 54594 74084
rect 54744 74070 55552 74084
rect 55702 74070 55842 74084
rect 55992 74070 56800 74084
rect 56950 74070 57090 74084
rect 57240 74070 58048 74084
rect 58198 74070 58338 74084
rect 58488 74070 58934 74084
rect 16418 74022 58934 74070
rect 16418 74008 16864 74022
rect 17014 74008 17154 74022
rect 17304 74008 18112 74022
rect 18262 74008 18402 74022
rect 18552 74008 19360 74022
rect 19510 74008 19650 74022
rect 19800 74008 20608 74022
rect 20758 74008 20898 74022
rect 21048 74008 21856 74022
rect 22006 74008 22146 74022
rect 22296 74008 23104 74022
rect 23254 74008 23394 74022
rect 23544 74008 24352 74022
rect 24502 74008 24642 74022
rect 24792 74008 25600 74022
rect 25750 74008 25890 74022
rect 26040 74008 26848 74022
rect 26998 74008 27138 74022
rect 27288 74008 28096 74022
rect 28246 74008 28386 74022
rect 28536 74008 29344 74022
rect 29494 74008 29634 74022
rect 29784 74008 30592 74022
rect 30742 74008 30882 74022
rect 31032 74008 31840 74022
rect 31990 74008 32130 74022
rect 32280 74008 33088 74022
rect 33238 74008 33378 74022
rect 33528 74008 34336 74022
rect 34486 74008 34626 74022
rect 34776 74008 35584 74022
rect 35734 74008 35874 74022
rect 36024 74008 36832 74022
rect 36982 74008 37122 74022
rect 37272 74008 38080 74022
rect 38230 74008 38370 74022
rect 38520 74008 39328 74022
rect 39478 74008 39618 74022
rect 39768 74008 40576 74022
rect 40726 74008 40866 74022
rect 41016 74008 41824 74022
rect 41974 74008 42114 74022
rect 42264 74008 43072 74022
rect 43222 74008 43362 74022
rect 43512 74008 44320 74022
rect 44470 74008 44610 74022
rect 44760 74008 45568 74022
rect 45718 74008 45858 74022
rect 46008 74008 46816 74022
rect 46966 74008 47106 74022
rect 47256 74008 48064 74022
rect 48214 74008 48354 74022
rect 48504 74008 49312 74022
rect 49462 74008 49602 74022
rect 49752 74008 50560 74022
rect 50710 74008 50850 74022
rect 51000 74008 51808 74022
rect 51958 74008 52098 74022
rect 52248 74008 53056 74022
rect 53206 74008 53346 74022
rect 53496 74008 54304 74022
rect 54454 74008 54594 74022
rect 54744 74008 55552 74022
rect 55702 74008 55842 74022
rect 55992 74008 56800 74022
rect 56950 74008 57090 74022
rect 57240 74008 58048 74022
rect 58198 74008 58338 74022
rect 58488 74008 58934 74022
rect 16898 73960 16980 73974
rect 17188 73960 17270 73974
rect 18146 73960 18228 73974
rect 18436 73960 18518 73974
rect 19394 73960 19476 73974
rect 19684 73960 19766 73974
rect 20642 73960 20724 73974
rect 20932 73960 21014 73974
rect 21890 73960 21972 73974
rect 22180 73960 22262 73974
rect 23138 73960 23220 73974
rect 23428 73960 23510 73974
rect 24386 73960 24468 73974
rect 24676 73960 24758 73974
rect 25634 73960 25716 73974
rect 25924 73960 26006 73974
rect 26882 73960 26964 73974
rect 27172 73960 27254 73974
rect 28130 73960 28212 73974
rect 28420 73960 28502 73974
rect 29378 73960 29460 73974
rect 29668 73960 29750 73974
rect 30626 73960 30708 73974
rect 30916 73960 30998 73974
rect 31874 73960 31956 73974
rect 32164 73960 32246 73974
rect 33122 73960 33204 73974
rect 33412 73960 33494 73974
rect 34370 73960 34452 73974
rect 34660 73960 34742 73974
rect 35618 73960 35700 73974
rect 35908 73960 35990 73974
rect 36866 73960 36948 73974
rect 37156 73960 37238 73974
rect 38114 73960 38196 73974
rect 38404 73960 38486 73974
rect 39362 73960 39444 73974
rect 39652 73960 39734 73974
rect 40610 73960 40692 73974
rect 40900 73960 40982 73974
rect 41858 73960 41940 73974
rect 42148 73960 42230 73974
rect 43106 73960 43188 73974
rect 43396 73960 43478 73974
rect 44354 73960 44436 73974
rect 44644 73960 44726 73974
rect 45602 73960 45684 73974
rect 45892 73960 45974 73974
rect 46850 73960 46932 73974
rect 47140 73960 47222 73974
rect 48098 73960 48180 73974
rect 48388 73960 48470 73974
rect 49346 73960 49428 73974
rect 49636 73960 49718 73974
rect 50594 73960 50676 73974
rect 50884 73960 50966 73974
rect 51842 73960 51924 73974
rect 52132 73960 52214 73974
rect 53090 73960 53172 73974
rect 53380 73960 53462 73974
rect 54338 73960 54420 73974
rect 54628 73960 54710 73974
rect 55586 73960 55668 73974
rect 55876 73960 55958 73974
rect 56834 73960 56916 73974
rect 57124 73960 57206 73974
rect 58082 73960 58164 73974
rect 58372 73960 58454 73974
rect 16418 73912 58934 73960
rect 16418 73816 58934 73864
rect 16898 73802 16980 73816
rect 17188 73802 17270 73816
rect 18146 73802 18228 73816
rect 18436 73802 18518 73816
rect 19394 73802 19476 73816
rect 19684 73802 19766 73816
rect 20642 73802 20724 73816
rect 20932 73802 21014 73816
rect 21890 73802 21972 73816
rect 22180 73802 22262 73816
rect 23138 73802 23220 73816
rect 23428 73802 23510 73816
rect 24386 73802 24468 73816
rect 24676 73802 24758 73816
rect 25634 73802 25716 73816
rect 25924 73802 26006 73816
rect 26882 73802 26964 73816
rect 27172 73802 27254 73816
rect 28130 73802 28212 73816
rect 28420 73802 28502 73816
rect 29378 73802 29460 73816
rect 29668 73802 29750 73816
rect 30626 73802 30708 73816
rect 30916 73802 30998 73816
rect 31874 73802 31956 73816
rect 32164 73802 32246 73816
rect 33122 73802 33204 73816
rect 33412 73802 33494 73816
rect 34370 73802 34452 73816
rect 34660 73802 34742 73816
rect 35618 73802 35700 73816
rect 35908 73802 35990 73816
rect 36866 73802 36948 73816
rect 37156 73802 37238 73816
rect 38114 73802 38196 73816
rect 38404 73802 38486 73816
rect 39362 73802 39444 73816
rect 39652 73802 39734 73816
rect 40610 73802 40692 73816
rect 40900 73802 40982 73816
rect 41858 73802 41940 73816
rect 42148 73802 42230 73816
rect 43106 73802 43188 73816
rect 43396 73802 43478 73816
rect 44354 73802 44436 73816
rect 44644 73802 44726 73816
rect 45602 73802 45684 73816
rect 45892 73802 45974 73816
rect 46850 73802 46932 73816
rect 47140 73802 47222 73816
rect 48098 73802 48180 73816
rect 48388 73802 48470 73816
rect 49346 73802 49428 73816
rect 49636 73802 49718 73816
rect 50594 73802 50676 73816
rect 50884 73802 50966 73816
rect 51842 73802 51924 73816
rect 52132 73802 52214 73816
rect 53090 73802 53172 73816
rect 53380 73802 53462 73816
rect 54338 73802 54420 73816
rect 54628 73802 54710 73816
rect 55586 73802 55668 73816
rect 55876 73802 55958 73816
rect 56834 73802 56916 73816
rect 57124 73802 57206 73816
rect 58082 73802 58164 73816
rect 58372 73802 58454 73816
rect 16418 73754 16864 73768
rect 17014 73754 17154 73768
rect 17304 73754 18112 73768
rect 18262 73754 18402 73768
rect 18552 73754 19360 73768
rect 19510 73754 19650 73768
rect 19800 73754 20608 73768
rect 20758 73754 20898 73768
rect 21048 73754 21856 73768
rect 22006 73754 22146 73768
rect 22296 73754 23104 73768
rect 23254 73754 23394 73768
rect 23544 73754 24352 73768
rect 24502 73754 24642 73768
rect 24792 73754 25600 73768
rect 25750 73754 25890 73768
rect 26040 73754 26848 73768
rect 26998 73754 27138 73768
rect 27288 73754 28096 73768
rect 28246 73754 28386 73768
rect 28536 73754 29344 73768
rect 29494 73754 29634 73768
rect 29784 73754 30592 73768
rect 30742 73754 30882 73768
rect 31032 73754 31840 73768
rect 31990 73754 32130 73768
rect 32280 73754 33088 73768
rect 33238 73754 33378 73768
rect 33528 73754 34336 73768
rect 34486 73754 34626 73768
rect 34776 73754 35584 73768
rect 35734 73754 35874 73768
rect 36024 73754 36832 73768
rect 36982 73754 37122 73768
rect 37272 73754 38080 73768
rect 38230 73754 38370 73768
rect 38520 73754 39328 73768
rect 39478 73754 39618 73768
rect 39768 73754 40576 73768
rect 40726 73754 40866 73768
rect 41016 73754 41824 73768
rect 41974 73754 42114 73768
rect 42264 73754 43072 73768
rect 43222 73754 43362 73768
rect 43512 73754 44320 73768
rect 44470 73754 44610 73768
rect 44760 73754 45568 73768
rect 45718 73754 45858 73768
rect 46008 73754 46816 73768
rect 46966 73754 47106 73768
rect 47256 73754 48064 73768
rect 48214 73754 48354 73768
rect 48504 73754 49312 73768
rect 49462 73754 49602 73768
rect 49752 73754 50560 73768
rect 50710 73754 50850 73768
rect 51000 73754 51808 73768
rect 51958 73754 52098 73768
rect 52248 73754 53056 73768
rect 53206 73754 53346 73768
rect 53496 73754 54304 73768
rect 54454 73754 54594 73768
rect 54744 73754 55552 73768
rect 55702 73754 55842 73768
rect 55992 73754 56800 73768
rect 56950 73754 57090 73768
rect 57240 73754 58048 73768
rect 58198 73754 58338 73768
rect 58488 73754 58934 73768
rect 16418 73706 58934 73754
rect 16418 73692 16864 73706
rect 17014 73692 17154 73706
rect 17304 73692 18112 73706
rect 18262 73692 18402 73706
rect 18552 73692 19360 73706
rect 19510 73692 19650 73706
rect 19800 73692 20608 73706
rect 20758 73692 20898 73706
rect 21048 73692 21856 73706
rect 22006 73692 22146 73706
rect 22296 73692 23104 73706
rect 23254 73692 23394 73706
rect 23544 73692 24352 73706
rect 24502 73692 24642 73706
rect 24792 73692 25600 73706
rect 25750 73692 25890 73706
rect 26040 73692 26848 73706
rect 26998 73692 27138 73706
rect 27288 73692 28096 73706
rect 28246 73692 28386 73706
rect 28536 73692 29344 73706
rect 29494 73692 29634 73706
rect 29784 73692 30592 73706
rect 30742 73692 30882 73706
rect 31032 73692 31840 73706
rect 31990 73692 32130 73706
rect 32280 73692 33088 73706
rect 33238 73692 33378 73706
rect 33528 73692 34336 73706
rect 34486 73692 34626 73706
rect 34776 73692 35584 73706
rect 35734 73692 35874 73706
rect 36024 73692 36832 73706
rect 36982 73692 37122 73706
rect 37272 73692 38080 73706
rect 38230 73692 38370 73706
rect 38520 73692 39328 73706
rect 39478 73692 39618 73706
rect 39768 73692 40576 73706
rect 40726 73692 40866 73706
rect 41016 73692 41824 73706
rect 41974 73692 42114 73706
rect 42264 73692 43072 73706
rect 43222 73692 43362 73706
rect 43512 73692 44320 73706
rect 44470 73692 44610 73706
rect 44760 73692 45568 73706
rect 45718 73692 45858 73706
rect 46008 73692 46816 73706
rect 46966 73692 47106 73706
rect 47256 73692 48064 73706
rect 48214 73692 48354 73706
rect 48504 73692 49312 73706
rect 49462 73692 49602 73706
rect 49752 73692 50560 73706
rect 50710 73692 50850 73706
rect 51000 73692 51808 73706
rect 51958 73692 52098 73706
rect 52248 73692 53056 73706
rect 53206 73692 53346 73706
rect 53496 73692 54304 73706
rect 54454 73692 54594 73706
rect 54744 73692 55552 73706
rect 55702 73692 55842 73706
rect 55992 73692 56800 73706
rect 56950 73692 57090 73706
rect 57240 73692 58048 73706
rect 58198 73692 58338 73706
rect 58488 73692 58934 73706
rect 16898 73644 16980 73658
rect 17188 73644 17270 73658
rect 18146 73644 18228 73658
rect 18436 73644 18518 73658
rect 19394 73644 19476 73658
rect 19684 73644 19766 73658
rect 20642 73644 20724 73658
rect 20932 73644 21014 73658
rect 21890 73644 21972 73658
rect 22180 73644 22262 73658
rect 23138 73644 23220 73658
rect 23428 73644 23510 73658
rect 24386 73644 24468 73658
rect 24676 73644 24758 73658
rect 25634 73644 25716 73658
rect 25924 73644 26006 73658
rect 26882 73644 26964 73658
rect 27172 73644 27254 73658
rect 28130 73644 28212 73658
rect 28420 73644 28502 73658
rect 29378 73644 29460 73658
rect 29668 73644 29750 73658
rect 30626 73644 30708 73658
rect 30916 73644 30998 73658
rect 31874 73644 31956 73658
rect 32164 73644 32246 73658
rect 33122 73644 33204 73658
rect 33412 73644 33494 73658
rect 34370 73644 34452 73658
rect 34660 73644 34742 73658
rect 35618 73644 35700 73658
rect 35908 73644 35990 73658
rect 36866 73644 36948 73658
rect 37156 73644 37238 73658
rect 38114 73644 38196 73658
rect 38404 73644 38486 73658
rect 39362 73644 39444 73658
rect 39652 73644 39734 73658
rect 40610 73644 40692 73658
rect 40900 73644 40982 73658
rect 41858 73644 41940 73658
rect 42148 73644 42230 73658
rect 43106 73644 43188 73658
rect 43396 73644 43478 73658
rect 44354 73644 44436 73658
rect 44644 73644 44726 73658
rect 45602 73644 45684 73658
rect 45892 73644 45974 73658
rect 46850 73644 46932 73658
rect 47140 73644 47222 73658
rect 48098 73644 48180 73658
rect 48388 73644 48470 73658
rect 49346 73644 49428 73658
rect 49636 73644 49718 73658
rect 50594 73644 50676 73658
rect 50884 73644 50966 73658
rect 51842 73644 51924 73658
rect 52132 73644 52214 73658
rect 53090 73644 53172 73658
rect 53380 73644 53462 73658
rect 54338 73644 54420 73658
rect 54628 73644 54710 73658
rect 55586 73644 55668 73658
rect 55876 73644 55958 73658
rect 56834 73644 56916 73658
rect 57124 73644 57206 73658
rect 58082 73644 58164 73658
rect 58372 73644 58454 73658
rect 16418 73596 58934 73644
rect 16418 73438 58934 73548
rect 16418 73342 58934 73390
rect 16898 73328 16980 73342
rect 17188 73328 17270 73342
rect 18146 73328 18228 73342
rect 18436 73328 18518 73342
rect 19394 73328 19476 73342
rect 19684 73328 19766 73342
rect 20642 73328 20724 73342
rect 20932 73328 21014 73342
rect 21890 73328 21972 73342
rect 22180 73328 22262 73342
rect 23138 73328 23220 73342
rect 23428 73328 23510 73342
rect 24386 73328 24468 73342
rect 24676 73328 24758 73342
rect 25634 73328 25716 73342
rect 25924 73328 26006 73342
rect 26882 73328 26964 73342
rect 27172 73328 27254 73342
rect 28130 73328 28212 73342
rect 28420 73328 28502 73342
rect 29378 73328 29460 73342
rect 29668 73328 29750 73342
rect 30626 73328 30708 73342
rect 30916 73328 30998 73342
rect 31874 73328 31956 73342
rect 32164 73328 32246 73342
rect 33122 73328 33204 73342
rect 33412 73328 33494 73342
rect 34370 73328 34452 73342
rect 34660 73328 34742 73342
rect 35618 73328 35700 73342
rect 35908 73328 35990 73342
rect 36866 73328 36948 73342
rect 37156 73328 37238 73342
rect 38114 73328 38196 73342
rect 38404 73328 38486 73342
rect 39362 73328 39444 73342
rect 39652 73328 39734 73342
rect 40610 73328 40692 73342
rect 40900 73328 40982 73342
rect 41858 73328 41940 73342
rect 42148 73328 42230 73342
rect 43106 73328 43188 73342
rect 43396 73328 43478 73342
rect 44354 73328 44436 73342
rect 44644 73328 44726 73342
rect 45602 73328 45684 73342
rect 45892 73328 45974 73342
rect 46850 73328 46932 73342
rect 47140 73328 47222 73342
rect 48098 73328 48180 73342
rect 48388 73328 48470 73342
rect 49346 73328 49428 73342
rect 49636 73328 49718 73342
rect 50594 73328 50676 73342
rect 50884 73328 50966 73342
rect 51842 73328 51924 73342
rect 52132 73328 52214 73342
rect 53090 73328 53172 73342
rect 53380 73328 53462 73342
rect 54338 73328 54420 73342
rect 54628 73328 54710 73342
rect 55586 73328 55668 73342
rect 55876 73328 55958 73342
rect 56834 73328 56916 73342
rect 57124 73328 57206 73342
rect 58082 73328 58164 73342
rect 58372 73328 58454 73342
rect 16418 73280 16864 73294
rect 17014 73280 17154 73294
rect 17304 73280 18112 73294
rect 18262 73280 18402 73294
rect 18552 73280 19360 73294
rect 19510 73280 19650 73294
rect 19800 73280 20608 73294
rect 20758 73280 20898 73294
rect 21048 73280 21856 73294
rect 22006 73280 22146 73294
rect 22296 73280 23104 73294
rect 23254 73280 23394 73294
rect 23544 73280 24352 73294
rect 24502 73280 24642 73294
rect 24792 73280 25600 73294
rect 25750 73280 25890 73294
rect 26040 73280 26848 73294
rect 26998 73280 27138 73294
rect 27288 73280 28096 73294
rect 28246 73280 28386 73294
rect 28536 73280 29344 73294
rect 29494 73280 29634 73294
rect 29784 73280 30592 73294
rect 30742 73280 30882 73294
rect 31032 73280 31840 73294
rect 31990 73280 32130 73294
rect 32280 73280 33088 73294
rect 33238 73280 33378 73294
rect 33528 73280 34336 73294
rect 34486 73280 34626 73294
rect 34776 73280 35584 73294
rect 35734 73280 35874 73294
rect 36024 73280 36832 73294
rect 36982 73280 37122 73294
rect 37272 73280 38080 73294
rect 38230 73280 38370 73294
rect 38520 73280 39328 73294
rect 39478 73280 39618 73294
rect 39768 73280 40576 73294
rect 40726 73280 40866 73294
rect 41016 73280 41824 73294
rect 41974 73280 42114 73294
rect 42264 73280 43072 73294
rect 43222 73280 43362 73294
rect 43512 73280 44320 73294
rect 44470 73280 44610 73294
rect 44760 73280 45568 73294
rect 45718 73280 45858 73294
rect 46008 73280 46816 73294
rect 46966 73280 47106 73294
rect 47256 73280 48064 73294
rect 48214 73280 48354 73294
rect 48504 73280 49312 73294
rect 49462 73280 49602 73294
rect 49752 73280 50560 73294
rect 50710 73280 50850 73294
rect 51000 73280 51808 73294
rect 51958 73280 52098 73294
rect 52248 73280 53056 73294
rect 53206 73280 53346 73294
rect 53496 73280 54304 73294
rect 54454 73280 54594 73294
rect 54744 73280 55552 73294
rect 55702 73280 55842 73294
rect 55992 73280 56800 73294
rect 56950 73280 57090 73294
rect 57240 73280 58048 73294
rect 58198 73280 58338 73294
rect 58488 73280 58934 73294
rect 16418 73232 58934 73280
rect 16418 73218 16864 73232
rect 17014 73218 17154 73232
rect 17304 73218 18112 73232
rect 18262 73218 18402 73232
rect 18552 73218 19360 73232
rect 19510 73218 19650 73232
rect 19800 73218 20608 73232
rect 20758 73218 20898 73232
rect 21048 73218 21856 73232
rect 22006 73218 22146 73232
rect 22296 73218 23104 73232
rect 23254 73218 23394 73232
rect 23544 73218 24352 73232
rect 24502 73218 24642 73232
rect 24792 73218 25600 73232
rect 25750 73218 25890 73232
rect 26040 73218 26848 73232
rect 26998 73218 27138 73232
rect 27288 73218 28096 73232
rect 28246 73218 28386 73232
rect 28536 73218 29344 73232
rect 29494 73218 29634 73232
rect 29784 73218 30592 73232
rect 30742 73218 30882 73232
rect 31032 73218 31840 73232
rect 31990 73218 32130 73232
rect 32280 73218 33088 73232
rect 33238 73218 33378 73232
rect 33528 73218 34336 73232
rect 34486 73218 34626 73232
rect 34776 73218 35584 73232
rect 35734 73218 35874 73232
rect 36024 73218 36832 73232
rect 36982 73218 37122 73232
rect 37272 73218 38080 73232
rect 38230 73218 38370 73232
rect 38520 73218 39328 73232
rect 39478 73218 39618 73232
rect 39768 73218 40576 73232
rect 40726 73218 40866 73232
rect 41016 73218 41824 73232
rect 41974 73218 42114 73232
rect 42264 73218 43072 73232
rect 43222 73218 43362 73232
rect 43512 73218 44320 73232
rect 44470 73218 44610 73232
rect 44760 73218 45568 73232
rect 45718 73218 45858 73232
rect 46008 73218 46816 73232
rect 46966 73218 47106 73232
rect 47256 73218 48064 73232
rect 48214 73218 48354 73232
rect 48504 73218 49312 73232
rect 49462 73218 49602 73232
rect 49752 73218 50560 73232
rect 50710 73218 50850 73232
rect 51000 73218 51808 73232
rect 51958 73218 52098 73232
rect 52248 73218 53056 73232
rect 53206 73218 53346 73232
rect 53496 73218 54304 73232
rect 54454 73218 54594 73232
rect 54744 73218 55552 73232
rect 55702 73218 55842 73232
rect 55992 73218 56800 73232
rect 56950 73218 57090 73232
rect 57240 73218 58048 73232
rect 58198 73218 58338 73232
rect 58488 73218 58934 73232
rect 16898 73170 16980 73184
rect 17188 73170 17270 73184
rect 18146 73170 18228 73184
rect 18436 73170 18518 73184
rect 19394 73170 19476 73184
rect 19684 73170 19766 73184
rect 20642 73170 20724 73184
rect 20932 73170 21014 73184
rect 21890 73170 21972 73184
rect 22180 73170 22262 73184
rect 23138 73170 23220 73184
rect 23428 73170 23510 73184
rect 24386 73170 24468 73184
rect 24676 73170 24758 73184
rect 25634 73170 25716 73184
rect 25924 73170 26006 73184
rect 26882 73170 26964 73184
rect 27172 73170 27254 73184
rect 28130 73170 28212 73184
rect 28420 73170 28502 73184
rect 29378 73170 29460 73184
rect 29668 73170 29750 73184
rect 30626 73170 30708 73184
rect 30916 73170 30998 73184
rect 31874 73170 31956 73184
rect 32164 73170 32246 73184
rect 33122 73170 33204 73184
rect 33412 73170 33494 73184
rect 34370 73170 34452 73184
rect 34660 73170 34742 73184
rect 35618 73170 35700 73184
rect 35908 73170 35990 73184
rect 36866 73170 36948 73184
rect 37156 73170 37238 73184
rect 38114 73170 38196 73184
rect 38404 73170 38486 73184
rect 39362 73170 39444 73184
rect 39652 73170 39734 73184
rect 40610 73170 40692 73184
rect 40900 73170 40982 73184
rect 41858 73170 41940 73184
rect 42148 73170 42230 73184
rect 43106 73170 43188 73184
rect 43396 73170 43478 73184
rect 44354 73170 44436 73184
rect 44644 73170 44726 73184
rect 45602 73170 45684 73184
rect 45892 73170 45974 73184
rect 46850 73170 46932 73184
rect 47140 73170 47222 73184
rect 48098 73170 48180 73184
rect 48388 73170 48470 73184
rect 49346 73170 49428 73184
rect 49636 73170 49718 73184
rect 50594 73170 50676 73184
rect 50884 73170 50966 73184
rect 51842 73170 51924 73184
rect 52132 73170 52214 73184
rect 53090 73170 53172 73184
rect 53380 73170 53462 73184
rect 54338 73170 54420 73184
rect 54628 73170 54710 73184
rect 55586 73170 55668 73184
rect 55876 73170 55958 73184
rect 56834 73170 56916 73184
rect 57124 73170 57206 73184
rect 58082 73170 58164 73184
rect 58372 73170 58454 73184
rect 16418 73122 58934 73170
rect 16418 73026 58934 73074
rect 16898 73012 16980 73026
rect 17188 73012 17270 73026
rect 18146 73012 18228 73026
rect 18436 73012 18518 73026
rect 19394 73012 19476 73026
rect 19684 73012 19766 73026
rect 20642 73012 20724 73026
rect 20932 73012 21014 73026
rect 21890 73012 21972 73026
rect 22180 73012 22262 73026
rect 23138 73012 23220 73026
rect 23428 73012 23510 73026
rect 24386 73012 24468 73026
rect 24676 73012 24758 73026
rect 25634 73012 25716 73026
rect 25924 73012 26006 73026
rect 26882 73012 26964 73026
rect 27172 73012 27254 73026
rect 28130 73012 28212 73026
rect 28420 73012 28502 73026
rect 29378 73012 29460 73026
rect 29668 73012 29750 73026
rect 30626 73012 30708 73026
rect 30916 73012 30998 73026
rect 31874 73012 31956 73026
rect 32164 73012 32246 73026
rect 33122 73012 33204 73026
rect 33412 73012 33494 73026
rect 34370 73012 34452 73026
rect 34660 73012 34742 73026
rect 35618 73012 35700 73026
rect 35908 73012 35990 73026
rect 36866 73012 36948 73026
rect 37156 73012 37238 73026
rect 38114 73012 38196 73026
rect 38404 73012 38486 73026
rect 39362 73012 39444 73026
rect 39652 73012 39734 73026
rect 40610 73012 40692 73026
rect 40900 73012 40982 73026
rect 41858 73012 41940 73026
rect 42148 73012 42230 73026
rect 43106 73012 43188 73026
rect 43396 73012 43478 73026
rect 44354 73012 44436 73026
rect 44644 73012 44726 73026
rect 45602 73012 45684 73026
rect 45892 73012 45974 73026
rect 46850 73012 46932 73026
rect 47140 73012 47222 73026
rect 48098 73012 48180 73026
rect 48388 73012 48470 73026
rect 49346 73012 49428 73026
rect 49636 73012 49718 73026
rect 50594 73012 50676 73026
rect 50884 73012 50966 73026
rect 51842 73012 51924 73026
rect 52132 73012 52214 73026
rect 53090 73012 53172 73026
rect 53380 73012 53462 73026
rect 54338 73012 54420 73026
rect 54628 73012 54710 73026
rect 55586 73012 55668 73026
rect 55876 73012 55958 73026
rect 56834 73012 56916 73026
rect 57124 73012 57206 73026
rect 58082 73012 58164 73026
rect 58372 73012 58454 73026
rect 16418 72964 16864 72978
rect 17014 72964 17154 72978
rect 17304 72964 18112 72978
rect 18262 72964 18402 72978
rect 18552 72964 19360 72978
rect 19510 72964 19650 72978
rect 19800 72964 20608 72978
rect 20758 72964 20898 72978
rect 21048 72964 21856 72978
rect 22006 72964 22146 72978
rect 22296 72964 23104 72978
rect 23254 72964 23394 72978
rect 23544 72964 24352 72978
rect 24502 72964 24642 72978
rect 24792 72964 25600 72978
rect 25750 72964 25890 72978
rect 26040 72964 26848 72978
rect 26998 72964 27138 72978
rect 27288 72964 28096 72978
rect 28246 72964 28386 72978
rect 28536 72964 29344 72978
rect 29494 72964 29634 72978
rect 29784 72964 30592 72978
rect 30742 72964 30882 72978
rect 31032 72964 31840 72978
rect 31990 72964 32130 72978
rect 32280 72964 33088 72978
rect 33238 72964 33378 72978
rect 33528 72964 34336 72978
rect 34486 72964 34626 72978
rect 34776 72964 35584 72978
rect 35734 72964 35874 72978
rect 36024 72964 36832 72978
rect 36982 72964 37122 72978
rect 37272 72964 38080 72978
rect 38230 72964 38370 72978
rect 38520 72964 39328 72978
rect 39478 72964 39618 72978
rect 39768 72964 40576 72978
rect 40726 72964 40866 72978
rect 41016 72964 41824 72978
rect 41974 72964 42114 72978
rect 42264 72964 43072 72978
rect 43222 72964 43362 72978
rect 43512 72964 44320 72978
rect 44470 72964 44610 72978
rect 44760 72964 45568 72978
rect 45718 72964 45858 72978
rect 46008 72964 46816 72978
rect 46966 72964 47106 72978
rect 47256 72964 48064 72978
rect 48214 72964 48354 72978
rect 48504 72964 49312 72978
rect 49462 72964 49602 72978
rect 49752 72964 50560 72978
rect 50710 72964 50850 72978
rect 51000 72964 51808 72978
rect 51958 72964 52098 72978
rect 52248 72964 53056 72978
rect 53206 72964 53346 72978
rect 53496 72964 54304 72978
rect 54454 72964 54594 72978
rect 54744 72964 55552 72978
rect 55702 72964 55842 72978
rect 55992 72964 56800 72978
rect 56950 72964 57090 72978
rect 57240 72964 58048 72978
rect 58198 72964 58338 72978
rect 58488 72964 58934 72978
rect 16418 72916 58934 72964
rect 16418 72902 16864 72916
rect 17014 72902 17154 72916
rect 17304 72902 18112 72916
rect 18262 72902 18402 72916
rect 18552 72902 19360 72916
rect 19510 72902 19650 72916
rect 19800 72902 20608 72916
rect 20758 72902 20898 72916
rect 21048 72902 21856 72916
rect 22006 72902 22146 72916
rect 22296 72902 23104 72916
rect 23254 72902 23394 72916
rect 23544 72902 24352 72916
rect 24502 72902 24642 72916
rect 24792 72902 25600 72916
rect 25750 72902 25890 72916
rect 26040 72902 26848 72916
rect 26998 72902 27138 72916
rect 27288 72902 28096 72916
rect 28246 72902 28386 72916
rect 28536 72902 29344 72916
rect 29494 72902 29634 72916
rect 29784 72902 30592 72916
rect 30742 72902 30882 72916
rect 31032 72902 31840 72916
rect 31990 72902 32130 72916
rect 32280 72902 33088 72916
rect 33238 72902 33378 72916
rect 33528 72902 34336 72916
rect 34486 72902 34626 72916
rect 34776 72902 35584 72916
rect 35734 72902 35874 72916
rect 36024 72902 36832 72916
rect 36982 72902 37122 72916
rect 37272 72902 38080 72916
rect 38230 72902 38370 72916
rect 38520 72902 39328 72916
rect 39478 72902 39618 72916
rect 39768 72902 40576 72916
rect 40726 72902 40866 72916
rect 41016 72902 41824 72916
rect 41974 72902 42114 72916
rect 42264 72902 43072 72916
rect 43222 72902 43362 72916
rect 43512 72902 44320 72916
rect 44470 72902 44610 72916
rect 44760 72902 45568 72916
rect 45718 72902 45858 72916
rect 46008 72902 46816 72916
rect 46966 72902 47106 72916
rect 47256 72902 48064 72916
rect 48214 72902 48354 72916
rect 48504 72902 49312 72916
rect 49462 72902 49602 72916
rect 49752 72902 50560 72916
rect 50710 72902 50850 72916
rect 51000 72902 51808 72916
rect 51958 72902 52098 72916
rect 52248 72902 53056 72916
rect 53206 72902 53346 72916
rect 53496 72902 54304 72916
rect 54454 72902 54594 72916
rect 54744 72902 55552 72916
rect 55702 72902 55842 72916
rect 55992 72902 56800 72916
rect 56950 72902 57090 72916
rect 57240 72902 58048 72916
rect 58198 72902 58338 72916
rect 58488 72902 58934 72916
rect 16898 72854 16980 72868
rect 17188 72854 17270 72868
rect 18146 72854 18228 72868
rect 18436 72854 18518 72868
rect 19394 72854 19476 72868
rect 19684 72854 19766 72868
rect 20642 72854 20724 72868
rect 20932 72854 21014 72868
rect 21890 72854 21972 72868
rect 22180 72854 22262 72868
rect 23138 72854 23220 72868
rect 23428 72854 23510 72868
rect 24386 72854 24468 72868
rect 24676 72854 24758 72868
rect 25634 72854 25716 72868
rect 25924 72854 26006 72868
rect 26882 72854 26964 72868
rect 27172 72854 27254 72868
rect 28130 72854 28212 72868
rect 28420 72854 28502 72868
rect 29378 72854 29460 72868
rect 29668 72854 29750 72868
rect 30626 72854 30708 72868
rect 30916 72854 30998 72868
rect 31874 72854 31956 72868
rect 32164 72854 32246 72868
rect 33122 72854 33204 72868
rect 33412 72854 33494 72868
rect 34370 72854 34452 72868
rect 34660 72854 34742 72868
rect 35618 72854 35700 72868
rect 35908 72854 35990 72868
rect 36866 72854 36948 72868
rect 37156 72854 37238 72868
rect 38114 72854 38196 72868
rect 38404 72854 38486 72868
rect 39362 72854 39444 72868
rect 39652 72854 39734 72868
rect 40610 72854 40692 72868
rect 40900 72854 40982 72868
rect 41858 72854 41940 72868
rect 42148 72854 42230 72868
rect 43106 72854 43188 72868
rect 43396 72854 43478 72868
rect 44354 72854 44436 72868
rect 44644 72854 44726 72868
rect 45602 72854 45684 72868
rect 45892 72854 45974 72868
rect 46850 72854 46932 72868
rect 47140 72854 47222 72868
rect 48098 72854 48180 72868
rect 48388 72854 48470 72868
rect 49346 72854 49428 72868
rect 49636 72854 49718 72868
rect 50594 72854 50676 72868
rect 50884 72854 50966 72868
rect 51842 72854 51924 72868
rect 52132 72854 52214 72868
rect 53090 72854 53172 72868
rect 53380 72854 53462 72868
rect 54338 72854 54420 72868
rect 54628 72854 54710 72868
rect 55586 72854 55668 72868
rect 55876 72854 55958 72868
rect 56834 72854 56916 72868
rect 57124 72854 57206 72868
rect 58082 72854 58164 72868
rect 58372 72854 58454 72868
rect 16418 72806 58934 72854
rect 16418 72648 58934 72758
rect 16418 72552 58934 72600
rect 16898 72538 16980 72552
rect 17188 72538 17270 72552
rect 18146 72538 18228 72552
rect 18436 72538 18518 72552
rect 19394 72538 19476 72552
rect 19684 72538 19766 72552
rect 20642 72538 20724 72552
rect 20932 72538 21014 72552
rect 21890 72538 21972 72552
rect 22180 72538 22262 72552
rect 23138 72538 23220 72552
rect 23428 72538 23510 72552
rect 24386 72538 24468 72552
rect 24676 72538 24758 72552
rect 25634 72538 25716 72552
rect 25924 72538 26006 72552
rect 26882 72538 26964 72552
rect 27172 72538 27254 72552
rect 28130 72538 28212 72552
rect 28420 72538 28502 72552
rect 29378 72538 29460 72552
rect 29668 72538 29750 72552
rect 30626 72538 30708 72552
rect 30916 72538 30998 72552
rect 31874 72538 31956 72552
rect 32164 72538 32246 72552
rect 33122 72538 33204 72552
rect 33412 72538 33494 72552
rect 34370 72538 34452 72552
rect 34660 72538 34742 72552
rect 35618 72538 35700 72552
rect 35908 72538 35990 72552
rect 36866 72538 36948 72552
rect 37156 72538 37238 72552
rect 38114 72538 38196 72552
rect 38404 72538 38486 72552
rect 39362 72538 39444 72552
rect 39652 72538 39734 72552
rect 40610 72538 40692 72552
rect 40900 72538 40982 72552
rect 41858 72538 41940 72552
rect 42148 72538 42230 72552
rect 43106 72538 43188 72552
rect 43396 72538 43478 72552
rect 44354 72538 44436 72552
rect 44644 72538 44726 72552
rect 45602 72538 45684 72552
rect 45892 72538 45974 72552
rect 46850 72538 46932 72552
rect 47140 72538 47222 72552
rect 48098 72538 48180 72552
rect 48388 72538 48470 72552
rect 49346 72538 49428 72552
rect 49636 72538 49718 72552
rect 50594 72538 50676 72552
rect 50884 72538 50966 72552
rect 51842 72538 51924 72552
rect 52132 72538 52214 72552
rect 53090 72538 53172 72552
rect 53380 72538 53462 72552
rect 54338 72538 54420 72552
rect 54628 72538 54710 72552
rect 55586 72538 55668 72552
rect 55876 72538 55958 72552
rect 56834 72538 56916 72552
rect 57124 72538 57206 72552
rect 58082 72538 58164 72552
rect 58372 72538 58454 72552
rect 16418 72490 16864 72504
rect 17014 72490 17154 72504
rect 17304 72490 18112 72504
rect 18262 72490 18402 72504
rect 18552 72490 19360 72504
rect 19510 72490 19650 72504
rect 19800 72490 20608 72504
rect 20758 72490 20898 72504
rect 21048 72490 21856 72504
rect 22006 72490 22146 72504
rect 22296 72490 23104 72504
rect 23254 72490 23394 72504
rect 23544 72490 24352 72504
rect 24502 72490 24642 72504
rect 24792 72490 25600 72504
rect 25750 72490 25890 72504
rect 26040 72490 26848 72504
rect 26998 72490 27138 72504
rect 27288 72490 28096 72504
rect 28246 72490 28386 72504
rect 28536 72490 29344 72504
rect 29494 72490 29634 72504
rect 29784 72490 30592 72504
rect 30742 72490 30882 72504
rect 31032 72490 31840 72504
rect 31990 72490 32130 72504
rect 32280 72490 33088 72504
rect 33238 72490 33378 72504
rect 33528 72490 34336 72504
rect 34486 72490 34626 72504
rect 34776 72490 35584 72504
rect 35734 72490 35874 72504
rect 36024 72490 36832 72504
rect 36982 72490 37122 72504
rect 37272 72490 38080 72504
rect 38230 72490 38370 72504
rect 38520 72490 39328 72504
rect 39478 72490 39618 72504
rect 39768 72490 40576 72504
rect 40726 72490 40866 72504
rect 41016 72490 41824 72504
rect 41974 72490 42114 72504
rect 42264 72490 43072 72504
rect 43222 72490 43362 72504
rect 43512 72490 44320 72504
rect 44470 72490 44610 72504
rect 44760 72490 45568 72504
rect 45718 72490 45858 72504
rect 46008 72490 46816 72504
rect 46966 72490 47106 72504
rect 47256 72490 48064 72504
rect 48214 72490 48354 72504
rect 48504 72490 49312 72504
rect 49462 72490 49602 72504
rect 49752 72490 50560 72504
rect 50710 72490 50850 72504
rect 51000 72490 51808 72504
rect 51958 72490 52098 72504
rect 52248 72490 53056 72504
rect 53206 72490 53346 72504
rect 53496 72490 54304 72504
rect 54454 72490 54594 72504
rect 54744 72490 55552 72504
rect 55702 72490 55842 72504
rect 55992 72490 56800 72504
rect 56950 72490 57090 72504
rect 57240 72490 58048 72504
rect 58198 72490 58338 72504
rect 58488 72490 58934 72504
rect 16418 72442 58934 72490
rect 16418 72428 16864 72442
rect 17014 72428 17154 72442
rect 17304 72428 18112 72442
rect 18262 72428 18402 72442
rect 18552 72428 19360 72442
rect 19510 72428 19650 72442
rect 19800 72428 20608 72442
rect 20758 72428 20898 72442
rect 21048 72428 21856 72442
rect 22006 72428 22146 72442
rect 22296 72428 23104 72442
rect 23254 72428 23394 72442
rect 23544 72428 24352 72442
rect 24502 72428 24642 72442
rect 24792 72428 25600 72442
rect 25750 72428 25890 72442
rect 26040 72428 26848 72442
rect 26998 72428 27138 72442
rect 27288 72428 28096 72442
rect 28246 72428 28386 72442
rect 28536 72428 29344 72442
rect 29494 72428 29634 72442
rect 29784 72428 30592 72442
rect 30742 72428 30882 72442
rect 31032 72428 31840 72442
rect 31990 72428 32130 72442
rect 32280 72428 33088 72442
rect 33238 72428 33378 72442
rect 33528 72428 34336 72442
rect 34486 72428 34626 72442
rect 34776 72428 35584 72442
rect 35734 72428 35874 72442
rect 36024 72428 36832 72442
rect 36982 72428 37122 72442
rect 37272 72428 38080 72442
rect 38230 72428 38370 72442
rect 38520 72428 39328 72442
rect 39478 72428 39618 72442
rect 39768 72428 40576 72442
rect 40726 72428 40866 72442
rect 41016 72428 41824 72442
rect 41974 72428 42114 72442
rect 42264 72428 43072 72442
rect 43222 72428 43362 72442
rect 43512 72428 44320 72442
rect 44470 72428 44610 72442
rect 44760 72428 45568 72442
rect 45718 72428 45858 72442
rect 46008 72428 46816 72442
rect 46966 72428 47106 72442
rect 47256 72428 48064 72442
rect 48214 72428 48354 72442
rect 48504 72428 49312 72442
rect 49462 72428 49602 72442
rect 49752 72428 50560 72442
rect 50710 72428 50850 72442
rect 51000 72428 51808 72442
rect 51958 72428 52098 72442
rect 52248 72428 53056 72442
rect 53206 72428 53346 72442
rect 53496 72428 54304 72442
rect 54454 72428 54594 72442
rect 54744 72428 55552 72442
rect 55702 72428 55842 72442
rect 55992 72428 56800 72442
rect 56950 72428 57090 72442
rect 57240 72428 58048 72442
rect 58198 72428 58338 72442
rect 58488 72428 58934 72442
rect 16898 72380 16980 72394
rect 17188 72380 17270 72394
rect 18146 72380 18228 72394
rect 18436 72380 18518 72394
rect 19394 72380 19476 72394
rect 19684 72380 19766 72394
rect 20642 72380 20724 72394
rect 20932 72380 21014 72394
rect 21890 72380 21972 72394
rect 22180 72380 22262 72394
rect 23138 72380 23220 72394
rect 23428 72380 23510 72394
rect 24386 72380 24468 72394
rect 24676 72380 24758 72394
rect 25634 72380 25716 72394
rect 25924 72380 26006 72394
rect 26882 72380 26964 72394
rect 27172 72380 27254 72394
rect 28130 72380 28212 72394
rect 28420 72380 28502 72394
rect 29378 72380 29460 72394
rect 29668 72380 29750 72394
rect 30626 72380 30708 72394
rect 30916 72380 30998 72394
rect 31874 72380 31956 72394
rect 32164 72380 32246 72394
rect 33122 72380 33204 72394
rect 33412 72380 33494 72394
rect 34370 72380 34452 72394
rect 34660 72380 34742 72394
rect 35618 72380 35700 72394
rect 35908 72380 35990 72394
rect 36866 72380 36948 72394
rect 37156 72380 37238 72394
rect 38114 72380 38196 72394
rect 38404 72380 38486 72394
rect 39362 72380 39444 72394
rect 39652 72380 39734 72394
rect 40610 72380 40692 72394
rect 40900 72380 40982 72394
rect 41858 72380 41940 72394
rect 42148 72380 42230 72394
rect 43106 72380 43188 72394
rect 43396 72380 43478 72394
rect 44354 72380 44436 72394
rect 44644 72380 44726 72394
rect 45602 72380 45684 72394
rect 45892 72380 45974 72394
rect 46850 72380 46932 72394
rect 47140 72380 47222 72394
rect 48098 72380 48180 72394
rect 48388 72380 48470 72394
rect 49346 72380 49428 72394
rect 49636 72380 49718 72394
rect 50594 72380 50676 72394
rect 50884 72380 50966 72394
rect 51842 72380 51924 72394
rect 52132 72380 52214 72394
rect 53090 72380 53172 72394
rect 53380 72380 53462 72394
rect 54338 72380 54420 72394
rect 54628 72380 54710 72394
rect 55586 72380 55668 72394
rect 55876 72380 55958 72394
rect 56834 72380 56916 72394
rect 57124 72380 57206 72394
rect 58082 72380 58164 72394
rect 58372 72380 58454 72394
rect 16418 72332 58934 72380
rect 16418 72236 58934 72284
rect 16898 72222 16980 72236
rect 17188 72222 17270 72236
rect 18146 72222 18228 72236
rect 18436 72222 18518 72236
rect 19394 72222 19476 72236
rect 19684 72222 19766 72236
rect 20642 72222 20724 72236
rect 20932 72222 21014 72236
rect 21890 72222 21972 72236
rect 22180 72222 22262 72236
rect 23138 72222 23220 72236
rect 23428 72222 23510 72236
rect 24386 72222 24468 72236
rect 24676 72222 24758 72236
rect 25634 72222 25716 72236
rect 25924 72222 26006 72236
rect 26882 72222 26964 72236
rect 27172 72222 27254 72236
rect 28130 72222 28212 72236
rect 28420 72222 28502 72236
rect 29378 72222 29460 72236
rect 29668 72222 29750 72236
rect 30626 72222 30708 72236
rect 30916 72222 30998 72236
rect 31874 72222 31956 72236
rect 32164 72222 32246 72236
rect 33122 72222 33204 72236
rect 33412 72222 33494 72236
rect 34370 72222 34452 72236
rect 34660 72222 34742 72236
rect 35618 72222 35700 72236
rect 35908 72222 35990 72236
rect 36866 72222 36948 72236
rect 37156 72222 37238 72236
rect 38114 72222 38196 72236
rect 38404 72222 38486 72236
rect 39362 72222 39444 72236
rect 39652 72222 39734 72236
rect 40610 72222 40692 72236
rect 40900 72222 40982 72236
rect 41858 72222 41940 72236
rect 42148 72222 42230 72236
rect 43106 72222 43188 72236
rect 43396 72222 43478 72236
rect 44354 72222 44436 72236
rect 44644 72222 44726 72236
rect 45602 72222 45684 72236
rect 45892 72222 45974 72236
rect 46850 72222 46932 72236
rect 47140 72222 47222 72236
rect 48098 72222 48180 72236
rect 48388 72222 48470 72236
rect 49346 72222 49428 72236
rect 49636 72222 49718 72236
rect 50594 72222 50676 72236
rect 50884 72222 50966 72236
rect 51842 72222 51924 72236
rect 52132 72222 52214 72236
rect 53090 72222 53172 72236
rect 53380 72222 53462 72236
rect 54338 72222 54420 72236
rect 54628 72222 54710 72236
rect 55586 72222 55668 72236
rect 55876 72222 55958 72236
rect 56834 72222 56916 72236
rect 57124 72222 57206 72236
rect 58082 72222 58164 72236
rect 58372 72222 58454 72236
rect 16418 72174 16864 72188
rect 17014 72174 17154 72188
rect 17304 72174 18112 72188
rect 18262 72174 18402 72188
rect 18552 72174 19360 72188
rect 19510 72174 19650 72188
rect 19800 72174 20608 72188
rect 20758 72174 20898 72188
rect 21048 72174 21856 72188
rect 22006 72174 22146 72188
rect 22296 72174 23104 72188
rect 23254 72174 23394 72188
rect 23544 72174 24352 72188
rect 24502 72174 24642 72188
rect 24792 72174 25600 72188
rect 25750 72174 25890 72188
rect 26040 72174 26848 72188
rect 26998 72174 27138 72188
rect 27288 72174 28096 72188
rect 28246 72174 28386 72188
rect 28536 72174 29344 72188
rect 29494 72174 29634 72188
rect 29784 72174 30592 72188
rect 30742 72174 30882 72188
rect 31032 72174 31840 72188
rect 31990 72174 32130 72188
rect 32280 72174 33088 72188
rect 33238 72174 33378 72188
rect 33528 72174 34336 72188
rect 34486 72174 34626 72188
rect 34776 72174 35584 72188
rect 35734 72174 35874 72188
rect 36024 72174 36832 72188
rect 36982 72174 37122 72188
rect 37272 72174 38080 72188
rect 38230 72174 38370 72188
rect 38520 72174 39328 72188
rect 39478 72174 39618 72188
rect 39768 72174 40576 72188
rect 40726 72174 40866 72188
rect 41016 72174 41824 72188
rect 41974 72174 42114 72188
rect 42264 72174 43072 72188
rect 43222 72174 43362 72188
rect 43512 72174 44320 72188
rect 44470 72174 44610 72188
rect 44760 72174 45568 72188
rect 45718 72174 45858 72188
rect 46008 72174 46816 72188
rect 46966 72174 47106 72188
rect 47256 72174 48064 72188
rect 48214 72174 48354 72188
rect 48504 72174 49312 72188
rect 49462 72174 49602 72188
rect 49752 72174 50560 72188
rect 50710 72174 50850 72188
rect 51000 72174 51808 72188
rect 51958 72174 52098 72188
rect 52248 72174 53056 72188
rect 53206 72174 53346 72188
rect 53496 72174 54304 72188
rect 54454 72174 54594 72188
rect 54744 72174 55552 72188
rect 55702 72174 55842 72188
rect 55992 72174 56800 72188
rect 56950 72174 57090 72188
rect 57240 72174 58048 72188
rect 58198 72174 58338 72188
rect 58488 72174 58934 72188
rect 16418 72126 58934 72174
rect 16418 72112 16864 72126
rect 17014 72112 17154 72126
rect 17304 72112 18112 72126
rect 18262 72112 18402 72126
rect 18552 72112 19360 72126
rect 19510 72112 19650 72126
rect 19800 72112 20608 72126
rect 20758 72112 20898 72126
rect 21048 72112 21856 72126
rect 22006 72112 22146 72126
rect 22296 72112 23104 72126
rect 23254 72112 23394 72126
rect 23544 72112 24352 72126
rect 24502 72112 24642 72126
rect 24792 72112 25600 72126
rect 25750 72112 25890 72126
rect 26040 72112 26848 72126
rect 26998 72112 27138 72126
rect 27288 72112 28096 72126
rect 28246 72112 28386 72126
rect 28536 72112 29344 72126
rect 29494 72112 29634 72126
rect 29784 72112 30592 72126
rect 30742 72112 30882 72126
rect 31032 72112 31840 72126
rect 31990 72112 32130 72126
rect 32280 72112 33088 72126
rect 33238 72112 33378 72126
rect 33528 72112 34336 72126
rect 34486 72112 34626 72126
rect 34776 72112 35584 72126
rect 35734 72112 35874 72126
rect 36024 72112 36832 72126
rect 36982 72112 37122 72126
rect 37272 72112 38080 72126
rect 38230 72112 38370 72126
rect 38520 72112 39328 72126
rect 39478 72112 39618 72126
rect 39768 72112 40576 72126
rect 40726 72112 40866 72126
rect 41016 72112 41824 72126
rect 41974 72112 42114 72126
rect 42264 72112 43072 72126
rect 43222 72112 43362 72126
rect 43512 72112 44320 72126
rect 44470 72112 44610 72126
rect 44760 72112 45568 72126
rect 45718 72112 45858 72126
rect 46008 72112 46816 72126
rect 46966 72112 47106 72126
rect 47256 72112 48064 72126
rect 48214 72112 48354 72126
rect 48504 72112 49312 72126
rect 49462 72112 49602 72126
rect 49752 72112 50560 72126
rect 50710 72112 50850 72126
rect 51000 72112 51808 72126
rect 51958 72112 52098 72126
rect 52248 72112 53056 72126
rect 53206 72112 53346 72126
rect 53496 72112 54304 72126
rect 54454 72112 54594 72126
rect 54744 72112 55552 72126
rect 55702 72112 55842 72126
rect 55992 72112 56800 72126
rect 56950 72112 57090 72126
rect 57240 72112 58048 72126
rect 58198 72112 58338 72126
rect 58488 72112 58934 72126
rect 16898 72064 16980 72078
rect 17188 72064 17270 72078
rect 18146 72064 18228 72078
rect 18436 72064 18518 72078
rect 19394 72064 19476 72078
rect 19684 72064 19766 72078
rect 20642 72064 20724 72078
rect 20932 72064 21014 72078
rect 21890 72064 21972 72078
rect 22180 72064 22262 72078
rect 23138 72064 23220 72078
rect 23428 72064 23510 72078
rect 24386 72064 24468 72078
rect 24676 72064 24758 72078
rect 25634 72064 25716 72078
rect 25924 72064 26006 72078
rect 26882 72064 26964 72078
rect 27172 72064 27254 72078
rect 28130 72064 28212 72078
rect 28420 72064 28502 72078
rect 29378 72064 29460 72078
rect 29668 72064 29750 72078
rect 30626 72064 30708 72078
rect 30916 72064 30998 72078
rect 31874 72064 31956 72078
rect 32164 72064 32246 72078
rect 33122 72064 33204 72078
rect 33412 72064 33494 72078
rect 34370 72064 34452 72078
rect 34660 72064 34742 72078
rect 35618 72064 35700 72078
rect 35908 72064 35990 72078
rect 36866 72064 36948 72078
rect 37156 72064 37238 72078
rect 38114 72064 38196 72078
rect 38404 72064 38486 72078
rect 39362 72064 39444 72078
rect 39652 72064 39734 72078
rect 40610 72064 40692 72078
rect 40900 72064 40982 72078
rect 41858 72064 41940 72078
rect 42148 72064 42230 72078
rect 43106 72064 43188 72078
rect 43396 72064 43478 72078
rect 44354 72064 44436 72078
rect 44644 72064 44726 72078
rect 45602 72064 45684 72078
rect 45892 72064 45974 72078
rect 46850 72064 46932 72078
rect 47140 72064 47222 72078
rect 48098 72064 48180 72078
rect 48388 72064 48470 72078
rect 49346 72064 49428 72078
rect 49636 72064 49718 72078
rect 50594 72064 50676 72078
rect 50884 72064 50966 72078
rect 51842 72064 51924 72078
rect 52132 72064 52214 72078
rect 53090 72064 53172 72078
rect 53380 72064 53462 72078
rect 54338 72064 54420 72078
rect 54628 72064 54710 72078
rect 55586 72064 55668 72078
rect 55876 72064 55958 72078
rect 56834 72064 56916 72078
rect 57124 72064 57206 72078
rect 58082 72064 58164 72078
rect 58372 72064 58454 72078
rect 16418 72016 58934 72064
rect 16418 71858 58934 71968
rect 16418 71762 58934 71810
rect 16898 71748 16980 71762
rect 17188 71748 17270 71762
rect 18146 71748 18228 71762
rect 18436 71748 18518 71762
rect 19394 71748 19476 71762
rect 19684 71748 19766 71762
rect 20642 71748 20724 71762
rect 20932 71748 21014 71762
rect 21890 71748 21972 71762
rect 22180 71748 22262 71762
rect 23138 71748 23220 71762
rect 23428 71748 23510 71762
rect 24386 71748 24468 71762
rect 24676 71748 24758 71762
rect 25634 71748 25716 71762
rect 25924 71748 26006 71762
rect 26882 71748 26964 71762
rect 27172 71748 27254 71762
rect 28130 71748 28212 71762
rect 28420 71748 28502 71762
rect 29378 71748 29460 71762
rect 29668 71748 29750 71762
rect 30626 71748 30708 71762
rect 30916 71748 30998 71762
rect 31874 71748 31956 71762
rect 32164 71748 32246 71762
rect 33122 71748 33204 71762
rect 33412 71748 33494 71762
rect 34370 71748 34452 71762
rect 34660 71748 34742 71762
rect 35618 71748 35700 71762
rect 35908 71748 35990 71762
rect 36866 71748 36948 71762
rect 37156 71748 37238 71762
rect 38114 71748 38196 71762
rect 38404 71748 38486 71762
rect 39362 71748 39444 71762
rect 39652 71748 39734 71762
rect 40610 71748 40692 71762
rect 40900 71748 40982 71762
rect 41858 71748 41940 71762
rect 42148 71748 42230 71762
rect 43106 71748 43188 71762
rect 43396 71748 43478 71762
rect 44354 71748 44436 71762
rect 44644 71748 44726 71762
rect 45602 71748 45684 71762
rect 45892 71748 45974 71762
rect 46850 71748 46932 71762
rect 47140 71748 47222 71762
rect 48098 71748 48180 71762
rect 48388 71748 48470 71762
rect 49346 71748 49428 71762
rect 49636 71748 49718 71762
rect 50594 71748 50676 71762
rect 50884 71748 50966 71762
rect 51842 71748 51924 71762
rect 52132 71748 52214 71762
rect 53090 71748 53172 71762
rect 53380 71748 53462 71762
rect 54338 71748 54420 71762
rect 54628 71748 54710 71762
rect 55586 71748 55668 71762
rect 55876 71748 55958 71762
rect 56834 71748 56916 71762
rect 57124 71748 57206 71762
rect 58082 71748 58164 71762
rect 58372 71748 58454 71762
rect 16418 71700 16864 71714
rect 17014 71700 17154 71714
rect 17304 71700 18112 71714
rect 18262 71700 18402 71714
rect 18552 71700 19360 71714
rect 19510 71700 19650 71714
rect 19800 71700 20608 71714
rect 20758 71700 20898 71714
rect 21048 71700 21856 71714
rect 22006 71700 22146 71714
rect 22296 71700 23104 71714
rect 23254 71700 23394 71714
rect 23544 71700 24352 71714
rect 24502 71700 24642 71714
rect 24792 71700 25600 71714
rect 25750 71700 25890 71714
rect 26040 71700 26848 71714
rect 26998 71700 27138 71714
rect 27288 71700 28096 71714
rect 28246 71700 28386 71714
rect 28536 71700 29344 71714
rect 29494 71700 29634 71714
rect 29784 71700 30592 71714
rect 30742 71700 30882 71714
rect 31032 71700 31840 71714
rect 31990 71700 32130 71714
rect 32280 71700 33088 71714
rect 33238 71700 33378 71714
rect 33528 71700 34336 71714
rect 34486 71700 34626 71714
rect 34776 71700 35584 71714
rect 35734 71700 35874 71714
rect 36024 71700 36832 71714
rect 36982 71700 37122 71714
rect 37272 71700 38080 71714
rect 38230 71700 38370 71714
rect 38520 71700 39328 71714
rect 39478 71700 39618 71714
rect 39768 71700 40576 71714
rect 40726 71700 40866 71714
rect 41016 71700 41824 71714
rect 41974 71700 42114 71714
rect 42264 71700 43072 71714
rect 43222 71700 43362 71714
rect 43512 71700 44320 71714
rect 44470 71700 44610 71714
rect 44760 71700 45568 71714
rect 45718 71700 45858 71714
rect 46008 71700 46816 71714
rect 46966 71700 47106 71714
rect 47256 71700 48064 71714
rect 48214 71700 48354 71714
rect 48504 71700 49312 71714
rect 49462 71700 49602 71714
rect 49752 71700 50560 71714
rect 50710 71700 50850 71714
rect 51000 71700 51808 71714
rect 51958 71700 52098 71714
rect 52248 71700 53056 71714
rect 53206 71700 53346 71714
rect 53496 71700 54304 71714
rect 54454 71700 54594 71714
rect 54744 71700 55552 71714
rect 55702 71700 55842 71714
rect 55992 71700 56800 71714
rect 56950 71700 57090 71714
rect 57240 71700 58048 71714
rect 58198 71700 58338 71714
rect 58488 71700 58934 71714
rect 16418 71652 58934 71700
rect 16418 71638 16864 71652
rect 17014 71638 17154 71652
rect 17304 71638 18112 71652
rect 18262 71638 18402 71652
rect 18552 71638 19360 71652
rect 19510 71638 19650 71652
rect 19800 71638 20608 71652
rect 20758 71638 20898 71652
rect 21048 71638 21856 71652
rect 22006 71638 22146 71652
rect 22296 71638 23104 71652
rect 23254 71638 23394 71652
rect 23544 71638 24352 71652
rect 24502 71638 24642 71652
rect 24792 71638 25600 71652
rect 25750 71638 25890 71652
rect 26040 71638 26848 71652
rect 26998 71638 27138 71652
rect 27288 71638 28096 71652
rect 28246 71638 28386 71652
rect 28536 71638 29344 71652
rect 29494 71638 29634 71652
rect 29784 71638 30592 71652
rect 30742 71638 30882 71652
rect 31032 71638 31840 71652
rect 31990 71638 32130 71652
rect 32280 71638 33088 71652
rect 33238 71638 33378 71652
rect 33528 71638 34336 71652
rect 34486 71638 34626 71652
rect 34776 71638 35584 71652
rect 35734 71638 35874 71652
rect 36024 71638 36832 71652
rect 36982 71638 37122 71652
rect 37272 71638 38080 71652
rect 38230 71638 38370 71652
rect 38520 71638 39328 71652
rect 39478 71638 39618 71652
rect 39768 71638 40576 71652
rect 40726 71638 40866 71652
rect 41016 71638 41824 71652
rect 41974 71638 42114 71652
rect 42264 71638 43072 71652
rect 43222 71638 43362 71652
rect 43512 71638 44320 71652
rect 44470 71638 44610 71652
rect 44760 71638 45568 71652
rect 45718 71638 45858 71652
rect 46008 71638 46816 71652
rect 46966 71638 47106 71652
rect 47256 71638 48064 71652
rect 48214 71638 48354 71652
rect 48504 71638 49312 71652
rect 49462 71638 49602 71652
rect 49752 71638 50560 71652
rect 50710 71638 50850 71652
rect 51000 71638 51808 71652
rect 51958 71638 52098 71652
rect 52248 71638 53056 71652
rect 53206 71638 53346 71652
rect 53496 71638 54304 71652
rect 54454 71638 54594 71652
rect 54744 71638 55552 71652
rect 55702 71638 55842 71652
rect 55992 71638 56800 71652
rect 56950 71638 57090 71652
rect 57240 71638 58048 71652
rect 58198 71638 58338 71652
rect 58488 71638 58934 71652
rect 16898 71590 16980 71604
rect 17188 71590 17270 71604
rect 18146 71590 18228 71604
rect 18436 71590 18518 71604
rect 19394 71590 19476 71604
rect 19684 71590 19766 71604
rect 20642 71590 20724 71604
rect 20932 71590 21014 71604
rect 21890 71590 21972 71604
rect 22180 71590 22262 71604
rect 23138 71590 23220 71604
rect 23428 71590 23510 71604
rect 24386 71590 24468 71604
rect 24676 71590 24758 71604
rect 25634 71590 25716 71604
rect 25924 71590 26006 71604
rect 26882 71590 26964 71604
rect 27172 71590 27254 71604
rect 28130 71590 28212 71604
rect 28420 71590 28502 71604
rect 29378 71590 29460 71604
rect 29668 71590 29750 71604
rect 30626 71590 30708 71604
rect 30916 71590 30998 71604
rect 31874 71590 31956 71604
rect 32164 71590 32246 71604
rect 33122 71590 33204 71604
rect 33412 71590 33494 71604
rect 34370 71590 34452 71604
rect 34660 71590 34742 71604
rect 35618 71590 35700 71604
rect 35908 71590 35990 71604
rect 36866 71590 36948 71604
rect 37156 71590 37238 71604
rect 38114 71590 38196 71604
rect 38404 71590 38486 71604
rect 39362 71590 39444 71604
rect 39652 71590 39734 71604
rect 40610 71590 40692 71604
rect 40900 71590 40982 71604
rect 41858 71590 41940 71604
rect 42148 71590 42230 71604
rect 43106 71590 43188 71604
rect 43396 71590 43478 71604
rect 44354 71590 44436 71604
rect 44644 71590 44726 71604
rect 45602 71590 45684 71604
rect 45892 71590 45974 71604
rect 46850 71590 46932 71604
rect 47140 71590 47222 71604
rect 48098 71590 48180 71604
rect 48388 71590 48470 71604
rect 49346 71590 49428 71604
rect 49636 71590 49718 71604
rect 50594 71590 50676 71604
rect 50884 71590 50966 71604
rect 51842 71590 51924 71604
rect 52132 71590 52214 71604
rect 53090 71590 53172 71604
rect 53380 71590 53462 71604
rect 54338 71590 54420 71604
rect 54628 71590 54710 71604
rect 55586 71590 55668 71604
rect 55876 71590 55958 71604
rect 56834 71590 56916 71604
rect 57124 71590 57206 71604
rect 58082 71590 58164 71604
rect 58372 71590 58454 71604
rect 16418 71542 58934 71590
rect 16418 71446 58934 71494
rect 16898 71432 16980 71446
rect 17188 71432 17270 71446
rect 18146 71432 18228 71446
rect 18436 71432 18518 71446
rect 19394 71432 19476 71446
rect 19684 71432 19766 71446
rect 20642 71432 20724 71446
rect 20932 71432 21014 71446
rect 21890 71432 21972 71446
rect 22180 71432 22262 71446
rect 23138 71432 23220 71446
rect 23428 71432 23510 71446
rect 24386 71432 24468 71446
rect 24676 71432 24758 71446
rect 25634 71432 25716 71446
rect 25924 71432 26006 71446
rect 26882 71432 26964 71446
rect 27172 71432 27254 71446
rect 28130 71432 28212 71446
rect 28420 71432 28502 71446
rect 29378 71432 29460 71446
rect 29668 71432 29750 71446
rect 30626 71432 30708 71446
rect 30916 71432 30998 71446
rect 31874 71432 31956 71446
rect 32164 71432 32246 71446
rect 33122 71432 33204 71446
rect 33412 71432 33494 71446
rect 34370 71432 34452 71446
rect 34660 71432 34742 71446
rect 35618 71432 35700 71446
rect 35908 71432 35990 71446
rect 36866 71432 36948 71446
rect 37156 71432 37238 71446
rect 38114 71432 38196 71446
rect 38404 71432 38486 71446
rect 39362 71432 39444 71446
rect 39652 71432 39734 71446
rect 40610 71432 40692 71446
rect 40900 71432 40982 71446
rect 41858 71432 41940 71446
rect 42148 71432 42230 71446
rect 43106 71432 43188 71446
rect 43396 71432 43478 71446
rect 44354 71432 44436 71446
rect 44644 71432 44726 71446
rect 45602 71432 45684 71446
rect 45892 71432 45974 71446
rect 46850 71432 46932 71446
rect 47140 71432 47222 71446
rect 48098 71432 48180 71446
rect 48388 71432 48470 71446
rect 49346 71432 49428 71446
rect 49636 71432 49718 71446
rect 50594 71432 50676 71446
rect 50884 71432 50966 71446
rect 51842 71432 51924 71446
rect 52132 71432 52214 71446
rect 53090 71432 53172 71446
rect 53380 71432 53462 71446
rect 54338 71432 54420 71446
rect 54628 71432 54710 71446
rect 55586 71432 55668 71446
rect 55876 71432 55958 71446
rect 56834 71432 56916 71446
rect 57124 71432 57206 71446
rect 58082 71432 58164 71446
rect 58372 71432 58454 71446
rect 16418 71384 16864 71398
rect 17014 71384 17154 71398
rect 17304 71384 18112 71398
rect 18262 71384 18402 71398
rect 18552 71384 19360 71398
rect 19510 71384 19650 71398
rect 19800 71384 20608 71398
rect 20758 71384 20898 71398
rect 21048 71384 21856 71398
rect 22006 71384 22146 71398
rect 22296 71384 23104 71398
rect 23254 71384 23394 71398
rect 23544 71384 24352 71398
rect 24502 71384 24642 71398
rect 24792 71384 25600 71398
rect 25750 71384 25890 71398
rect 26040 71384 26848 71398
rect 26998 71384 27138 71398
rect 27288 71384 28096 71398
rect 28246 71384 28386 71398
rect 28536 71384 29344 71398
rect 29494 71384 29634 71398
rect 29784 71384 30592 71398
rect 30742 71384 30882 71398
rect 31032 71384 31840 71398
rect 31990 71384 32130 71398
rect 32280 71384 33088 71398
rect 33238 71384 33378 71398
rect 33528 71384 34336 71398
rect 34486 71384 34626 71398
rect 34776 71384 35584 71398
rect 35734 71384 35874 71398
rect 36024 71384 36832 71398
rect 36982 71384 37122 71398
rect 37272 71384 38080 71398
rect 38230 71384 38370 71398
rect 38520 71384 39328 71398
rect 39478 71384 39618 71398
rect 39768 71384 40576 71398
rect 40726 71384 40866 71398
rect 41016 71384 41824 71398
rect 41974 71384 42114 71398
rect 42264 71384 43072 71398
rect 43222 71384 43362 71398
rect 43512 71384 44320 71398
rect 44470 71384 44610 71398
rect 44760 71384 45568 71398
rect 45718 71384 45858 71398
rect 46008 71384 46816 71398
rect 46966 71384 47106 71398
rect 47256 71384 48064 71398
rect 48214 71384 48354 71398
rect 48504 71384 49312 71398
rect 49462 71384 49602 71398
rect 49752 71384 50560 71398
rect 50710 71384 50850 71398
rect 51000 71384 51808 71398
rect 51958 71384 52098 71398
rect 52248 71384 53056 71398
rect 53206 71384 53346 71398
rect 53496 71384 54304 71398
rect 54454 71384 54594 71398
rect 54744 71384 55552 71398
rect 55702 71384 55842 71398
rect 55992 71384 56800 71398
rect 56950 71384 57090 71398
rect 57240 71384 58048 71398
rect 58198 71384 58338 71398
rect 58488 71384 58934 71398
rect 16418 71336 58934 71384
rect 16418 71322 16864 71336
rect 17014 71322 17154 71336
rect 17304 71322 18112 71336
rect 18262 71322 18402 71336
rect 18552 71322 19360 71336
rect 19510 71322 19650 71336
rect 19800 71322 20608 71336
rect 20758 71322 20898 71336
rect 21048 71322 21856 71336
rect 22006 71322 22146 71336
rect 22296 71322 23104 71336
rect 23254 71322 23394 71336
rect 23544 71322 24352 71336
rect 24502 71322 24642 71336
rect 24792 71322 25600 71336
rect 25750 71322 25890 71336
rect 26040 71322 26848 71336
rect 26998 71322 27138 71336
rect 27288 71322 28096 71336
rect 28246 71322 28386 71336
rect 28536 71322 29344 71336
rect 29494 71322 29634 71336
rect 29784 71322 30592 71336
rect 30742 71322 30882 71336
rect 31032 71322 31840 71336
rect 31990 71322 32130 71336
rect 32280 71322 33088 71336
rect 33238 71322 33378 71336
rect 33528 71322 34336 71336
rect 34486 71322 34626 71336
rect 34776 71322 35584 71336
rect 35734 71322 35874 71336
rect 36024 71322 36832 71336
rect 36982 71322 37122 71336
rect 37272 71322 38080 71336
rect 38230 71322 38370 71336
rect 38520 71322 39328 71336
rect 39478 71322 39618 71336
rect 39768 71322 40576 71336
rect 40726 71322 40866 71336
rect 41016 71322 41824 71336
rect 41974 71322 42114 71336
rect 42264 71322 43072 71336
rect 43222 71322 43362 71336
rect 43512 71322 44320 71336
rect 44470 71322 44610 71336
rect 44760 71322 45568 71336
rect 45718 71322 45858 71336
rect 46008 71322 46816 71336
rect 46966 71322 47106 71336
rect 47256 71322 48064 71336
rect 48214 71322 48354 71336
rect 48504 71322 49312 71336
rect 49462 71322 49602 71336
rect 49752 71322 50560 71336
rect 50710 71322 50850 71336
rect 51000 71322 51808 71336
rect 51958 71322 52098 71336
rect 52248 71322 53056 71336
rect 53206 71322 53346 71336
rect 53496 71322 54304 71336
rect 54454 71322 54594 71336
rect 54744 71322 55552 71336
rect 55702 71322 55842 71336
rect 55992 71322 56800 71336
rect 56950 71322 57090 71336
rect 57240 71322 58048 71336
rect 58198 71322 58338 71336
rect 58488 71322 58934 71336
rect 16898 71274 16980 71288
rect 17188 71274 17270 71288
rect 18146 71274 18228 71288
rect 18436 71274 18518 71288
rect 19394 71274 19476 71288
rect 19684 71274 19766 71288
rect 20642 71274 20724 71288
rect 20932 71274 21014 71288
rect 21890 71274 21972 71288
rect 22180 71274 22262 71288
rect 23138 71274 23220 71288
rect 23428 71274 23510 71288
rect 24386 71274 24468 71288
rect 24676 71274 24758 71288
rect 25634 71274 25716 71288
rect 25924 71274 26006 71288
rect 26882 71274 26964 71288
rect 27172 71274 27254 71288
rect 28130 71274 28212 71288
rect 28420 71274 28502 71288
rect 29378 71274 29460 71288
rect 29668 71274 29750 71288
rect 30626 71274 30708 71288
rect 30916 71274 30998 71288
rect 31874 71274 31956 71288
rect 32164 71274 32246 71288
rect 33122 71274 33204 71288
rect 33412 71274 33494 71288
rect 34370 71274 34452 71288
rect 34660 71274 34742 71288
rect 35618 71274 35700 71288
rect 35908 71274 35990 71288
rect 36866 71274 36948 71288
rect 37156 71274 37238 71288
rect 38114 71274 38196 71288
rect 38404 71274 38486 71288
rect 39362 71274 39444 71288
rect 39652 71274 39734 71288
rect 40610 71274 40692 71288
rect 40900 71274 40982 71288
rect 41858 71274 41940 71288
rect 42148 71274 42230 71288
rect 43106 71274 43188 71288
rect 43396 71274 43478 71288
rect 44354 71274 44436 71288
rect 44644 71274 44726 71288
rect 45602 71274 45684 71288
rect 45892 71274 45974 71288
rect 46850 71274 46932 71288
rect 47140 71274 47222 71288
rect 48098 71274 48180 71288
rect 48388 71274 48470 71288
rect 49346 71274 49428 71288
rect 49636 71274 49718 71288
rect 50594 71274 50676 71288
rect 50884 71274 50966 71288
rect 51842 71274 51924 71288
rect 52132 71274 52214 71288
rect 53090 71274 53172 71288
rect 53380 71274 53462 71288
rect 54338 71274 54420 71288
rect 54628 71274 54710 71288
rect 55586 71274 55668 71288
rect 55876 71274 55958 71288
rect 56834 71274 56916 71288
rect 57124 71274 57206 71288
rect 58082 71274 58164 71288
rect 58372 71274 58454 71288
rect 16418 71226 58934 71274
rect 16418 71068 58934 71178
rect 16418 70972 58934 71020
rect 16898 70958 16980 70972
rect 17188 70958 17270 70972
rect 18146 70958 18228 70972
rect 18436 70958 18518 70972
rect 19394 70958 19476 70972
rect 19684 70958 19766 70972
rect 20642 70958 20724 70972
rect 20932 70958 21014 70972
rect 21890 70958 21972 70972
rect 22180 70958 22262 70972
rect 23138 70958 23220 70972
rect 23428 70958 23510 70972
rect 24386 70958 24468 70972
rect 24676 70958 24758 70972
rect 25634 70958 25716 70972
rect 25924 70958 26006 70972
rect 26882 70958 26964 70972
rect 27172 70958 27254 70972
rect 28130 70958 28212 70972
rect 28420 70958 28502 70972
rect 29378 70958 29460 70972
rect 29668 70958 29750 70972
rect 30626 70958 30708 70972
rect 30916 70958 30998 70972
rect 31874 70958 31956 70972
rect 32164 70958 32246 70972
rect 33122 70958 33204 70972
rect 33412 70958 33494 70972
rect 34370 70958 34452 70972
rect 34660 70958 34742 70972
rect 35618 70958 35700 70972
rect 35908 70958 35990 70972
rect 36866 70958 36948 70972
rect 37156 70958 37238 70972
rect 38114 70958 38196 70972
rect 38404 70958 38486 70972
rect 39362 70958 39444 70972
rect 39652 70958 39734 70972
rect 40610 70958 40692 70972
rect 40900 70958 40982 70972
rect 41858 70958 41940 70972
rect 42148 70958 42230 70972
rect 43106 70958 43188 70972
rect 43396 70958 43478 70972
rect 44354 70958 44436 70972
rect 44644 70958 44726 70972
rect 45602 70958 45684 70972
rect 45892 70958 45974 70972
rect 46850 70958 46932 70972
rect 47140 70958 47222 70972
rect 48098 70958 48180 70972
rect 48388 70958 48470 70972
rect 49346 70958 49428 70972
rect 49636 70958 49718 70972
rect 50594 70958 50676 70972
rect 50884 70958 50966 70972
rect 51842 70958 51924 70972
rect 52132 70958 52214 70972
rect 53090 70958 53172 70972
rect 53380 70958 53462 70972
rect 54338 70958 54420 70972
rect 54628 70958 54710 70972
rect 55586 70958 55668 70972
rect 55876 70958 55958 70972
rect 56834 70958 56916 70972
rect 57124 70958 57206 70972
rect 58082 70958 58164 70972
rect 58372 70958 58454 70972
rect 16418 70910 16864 70924
rect 17014 70910 17154 70924
rect 17304 70910 18112 70924
rect 18262 70910 18402 70924
rect 18552 70910 19360 70924
rect 19510 70910 19650 70924
rect 19800 70910 20608 70924
rect 20758 70910 20898 70924
rect 21048 70910 21856 70924
rect 22006 70910 22146 70924
rect 22296 70910 23104 70924
rect 23254 70910 23394 70924
rect 23544 70910 24352 70924
rect 24502 70910 24642 70924
rect 24792 70910 25600 70924
rect 25750 70910 25890 70924
rect 26040 70910 26848 70924
rect 26998 70910 27138 70924
rect 27288 70910 28096 70924
rect 28246 70910 28386 70924
rect 28536 70910 29344 70924
rect 29494 70910 29634 70924
rect 29784 70910 30592 70924
rect 30742 70910 30882 70924
rect 31032 70910 31840 70924
rect 31990 70910 32130 70924
rect 32280 70910 33088 70924
rect 33238 70910 33378 70924
rect 33528 70910 34336 70924
rect 34486 70910 34626 70924
rect 34776 70910 35584 70924
rect 35734 70910 35874 70924
rect 36024 70910 36832 70924
rect 36982 70910 37122 70924
rect 37272 70910 38080 70924
rect 38230 70910 38370 70924
rect 38520 70910 39328 70924
rect 39478 70910 39618 70924
rect 39768 70910 40576 70924
rect 40726 70910 40866 70924
rect 41016 70910 41824 70924
rect 41974 70910 42114 70924
rect 42264 70910 43072 70924
rect 43222 70910 43362 70924
rect 43512 70910 44320 70924
rect 44470 70910 44610 70924
rect 44760 70910 45568 70924
rect 45718 70910 45858 70924
rect 46008 70910 46816 70924
rect 46966 70910 47106 70924
rect 47256 70910 48064 70924
rect 48214 70910 48354 70924
rect 48504 70910 49312 70924
rect 49462 70910 49602 70924
rect 49752 70910 50560 70924
rect 50710 70910 50850 70924
rect 51000 70910 51808 70924
rect 51958 70910 52098 70924
rect 52248 70910 53056 70924
rect 53206 70910 53346 70924
rect 53496 70910 54304 70924
rect 54454 70910 54594 70924
rect 54744 70910 55552 70924
rect 55702 70910 55842 70924
rect 55992 70910 56800 70924
rect 56950 70910 57090 70924
rect 57240 70910 58048 70924
rect 58198 70910 58338 70924
rect 58488 70910 58934 70924
rect 16418 70862 58934 70910
rect 16418 70848 16864 70862
rect 17014 70848 17154 70862
rect 17304 70848 18112 70862
rect 18262 70848 18402 70862
rect 18552 70848 19360 70862
rect 19510 70848 19650 70862
rect 19800 70848 20608 70862
rect 20758 70848 20898 70862
rect 21048 70848 21856 70862
rect 22006 70848 22146 70862
rect 22296 70848 23104 70862
rect 23254 70848 23394 70862
rect 23544 70848 24352 70862
rect 24502 70848 24642 70862
rect 24792 70848 25600 70862
rect 25750 70848 25890 70862
rect 26040 70848 26848 70862
rect 26998 70848 27138 70862
rect 27288 70848 28096 70862
rect 28246 70848 28386 70862
rect 28536 70848 29344 70862
rect 29494 70848 29634 70862
rect 29784 70848 30592 70862
rect 30742 70848 30882 70862
rect 31032 70848 31840 70862
rect 31990 70848 32130 70862
rect 32280 70848 33088 70862
rect 33238 70848 33378 70862
rect 33528 70848 34336 70862
rect 34486 70848 34626 70862
rect 34776 70848 35584 70862
rect 35734 70848 35874 70862
rect 36024 70848 36832 70862
rect 36982 70848 37122 70862
rect 37272 70848 38080 70862
rect 38230 70848 38370 70862
rect 38520 70848 39328 70862
rect 39478 70848 39618 70862
rect 39768 70848 40576 70862
rect 40726 70848 40866 70862
rect 41016 70848 41824 70862
rect 41974 70848 42114 70862
rect 42264 70848 43072 70862
rect 43222 70848 43362 70862
rect 43512 70848 44320 70862
rect 44470 70848 44610 70862
rect 44760 70848 45568 70862
rect 45718 70848 45858 70862
rect 46008 70848 46816 70862
rect 46966 70848 47106 70862
rect 47256 70848 48064 70862
rect 48214 70848 48354 70862
rect 48504 70848 49312 70862
rect 49462 70848 49602 70862
rect 49752 70848 50560 70862
rect 50710 70848 50850 70862
rect 51000 70848 51808 70862
rect 51958 70848 52098 70862
rect 52248 70848 53056 70862
rect 53206 70848 53346 70862
rect 53496 70848 54304 70862
rect 54454 70848 54594 70862
rect 54744 70848 55552 70862
rect 55702 70848 55842 70862
rect 55992 70848 56800 70862
rect 56950 70848 57090 70862
rect 57240 70848 58048 70862
rect 58198 70848 58338 70862
rect 58488 70848 58934 70862
rect 16898 70800 16980 70814
rect 17188 70800 17270 70814
rect 18146 70800 18228 70814
rect 18436 70800 18518 70814
rect 19394 70800 19476 70814
rect 19684 70800 19766 70814
rect 20642 70800 20724 70814
rect 20932 70800 21014 70814
rect 21890 70800 21972 70814
rect 22180 70800 22262 70814
rect 23138 70800 23220 70814
rect 23428 70800 23510 70814
rect 24386 70800 24468 70814
rect 24676 70800 24758 70814
rect 25634 70800 25716 70814
rect 25924 70800 26006 70814
rect 26882 70800 26964 70814
rect 27172 70800 27254 70814
rect 28130 70800 28212 70814
rect 28420 70800 28502 70814
rect 29378 70800 29460 70814
rect 29668 70800 29750 70814
rect 30626 70800 30708 70814
rect 30916 70800 30998 70814
rect 31874 70800 31956 70814
rect 32164 70800 32246 70814
rect 33122 70800 33204 70814
rect 33412 70800 33494 70814
rect 34370 70800 34452 70814
rect 34660 70800 34742 70814
rect 35618 70800 35700 70814
rect 35908 70800 35990 70814
rect 36866 70800 36948 70814
rect 37156 70800 37238 70814
rect 38114 70800 38196 70814
rect 38404 70800 38486 70814
rect 39362 70800 39444 70814
rect 39652 70800 39734 70814
rect 40610 70800 40692 70814
rect 40900 70800 40982 70814
rect 41858 70800 41940 70814
rect 42148 70800 42230 70814
rect 43106 70800 43188 70814
rect 43396 70800 43478 70814
rect 44354 70800 44436 70814
rect 44644 70800 44726 70814
rect 45602 70800 45684 70814
rect 45892 70800 45974 70814
rect 46850 70800 46932 70814
rect 47140 70800 47222 70814
rect 48098 70800 48180 70814
rect 48388 70800 48470 70814
rect 49346 70800 49428 70814
rect 49636 70800 49718 70814
rect 50594 70800 50676 70814
rect 50884 70800 50966 70814
rect 51842 70800 51924 70814
rect 52132 70800 52214 70814
rect 53090 70800 53172 70814
rect 53380 70800 53462 70814
rect 54338 70800 54420 70814
rect 54628 70800 54710 70814
rect 55586 70800 55668 70814
rect 55876 70800 55958 70814
rect 56834 70800 56916 70814
rect 57124 70800 57206 70814
rect 58082 70800 58164 70814
rect 58372 70800 58454 70814
rect 16418 70752 58934 70800
rect 16418 70656 58934 70704
rect 16898 70642 16980 70656
rect 17188 70642 17270 70656
rect 18146 70642 18228 70656
rect 18436 70642 18518 70656
rect 19394 70642 19476 70656
rect 19684 70642 19766 70656
rect 20642 70642 20724 70656
rect 20932 70642 21014 70656
rect 21890 70642 21972 70656
rect 22180 70642 22262 70656
rect 23138 70642 23220 70656
rect 23428 70642 23510 70656
rect 24386 70642 24468 70656
rect 24676 70642 24758 70656
rect 25634 70642 25716 70656
rect 25924 70642 26006 70656
rect 26882 70642 26964 70656
rect 27172 70642 27254 70656
rect 28130 70642 28212 70656
rect 28420 70642 28502 70656
rect 29378 70642 29460 70656
rect 29668 70642 29750 70656
rect 30626 70642 30708 70656
rect 30916 70642 30998 70656
rect 31874 70642 31956 70656
rect 32164 70642 32246 70656
rect 33122 70642 33204 70656
rect 33412 70642 33494 70656
rect 34370 70642 34452 70656
rect 34660 70642 34742 70656
rect 35618 70642 35700 70656
rect 35908 70642 35990 70656
rect 36866 70642 36948 70656
rect 37156 70642 37238 70656
rect 38114 70642 38196 70656
rect 38404 70642 38486 70656
rect 39362 70642 39444 70656
rect 39652 70642 39734 70656
rect 40610 70642 40692 70656
rect 40900 70642 40982 70656
rect 41858 70642 41940 70656
rect 42148 70642 42230 70656
rect 43106 70642 43188 70656
rect 43396 70642 43478 70656
rect 44354 70642 44436 70656
rect 44644 70642 44726 70656
rect 45602 70642 45684 70656
rect 45892 70642 45974 70656
rect 46850 70642 46932 70656
rect 47140 70642 47222 70656
rect 48098 70642 48180 70656
rect 48388 70642 48470 70656
rect 49346 70642 49428 70656
rect 49636 70642 49718 70656
rect 50594 70642 50676 70656
rect 50884 70642 50966 70656
rect 51842 70642 51924 70656
rect 52132 70642 52214 70656
rect 53090 70642 53172 70656
rect 53380 70642 53462 70656
rect 54338 70642 54420 70656
rect 54628 70642 54710 70656
rect 55586 70642 55668 70656
rect 55876 70642 55958 70656
rect 56834 70642 56916 70656
rect 57124 70642 57206 70656
rect 58082 70642 58164 70656
rect 58372 70642 58454 70656
rect 16418 70594 16864 70608
rect 17014 70594 17154 70608
rect 17304 70594 18112 70608
rect 18262 70594 18402 70608
rect 18552 70594 19360 70608
rect 19510 70594 19650 70608
rect 19800 70594 20608 70608
rect 20758 70594 20898 70608
rect 21048 70594 21856 70608
rect 22006 70594 22146 70608
rect 22296 70594 23104 70608
rect 23254 70594 23394 70608
rect 23544 70594 24352 70608
rect 24502 70594 24642 70608
rect 24792 70594 25600 70608
rect 25750 70594 25890 70608
rect 26040 70594 26848 70608
rect 26998 70594 27138 70608
rect 27288 70594 28096 70608
rect 28246 70594 28386 70608
rect 28536 70594 29344 70608
rect 29494 70594 29634 70608
rect 29784 70594 30592 70608
rect 30742 70594 30882 70608
rect 31032 70594 31840 70608
rect 31990 70594 32130 70608
rect 32280 70594 33088 70608
rect 33238 70594 33378 70608
rect 33528 70594 34336 70608
rect 34486 70594 34626 70608
rect 34776 70594 35584 70608
rect 35734 70594 35874 70608
rect 36024 70594 36832 70608
rect 36982 70594 37122 70608
rect 37272 70594 38080 70608
rect 38230 70594 38370 70608
rect 38520 70594 39328 70608
rect 39478 70594 39618 70608
rect 39768 70594 40576 70608
rect 40726 70594 40866 70608
rect 41016 70594 41824 70608
rect 41974 70594 42114 70608
rect 42264 70594 43072 70608
rect 43222 70594 43362 70608
rect 43512 70594 44320 70608
rect 44470 70594 44610 70608
rect 44760 70594 45568 70608
rect 45718 70594 45858 70608
rect 46008 70594 46816 70608
rect 46966 70594 47106 70608
rect 47256 70594 48064 70608
rect 48214 70594 48354 70608
rect 48504 70594 49312 70608
rect 49462 70594 49602 70608
rect 49752 70594 50560 70608
rect 50710 70594 50850 70608
rect 51000 70594 51808 70608
rect 51958 70594 52098 70608
rect 52248 70594 53056 70608
rect 53206 70594 53346 70608
rect 53496 70594 54304 70608
rect 54454 70594 54594 70608
rect 54744 70594 55552 70608
rect 55702 70594 55842 70608
rect 55992 70594 56800 70608
rect 56950 70594 57090 70608
rect 57240 70594 58048 70608
rect 58198 70594 58338 70608
rect 58488 70594 58934 70608
rect 16418 70546 58934 70594
rect 16418 70532 16864 70546
rect 17014 70532 17154 70546
rect 17304 70532 18112 70546
rect 18262 70532 18402 70546
rect 18552 70532 19360 70546
rect 19510 70532 19650 70546
rect 19800 70532 20608 70546
rect 20758 70532 20898 70546
rect 21048 70532 21856 70546
rect 22006 70532 22146 70546
rect 22296 70532 23104 70546
rect 23254 70532 23394 70546
rect 23544 70532 24352 70546
rect 24502 70532 24642 70546
rect 24792 70532 25600 70546
rect 25750 70532 25890 70546
rect 26040 70532 26848 70546
rect 26998 70532 27138 70546
rect 27288 70532 28096 70546
rect 28246 70532 28386 70546
rect 28536 70532 29344 70546
rect 29494 70532 29634 70546
rect 29784 70532 30592 70546
rect 30742 70532 30882 70546
rect 31032 70532 31840 70546
rect 31990 70532 32130 70546
rect 32280 70532 33088 70546
rect 33238 70532 33378 70546
rect 33528 70532 34336 70546
rect 34486 70532 34626 70546
rect 34776 70532 35584 70546
rect 35734 70532 35874 70546
rect 36024 70532 36832 70546
rect 36982 70532 37122 70546
rect 37272 70532 38080 70546
rect 38230 70532 38370 70546
rect 38520 70532 39328 70546
rect 39478 70532 39618 70546
rect 39768 70532 40576 70546
rect 40726 70532 40866 70546
rect 41016 70532 41824 70546
rect 41974 70532 42114 70546
rect 42264 70532 43072 70546
rect 43222 70532 43362 70546
rect 43512 70532 44320 70546
rect 44470 70532 44610 70546
rect 44760 70532 45568 70546
rect 45718 70532 45858 70546
rect 46008 70532 46816 70546
rect 46966 70532 47106 70546
rect 47256 70532 48064 70546
rect 48214 70532 48354 70546
rect 48504 70532 49312 70546
rect 49462 70532 49602 70546
rect 49752 70532 50560 70546
rect 50710 70532 50850 70546
rect 51000 70532 51808 70546
rect 51958 70532 52098 70546
rect 52248 70532 53056 70546
rect 53206 70532 53346 70546
rect 53496 70532 54304 70546
rect 54454 70532 54594 70546
rect 54744 70532 55552 70546
rect 55702 70532 55842 70546
rect 55992 70532 56800 70546
rect 56950 70532 57090 70546
rect 57240 70532 58048 70546
rect 58198 70532 58338 70546
rect 58488 70532 58934 70546
rect 16898 70484 16980 70498
rect 17188 70484 17270 70498
rect 18146 70484 18228 70498
rect 18436 70484 18518 70498
rect 19394 70484 19476 70498
rect 19684 70484 19766 70498
rect 20642 70484 20724 70498
rect 20932 70484 21014 70498
rect 21890 70484 21972 70498
rect 22180 70484 22262 70498
rect 23138 70484 23220 70498
rect 23428 70484 23510 70498
rect 24386 70484 24468 70498
rect 24676 70484 24758 70498
rect 25634 70484 25716 70498
rect 25924 70484 26006 70498
rect 26882 70484 26964 70498
rect 27172 70484 27254 70498
rect 28130 70484 28212 70498
rect 28420 70484 28502 70498
rect 29378 70484 29460 70498
rect 29668 70484 29750 70498
rect 30626 70484 30708 70498
rect 30916 70484 30998 70498
rect 31874 70484 31956 70498
rect 32164 70484 32246 70498
rect 33122 70484 33204 70498
rect 33412 70484 33494 70498
rect 34370 70484 34452 70498
rect 34660 70484 34742 70498
rect 35618 70484 35700 70498
rect 35908 70484 35990 70498
rect 36866 70484 36948 70498
rect 37156 70484 37238 70498
rect 38114 70484 38196 70498
rect 38404 70484 38486 70498
rect 39362 70484 39444 70498
rect 39652 70484 39734 70498
rect 40610 70484 40692 70498
rect 40900 70484 40982 70498
rect 41858 70484 41940 70498
rect 42148 70484 42230 70498
rect 43106 70484 43188 70498
rect 43396 70484 43478 70498
rect 44354 70484 44436 70498
rect 44644 70484 44726 70498
rect 45602 70484 45684 70498
rect 45892 70484 45974 70498
rect 46850 70484 46932 70498
rect 47140 70484 47222 70498
rect 48098 70484 48180 70498
rect 48388 70484 48470 70498
rect 49346 70484 49428 70498
rect 49636 70484 49718 70498
rect 50594 70484 50676 70498
rect 50884 70484 50966 70498
rect 51842 70484 51924 70498
rect 52132 70484 52214 70498
rect 53090 70484 53172 70498
rect 53380 70484 53462 70498
rect 54338 70484 54420 70498
rect 54628 70484 54710 70498
rect 55586 70484 55668 70498
rect 55876 70484 55958 70498
rect 56834 70484 56916 70498
rect 57124 70484 57206 70498
rect 58082 70484 58164 70498
rect 58372 70484 58454 70498
rect 16418 70436 58934 70484
rect 16418 70278 58934 70388
rect 16418 70182 58934 70230
rect 16898 70168 16980 70182
rect 17188 70168 17270 70182
rect 18146 70168 18228 70182
rect 18436 70168 18518 70182
rect 19394 70168 19476 70182
rect 19684 70168 19766 70182
rect 20642 70168 20724 70182
rect 20932 70168 21014 70182
rect 21890 70168 21972 70182
rect 22180 70168 22262 70182
rect 23138 70168 23220 70182
rect 23428 70168 23510 70182
rect 24386 70168 24468 70182
rect 24676 70168 24758 70182
rect 25634 70168 25716 70182
rect 25924 70168 26006 70182
rect 26882 70168 26964 70182
rect 27172 70168 27254 70182
rect 28130 70168 28212 70182
rect 28420 70168 28502 70182
rect 29378 70168 29460 70182
rect 29668 70168 29750 70182
rect 30626 70168 30708 70182
rect 30916 70168 30998 70182
rect 31874 70168 31956 70182
rect 32164 70168 32246 70182
rect 33122 70168 33204 70182
rect 33412 70168 33494 70182
rect 34370 70168 34452 70182
rect 34660 70168 34742 70182
rect 35618 70168 35700 70182
rect 35908 70168 35990 70182
rect 36866 70168 36948 70182
rect 37156 70168 37238 70182
rect 38114 70168 38196 70182
rect 38404 70168 38486 70182
rect 39362 70168 39444 70182
rect 39652 70168 39734 70182
rect 40610 70168 40692 70182
rect 40900 70168 40982 70182
rect 41858 70168 41940 70182
rect 42148 70168 42230 70182
rect 43106 70168 43188 70182
rect 43396 70168 43478 70182
rect 44354 70168 44436 70182
rect 44644 70168 44726 70182
rect 45602 70168 45684 70182
rect 45892 70168 45974 70182
rect 46850 70168 46932 70182
rect 47140 70168 47222 70182
rect 48098 70168 48180 70182
rect 48388 70168 48470 70182
rect 49346 70168 49428 70182
rect 49636 70168 49718 70182
rect 50594 70168 50676 70182
rect 50884 70168 50966 70182
rect 51842 70168 51924 70182
rect 52132 70168 52214 70182
rect 53090 70168 53172 70182
rect 53380 70168 53462 70182
rect 54338 70168 54420 70182
rect 54628 70168 54710 70182
rect 55586 70168 55668 70182
rect 55876 70168 55958 70182
rect 56834 70168 56916 70182
rect 57124 70168 57206 70182
rect 58082 70168 58164 70182
rect 58372 70168 58454 70182
rect 16418 70120 16864 70134
rect 17014 70120 17154 70134
rect 17304 70120 18112 70134
rect 18262 70120 18402 70134
rect 18552 70120 19360 70134
rect 19510 70120 19650 70134
rect 19800 70120 20608 70134
rect 20758 70120 20898 70134
rect 21048 70120 21856 70134
rect 22006 70120 22146 70134
rect 22296 70120 23104 70134
rect 23254 70120 23394 70134
rect 23544 70120 24352 70134
rect 24502 70120 24642 70134
rect 24792 70120 25600 70134
rect 25750 70120 25890 70134
rect 26040 70120 26848 70134
rect 26998 70120 27138 70134
rect 27288 70120 28096 70134
rect 28246 70120 28386 70134
rect 28536 70120 29344 70134
rect 29494 70120 29634 70134
rect 29784 70120 30592 70134
rect 30742 70120 30882 70134
rect 31032 70120 31840 70134
rect 31990 70120 32130 70134
rect 32280 70120 33088 70134
rect 33238 70120 33378 70134
rect 33528 70120 34336 70134
rect 34486 70120 34626 70134
rect 34776 70120 35584 70134
rect 35734 70120 35874 70134
rect 36024 70120 36832 70134
rect 36982 70120 37122 70134
rect 37272 70120 38080 70134
rect 38230 70120 38370 70134
rect 38520 70120 39328 70134
rect 39478 70120 39618 70134
rect 39768 70120 40576 70134
rect 40726 70120 40866 70134
rect 41016 70120 41824 70134
rect 41974 70120 42114 70134
rect 42264 70120 43072 70134
rect 43222 70120 43362 70134
rect 43512 70120 44320 70134
rect 44470 70120 44610 70134
rect 44760 70120 45568 70134
rect 45718 70120 45858 70134
rect 46008 70120 46816 70134
rect 46966 70120 47106 70134
rect 47256 70120 48064 70134
rect 48214 70120 48354 70134
rect 48504 70120 49312 70134
rect 49462 70120 49602 70134
rect 49752 70120 50560 70134
rect 50710 70120 50850 70134
rect 51000 70120 51808 70134
rect 51958 70120 52098 70134
rect 52248 70120 53056 70134
rect 53206 70120 53346 70134
rect 53496 70120 54304 70134
rect 54454 70120 54594 70134
rect 54744 70120 55552 70134
rect 55702 70120 55842 70134
rect 55992 70120 56800 70134
rect 56950 70120 57090 70134
rect 57240 70120 58048 70134
rect 58198 70120 58338 70134
rect 58488 70120 58934 70134
rect 16418 70072 58934 70120
rect 16418 70058 16864 70072
rect 17014 70058 17154 70072
rect 17304 70058 18112 70072
rect 18262 70058 18402 70072
rect 18552 70058 19360 70072
rect 19510 70058 19650 70072
rect 19800 70058 20608 70072
rect 20758 70058 20898 70072
rect 21048 70058 21856 70072
rect 22006 70058 22146 70072
rect 22296 70058 23104 70072
rect 23254 70058 23394 70072
rect 23544 70058 24352 70072
rect 24502 70058 24642 70072
rect 24792 70058 25600 70072
rect 25750 70058 25890 70072
rect 26040 70058 26848 70072
rect 26998 70058 27138 70072
rect 27288 70058 28096 70072
rect 28246 70058 28386 70072
rect 28536 70058 29344 70072
rect 29494 70058 29634 70072
rect 29784 70058 30592 70072
rect 30742 70058 30882 70072
rect 31032 70058 31840 70072
rect 31990 70058 32130 70072
rect 32280 70058 33088 70072
rect 33238 70058 33378 70072
rect 33528 70058 34336 70072
rect 34486 70058 34626 70072
rect 34776 70058 35584 70072
rect 35734 70058 35874 70072
rect 36024 70058 36832 70072
rect 36982 70058 37122 70072
rect 37272 70058 38080 70072
rect 38230 70058 38370 70072
rect 38520 70058 39328 70072
rect 39478 70058 39618 70072
rect 39768 70058 40576 70072
rect 40726 70058 40866 70072
rect 41016 70058 41824 70072
rect 41974 70058 42114 70072
rect 42264 70058 43072 70072
rect 43222 70058 43362 70072
rect 43512 70058 44320 70072
rect 44470 70058 44610 70072
rect 44760 70058 45568 70072
rect 45718 70058 45858 70072
rect 46008 70058 46816 70072
rect 46966 70058 47106 70072
rect 47256 70058 48064 70072
rect 48214 70058 48354 70072
rect 48504 70058 49312 70072
rect 49462 70058 49602 70072
rect 49752 70058 50560 70072
rect 50710 70058 50850 70072
rect 51000 70058 51808 70072
rect 51958 70058 52098 70072
rect 52248 70058 53056 70072
rect 53206 70058 53346 70072
rect 53496 70058 54304 70072
rect 54454 70058 54594 70072
rect 54744 70058 55552 70072
rect 55702 70058 55842 70072
rect 55992 70058 56800 70072
rect 56950 70058 57090 70072
rect 57240 70058 58048 70072
rect 58198 70058 58338 70072
rect 58488 70058 58934 70072
rect 16898 70010 16980 70024
rect 17188 70010 17270 70024
rect 18146 70010 18228 70024
rect 18436 70010 18518 70024
rect 19394 70010 19476 70024
rect 19684 70010 19766 70024
rect 20642 70010 20724 70024
rect 20932 70010 21014 70024
rect 21890 70010 21972 70024
rect 22180 70010 22262 70024
rect 23138 70010 23220 70024
rect 23428 70010 23510 70024
rect 24386 70010 24468 70024
rect 24676 70010 24758 70024
rect 25634 70010 25716 70024
rect 25924 70010 26006 70024
rect 26882 70010 26964 70024
rect 27172 70010 27254 70024
rect 28130 70010 28212 70024
rect 28420 70010 28502 70024
rect 29378 70010 29460 70024
rect 29668 70010 29750 70024
rect 30626 70010 30708 70024
rect 30916 70010 30998 70024
rect 31874 70010 31956 70024
rect 32164 70010 32246 70024
rect 33122 70010 33204 70024
rect 33412 70010 33494 70024
rect 34370 70010 34452 70024
rect 34660 70010 34742 70024
rect 35618 70010 35700 70024
rect 35908 70010 35990 70024
rect 36866 70010 36948 70024
rect 37156 70010 37238 70024
rect 38114 70010 38196 70024
rect 38404 70010 38486 70024
rect 39362 70010 39444 70024
rect 39652 70010 39734 70024
rect 40610 70010 40692 70024
rect 40900 70010 40982 70024
rect 41858 70010 41940 70024
rect 42148 70010 42230 70024
rect 43106 70010 43188 70024
rect 43396 70010 43478 70024
rect 44354 70010 44436 70024
rect 44644 70010 44726 70024
rect 45602 70010 45684 70024
rect 45892 70010 45974 70024
rect 46850 70010 46932 70024
rect 47140 70010 47222 70024
rect 48098 70010 48180 70024
rect 48388 70010 48470 70024
rect 49346 70010 49428 70024
rect 49636 70010 49718 70024
rect 50594 70010 50676 70024
rect 50884 70010 50966 70024
rect 51842 70010 51924 70024
rect 52132 70010 52214 70024
rect 53090 70010 53172 70024
rect 53380 70010 53462 70024
rect 54338 70010 54420 70024
rect 54628 70010 54710 70024
rect 55586 70010 55668 70024
rect 55876 70010 55958 70024
rect 56834 70010 56916 70024
rect 57124 70010 57206 70024
rect 58082 70010 58164 70024
rect 58372 70010 58454 70024
rect 16418 69962 58934 70010
rect 16418 69866 58934 69914
rect 16898 69852 16980 69866
rect 17188 69852 17270 69866
rect 18146 69852 18228 69866
rect 18436 69852 18518 69866
rect 19394 69852 19476 69866
rect 19684 69852 19766 69866
rect 20642 69852 20724 69866
rect 20932 69852 21014 69866
rect 21890 69852 21972 69866
rect 22180 69852 22262 69866
rect 23138 69852 23220 69866
rect 23428 69852 23510 69866
rect 24386 69852 24468 69866
rect 24676 69852 24758 69866
rect 25634 69852 25716 69866
rect 25924 69852 26006 69866
rect 26882 69852 26964 69866
rect 27172 69852 27254 69866
rect 28130 69852 28212 69866
rect 28420 69852 28502 69866
rect 29378 69852 29460 69866
rect 29668 69852 29750 69866
rect 30626 69852 30708 69866
rect 30916 69852 30998 69866
rect 31874 69852 31956 69866
rect 32164 69852 32246 69866
rect 33122 69852 33204 69866
rect 33412 69852 33494 69866
rect 34370 69852 34452 69866
rect 34660 69852 34742 69866
rect 35618 69852 35700 69866
rect 35908 69852 35990 69866
rect 36866 69852 36948 69866
rect 37156 69852 37238 69866
rect 38114 69852 38196 69866
rect 38404 69852 38486 69866
rect 39362 69852 39444 69866
rect 39652 69852 39734 69866
rect 40610 69852 40692 69866
rect 40900 69852 40982 69866
rect 41858 69852 41940 69866
rect 42148 69852 42230 69866
rect 43106 69852 43188 69866
rect 43396 69852 43478 69866
rect 44354 69852 44436 69866
rect 44644 69852 44726 69866
rect 45602 69852 45684 69866
rect 45892 69852 45974 69866
rect 46850 69852 46932 69866
rect 47140 69852 47222 69866
rect 48098 69852 48180 69866
rect 48388 69852 48470 69866
rect 49346 69852 49428 69866
rect 49636 69852 49718 69866
rect 50594 69852 50676 69866
rect 50884 69852 50966 69866
rect 51842 69852 51924 69866
rect 52132 69852 52214 69866
rect 53090 69852 53172 69866
rect 53380 69852 53462 69866
rect 54338 69852 54420 69866
rect 54628 69852 54710 69866
rect 55586 69852 55668 69866
rect 55876 69852 55958 69866
rect 56834 69852 56916 69866
rect 57124 69852 57206 69866
rect 58082 69852 58164 69866
rect 58372 69852 58454 69866
rect 16418 69804 16864 69818
rect 17014 69804 17154 69818
rect 17304 69804 18112 69818
rect 18262 69804 18402 69818
rect 18552 69804 19360 69818
rect 19510 69804 19650 69818
rect 19800 69804 20608 69818
rect 20758 69804 20898 69818
rect 21048 69804 21856 69818
rect 22006 69804 22146 69818
rect 22296 69804 23104 69818
rect 23254 69804 23394 69818
rect 23544 69804 24352 69818
rect 24502 69804 24642 69818
rect 24792 69804 25600 69818
rect 25750 69804 25890 69818
rect 26040 69804 26848 69818
rect 26998 69804 27138 69818
rect 27288 69804 28096 69818
rect 28246 69804 28386 69818
rect 28536 69804 29344 69818
rect 29494 69804 29634 69818
rect 29784 69804 30592 69818
rect 30742 69804 30882 69818
rect 31032 69804 31840 69818
rect 31990 69804 32130 69818
rect 32280 69804 33088 69818
rect 33238 69804 33378 69818
rect 33528 69804 34336 69818
rect 34486 69804 34626 69818
rect 34776 69804 35584 69818
rect 35734 69804 35874 69818
rect 36024 69804 36832 69818
rect 36982 69804 37122 69818
rect 37272 69804 38080 69818
rect 38230 69804 38370 69818
rect 38520 69804 39328 69818
rect 39478 69804 39618 69818
rect 39768 69804 40576 69818
rect 40726 69804 40866 69818
rect 41016 69804 41824 69818
rect 41974 69804 42114 69818
rect 42264 69804 43072 69818
rect 43222 69804 43362 69818
rect 43512 69804 44320 69818
rect 44470 69804 44610 69818
rect 44760 69804 45568 69818
rect 45718 69804 45858 69818
rect 46008 69804 46816 69818
rect 46966 69804 47106 69818
rect 47256 69804 48064 69818
rect 48214 69804 48354 69818
rect 48504 69804 49312 69818
rect 49462 69804 49602 69818
rect 49752 69804 50560 69818
rect 50710 69804 50850 69818
rect 51000 69804 51808 69818
rect 51958 69804 52098 69818
rect 52248 69804 53056 69818
rect 53206 69804 53346 69818
rect 53496 69804 54304 69818
rect 54454 69804 54594 69818
rect 54744 69804 55552 69818
rect 55702 69804 55842 69818
rect 55992 69804 56800 69818
rect 56950 69804 57090 69818
rect 57240 69804 58048 69818
rect 58198 69804 58338 69818
rect 58488 69804 58934 69818
rect 16418 69756 58934 69804
rect 16418 69742 16864 69756
rect 17014 69742 17154 69756
rect 17304 69742 18112 69756
rect 18262 69742 18402 69756
rect 18552 69742 19360 69756
rect 19510 69742 19650 69756
rect 19800 69742 20608 69756
rect 20758 69742 20898 69756
rect 21048 69742 21856 69756
rect 22006 69742 22146 69756
rect 22296 69742 23104 69756
rect 23254 69742 23394 69756
rect 23544 69742 24352 69756
rect 24502 69742 24642 69756
rect 24792 69742 25600 69756
rect 25750 69742 25890 69756
rect 26040 69742 26848 69756
rect 26998 69742 27138 69756
rect 27288 69742 28096 69756
rect 28246 69742 28386 69756
rect 28536 69742 29344 69756
rect 29494 69742 29634 69756
rect 29784 69742 30592 69756
rect 30742 69742 30882 69756
rect 31032 69742 31840 69756
rect 31990 69742 32130 69756
rect 32280 69742 33088 69756
rect 33238 69742 33378 69756
rect 33528 69742 34336 69756
rect 34486 69742 34626 69756
rect 34776 69742 35584 69756
rect 35734 69742 35874 69756
rect 36024 69742 36832 69756
rect 36982 69742 37122 69756
rect 37272 69742 38080 69756
rect 38230 69742 38370 69756
rect 38520 69742 39328 69756
rect 39478 69742 39618 69756
rect 39768 69742 40576 69756
rect 40726 69742 40866 69756
rect 41016 69742 41824 69756
rect 41974 69742 42114 69756
rect 42264 69742 43072 69756
rect 43222 69742 43362 69756
rect 43512 69742 44320 69756
rect 44470 69742 44610 69756
rect 44760 69742 45568 69756
rect 45718 69742 45858 69756
rect 46008 69742 46816 69756
rect 46966 69742 47106 69756
rect 47256 69742 48064 69756
rect 48214 69742 48354 69756
rect 48504 69742 49312 69756
rect 49462 69742 49602 69756
rect 49752 69742 50560 69756
rect 50710 69742 50850 69756
rect 51000 69742 51808 69756
rect 51958 69742 52098 69756
rect 52248 69742 53056 69756
rect 53206 69742 53346 69756
rect 53496 69742 54304 69756
rect 54454 69742 54594 69756
rect 54744 69742 55552 69756
rect 55702 69742 55842 69756
rect 55992 69742 56800 69756
rect 56950 69742 57090 69756
rect 57240 69742 58048 69756
rect 58198 69742 58338 69756
rect 58488 69742 58934 69756
rect 16898 69694 16980 69708
rect 17188 69694 17270 69708
rect 18146 69694 18228 69708
rect 18436 69694 18518 69708
rect 19394 69694 19476 69708
rect 19684 69694 19766 69708
rect 20642 69694 20724 69708
rect 20932 69694 21014 69708
rect 21890 69694 21972 69708
rect 22180 69694 22262 69708
rect 23138 69694 23220 69708
rect 23428 69694 23510 69708
rect 24386 69694 24468 69708
rect 24676 69694 24758 69708
rect 25634 69694 25716 69708
rect 25924 69694 26006 69708
rect 26882 69694 26964 69708
rect 27172 69694 27254 69708
rect 28130 69694 28212 69708
rect 28420 69694 28502 69708
rect 29378 69694 29460 69708
rect 29668 69694 29750 69708
rect 30626 69694 30708 69708
rect 30916 69694 30998 69708
rect 31874 69694 31956 69708
rect 32164 69694 32246 69708
rect 33122 69694 33204 69708
rect 33412 69694 33494 69708
rect 34370 69694 34452 69708
rect 34660 69694 34742 69708
rect 35618 69694 35700 69708
rect 35908 69694 35990 69708
rect 36866 69694 36948 69708
rect 37156 69694 37238 69708
rect 38114 69694 38196 69708
rect 38404 69694 38486 69708
rect 39362 69694 39444 69708
rect 39652 69694 39734 69708
rect 40610 69694 40692 69708
rect 40900 69694 40982 69708
rect 41858 69694 41940 69708
rect 42148 69694 42230 69708
rect 43106 69694 43188 69708
rect 43396 69694 43478 69708
rect 44354 69694 44436 69708
rect 44644 69694 44726 69708
rect 45602 69694 45684 69708
rect 45892 69694 45974 69708
rect 46850 69694 46932 69708
rect 47140 69694 47222 69708
rect 48098 69694 48180 69708
rect 48388 69694 48470 69708
rect 49346 69694 49428 69708
rect 49636 69694 49718 69708
rect 50594 69694 50676 69708
rect 50884 69694 50966 69708
rect 51842 69694 51924 69708
rect 52132 69694 52214 69708
rect 53090 69694 53172 69708
rect 53380 69694 53462 69708
rect 54338 69694 54420 69708
rect 54628 69694 54710 69708
rect 55586 69694 55668 69708
rect 55876 69694 55958 69708
rect 56834 69694 56916 69708
rect 57124 69694 57206 69708
rect 58082 69694 58164 69708
rect 58372 69694 58454 69708
rect 16418 69646 58934 69694
rect 16418 69488 58934 69598
rect 16418 69392 58934 69440
rect 16898 69378 16980 69392
rect 17188 69378 17270 69392
rect 18146 69378 18228 69392
rect 18436 69378 18518 69392
rect 19394 69378 19476 69392
rect 19684 69378 19766 69392
rect 20642 69378 20724 69392
rect 20932 69378 21014 69392
rect 21890 69378 21972 69392
rect 22180 69378 22262 69392
rect 23138 69378 23220 69392
rect 23428 69378 23510 69392
rect 24386 69378 24468 69392
rect 24676 69378 24758 69392
rect 25634 69378 25716 69392
rect 25924 69378 26006 69392
rect 26882 69378 26964 69392
rect 27172 69378 27254 69392
rect 28130 69378 28212 69392
rect 28420 69378 28502 69392
rect 29378 69378 29460 69392
rect 29668 69378 29750 69392
rect 30626 69378 30708 69392
rect 30916 69378 30998 69392
rect 31874 69378 31956 69392
rect 32164 69378 32246 69392
rect 33122 69378 33204 69392
rect 33412 69378 33494 69392
rect 34370 69378 34452 69392
rect 34660 69378 34742 69392
rect 35618 69378 35700 69392
rect 35908 69378 35990 69392
rect 36866 69378 36948 69392
rect 37156 69378 37238 69392
rect 38114 69378 38196 69392
rect 38404 69378 38486 69392
rect 39362 69378 39444 69392
rect 39652 69378 39734 69392
rect 40610 69378 40692 69392
rect 40900 69378 40982 69392
rect 41858 69378 41940 69392
rect 42148 69378 42230 69392
rect 43106 69378 43188 69392
rect 43396 69378 43478 69392
rect 44354 69378 44436 69392
rect 44644 69378 44726 69392
rect 45602 69378 45684 69392
rect 45892 69378 45974 69392
rect 46850 69378 46932 69392
rect 47140 69378 47222 69392
rect 48098 69378 48180 69392
rect 48388 69378 48470 69392
rect 49346 69378 49428 69392
rect 49636 69378 49718 69392
rect 50594 69378 50676 69392
rect 50884 69378 50966 69392
rect 51842 69378 51924 69392
rect 52132 69378 52214 69392
rect 53090 69378 53172 69392
rect 53380 69378 53462 69392
rect 54338 69378 54420 69392
rect 54628 69378 54710 69392
rect 55586 69378 55668 69392
rect 55876 69378 55958 69392
rect 56834 69378 56916 69392
rect 57124 69378 57206 69392
rect 58082 69378 58164 69392
rect 58372 69378 58454 69392
rect 16418 69330 16864 69344
rect 17014 69330 17154 69344
rect 17304 69330 18112 69344
rect 18262 69330 18402 69344
rect 18552 69330 19360 69344
rect 19510 69330 19650 69344
rect 19800 69330 20608 69344
rect 20758 69330 20898 69344
rect 21048 69330 21856 69344
rect 22006 69330 22146 69344
rect 22296 69330 23104 69344
rect 23254 69330 23394 69344
rect 23544 69330 24352 69344
rect 24502 69330 24642 69344
rect 24792 69330 25600 69344
rect 25750 69330 25890 69344
rect 26040 69330 26848 69344
rect 26998 69330 27138 69344
rect 27288 69330 28096 69344
rect 28246 69330 28386 69344
rect 28536 69330 29344 69344
rect 29494 69330 29634 69344
rect 29784 69330 30592 69344
rect 30742 69330 30882 69344
rect 31032 69330 31840 69344
rect 31990 69330 32130 69344
rect 32280 69330 33088 69344
rect 33238 69330 33378 69344
rect 33528 69330 34336 69344
rect 34486 69330 34626 69344
rect 34776 69330 35584 69344
rect 35734 69330 35874 69344
rect 36024 69330 36832 69344
rect 36982 69330 37122 69344
rect 37272 69330 38080 69344
rect 38230 69330 38370 69344
rect 38520 69330 39328 69344
rect 39478 69330 39618 69344
rect 39768 69330 40576 69344
rect 40726 69330 40866 69344
rect 41016 69330 41824 69344
rect 41974 69330 42114 69344
rect 42264 69330 43072 69344
rect 43222 69330 43362 69344
rect 43512 69330 44320 69344
rect 44470 69330 44610 69344
rect 44760 69330 45568 69344
rect 45718 69330 45858 69344
rect 46008 69330 46816 69344
rect 46966 69330 47106 69344
rect 47256 69330 48064 69344
rect 48214 69330 48354 69344
rect 48504 69330 49312 69344
rect 49462 69330 49602 69344
rect 49752 69330 50560 69344
rect 50710 69330 50850 69344
rect 51000 69330 51808 69344
rect 51958 69330 52098 69344
rect 52248 69330 53056 69344
rect 53206 69330 53346 69344
rect 53496 69330 54304 69344
rect 54454 69330 54594 69344
rect 54744 69330 55552 69344
rect 55702 69330 55842 69344
rect 55992 69330 56800 69344
rect 56950 69330 57090 69344
rect 57240 69330 58048 69344
rect 58198 69330 58338 69344
rect 58488 69330 58934 69344
rect 16418 69282 58934 69330
rect 16418 69268 16864 69282
rect 17014 69268 17154 69282
rect 17304 69268 18112 69282
rect 18262 69268 18402 69282
rect 18552 69268 19360 69282
rect 19510 69268 19650 69282
rect 19800 69268 20608 69282
rect 20758 69268 20898 69282
rect 21048 69268 21856 69282
rect 22006 69268 22146 69282
rect 22296 69268 23104 69282
rect 23254 69268 23394 69282
rect 23544 69268 24352 69282
rect 24502 69268 24642 69282
rect 24792 69268 25600 69282
rect 25750 69268 25890 69282
rect 26040 69268 26848 69282
rect 26998 69268 27138 69282
rect 27288 69268 28096 69282
rect 28246 69268 28386 69282
rect 28536 69268 29344 69282
rect 29494 69268 29634 69282
rect 29784 69268 30592 69282
rect 30742 69268 30882 69282
rect 31032 69268 31840 69282
rect 31990 69268 32130 69282
rect 32280 69268 33088 69282
rect 33238 69268 33378 69282
rect 33528 69268 34336 69282
rect 34486 69268 34626 69282
rect 34776 69268 35584 69282
rect 35734 69268 35874 69282
rect 36024 69268 36832 69282
rect 36982 69268 37122 69282
rect 37272 69268 38080 69282
rect 38230 69268 38370 69282
rect 38520 69268 39328 69282
rect 39478 69268 39618 69282
rect 39768 69268 40576 69282
rect 40726 69268 40866 69282
rect 41016 69268 41824 69282
rect 41974 69268 42114 69282
rect 42264 69268 43072 69282
rect 43222 69268 43362 69282
rect 43512 69268 44320 69282
rect 44470 69268 44610 69282
rect 44760 69268 45568 69282
rect 45718 69268 45858 69282
rect 46008 69268 46816 69282
rect 46966 69268 47106 69282
rect 47256 69268 48064 69282
rect 48214 69268 48354 69282
rect 48504 69268 49312 69282
rect 49462 69268 49602 69282
rect 49752 69268 50560 69282
rect 50710 69268 50850 69282
rect 51000 69268 51808 69282
rect 51958 69268 52098 69282
rect 52248 69268 53056 69282
rect 53206 69268 53346 69282
rect 53496 69268 54304 69282
rect 54454 69268 54594 69282
rect 54744 69268 55552 69282
rect 55702 69268 55842 69282
rect 55992 69268 56800 69282
rect 56950 69268 57090 69282
rect 57240 69268 58048 69282
rect 58198 69268 58338 69282
rect 58488 69268 58934 69282
rect 16898 69220 16980 69234
rect 17188 69220 17270 69234
rect 18146 69220 18228 69234
rect 18436 69220 18518 69234
rect 19394 69220 19476 69234
rect 19684 69220 19766 69234
rect 20642 69220 20724 69234
rect 20932 69220 21014 69234
rect 21890 69220 21972 69234
rect 22180 69220 22262 69234
rect 23138 69220 23220 69234
rect 23428 69220 23510 69234
rect 24386 69220 24468 69234
rect 24676 69220 24758 69234
rect 25634 69220 25716 69234
rect 25924 69220 26006 69234
rect 26882 69220 26964 69234
rect 27172 69220 27254 69234
rect 28130 69220 28212 69234
rect 28420 69220 28502 69234
rect 29378 69220 29460 69234
rect 29668 69220 29750 69234
rect 30626 69220 30708 69234
rect 30916 69220 30998 69234
rect 31874 69220 31956 69234
rect 32164 69220 32246 69234
rect 33122 69220 33204 69234
rect 33412 69220 33494 69234
rect 34370 69220 34452 69234
rect 34660 69220 34742 69234
rect 35618 69220 35700 69234
rect 35908 69220 35990 69234
rect 36866 69220 36948 69234
rect 37156 69220 37238 69234
rect 38114 69220 38196 69234
rect 38404 69220 38486 69234
rect 39362 69220 39444 69234
rect 39652 69220 39734 69234
rect 40610 69220 40692 69234
rect 40900 69220 40982 69234
rect 41858 69220 41940 69234
rect 42148 69220 42230 69234
rect 43106 69220 43188 69234
rect 43396 69220 43478 69234
rect 44354 69220 44436 69234
rect 44644 69220 44726 69234
rect 45602 69220 45684 69234
rect 45892 69220 45974 69234
rect 46850 69220 46932 69234
rect 47140 69220 47222 69234
rect 48098 69220 48180 69234
rect 48388 69220 48470 69234
rect 49346 69220 49428 69234
rect 49636 69220 49718 69234
rect 50594 69220 50676 69234
rect 50884 69220 50966 69234
rect 51842 69220 51924 69234
rect 52132 69220 52214 69234
rect 53090 69220 53172 69234
rect 53380 69220 53462 69234
rect 54338 69220 54420 69234
rect 54628 69220 54710 69234
rect 55586 69220 55668 69234
rect 55876 69220 55958 69234
rect 56834 69220 56916 69234
rect 57124 69220 57206 69234
rect 58082 69220 58164 69234
rect 58372 69220 58454 69234
rect 16418 69172 58934 69220
rect 16418 69076 58934 69124
rect 16898 69062 16980 69076
rect 17188 69062 17270 69076
rect 18146 69062 18228 69076
rect 18436 69062 18518 69076
rect 19394 69062 19476 69076
rect 19684 69062 19766 69076
rect 20642 69062 20724 69076
rect 20932 69062 21014 69076
rect 21890 69062 21972 69076
rect 22180 69062 22262 69076
rect 23138 69062 23220 69076
rect 23428 69062 23510 69076
rect 24386 69062 24468 69076
rect 24676 69062 24758 69076
rect 25634 69062 25716 69076
rect 25924 69062 26006 69076
rect 26882 69062 26964 69076
rect 27172 69062 27254 69076
rect 28130 69062 28212 69076
rect 28420 69062 28502 69076
rect 29378 69062 29460 69076
rect 29668 69062 29750 69076
rect 30626 69062 30708 69076
rect 30916 69062 30998 69076
rect 31874 69062 31956 69076
rect 32164 69062 32246 69076
rect 33122 69062 33204 69076
rect 33412 69062 33494 69076
rect 34370 69062 34452 69076
rect 34660 69062 34742 69076
rect 35618 69062 35700 69076
rect 35908 69062 35990 69076
rect 36866 69062 36948 69076
rect 37156 69062 37238 69076
rect 38114 69062 38196 69076
rect 38404 69062 38486 69076
rect 39362 69062 39444 69076
rect 39652 69062 39734 69076
rect 40610 69062 40692 69076
rect 40900 69062 40982 69076
rect 41858 69062 41940 69076
rect 42148 69062 42230 69076
rect 43106 69062 43188 69076
rect 43396 69062 43478 69076
rect 44354 69062 44436 69076
rect 44644 69062 44726 69076
rect 45602 69062 45684 69076
rect 45892 69062 45974 69076
rect 46850 69062 46932 69076
rect 47140 69062 47222 69076
rect 48098 69062 48180 69076
rect 48388 69062 48470 69076
rect 49346 69062 49428 69076
rect 49636 69062 49718 69076
rect 50594 69062 50676 69076
rect 50884 69062 50966 69076
rect 51842 69062 51924 69076
rect 52132 69062 52214 69076
rect 53090 69062 53172 69076
rect 53380 69062 53462 69076
rect 54338 69062 54420 69076
rect 54628 69062 54710 69076
rect 55586 69062 55668 69076
rect 55876 69062 55958 69076
rect 56834 69062 56916 69076
rect 57124 69062 57206 69076
rect 58082 69062 58164 69076
rect 58372 69062 58454 69076
rect 16418 69014 16864 69028
rect 17014 69014 17154 69028
rect 17304 69014 18112 69028
rect 18262 69014 18402 69028
rect 18552 69014 19360 69028
rect 19510 69014 19650 69028
rect 19800 69014 20608 69028
rect 20758 69014 20898 69028
rect 21048 69014 21856 69028
rect 22006 69014 22146 69028
rect 22296 69014 23104 69028
rect 23254 69014 23394 69028
rect 23544 69014 24352 69028
rect 24502 69014 24642 69028
rect 24792 69014 25600 69028
rect 25750 69014 25890 69028
rect 26040 69014 26848 69028
rect 26998 69014 27138 69028
rect 27288 69014 28096 69028
rect 28246 69014 28386 69028
rect 28536 69014 29344 69028
rect 29494 69014 29634 69028
rect 29784 69014 30592 69028
rect 30742 69014 30882 69028
rect 31032 69014 31840 69028
rect 31990 69014 32130 69028
rect 32280 69014 33088 69028
rect 33238 69014 33378 69028
rect 33528 69014 34336 69028
rect 34486 69014 34626 69028
rect 34776 69014 35584 69028
rect 35734 69014 35874 69028
rect 36024 69014 36832 69028
rect 36982 69014 37122 69028
rect 37272 69014 38080 69028
rect 38230 69014 38370 69028
rect 38520 69014 39328 69028
rect 39478 69014 39618 69028
rect 39768 69014 40576 69028
rect 40726 69014 40866 69028
rect 41016 69014 41824 69028
rect 41974 69014 42114 69028
rect 42264 69014 43072 69028
rect 43222 69014 43362 69028
rect 43512 69014 44320 69028
rect 44470 69014 44610 69028
rect 44760 69014 45568 69028
rect 45718 69014 45858 69028
rect 46008 69014 46816 69028
rect 46966 69014 47106 69028
rect 47256 69014 48064 69028
rect 48214 69014 48354 69028
rect 48504 69014 49312 69028
rect 49462 69014 49602 69028
rect 49752 69014 50560 69028
rect 50710 69014 50850 69028
rect 51000 69014 51808 69028
rect 51958 69014 52098 69028
rect 52248 69014 53056 69028
rect 53206 69014 53346 69028
rect 53496 69014 54304 69028
rect 54454 69014 54594 69028
rect 54744 69014 55552 69028
rect 55702 69014 55842 69028
rect 55992 69014 56800 69028
rect 56950 69014 57090 69028
rect 57240 69014 58048 69028
rect 58198 69014 58338 69028
rect 58488 69014 58934 69028
rect 16418 68966 58934 69014
rect 16418 68952 16864 68966
rect 17014 68952 17154 68966
rect 17304 68952 18112 68966
rect 18262 68952 18402 68966
rect 18552 68952 19360 68966
rect 19510 68952 19650 68966
rect 19800 68952 20608 68966
rect 20758 68952 20898 68966
rect 21048 68952 21856 68966
rect 22006 68952 22146 68966
rect 22296 68952 23104 68966
rect 23254 68952 23394 68966
rect 23544 68952 24352 68966
rect 24502 68952 24642 68966
rect 24792 68952 25600 68966
rect 25750 68952 25890 68966
rect 26040 68952 26848 68966
rect 26998 68952 27138 68966
rect 27288 68952 28096 68966
rect 28246 68952 28386 68966
rect 28536 68952 29344 68966
rect 29494 68952 29634 68966
rect 29784 68952 30592 68966
rect 30742 68952 30882 68966
rect 31032 68952 31840 68966
rect 31990 68952 32130 68966
rect 32280 68952 33088 68966
rect 33238 68952 33378 68966
rect 33528 68952 34336 68966
rect 34486 68952 34626 68966
rect 34776 68952 35584 68966
rect 35734 68952 35874 68966
rect 36024 68952 36832 68966
rect 36982 68952 37122 68966
rect 37272 68952 38080 68966
rect 38230 68952 38370 68966
rect 38520 68952 39328 68966
rect 39478 68952 39618 68966
rect 39768 68952 40576 68966
rect 40726 68952 40866 68966
rect 41016 68952 41824 68966
rect 41974 68952 42114 68966
rect 42264 68952 43072 68966
rect 43222 68952 43362 68966
rect 43512 68952 44320 68966
rect 44470 68952 44610 68966
rect 44760 68952 45568 68966
rect 45718 68952 45858 68966
rect 46008 68952 46816 68966
rect 46966 68952 47106 68966
rect 47256 68952 48064 68966
rect 48214 68952 48354 68966
rect 48504 68952 49312 68966
rect 49462 68952 49602 68966
rect 49752 68952 50560 68966
rect 50710 68952 50850 68966
rect 51000 68952 51808 68966
rect 51958 68952 52098 68966
rect 52248 68952 53056 68966
rect 53206 68952 53346 68966
rect 53496 68952 54304 68966
rect 54454 68952 54594 68966
rect 54744 68952 55552 68966
rect 55702 68952 55842 68966
rect 55992 68952 56800 68966
rect 56950 68952 57090 68966
rect 57240 68952 58048 68966
rect 58198 68952 58338 68966
rect 58488 68952 58934 68966
rect 16898 68904 16980 68918
rect 17188 68904 17270 68918
rect 18146 68904 18228 68918
rect 18436 68904 18518 68918
rect 19394 68904 19476 68918
rect 19684 68904 19766 68918
rect 20642 68904 20724 68918
rect 20932 68904 21014 68918
rect 21890 68904 21972 68918
rect 22180 68904 22262 68918
rect 23138 68904 23220 68918
rect 23428 68904 23510 68918
rect 24386 68904 24468 68918
rect 24676 68904 24758 68918
rect 25634 68904 25716 68918
rect 25924 68904 26006 68918
rect 26882 68904 26964 68918
rect 27172 68904 27254 68918
rect 28130 68904 28212 68918
rect 28420 68904 28502 68918
rect 29378 68904 29460 68918
rect 29668 68904 29750 68918
rect 30626 68904 30708 68918
rect 30916 68904 30998 68918
rect 31874 68904 31956 68918
rect 32164 68904 32246 68918
rect 33122 68904 33204 68918
rect 33412 68904 33494 68918
rect 34370 68904 34452 68918
rect 34660 68904 34742 68918
rect 35618 68904 35700 68918
rect 35908 68904 35990 68918
rect 36866 68904 36948 68918
rect 37156 68904 37238 68918
rect 38114 68904 38196 68918
rect 38404 68904 38486 68918
rect 39362 68904 39444 68918
rect 39652 68904 39734 68918
rect 40610 68904 40692 68918
rect 40900 68904 40982 68918
rect 41858 68904 41940 68918
rect 42148 68904 42230 68918
rect 43106 68904 43188 68918
rect 43396 68904 43478 68918
rect 44354 68904 44436 68918
rect 44644 68904 44726 68918
rect 45602 68904 45684 68918
rect 45892 68904 45974 68918
rect 46850 68904 46932 68918
rect 47140 68904 47222 68918
rect 48098 68904 48180 68918
rect 48388 68904 48470 68918
rect 49346 68904 49428 68918
rect 49636 68904 49718 68918
rect 50594 68904 50676 68918
rect 50884 68904 50966 68918
rect 51842 68904 51924 68918
rect 52132 68904 52214 68918
rect 53090 68904 53172 68918
rect 53380 68904 53462 68918
rect 54338 68904 54420 68918
rect 54628 68904 54710 68918
rect 55586 68904 55668 68918
rect 55876 68904 55958 68918
rect 56834 68904 56916 68918
rect 57124 68904 57206 68918
rect 58082 68904 58164 68918
rect 58372 68904 58454 68918
rect 16418 68856 58934 68904
rect 16418 68698 58934 68808
rect 16418 68602 58934 68650
rect 16898 68588 16980 68602
rect 17188 68588 17270 68602
rect 18146 68588 18228 68602
rect 18436 68588 18518 68602
rect 19394 68588 19476 68602
rect 19684 68588 19766 68602
rect 20642 68588 20724 68602
rect 20932 68588 21014 68602
rect 21890 68588 21972 68602
rect 22180 68588 22262 68602
rect 23138 68588 23220 68602
rect 23428 68588 23510 68602
rect 24386 68588 24468 68602
rect 24676 68588 24758 68602
rect 25634 68588 25716 68602
rect 25924 68588 26006 68602
rect 26882 68588 26964 68602
rect 27172 68588 27254 68602
rect 28130 68588 28212 68602
rect 28420 68588 28502 68602
rect 29378 68588 29460 68602
rect 29668 68588 29750 68602
rect 30626 68588 30708 68602
rect 30916 68588 30998 68602
rect 31874 68588 31956 68602
rect 32164 68588 32246 68602
rect 33122 68588 33204 68602
rect 33412 68588 33494 68602
rect 34370 68588 34452 68602
rect 34660 68588 34742 68602
rect 35618 68588 35700 68602
rect 35908 68588 35990 68602
rect 36866 68588 36948 68602
rect 37156 68588 37238 68602
rect 38114 68588 38196 68602
rect 38404 68588 38486 68602
rect 39362 68588 39444 68602
rect 39652 68588 39734 68602
rect 40610 68588 40692 68602
rect 40900 68588 40982 68602
rect 41858 68588 41940 68602
rect 42148 68588 42230 68602
rect 43106 68588 43188 68602
rect 43396 68588 43478 68602
rect 44354 68588 44436 68602
rect 44644 68588 44726 68602
rect 45602 68588 45684 68602
rect 45892 68588 45974 68602
rect 46850 68588 46932 68602
rect 47140 68588 47222 68602
rect 48098 68588 48180 68602
rect 48388 68588 48470 68602
rect 49346 68588 49428 68602
rect 49636 68588 49718 68602
rect 50594 68588 50676 68602
rect 50884 68588 50966 68602
rect 51842 68588 51924 68602
rect 52132 68588 52214 68602
rect 53090 68588 53172 68602
rect 53380 68588 53462 68602
rect 54338 68588 54420 68602
rect 54628 68588 54710 68602
rect 55586 68588 55668 68602
rect 55876 68588 55958 68602
rect 56834 68588 56916 68602
rect 57124 68588 57206 68602
rect 58082 68588 58164 68602
rect 58372 68588 58454 68602
rect 16418 68540 16864 68554
rect 17014 68540 17154 68554
rect 17304 68540 18112 68554
rect 18262 68540 18402 68554
rect 18552 68540 19360 68554
rect 19510 68540 19650 68554
rect 19800 68540 20608 68554
rect 20758 68540 20898 68554
rect 21048 68540 21856 68554
rect 22006 68540 22146 68554
rect 22296 68540 23104 68554
rect 23254 68540 23394 68554
rect 23544 68540 24352 68554
rect 24502 68540 24642 68554
rect 24792 68540 25600 68554
rect 25750 68540 25890 68554
rect 26040 68540 26848 68554
rect 26998 68540 27138 68554
rect 27288 68540 28096 68554
rect 28246 68540 28386 68554
rect 28536 68540 29344 68554
rect 29494 68540 29634 68554
rect 29784 68540 30592 68554
rect 30742 68540 30882 68554
rect 31032 68540 31840 68554
rect 31990 68540 32130 68554
rect 32280 68540 33088 68554
rect 33238 68540 33378 68554
rect 33528 68540 34336 68554
rect 34486 68540 34626 68554
rect 34776 68540 35584 68554
rect 35734 68540 35874 68554
rect 36024 68540 36832 68554
rect 36982 68540 37122 68554
rect 37272 68540 38080 68554
rect 38230 68540 38370 68554
rect 38520 68540 39328 68554
rect 39478 68540 39618 68554
rect 39768 68540 40576 68554
rect 40726 68540 40866 68554
rect 41016 68540 41824 68554
rect 41974 68540 42114 68554
rect 42264 68540 43072 68554
rect 43222 68540 43362 68554
rect 43512 68540 44320 68554
rect 44470 68540 44610 68554
rect 44760 68540 45568 68554
rect 45718 68540 45858 68554
rect 46008 68540 46816 68554
rect 46966 68540 47106 68554
rect 47256 68540 48064 68554
rect 48214 68540 48354 68554
rect 48504 68540 49312 68554
rect 49462 68540 49602 68554
rect 49752 68540 50560 68554
rect 50710 68540 50850 68554
rect 51000 68540 51808 68554
rect 51958 68540 52098 68554
rect 52248 68540 53056 68554
rect 53206 68540 53346 68554
rect 53496 68540 54304 68554
rect 54454 68540 54594 68554
rect 54744 68540 55552 68554
rect 55702 68540 55842 68554
rect 55992 68540 56800 68554
rect 56950 68540 57090 68554
rect 57240 68540 58048 68554
rect 58198 68540 58338 68554
rect 58488 68540 58934 68554
rect 16418 68492 58934 68540
rect 16418 68478 16864 68492
rect 17014 68478 17154 68492
rect 17304 68478 18112 68492
rect 18262 68478 18402 68492
rect 18552 68478 19360 68492
rect 19510 68478 19650 68492
rect 19800 68478 20608 68492
rect 20758 68478 20898 68492
rect 21048 68478 21856 68492
rect 22006 68478 22146 68492
rect 22296 68478 23104 68492
rect 23254 68478 23394 68492
rect 23544 68478 24352 68492
rect 24502 68478 24642 68492
rect 24792 68478 25600 68492
rect 25750 68478 25890 68492
rect 26040 68478 26848 68492
rect 26998 68478 27138 68492
rect 27288 68478 28096 68492
rect 28246 68478 28386 68492
rect 28536 68478 29344 68492
rect 29494 68478 29634 68492
rect 29784 68478 30592 68492
rect 30742 68478 30882 68492
rect 31032 68478 31840 68492
rect 31990 68478 32130 68492
rect 32280 68478 33088 68492
rect 33238 68478 33378 68492
rect 33528 68478 34336 68492
rect 34486 68478 34626 68492
rect 34776 68478 35584 68492
rect 35734 68478 35874 68492
rect 36024 68478 36832 68492
rect 36982 68478 37122 68492
rect 37272 68478 38080 68492
rect 38230 68478 38370 68492
rect 38520 68478 39328 68492
rect 39478 68478 39618 68492
rect 39768 68478 40576 68492
rect 40726 68478 40866 68492
rect 41016 68478 41824 68492
rect 41974 68478 42114 68492
rect 42264 68478 43072 68492
rect 43222 68478 43362 68492
rect 43512 68478 44320 68492
rect 44470 68478 44610 68492
rect 44760 68478 45568 68492
rect 45718 68478 45858 68492
rect 46008 68478 46816 68492
rect 46966 68478 47106 68492
rect 47256 68478 48064 68492
rect 48214 68478 48354 68492
rect 48504 68478 49312 68492
rect 49462 68478 49602 68492
rect 49752 68478 50560 68492
rect 50710 68478 50850 68492
rect 51000 68478 51808 68492
rect 51958 68478 52098 68492
rect 52248 68478 53056 68492
rect 53206 68478 53346 68492
rect 53496 68478 54304 68492
rect 54454 68478 54594 68492
rect 54744 68478 55552 68492
rect 55702 68478 55842 68492
rect 55992 68478 56800 68492
rect 56950 68478 57090 68492
rect 57240 68478 58048 68492
rect 58198 68478 58338 68492
rect 58488 68478 58934 68492
rect 16898 68430 16980 68444
rect 17188 68430 17270 68444
rect 18146 68430 18228 68444
rect 18436 68430 18518 68444
rect 19394 68430 19476 68444
rect 19684 68430 19766 68444
rect 20642 68430 20724 68444
rect 20932 68430 21014 68444
rect 21890 68430 21972 68444
rect 22180 68430 22262 68444
rect 23138 68430 23220 68444
rect 23428 68430 23510 68444
rect 24386 68430 24468 68444
rect 24676 68430 24758 68444
rect 25634 68430 25716 68444
rect 25924 68430 26006 68444
rect 26882 68430 26964 68444
rect 27172 68430 27254 68444
rect 28130 68430 28212 68444
rect 28420 68430 28502 68444
rect 29378 68430 29460 68444
rect 29668 68430 29750 68444
rect 30626 68430 30708 68444
rect 30916 68430 30998 68444
rect 31874 68430 31956 68444
rect 32164 68430 32246 68444
rect 33122 68430 33204 68444
rect 33412 68430 33494 68444
rect 34370 68430 34452 68444
rect 34660 68430 34742 68444
rect 35618 68430 35700 68444
rect 35908 68430 35990 68444
rect 36866 68430 36948 68444
rect 37156 68430 37238 68444
rect 38114 68430 38196 68444
rect 38404 68430 38486 68444
rect 39362 68430 39444 68444
rect 39652 68430 39734 68444
rect 40610 68430 40692 68444
rect 40900 68430 40982 68444
rect 41858 68430 41940 68444
rect 42148 68430 42230 68444
rect 43106 68430 43188 68444
rect 43396 68430 43478 68444
rect 44354 68430 44436 68444
rect 44644 68430 44726 68444
rect 45602 68430 45684 68444
rect 45892 68430 45974 68444
rect 46850 68430 46932 68444
rect 47140 68430 47222 68444
rect 48098 68430 48180 68444
rect 48388 68430 48470 68444
rect 49346 68430 49428 68444
rect 49636 68430 49718 68444
rect 50594 68430 50676 68444
rect 50884 68430 50966 68444
rect 51842 68430 51924 68444
rect 52132 68430 52214 68444
rect 53090 68430 53172 68444
rect 53380 68430 53462 68444
rect 54338 68430 54420 68444
rect 54628 68430 54710 68444
rect 55586 68430 55668 68444
rect 55876 68430 55958 68444
rect 56834 68430 56916 68444
rect 57124 68430 57206 68444
rect 58082 68430 58164 68444
rect 58372 68430 58454 68444
rect 16418 68382 58934 68430
rect 16418 68286 58934 68334
rect 16898 68272 16980 68286
rect 17188 68272 17270 68286
rect 18146 68272 18228 68286
rect 18436 68272 18518 68286
rect 19394 68272 19476 68286
rect 19684 68272 19766 68286
rect 20642 68272 20724 68286
rect 20932 68272 21014 68286
rect 21890 68272 21972 68286
rect 22180 68272 22262 68286
rect 23138 68272 23220 68286
rect 23428 68272 23510 68286
rect 24386 68272 24468 68286
rect 24676 68272 24758 68286
rect 25634 68272 25716 68286
rect 25924 68272 26006 68286
rect 26882 68272 26964 68286
rect 27172 68272 27254 68286
rect 28130 68272 28212 68286
rect 28420 68272 28502 68286
rect 29378 68272 29460 68286
rect 29668 68272 29750 68286
rect 30626 68272 30708 68286
rect 30916 68272 30998 68286
rect 31874 68272 31956 68286
rect 32164 68272 32246 68286
rect 33122 68272 33204 68286
rect 33412 68272 33494 68286
rect 34370 68272 34452 68286
rect 34660 68272 34742 68286
rect 35618 68272 35700 68286
rect 35908 68272 35990 68286
rect 36866 68272 36948 68286
rect 37156 68272 37238 68286
rect 38114 68272 38196 68286
rect 38404 68272 38486 68286
rect 39362 68272 39444 68286
rect 39652 68272 39734 68286
rect 40610 68272 40692 68286
rect 40900 68272 40982 68286
rect 41858 68272 41940 68286
rect 42148 68272 42230 68286
rect 43106 68272 43188 68286
rect 43396 68272 43478 68286
rect 44354 68272 44436 68286
rect 44644 68272 44726 68286
rect 45602 68272 45684 68286
rect 45892 68272 45974 68286
rect 46850 68272 46932 68286
rect 47140 68272 47222 68286
rect 48098 68272 48180 68286
rect 48388 68272 48470 68286
rect 49346 68272 49428 68286
rect 49636 68272 49718 68286
rect 50594 68272 50676 68286
rect 50884 68272 50966 68286
rect 51842 68272 51924 68286
rect 52132 68272 52214 68286
rect 53090 68272 53172 68286
rect 53380 68272 53462 68286
rect 54338 68272 54420 68286
rect 54628 68272 54710 68286
rect 55586 68272 55668 68286
rect 55876 68272 55958 68286
rect 56834 68272 56916 68286
rect 57124 68272 57206 68286
rect 58082 68272 58164 68286
rect 58372 68272 58454 68286
rect 16418 68224 16864 68238
rect 17014 68224 17154 68238
rect 17304 68224 18112 68238
rect 18262 68224 18402 68238
rect 18552 68224 19360 68238
rect 19510 68224 19650 68238
rect 19800 68224 20608 68238
rect 20758 68224 20898 68238
rect 21048 68224 21856 68238
rect 22006 68224 22146 68238
rect 22296 68224 23104 68238
rect 23254 68224 23394 68238
rect 23544 68224 24352 68238
rect 24502 68224 24642 68238
rect 24792 68224 25600 68238
rect 25750 68224 25890 68238
rect 26040 68224 26848 68238
rect 26998 68224 27138 68238
rect 27288 68224 28096 68238
rect 28246 68224 28386 68238
rect 28536 68224 29344 68238
rect 29494 68224 29634 68238
rect 29784 68224 30592 68238
rect 30742 68224 30882 68238
rect 31032 68224 31840 68238
rect 31990 68224 32130 68238
rect 32280 68224 33088 68238
rect 33238 68224 33378 68238
rect 33528 68224 34336 68238
rect 34486 68224 34626 68238
rect 34776 68224 35584 68238
rect 35734 68224 35874 68238
rect 36024 68224 36832 68238
rect 36982 68224 37122 68238
rect 37272 68224 38080 68238
rect 38230 68224 38370 68238
rect 38520 68224 39328 68238
rect 39478 68224 39618 68238
rect 39768 68224 40576 68238
rect 40726 68224 40866 68238
rect 41016 68224 41824 68238
rect 41974 68224 42114 68238
rect 42264 68224 43072 68238
rect 43222 68224 43362 68238
rect 43512 68224 44320 68238
rect 44470 68224 44610 68238
rect 44760 68224 45568 68238
rect 45718 68224 45858 68238
rect 46008 68224 46816 68238
rect 46966 68224 47106 68238
rect 47256 68224 48064 68238
rect 48214 68224 48354 68238
rect 48504 68224 49312 68238
rect 49462 68224 49602 68238
rect 49752 68224 50560 68238
rect 50710 68224 50850 68238
rect 51000 68224 51808 68238
rect 51958 68224 52098 68238
rect 52248 68224 53056 68238
rect 53206 68224 53346 68238
rect 53496 68224 54304 68238
rect 54454 68224 54594 68238
rect 54744 68224 55552 68238
rect 55702 68224 55842 68238
rect 55992 68224 56800 68238
rect 56950 68224 57090 68238
rect 57240 68224 58048 68238
rect 58198 68224 58338 68238
rect 58488 68224 58934 68238
rect 16418 68176 58934 68224
rect 16418 68162 16864 68176
rect 17014 68162 17154 68176
rect 17304 68162 18112 68176
rect 18262 68162 18402 68176
rect 18552 68162 19360 68176
rect 19510 68162 19650 68176
rect 19800 68162 20608 68176
rect 20758 68162 20898 68176
rect 21048 68162 21856 68176
rect 22006 68162 22146 68176
rect 22296 68162 23104 68176
rect 23254 68162 23394 68176
rect 23544 68162 24352 68176
rect 24502 68162 24642 68176
rect 24792 68162 25600 68176
rect 25750 68162 25890 68176
rect 26040 68162 26848 68176
rect 26998 68162 27138 68176
rect 27288 68162 28096 68176
rect 28246 68162 28386 68176
rect 28536 68162 29344 68176
rect 29494 68162 29634 68176
rect 29784 68162 30592 68176
rect 30742 68162 30882 68176
rect 31032 68162 31840 68176
rect 31990 68162 32130 68176
rect 32280 68162 33088 68176
rect 33238 68162 33378 68176
rect 33528 68162 34336 68176
rect 34486 68162 34626 68176
rect 34776 68162 35584 68176
rect 35734 68162 35874 68176
rect 36024 68162 36832 68176
rect 36982 68162 37122 68176
rect 37272 68162 38080 68176
rect 38230 68162 38370 68176
rect 38520 68162 39328 68176
rect 39478 68162 39618 68176
rect 39768 68162 40576 68176
rect 40726 68162 40866 68176
rect 41016 68162 41824 68176
rect 41974 68162 42114 68176
rect 42264 68162 43072 68176
rect 43222 68162 43362 68176
rect 43512 68162 44320 68176
rect 44470 68162 44610 68176
rect 44760 68162 45568 68176
rect 45718 68162 45858 68176
rect 46008 68162 46816 68176
rect 46966 68162 47106 68176
rect 47256 68162 48064 68176
rect 48214 68162 48354 68176
rect 48504 68162 49312 68176
rect 49462 68162 49602 68176
rect 49752 68162 50560 68176
rect 50710 68162 50850 68176
rect 51000 68162 51808 68176
rect 51958 68162 52098 68176
rect 52248 68162 53056 68176
rect 53206 68162 53346 68176
rect 53496 68162 54304 68176
rect 54454 68162 54594 68176
rect 54744 68162 55552 68176
rect 55702 68162 55842 68176
rect 55992 68162 56800 68176
rect 56950 68162 57090 68176
rect 57240 68162 58048 68176
rect 58198 68162 58338 68176
rect 58488 68162 58934 68176
rect 16898 68114 16980 68128
rect 17188 68114 17270 68128
rect 18146 68114 18228 68128
rect 18436 68114 18518 68128
rect 19394 68114 19476 68128
rect 19684 68114 19766 68128
rect 20642 68114 20724 68128
rect 20932 68114 21014 68128
rect 21890 68114 21972 68128
rect 22180 68114 22262 68128
rect 23138 68114 23220 68128
rect 23428 68114 23510 68128
rect 24386 68114 24468 68128
rect 24676 68114 24758 68128
rect 25634 68114 25716 68128
rect 25924 68114 26006 68128
rect 26882 68114 26964 68128
rect 27172 68114 27254 68128
rect 28130 68114 28212 68128
rect 28420 68114 28502 68128
rect 29378 68114 29460 68128
rect 29668 68114 29750 68128
rect 30626 68114 30708 68128
rect 30916 68114 30998 68128
rect 31874 68114 31956 68128
rect 32164 68114 32246 68128
rect 33122 68114 33204 68128
rect 33412 68114 33494 68128
rect 34370 68114 34452 68128
rect 34660 68114 34742 68128
rect 35618 68114 35700 68128
rect 35908 68114 35990 68128
rect 36866 68114 36948 68128
rect 37156 68114 37238 68128
rect 38114 68114 38196 68128
rect 38404 68114 38486 68128
rect 39362 68114 39444 68128
rect 39652 68114 39734 68128
rect 40610 68114 40692 68128
rect 40900 68114 40982 68128
rect 41858 68114 41940 68128
rect 42148 68114 42230 68128
rect 43106 68114 43188 68128
rect 43396 68114 43478 68128
rect 44354 68114 44436 68128
rect 44644 68114 44726 68128
rect 45602 68114 45684 68128
rect 45892 68114 45974 68128
rect 46850 68114 46932 68128
rect 47140 68114 47222 68128
rect 48098 68114 48180 68128
rect 48388 68114 48470 68128
rect 49346 68114 49428 68128
rect 49636 68114 49718 68128
rect 50594 68114 50676 68128
rect 50884 68114 50966 68128
rect 51842 68114 51924 68128
rect 52132 68114 52214 68128
rect 53090 68114 53172 68128
rect 53380 68114 53462 68128
rect 54338 68114 54420 68128
rect 54628 68114 54710 68128
rect 55586 68114 55668 68128
rect 55876 68114 55958 68128
rect 56834 68114 56916 68128
rect 57124 68114 57206 68128
rect 58082 68114 58164 68128
rect 58372 68114 58454 68128
rect 16418 68066 58934 68114
rect 16418 67908 58934 68018
rect 16418 67812 58934 67860
rect 16898 67798 16980 67812
rect 17188 67798 17270 67812
rect 18146 67798 18228 67812
rect 18436 67798 18518 67812
rect 19394 67798 19476 67812
rect 19684 67798 19766 67812
rect 20642 67798 20724 67812
rect 20932 67798 21014 67812
rect 21890 67798 21972 67812
rect 22180 67798 22262 67812
rect 23138 67798 23220 67812
rect 23428 67798 23510 67812
rect 24386 67798 24468 67812
rect 24676 67798 24758 67812
rect 25634 67798 25716 67812
rect 25924 67798 26006 67812
rect 26882 67798 26964 67812
rect 27172 67798 27254 67812
rect 28130 67798 28212 67812
rect 28420 67798 28502 67812
rect 29378 67798 29460 67812
rect 29668 67798 29750 67812
rect 30626 67798 30708 67812
rect 30916 67798 30998 67812
rect 31874 67798 31956 67812
rect 32164 67798 32246 67812
rect 33122 67798 33204 67812
rect 33412 67798 33494 67812
rect 34370 67798 34452 67812
rect 34660 67798 34742 67812
rect 35618 67798 35700 67812
rect 35908 67798 35990 67812
rect 36866 67798 36948 67812
rect 37156 67798 37238 67812
rect 38114 67798 38196 67812
rect 38404 67798 38486 67812
rect 39362 67798 39444 67812
rect 39652 67798 39734 67812
rect 40610 67798 40692 67812
rect 40900 67798 40982 67812
rect 41858 67798 41940 67812
rect 42148 67798 42230 67812
rect 43106 67798 43188 67812
rect 43396 67798 43478 67812
rect 44354 67798 44436 67812
rect 44644 67798 44726 67812
rect 45602 67798 45684 67812
rect 45892 67798 45974 67812
rect 46850 67798 46932 67812
rect 47140 67798 47222 67812
rect 48098 67798 48180 67812
rect 48388 67798 48470 67812
rect 49346 67798 49428 67812
rect 49636 67798 49718 67812
rect 50594 67798 50676 67812
rect 50884 67798 50966 67812
rect 51842 67798 51924 67812
rect 52132 67798 52214 67812
rect 53090 67798 53172 67812
rect 53380 67798 53462 67812
rect 54338 67798 54420 67812
rect 54628 67798 54710 67812
rect 55586 67798 55668 67812
rect 55876 67798 55958 67812
rect 56834 67798 56916 67812
rect 57124 67798 57206 67812
rect 58082 67798 58164 67812
rect 58372 67798 58454 67812
rect 16418 67750 16864 67764
rect 17014 67750 17154 67764
rect 17304 67750 18112 67764
rect 18262 67750 18402 67764
rect 18552 67750 19360 67764
rect 19510 67750 19650 67764
rect 19800 67750 20608 67764
rect 20758 67750 20898 67764
rect 21048 67750 21856 67764
rect 22006 67750 22146 67764
rect 22296 67750 23104 67764
rect 23254 67750 23394 67764
rect 23544 67750 24352 67764
rect 24502 67750 24642 67764
rect 24792 67750 25600 67764
rect 25750 67750 25890 67764
rect 26040 67750 26848 67764
rect 26998 67750 27138 67764
rect 27288 67750 28096 67764
rect 28246 67750 28386 67764
rect 28536 67750 29344 67764
rect 29494 67750 29634 67764
rect 29784 67750 30592 67764
rect 30742 67750 30882 67764
rect 31032 67750 31840 67764
rect 31990 67750 32130 67764
rect 32280 67750 33088 67764
rect 33238 67750 33378 67764
rect 33528 67750 34336 67764
rect 34486 67750 34626 67764
rect 34776 67750 35584 67764
rect 35734 67750 35874 67764
rect 36024 67750 36832 67764
rect 36982 67750 37122 67764
rect 37272 67750 38080 67764
rect 38230 67750 38370 67764
rect 38520 67750 39328 67764
rect 39478 67750 39618 67764
rect 39768 67750 40576 67764
rect 40726 67750 40866 67764
rect 41016 67750 41824 67764
rect 41974 67750 42114 67764
rect 42264 67750 43072 67764
rect 43222 67750 43362 67764
rect 43512 67750 44320 67764
rect 44470 67750 44610 67764
rect 44760 67750 45568 67764
rect 45718 67750 45858 67764
rect 46008 67750 46816 67764
rect 46966 67750 47106 67764
rect 47256 67750 48064 67764
rect 48214 67750 48354 67764
rect 48504 67750 49312 67764
rect 49462 67750 49602 67764
rect 49752 67750 50560 67764
rect 50710 67750 50850 67764
rect 51000 67750 51808 67764
rect 51958 67750 52098 67764
rect 52248 67750 53056 67764
rect 53206 67750 53346 67764
rect 53496 67750 54304 67764
rect 54454 67750 54594 67764
rect 54744 67750 55552 67764
rect 55702 67750 55842 67764
rect 55992 67750 56800 67764
rect 56950 67750 57090 67764
rect 57240 67750 58048 67764
rect 58198 67750 58338 67764
rect 58488 67750 58934 67764
rect 16418 67702 58934 67750
rect 16418 67688 16864 67702
rect 17014 67688 17154 67702
rect 17304 67688 18112 67702
rect 18262 67688 18402 67702
rect 18552 67688 19360 67702
rect 19510 67688 19650 67702
rect 19800 67688 20608 67702
rect 20758 67688 20898 67702
rect 21048 67688 21856 67702
rect 22006 67688 22146 67702
rect 22296 67688 23104 67702
rect 23254 67688 23394 67702
rect 23544 67688 24352 67702
rect 24502 67688 24642 67702
rect 24792 67688 25600 67702
rect 25750 67688 25890 67702
rect 26040 67688 26848 67702
rect 26998 67688 27138 67702
rect 27288 67688 28096 67702
rect 28246 67688 28386 67702
rect 28536 67688 29344 67702
rect 29494 67688 29634 67702
rect 29784 67688 30592 67702
rect 30742 67688 30882 67702
rect 31032 67688 31840 67702
rect 31990 67688 32130 67702
rect 32280 67688 33088 67702
rect 33238 67688 33378 67702
rect 33528 67688 34336 67702
rect 34486 67688 34626 67702
rect 34776 67688 35584 67702
rect 35734 67688 35874 67702
rect 36024 67688 36832 67702
rect 36982 67688 37122 67702
rect 37272 67688 38080 67702
rect 38230 67688 38370 67702
rect 38520 67688 39328 67702
rect 39478 67688 39618 67702
rect 39768 67688 40576 67702
rect 40726 67688 40866 67702
rect 41016 67688 41824 67702
rect 41974 67688 42114 67702
rect 42264 67688 43072 67702
rect 43222 67688 43362 67702
rect 43512 67688 44320 67702
rect 44470 67688 44610 67702
rect 44760 67688 45568 67702
rect 45718 67688 45858 67702
rect 46008 67688 46816 67702
rect 46966 67688 47106 67702
rect 47256 67688 48064 67702
rect 48214 67688 48354 67702
rect 48504 67688 49312 67702
rect 49462 67688 49602 67702
rect 49752 67688 50560 67702
rect 50710 67688 50850 67702
rect 51000 67688 51808 67702
rect 51958 67688 52098 67702
rect 52248 67688 53056 67702
rect 53206 67688 53346 67702
rect 53496 67688 54304 67702
rect 54454 67688 54594 67702
rect 54744 67688 55552 67702
rect 55702 67688 55842 67702
rect 55992 67688 56800 67702
rect 56950 67688 57090 67702
rect 57240 67688 58048 67702
rect 58198 67688 58338 67702
rect 58488 67688 58934 67702
rect 16898 67640 16980 67654
rect 17188 67640 17270 67654
rect 18146 67640 18228 67654
rect 18436 67640 18518 67654
rect 19394 67640 19476 67654
rect 19684 67640 19766 67654
rect 20642 67640 20724 67654
rect 20932 67640 21014 67654
rect 21890 67640 21972 67654
rect 22180 67640 22262 67654
rect 23138 67640 23220 67654
rect 23428 67640 23510 67654
rect 24386 67640 24468 67654
rect 24676 67640 24758 67654
rect 25634 67640 25716 67654
rect 25924 67640 26006 67654
rect 26882 67640 26964 67654
rect 27172 67640 27254 67654
rect 28130 67640 28212 67654
rect 28420 67640 28502 67654
rect 29378 67640 29460 67654
rect 29668 67640 29750 67654
rect 30626 67640 30708 67654
rect 30916 67640 30998 67654
rect 31874 67640 31956 67654
rect 32164 67640 32246 67654
rect 33122 67640 33204 67654
rect 33412 67640 33494 67654
rect 34370 67640 34452 67654
rect 34660 67640 34742 67654
rect 35618 67640 35700 67654
rect 35908 67640 35990 67654
rect 36866 67640 36948 67654
rect 37156 67640 37238 67654
rect 38114 67640 38196 67654
rect 38404 67640 38486 67654
rect 39362 67640 39444 67654
rect 39652 67640 39734 67654
rect 40610 67640 40692 67654
rect 40900 67640 40982 67654
rect 41858 67640 41940 67654
rect 42148 67640 42230 67654
rect 43106 67640 43188 67654
rect 43396 67640 43478 67654
rect 44354 67640 44436 67654
rect 44644 67640 44726 67654
rect 45602 67640 45684 67654
rect 45892 67640 45974 67654
rect 46850 67640 46932 67654
rect 47140 67640 47222 67654
rect 48098 67640 48180 67654
rect 48388 67640 48470 67654
rect 49346 67640 49428 67654
rect 49636 67640 49718 67654
rect 50594 67640 50676 67654
rect 50884 67640 50966 67654
rect 51842 67640 51924 67654
rect 52132 67640 52214 67654
rect 53090 67640 53172 67654
rect 53380 67640 53462 67654
rect 54338 67640 54420 67654
rect 54628 67640 54710 67654
rect 55586 67640 55668 67654
rect 55876 67640 55958 67654
rect 56834 67640 56916 67654
rect 57124 67640 57206 67654
rect 58082 67640 58164 67654
rect 58372 67640 58454 67654
rect 16418 67592 58934 67640
rect 16418 67496 58934 67544
rect 16898 67482 16980 67496
rect 17188 67482 17270 67496
rect 18146 67482 18228 67496
rect 18436 67482 18518 67496
rect 19394 67482 19476 67496
rect 19684 67482 19766 67496
rect 20642 67482 20724 67496
rect 20932 67482 21014 67496
rect 21890 67482 21972 67496
rect 22180 67482 22262 67496
rect 23138 67482 23220 67496
rect 23428 67482 23510 67496
rect 24386 67482 24468 67496
rect 24676 67482 24758 67496
rect 25634 67482 25716 67496
rect 25924 67482 26006 67496
rect 26882 67482 26964 67496
rect 27172 67482 27254 67496
rect 28130 67482 28212 67496
rect 28420 67482 28502 67496
rect 29378 67482 29460 67496
rect 29668 67482 29750 67496
rect 30626 67482 30708 67496
rect 30916 67482 30998 67496
rect 31874 67482 31956 67496
rect 32164 67482 32246 67496
rect 33122 67482 33204 67496
rect 33412 67482 33494 67496
rect 34370 67482 34452 67496
rect 34660 67482 34742 67496
rect 35618 67482 35700 67496
rect 35908 67482 35990 67496
rect 36866 67482 36948 67496
rect 37156 67482 37238 67496
rect 38114 67482 38196 67496
rect 38404 67482 38486 67496
rect 39362 67482 39444 67496
rect 39652 67482 39734 67496
rect 40610 67482 40692 67496
rect 40900 67482 40982 67496
rect 41858 67482 41940 67496
rect 42148 67482 42230 67496
rect 43106 67482 43188 67496
rect 43396 67482 43478 67496
rect 44354 67482 44436 67496
rect 44644 67482 44726 67496
rect 45602 67482 45684 67496
rect 45892 67482 45974 67496
rect 46850 67482 46932 67496
rect 47140 67482 47222 67496
rect 48098 67482 48180 67496
rect 48388 67482 48470 67496
rect 49346 67482 49428 67496
rect 49636 67482 49718 67496
rect 50594 67482 50676 67496
rect 50884 67482 50966 67496
rect 51842 67482 51924 67496
rect 52132 67482 52214 67496
rect 53090 67482 53172 67496
rect 53380 67482 53462 67496
rect 54338 67482 54420 67496
rect 54628 67482 54710 67496
rect 55586 67482 55668 67496
rect 55876 67482 55958 67496
rect 56834 67482 56916 67496
rect 57124 67482 57206 67496
rect 58082 67482 58164 67496
rect 58372 67482 58454 67496
rect 16418 67434 16864 67448
rect 17014 67434 17154 67448
rect 17304 67434 18112 67448
rect 18262 67434 18402 67448
rect 18552 67434 19360 67448
rect 19510 67434 19650 67448
rect 19800 67434 20608 67448
rect 20758 67434 20898 67448
rect 21048 67434 21856 67448
rect 22006 67434 22146 67448
rect 22296 67434 23104 67448
rect 23254 67434 23394 67448
rect 23544 67434 24352 67448
rect 24502 67434 24642 67448
rect 24792 67434 25600 67448
rect 25750 67434 25890 67448
rect 26040 67434 26848 67448
rect 26998 67434 27138 67448
rect 27288 67434 28096 67448
rect 28246 67434 28386 67448
rect 28536 67434 29344 67448
rect 29494 67434 29634 67448
rect 29784 67434 30592 67448
rect 30742 67434 30882 67448
rect 31032 67434 31840 67448
rect 31990 67434 32130 67448
rect 32280 67434 33088 67448
rect 33238 67434 33378 67448
rect 33528 67434 34336 67448
rect 34486 67434 34626 67448
rect 34776 67434 35584 67448
rect 35734 67434 35874 67448
rect 36024 67434 36832 67448
rect 36982 67434 37122 67448
rect 37272 67434 38080 67448
rect 38230 67434 38370 67448
rect 38520 67434 39328 67448
rect 39478 67434 39618 67448
rect 39768 67434 40576 67448
rect 40726 67434 40866 67448
rect 41016 67434 41824 67448
rect 41974 67434 42114 67448
rect 42264 67434 43072 67448
rect 43222 67434 43362 67448
rect 43512 67434 44320 67448
rect 44470 67434 44610 67448
rect 44760 67434 45568 67448
rect 45718 67434 45858 67448
rect 46008 67434 46816 67448
rect 46966 67434 47106 67448
rect 47256 67434 48064 67448
rect 48214 67434 48354 67448
rect 48504 67434 49312 67448
rect 49462 67434 49602 67448
rect 49752 67434 50560 67448
rect 50710 67434 50850 67448
rect 51000 67434 51808 67448
rect 51958 67434 52098 67448
rect 52248 67434 53056 67448
rect 53206 67434 53346 67448
rect 53496 67434 54304 67448
rect 54454 67434 54594 67448
rect 54744 67434 55552 67448
rect 55702 67434 55842 67448
rect 55992 67434 56800 67448
rect 56950 67434 57090 67448
rect 57240 67434 58048 67448
rect 58198 67434 58338 67448
rect 58488 67434 58934 67448
rect 16418 67386 58934 67434
rect 16418 67372 16864 67386
rect 17014 67372 17154 67386
rect 17304 67372 18112 67386
rect 18262 67372 18402 67386
rect 18552 67372 19360 67386
rect 19510 67372 19650 67386
rect 19800 67372 20608 67386
rect 20758 67372 20898 67386
rect 21048 67372 21856 67386
rect 22006 67372 22146 67386
rect 22296 67372 23104 67386
rect 23254 67372 23394 67386
rect 23544 67372 24352 67386
rect 24502 67372 24642 67386
rect 24792 67372 25600 67386
rect 25750 67372 25890 67386
rect 26040 67372 26848 67386
rect 26998 67372 27138 67386
rect 27288 67372 28096 67386
rect 28246 67372 28386 67386
rect 28536 67372 29344 67386
rect 29494 67372 29634 67386
rect 29784 67372 30592 67386
rect 30742 67372 30882 67386
rect 31032 67372 31840 67386
rect 31990 67372 32130 67386
rect 32280 67372 33088 67386
rect 33238 67372 33378 67386
rect 33528 67372 34336 67386
rect 34486 67372 34626 67386
rect 34776 67372 35584 67386
rect 35734 67372 35874 67386
rect 36024 67372 36832 67386
rect 36982 67372 37122 67386
rect 37272 67372 38080 67386
rect 38230 67372 38370 67386
rect 38520 67372 39328 67386
rect 39478 67372 39618 67386
rect 39768 67372 40576 67386
rect 40726 67372 40866 67386
rect 41016 67372 41824 67386
rect 41974 67372 42114 67386
rect 42264 67372 43072 67386
rect 43222 67372 43362 67386
rect 43512 67372 44320 67386
rect 44470 67372 44610 67386
rect 44760 67372 45568 67386
rect 45718 67372 45858 67386
rect 46008 67372 46816 67386
rect 46966 67372 47106 67386
rect 47256 67372 48064 67386
rect 48214 67372 48354 67386
rect 48504 67372 49312 67386
rect 49462 67372 49602 67386
rect 49752 67372 50560 67386
rect 50710 67372 50850 67386
rect 51000 67372 51808 67386
rect 51958 67372 52098 67386
rect 52248 67372 53056 67386
rect 53206 67372 53346 67386
rect 53496 67372 54304 67386
rect 54454 67372 54594 67386
rect 54744 67372 55552 67386
rect 55702 67372 55842 67386
rect 55992 67372 56800 67386
rect 56950 67372 57090 67386
rect 57240 67372 58048 67386
rect 58198 67372 58338 67386
rect 58488 67372 58934 67386
rect 16898 67324 16980 67338
rect 17188 67324 17270 67338
rect 18146 67324 18228 67338
rect 18436 67324 18518 67338
rect 19394 67324 19476 67338
rect 19684 67324 19766 67338
rect 20642 67324 20724 67338
rect 20932 67324 21014 67338
rect 21890 67324 21972 67338
rect 22180 67324 22262 67338
rect 23138 67324 23220 67338
rect 23428 67324 23510 67338
rect 24386 67324 24468 67338
rect 24676 67324 24758 67338
rect 25634 67324 25716 67338
rect 25924 67324 26006 67338
rect 26882 67324 26964 67338
rect 27172 67324 27254 67338
rect 28130 67324 28212 67338
rect 28420 67324 28502 67338
rect 29378 67324 29460 67338
rect 29668 67324 29750 67338
rect 30626 67324 30708 67338
rect 30916 67324 30998 67338
rect 31874 67324 31956 67338
rect 32164 67324 32246 67338
rect 33122 67324 33204 67338
rect 33412 67324 33494 67338
rect 34370 67324 34452 67338
rect 34660 67324 34742 67338
rect 35618 67324 35700 67338
rect 35908 67324 35990 67338
rect 36866 67324 36948 67338
rect 37156 67324 37238 67338
rect 38114 67324 38196 67338
rect 38404 67324 38486 67338
rect 39362 67324 39444 67338
rect 39652 67324 39734 67338
rect 40610 67324 40692 67338
rect 40900 67324 40982 67338
rect 41858 67324 41940 67338
rect 42148 67324 42230 67338
rect 43106 67324 43188 67338
rect 43396 67324 43478 67338
rect 44354 67324 44436 67338
rect 44644 67324 44726 67338
rect 45602 67324 45684 67338
rect 45892 67324 45974 67338
rect 46850 67324 46932 67338
rect 47140 67324 47222 67338
rect 48098 67324 48180 67338
rect 48388 67324 48470 67338
rect 49346 67324 49428 67338
rect 49636 67324 49718 67338
rect 50594 67324 50676 67338
rect 50884 67324 50966 67338
rect 51842 67324 51924 67338
rect 52132 67324 52214 67338
rect 53090 67324 53172 67338
rect 53380 67324 53462 67338
rect 54338 67324 54420 67338
rect 54628 67324 54710 67338
rect 55586 67324 55668 67338
rect 55876 67324 55958 67338
rect 56834 67324 56916 67338
rect 57124 67324 57206 67338
rect 58082 67324 58164 67338
rect 58372 67324 58454 67338
rect 16418 67276 58934 67324
rect 16418 67118 58934 67228
rect 16418 67022 58934 67070
rect 16898 67008 16980 67022
rect 17188 67008 17270 67022
rect 18146 67008 18228 67022
rect 18436 67008 18518 67022
rect 19394 67008 19476 67022
rect 19684 67008 19766 67022
rect 20642 67008 20724 67022
rect 20932 67008 21014 67022
rect 21890 67008 21972 67022
rect 22180 67008 22262 67022
rect 23138 67008 23220 67022
rect 23428 67008 23510 67022
rect 24386 67008 24468 67022
rect 24676 67008 24758 67022
rect 25634 67008 25716 67022
rect 25924 67008 26006 67022
rect 26882 67008 26964 67022
rect 27172 67008 27254 67022
rect 28130 67008 28212 67022
rect 28420 67008 28502 67022
rect 29378 67008 29460 67022
rect 29668 67008 29750 67022
rect 30626 67008 30708 67022
rect 30916 67008 30998 67022
rect 31874 67008 31956 67022
rect 32164 67008 32246 67022
rect 33122 67008 33204 67022
rect 33412 67008 33494 67022
rect 34370 67008 34452 67022
rect 34660 67008 34742 67022
rect 35618 67008 35700 67022
rect 35908 67008 35990 67022
rect 36866 67008 36948 67022
rect 37156 67008 37238 67022
rect 38114 67008 38196 67022
rect 38404 67008 38486 67022
rect 39362 67008 39444 67022
rect 39652 67008 39734 67022
rect 40610 67008 40692 67022
rect 40900 67008 40982 67022
rect 41858 67008 41940 67022
rect 42148 67008 42230 67022
rect 43106 67008 43188 67022
rect 43396 67008 43478 67022
rect 44354 67008 44436 67022
rect 44644 67008 44726 67022
rect 45602 67008 45684 67022
rect 45892 67008 45974 67022
rect 46850 67008 46932 67022
rect 47140 67008 47222 67022
rect 48098 67008 48180 67022
rect 48388 67008 48470 67022
rect 49346 67008 49428 67022
rect 49636 67008 49718 67022
rect 50594 67008 50676 67022
rect 50884 67008 50966 67022
rect 51842 67008 51924 67022
rect 52132 67008 52214 67022
rect 53090 67008 53172 67022
rect 53380 67008 53462 67022
rect 54338 67008 54420 67022
rect 54628 67008 54710 67022
rect 55586 67008 55668 67022
rect 55876 67008 55958 67022
rect 56834 67008 56916 67022
rect 57124 67008 57206 67022
rect 58082 67008 58164 67022
rect 58372 67008 58454 67022
rect 16418 66960 16864 66974
rect 17014 66960 17154 66974
rect 17304 66960 18112 66974
rect 18262 66960 18402 66974
rect 18552 66960 19360 66974
rect 19510 66960 19650 66974
rect 19800 66960 20608 66974
rect 20758 66960 20898 66974
rect 21048 66960 21856 66974
rect 22006 66960 22146 66974
rect 22296 66960 23104 66974
rect 23254 66960 23394 66974
rect 23544 66960 24352 66974
rect 24502 66960 24642 66974
rect 24792 66960 25600 66974
rect 25750 66960 25890 66974
rect 26040 66960 26848 66974
rect 26998 66960 27138 66974
rect 27288 66960 28096 66974
rect 28246 66960 28386 66974
rect 28536 66960 29344 66974
rect 29494 66960 29634 66974
rect 29784 66960 30592 66974
rect 30742 66960 30882 66974
rect 31032 66960 31840 66974
rect 31990 66960 32130 66974
rect 32280 66960 33088 66974
rect 33238 66960 33378 66974
rect 33528 66960 34336 66974
rect 34486 66960 34626 66974
rect 34776 66960 35584 66974
rect 35734 66960 35874 66974
rect 36024 66960 36832 66974
rect 36982 66960 37122 66974
rect 37272 66960 38080 66974
rect 38230 66960 38370 66974
rect 38520 66960 39328 66974
rect 39478 66960 39618 66974
rect 39768 66960 40576 66974
rect 40726 66960 40866 66974
rect 41016 66960 41824 66974
rect 41974 66960 42114 66974
rect 42264 66960 43072 66974
rect 43222 66960 43362 66974
rect 43512 66960 44320 66974
rect 44470 66960 44610 66974
rect 44760 66960 45568 66974
rect 45718 66960 45858 66974
rect 46008 66960 46816 66974
rect 46966 66960 47106 66974
rect 47256 66960 48064 66974
rect 48214 66960 48354 66974
rect 48504 66960 49312 66974
rect 49462 66960 49602 66974
rect 49752 66960 50560 66974
rect 50710 66960 50850 66974
rect 51000 66960 51808 66974
rect 51958 66960 52098 66974
rect 52248 66960 53056 66974
rect 53206 66960 53346 66974
rect 53496 66960 54304 66974
rect 54454 66960 54594 66974
rect 54744 66960 55552 66974
rect 55702 66960 55842 66974
rect 55992 66960 56800 66974
rect 56950 66960 57090 66974
rect 57240 66960 58048 66974
rect 58198 66960 58338 66974
rect 58488 66960 58934 66974
rect 16418 66912 58934 66960
rect 16418 66898 16864 66912
rect 17014 66898 17154 66912
rect 17304 66898 18112 66912
rect 18262 66898 18402 66912
rect 18552 66898 19360 66912
rect 19510 66898 19650 66912
rect 19800 66898 20608 66912
rect 20758 66898 20898 66912
rect 21048 66898 21856 66912
rect 22006 66898 22146 66912
rect 22296 66898 23104 66912
rect 23254 66898 23394 66912
rect 23544 66898 24352 66912
rect 24502 66898 24642 66912
rect 24792 66898 25600 66912
rect 25750 66898 25890 66912
rect 26040 66898 26848 66912
rect 26998 66898 27138 66912
rect 27288 66898 28096 66912
rect 28246 66898 28386 66912
rect 28536 66898 29344 66912
rect 29494 66898 29634 66912
rect 29784 66898 30592 66912
rect 30742 66898 30882 66912
rect 31032 66898 31840 66912
rect 31990 66898 32130 66912
rect 32280 66898 33088 66912
rect 33238 66898 33378 66912
rect 33528 66898 34336 66912
rect 34486 66898 34626 66912
rect 34776 66898 35584 66912
rect 35734 66898 35874 66912
rect 36024 66898 36832 66912
rect 36982 66898 37122 66912
rect 37272 66898 38080 66912
rect 38230 66898 38370 66912
rect 38520 66898 39328 66912
rect 39478 66898 39618 66912
rect 39768 66898 40576 66912
rect 40726 66898 40866 66912
rect 41016 66898 41824 66912
rect 41974 66898 42114 66912
rect 42264 66898 43072 66912
rect 43222 66898 43362 66912
rect 43512 66898 44320 66912
rect 44470 66898 44610 66912
rect 44760 66898 45568 66912
rect 45718 66898 45858 66912
rect 46008 66898 46816 66912
rect 46966 66898 47106 66912
rect 47256 66898 48064 66912
rect 48214 66898 48354 66912
rect 48504 66898 49312 66912
rect 49462 66898 49602 66912
rect 49752 66898 50560 66912
rect 50710 66898 50850 66912
rect 51000 66898 51808 66912
rect 51958 66898 52098 66912
rect 52248 66898 53056 66912
rect 53206 66898 53346 66912
rect 53496 66898 54304 66912
rect 54454 66898 54594 66912
rect 54744 66898 55552 66912
rect 55702 66898 55842 66912
rect 55992 66898 56800 66912
rect 56950 66898 57090 66912
rect 57240 66898 58048 66912
rect 58198 66898 58338 66912
rect 58488 66898 58934 66912
rect 16898 66850 16980 66864
rect 17188 66850 17270 66864
rect 18146 66850 18228 66864
rect 18436 66850 18518 66864
rect 19394 66850 19476 66864
rect 19684 66850 19766 66864
rect 20642 66850 20724 66864
rect 20932 66850 21014 66864
rect 21890 66850 21972 66864
rect 22180 66850 22262 66864
rect 23138 66850 23220 66864
rect 23428 66850 23510 66864
rect 24386 66850 24468 66864
rect 24676 66850 24758 66864
rect 25634 66850 25716 66864
rect 25924 66850 26006 66864
rect 26882 66850 26964 66864
rect 27172 66850 27254 66864
rect 28130 66850 28212 66864
rect 28420 66850 28502 66864
rect 29378 66850 29460 66864
rect 29668 66850 29750 66864
rect 30626 66850 30708 66864
rect 30916 66850 30998 66864
rect 31874 66850 31956 66864
rect 32164 66850 32246 66864
rect 33122 66850 33204 66864
rect 33412 66850 33494 66864
rect 34370 66850 34452 66864
rect 34660 66850 34742 66864
rect 35618 66850 35700 66864
rect 35908 66850 35990 66864
rect 36866 66850 36948 66864
rect 37156 66850 37238 66864
rect 38114 66850 38196 66864
rect 38404 66850 38486 66864
rect 39362 66850 39444 66864
rect 39652 66850 39734 66864
rect 40610 66850 40692 66864
rect 40900 66850 40982 66864
rect 41858 66850 41940 66864
rect 42148 66850 42230 66864
rect 43106 66850 43188 66864
rect 43396 66850 43478 66864
rect 44354 66850 44436 66864
rect 44644 66850 44726 66864
rect 45602 66850 45684 66864
rect 45892 66850 45974 66864
rect 46850 66850 46932 66864
rect 47140 66850 47222 66864
rect 48098 66850 48180 66864
rect 48388 66850 48470 66864
rect 49346 66850 49428 66864
rect 49636 66850 49718 66864
rect 50594 66850 50676 66864
rect 50884 66850 50966 66864
rect 51842 66850 51924 66864
rect 52132 66850 52214 66864
rect 53090 66850 53172 66864
rect 53380 66850 53462 66864
rect 54338 66850 54420 66864
rect 54628 66850 54710 66864
rect 55586 66850 55668 66864
rect 55876 66850 55958 66864
rect 56834 66850 56916 66864
rect 57124 66850 57206 66864
rect 58082 66850 58164 66864
rect 58372 66850 58454 66864
rect 16418 66802 58934 66850
rect 16418 66706 58934 66754
rect 16898 66692 16980 66706
rect 17188 66692 17270 66706
rect 18146 66692 18228 66706
rect 18436 66692 18518 66706
rect 19394 66692 19476 66706
rect 19684 66692 19766 66706
rect 20642 66692 20724 66706
rect 20932 66692 21014 66706
rect 21890 66692 21972 66706
rect 22180 66692 22262 66706
rect 23138 66692 23220 66706
rect 23428 66692 23510 66706
rect 24386 66692 24468 66706
rect 24676 66692 24758 66706
rect 25634 66692 25716 66706
rect 25924 66692 26006 66706
rect 26882 66692 26964 66706
rect 27172 66692 27254 66706
rect 28130 66692 28212 66706
rect 28420 66692 28502 66706
rect 29378 66692 29460 66706
rect 29668 66692 29750 66706
rect 30626 66692 30708 66706
rect 30916 66692 30998 66706
rect 31874 66692 31956 66706
rect 32164 66692 32246 66706
rect 33122 66692 33204 66706
rect 33412 66692 33494 66706
rect 34370 66692 34452 66706
rect 34660 66692 34742 66706
rect 35618 66692 35700 66706
rect 35908 66692 35990 66706
rect 36866 66692 36948 66706
rect 37156 66692 37238 66706
rect 38114 66692 38196 66706
rect 38404 66692 38486 66706
rect 39362 66692 39444 66706
rect 39652 66692 39734 66706
rect 40610 66692 40692 66706
rect 40900 66692 40982 66706
rect 41858 66692 41940 66706
rect 42148 66692 42230 66706
rect 43106 66692 43188 66706
rect 43396 66692 43478 66706
rect 44354 66692 44436 66706
rect 44644 66692 44726 66706
rect 45602 66692 45684 66706
rect 45892 66692 45974 66706
rect 46850 66692 46932 66706
rect 47140 66692 47222 66706
rect 48098 66692 48180 66706
rect 48388 66692 48470 66706
rect 49346 66692 49428 66706
rect 49636 66692 49718 66706
rect 50594 66692 50676 66706
rect 50884 66692 50966 66706
rect 51842 66692 51924 66706
rect 52132 66692 52214 66706
rect 53090 66692 53172 66706
rect 53380 66692 53462 66706
rect 54338 66692 54420 66706
rect 54628 66692 54710 66706
rect 55586 66692 55668 66706
rect 55876 66692 55958 66706
rect 56834 66692 56916 66706
rect 57124 66692 57206 66706
rect 58082 66692 58164 66706
rect 58372 66692 58454 66706
rect 16418 66644 16864 66658
rect 17014 66644 17154 66658
rect 17304 66644 18112 66658
rect 18262 66644 18402 66658
rect 18552 66644 19360 66658
rect 19510 66644 19650 66658
rect 19800 66644 20608 66658
rect 20758 66644 20898 66658
rect 21048 66644 21856 66658
rect 22006 66644 22146 66658
rect 22296 66644 23104 66658
rect 23254 66644 23394 66658
rect 23544 66644 24352 66658
rect 24502 66644 24642 66658
rect 24792 66644 25600 66658
rect 25750 66644 25890 66658
rect 26040 66644 26848 66658
rect 26998 66644 27138 66658
rect 27288 66644 28096 66658
rect 28246 66644 28386 66658
rect 28536 66644 29344 66658
rect 29494 66644 29634 66658
rect 29784 66644 30592 66658
rect 30742 66644 30882 66658
rect 31032 66644 31840 66658
rect 31990 66644 32130 66658
rect 32280 66644 33088 66658
rect 33238 66644 33378 66658
rect 33528 66644 34336 66658
rect 34486 66644 34626 66658
rect 34776 66644 35584 66658
rect 35734 66644 35874 66658
rect 36024 66644 36832 66658
rect 36982 66644 37122 66658
rect 37272 66644 38080 66658
rect 38230 66644 38370 66658
rect 38520 66644 39328 66658
rect 39478 66644 39618 66658
rect 39768 66644 40576 66658
rect 40726 66644 40866 66658
rect 41016 66644 41824 66658
rect 41974 66644 42114 66658
rect 42264 66644 43072 66658
rect 43222 66644 43362 66658
rect 43512 66644 44320 66658
rect 44470 66644 44610 66658
rect 44760 66644 45568 66658
rect 45718 66644 45858 66658
rect 46008 66644 46816 66658
rect 46966 66644 47106 66658
rect 47256 66644 48064 66658
rect 48214 66644 48354 66658
rect 48504 66644 49312 66658
rect 49462 66644 49602 66658
rect 49752 66644 50560 66658
rect 50710 66644 50850 66658
rect 51000 66644 51808 66658
rect 51958 66644 52098 66658
rect 52248 66644 53056 66658
rect 53206 66644 53346 66658
rect 53496 66644 54304 66658
rect 54454 66644 54594 66658
rect 54744 66644 55552 66658
rect 55702 66644 55842 66658
rect 55992 66644 56800 66658
rect 56950 66644 57090 66658
rect 57240 66644 58048 66658
rect 58198 66644 58338 66658
rect 58488 66644 58934 66658
rect 16418 66596 58934 66644
rect 16418 66582 16864 66596
rect 17014 66582 17154 66596
rect 17304 66582 18112 66596
rect 18262 66582 18402 66596
rect 18552 66582 19360 66596
rect 19510 66582 19650 66596
rect 19800 66582 20608 66596
rect 20758 66582 20898 66596
rect 21048 66582 21856 66596
rect 22006 66582 22146 66596
rect 22296 66582 23104 66596
rect 23254 66582 23394 66596
rect 23544 66582 24352 66596
rect 24502 66582 24642 66596
rect 24792 66582 25600 66596
rect 25750 66582 25890 66596
rect 26040 66582 26848 66596
rect 26998 66582 27138 66596
rect 27288 66582 28096 66596
rect 28246 66582 28386 66596
rect 28536 66582 29344 66596
rect 29494 66582 29634 66596
rect 29784 66582 30592 66596
rect 30742 66582 30882 66596
rect 31032 66582 31840 66596
rect 31990 66582 32130 66596
rect 32280 66582 33088 66596
rect 33238 66582 33378 66596
rect 33528 66582 34336 66596
rect 34486 66582 34626 66596
rect 34776 66582 35584 66596
rect 35734 66582 35874 66596
rect 36024 66582 36832 66596
rect 36982 66582 37122 66596
rect 37272 66582 38080 66596
rect 38230 66582 38370 66596
rect 38520 66582 39328 66596
rect 39478 66582 39618 66596
rect 39768 66582 40576 66596
rect 40726 66582 40866 66596
rect 41016 66582 41824 66596
rect 41974 66582 42114 66596
rect 42264 66582 43072 66596
rect 43222 66582 43362 66596
rect 43512 66582 44320 66596
rect 44470 66582 44610 66596
rect 44760 66582 45568 66596
rect 45718 66582 45858 66596
rect 46008 66582 46816 66596
rect 46966 66582 47106 66596
rect 47256 66582 48064 66596
rect 48214 66582 48354 66596
rect 48504 66582 49312 66596
rect 49462 66582 49602 66596
rect 49752 66582 50560 66596
rect 50710 66582 50850 66596
rect 51000 66582 51808 66596
rect 51958 66582 52098 66596
rect 52248 66582 53056 66596
rect 53206 66582 53346 66596
rect 53496 66582 54304 66596
rect 54454 66582 54594 66596
rect 54744 66582 55552 66596
rect 55702 66582 55842 66596
rect 55992 66582 56800 66596
rect 56950 66582 57090 66596
rect 57240 66582 58048 66596
rect 58198 66582 58338 66596
rect 58488 66582 58934 66596
rect 16898 66534 16980 66548
rect 17188 66534 17270 66548
rect 18146 66534 18228 66548
rect 18436 66534 18518 66548
rect 19394 66534 19476 66548
rect 19684 66534 19766 66548
rect 20642 66534 20724 66548
rect 20932 66534 21014 66548
rect 21890 66534 21972 66548
rect 22180 66534 22262 66548
rect 23138 66534 23220 66548
rect 23428 66534 23510 66548
rect 24386 66534 24468 66548
rect 24676 66534 24758 66548
rect 25634 66534 25716 66548
rect 25924 66534 26006 66548
rect 26882 66534 26964 66548
rect 27172 66534 27254 66548
rect 28130 66534 28212 66548
rect 28420 66534 28502 66548
rect 29378 66534 29460 66548
rect 29668 66534 29750 66548
rect 30626 66534 30708 66548
rect 30916 66534 30998 66548
rect 31874 66534 31956 66548
rect 32164 66534 32246 66548
rect 33122 66534 33204 66548
rect 33412 66534 33494 66548
rect 34370 66534 34452 66548
rect 34660 66534 34742 66548
rect 35618 66534 35700 66548
rect 35908 66534 35990 66548
rect 36866 66534 36948 66548
rect 37156 66534 37238 66548
rect 38114 66534 38196 66548
rect 38404 66534 38486 66548
rect 39362 66534 39444 66548
rect 39652 66534 39734 66548
rect 40610 66534 40692 66548
rect 40900 66534 40982 66548
rect 41858 66534 41940 66548
rect 42148 66534 42230 66548
rect 43106 66534 43188 66548
rect 43396 66534 43478 66548
rect 44354 66534 44436 66548
rect 44644 66534 44726 66548
rect 45602 66534 45684 66548
rect 45892 66534 45974 66548
rect 46850 66534 46932 66548
rect 47140 66534 47222 66548
rect 48098 66534 48180 66548
rect 48388 66534 48470 66548
rect 49346 66534 49428 66548
rect 49636 66534 49718 66548
rect 50594 66534 50676 66548
rect 50884 66534 50966 66548
rect 51842 66534 51924 66548
rect 52132 66534 52214 66548
rect 53090 66534 53172 66548
rect 53380 66534 53462 66548
rect 54338 66534 54420 66548
rect 54628 66534 54710 66548
rect 55586 66534 55668 66548
rect 55876 66534 55958 66548
rect 56834 66534 56916 66548
rect 57124 66534 57206 66548
rect 58082 66534 58164 66548
rect 58372 66534 58454 66548
rect 16418 66486 58934 66534
rect 16418 66328 58934 66438
rect 16418 66232 58934 66280
rect 16898 66218 16980 66232
rect 17188 66218 17270 66232
rect 18146 66218 18228 66232
rect 18436 66218 18518 66232
rect 19394 66218 19476 66232
rect 19684 66218 19766 66232
rect 20642 66218 20724 66232
rect 20932 66218 21014 66232
rect 21890 66218 21972 66232
rect 22180 66218 22262 66232
rect 23138 66218 23220 66232
rect 23428 66218 23510 66232
rect 24386 66218 24468 66232
rect 24676 66218 24758 66232
rect 25634 66218 25716 66232
rect 25924 66218 26006 66232
rect 26882 66218 26964 66232
rect 27172 66218 27254 66232
rect 28130 66218 28212 66232
rect 28420 66218 28502 66232
rect 29378 66218 29460 66232
rect 29668 66218 29750 66232
rect 30626 66218 30708 66232
rect 30916 66218 30998 66232
rect 31874 66218 31956 66232
rect 32164 66218 32246 66232
rect 33122 66218 33204 66232
rect 33412 66218 33494 66232
rect 34370 66218 34452 66232
rect 34660 66218 34742 66232
rect 35618 66218 35700 66232
rect 35908 66218 35990 66232
rect 36866 66218 36948 66232
rect 37156 66218 37238 66232
rect 38114 66218 38196 66232
rect 38404 66218 38486 66232
rect 39362 66218 39444 66232
rect 39652 66218 39734 66232
rect 40610 66218 40692 66232
rect 40900 66218 40982 66232
rect 41858 66218 41940 66232
rect 42148 66218 42230 66232
rect 43106 66218 43188 66232
rect 43396 66218 43478 66232
rect 44354 66218 44436 66232
rect 44644 66218 44726 66232
rect 45602 66218 45684 66232
rect 45892 66218 45974 66232
rect 46850 66218 46932 66232
rect 47140 66218 47222 66232
rect 48098 66218 48180 66232
rect 48388 66218 48470 66232
rect 49346 66218 49428 66232
rect 49636 66218 49718 66232
rect 50594 66218 50676 66232
rect 50884 66218 50966 66232
rect 51842 66218 51924 66232
rect 52132 66218 52214 66232
rect 53090 66218 53172 66232
rect 53380 66218 53462 66232
rect 54338 66218 54420 66232
rect 54628 66218 54710 66232
rect 55586 66218 55668 66232
rect 55876 66218 55958 66232
rect 56834 66218 56916 66232
rect 57124 66218 57206 66232
rect 58082 66218 58164 66232
rect 58372 66218 58454 66232
rect 16418 66170 16864 66184
rect 17014 66170 17154 66184
rect 17304 66170 18112 66184
rect 18262 66170 18402 66184
rect 18552 66170 19360 66184
rect 19510 66170 19650 66184
rect 19800 66170 20608 66184
rect 20758 66170 20898 66184
rect 21048 66170 21856 66184
rect 22006 66170 22146 66184
rect 22296 66170 23104 66184
rect 23254 66170 23394 66184
rect 23544 66170 24352 66184
rect 24502 66170 24642 66184
rect 24792 66170 25600 66184
rect 25750 66170 25890 66184
rect 26040 66170 26848 66184
rect 26998 66170 27138 66184
rect 27288 66170 28096 66184
rect 28246 66170 28386 66184
rect 28536 66170 29344 66184
rect 29494 66170 29634 66184
rect 29784 66170 30592 66184
rect 30742 66170 30882 66184
rect 31032 66170 31840 66184
rect 31990 66170 32130 66184
rect 32280 66170 33088 66184
rect 33238 66170 33378 66184
rect 33528 66170 34336 66184
rect 34486 66170 34626 66184
rect 34776 66170 35584 66184
rect 35734 66170 35874 66184
rect 36024 66170 36832 66184
rect 36982 66170 37122 66184
rect 37272 66170 38080 66184
rect 38230 66170 38370 66184
rect 38520 66170 39328 66184
rect 39478 66170 39618 66184
rect 39768 66170 40576 66184
rect 40726 66170 40866 66184
rect 41016 66170 41824 66184
rect 41974 66170 42114 66184
rect 42264 66170 43072 66184
rect 43222 66170 43362 66184
rect 43512 66170 44320 66184
rect 44470 66170 44610 66184
rect 44760 66170 45568 66184
rect 45718 66170 45858 66184
rect 46008 66170 46816 66184
rect 46966 66170 47106 66184
rect 47256 66170 48064 66184
rect 48214 66170 48354 66184
rect 48504 66170 49312 66184
rect 49462 66170 49602 66184
rect 49752 66170 50560 66184
rect 50710 66170 50850 66184
rect 51000 66170 51808 66184
rect 51958 66170 52098 66184
rect 52248 66170 53056 66184
rect 53206 66170 53346 66184
rect 53496 66170 54304 66184
rect 54454 66170 54594 66184
rect 54744 66170 55552 66184
rect 55702 66170 55842 66184
rect 55992 66170 56800 66184
rect 56950 66170 57090 66184
rect 57240 66170 58048 66184
rect 58198 66170 58338 66184
rect 58488 66170 58934 66184
rect 16418 66122 58934 66170
rect 16418 66108 16864 66122
rect 17014 66108 17154 66122
rect 17304 66108 18112 66122
rect 18262 66108 18402 66122
rect 18552 66108 19360 66122
rect 19510 66108 19650 66122
rect 19800 66108 20608 66122
rect 20758 66108 20898 66122
rect 21048 66108 21856 66122
rect 22006 66108 22146 66122
rect 22296 66108 23104 66122
rect 23254 66108 23394 66122
rect 23544 66108 24352 66122
rect 24502 66108 24642 66122
rect 24792 66108 25600 66122
rect 25750 66108 25890 66122
rect 26040 66108 26848 66122
rect 26998 66108 27138 66122
rect 27288 66108 28096 66122
rect 28246 66108 28386 66122
rect 28536 66108 29344 66122
rect 29494 66108 29634 66122
rect 29784 66108 30592 66122
rect 30742 66108 30882 66122
rect 31032 66108 31840 66122
rect 31990 66108 32130 66122
rect 32280 66108 33088 66122
rect 33238 66108 33378 66122
rect 33528 66108 34336 66122
rect 34486 66108 34626 66122
rect 34776 66108 35584 66122
rect 35734 66108 35874 66122
rect 36024 66108 36832 66122
rect 36982 66108 37122 66122
rect 37272 66108 38080 66122
rect 38230 66108 38370 66122
rect 38520 66108 39328 66122
rect 39478 66108 39618 66122
rect 39768 66108 40576 66122
rect 40726 66108 40866 66122
rect 41016 66108 41824 66122
rect 41974 66108 42114 66122
rect 42264 66108 43072 66122
rect 43222 66108 43362 66122
rect 43512 66108 44320 66122
rect 44470 66108 44610 66122
rect 44760 66108 45568 66122
rect 45718 66108 45858 66122
rect 46008 66108 46816 66122
rect 46966 66108 47106 66122
rect 47256 66108 48064 66122
rect 48214 66108 48354 66122
rect 48504 66108 49312 66122
rect 49462 66108 49602 66122
rect 49752 66108 50560 66122
rect 50710 66108 50850 66122
rect 51000 66108 51808 66122
rect 51958 66108 52098 66122
rect 52248 66108 53056 66122
rect 53206 66108 53346 66122
rect 53496 66108 54304 66122
rect 54454 66108 54594 66122
rect 54744 66108 55552 66122
rect 55702 66108 55842 66122
rect 55992 66108 56800 66122
rect 56950 66108 57090 66122
rect 57240 66108 58048 66122
rect 58198 66108 58338 66122
rect 58488 66108 58934 66122
rect 16898 66060 16980 66074
rect 17188 66060 17270 66074
rect 18146 66060 18228 66074
rect 18436 66060 18518 66074
rect 19394 66060 19476 66074
rect 19684 66060 19766 66074
rect 20642 66060 20724 66074
rect 20932 66060 21014 66074
rect 21890 66060 21972 66074
rect 22180 66060 22262 66074
rect 23138 66060 23220 66074
rect 23428 66060 23510 66074
rect 24386 66060 24468 66074
rect 24676 66060 24758 66074
rect 25634 66060 25716 66074
rect 25924 66060 26006 66074
rect 26882 66060 26964 66074
rect 27172 66060 27254 66074
rect 28130 66060 28212 66074
rect 28420 66060 28502 66074
rect 29378 66060 29460 66074
rect 29668 66060 29750 66074
rect 30626 66060 30708 66074
rect 30916 66060 30998 66074
rect 31874 66060 31956 66074
rect 32164 66060 32246 66074
rect 33122 66060 33204 66074
rect 33412 66060 33494 66074
rect 34370 66060 34452 66074
rect 34660 66060 34742 66074
rect 35618 66060 35700 66074
rect 35908 66060 35990 66074
rect 36866 66060 36948 66074
rect 37156 66060 37238 66074
rect 38114 66060 38196 66074
rect 38404 66060 38486 66074
rect 39362 66060 39444 66074
rect 39652 66060 39734 66074
rect 40610 66060 40692 66074
rect 40900 66060 40982 66074
rect 41858 66060 41940 66074
rect 42148 66060 42230 66074
rect 43106 66060 43188 66074
rect 43396 66060 43478 66074
rect 44354 66060 44436 66074
rect 44644 66060 44726 66074
rect 45602 66060 45684 66074
rect 45892 66060 45974 66074
rect 46850 66060 46932 66074
rect 47140 66060 47222 66074
rect 48098 66060 48180 66074
rect 48388 66060 48470 66074
rect 49346 66060 49428 66074
rect 49636 66060 49718 66074
rect 50594 66060 50676 66074
rect 50884 66060 50966 66074
rect 51842 66060 51924 66074
rect 52132 66060 52214 66074
rect 53090 66060 53172 66074
rect 53380 66060 53462 66074
rect 54338 66060 54420 66074
rect 54628 66060 54710 66074
rect 55586 66060 55668 66074
rect 55876 66060 55958 66074
rect 56834 66060 56916 66074
rect 57124 66060 57206 66074
rect 58082 66060 58164 66074
rect 58372 66060 58454 66074
rect 16418 66012 58934 66060
rect 16418 65916 58934 65964
rect 16898 65902 16980 65916
rect 17188 65902 17270 65916
rect 18146 65902 18228 65916
rect 18436 65902 18518 65916
rect 19394 65902 19476 65916
rect 19684 65902 19766 65916
rect 20642 65902 20724 65916
rect 20932 65902 21014 65916
rect 21890 65902 21972 65916
rect 22180 65902 22262 65916
rect 23138 65902 23220 65916
rect 23428 65902 23510 65916
rect 24386 65902 24468 65916
rect 24676 65902 24758 65916
rect 25634 65902 25716 65916
rect 25924 65902 26006 65916
rect 26882 65902 26964 65916
rect 27172 65902 27254 65916
rect 28130 65902 28212 65916
rect 28420 65902 28502 65916
rect 29378 65902 29460 65916
rect 29668 65902 29750 65916
rect 30626 65902 30708 65916
rect 30916 65902 30998 65916
rect 31874 65902 31956 65916
rect 32164 65902 32246 65916
rect 33122 65902 33204 65916
rect 33412 65902 33494 65916
rect 34370 65902 34452 65916
rect 34660 65902 34742 65916
rect 35618 65902 35700 65916
rect 35908 65902 35990 65916
rect 36866 65902 36948 65916
rect 37156 65902 37238 65916
rect 38114 65902 38196 65916
rect 38404 65902 38486 65916
rect 39362 65902 39444 65916
rect 39652 65902 39734 65916
rect 40610 65902 40692 65916
rect 40900 65902 40982 65916
rect 41858 65902 41940 65916
rect 42148 65902 42230 65916
rect 43106 65902 43188 65916
rect 43396 65902 43478 65916
rect 44354 65902 44436 65916
rect 44644 65902 44726 65916
rect 45602 65902 45684 65916
rect 45892 65902 45974 65916
rect 46850 65902 46932 65916
rect 47140 65902 47222 65916
rect 48098 65902 48180 65916
rect 48388 65902 48470 65916
rect 49346 65902 49428 65916
rect 49636 65902 49718 65916
rect 50594 65902 50676 65916
rect 50884 65902 50966 65916
rect 51842 65902 51924 65916
rect 52132 65902 52214 65916
rect 53090 65902 53172 65916
rect 53380 65902 53462 65916
rect 54338 65902 54420 65916
rect 54628 65902 54710 65916
rect 55586 65902 55668 65916
rect 55876 65902 55958 65916
rect 56834 65902 56916 65916
rect 57124 65902 57206 65916
rect 58082 65902 58164 65916
rect 58372 65902 58454 65916
rect 16418 65854 16864 65868
rect 17014 65854 17154 65868
rect 17304 65854 18112 65868
rect 18262 65854 18402 65868
rect 18552 65854 19360 65868
rect 19510 65854 19650 65868
rect 19800 65854 20608 65868
rect 20758 65854 20898 65868
rect 21048 65854 21856 65868
rect 22006 65854 22146 65868
rect 22296 65854 23104 65868
rect 23254 65854 23394 65868
rect 23544 65854 24352 65868
rect 24502 65854 24642 65868
rect 24792 65854 25600 65868
rect 25750 65854 25890 65868
rect 26040 65854 26848 65868
rect 26998 65854 27138 65868
rect 27288 65854 28096 65868
rect 28246 65854 28386 65868
rect 28536 65854 29344 65868
rect 29494 65854 29634 65868
rect 29784 65854 30592 65868
rect 30742 65854 30882 65868
rect 31032 65854 31840 65868
rect 31990 65854 32130 65868
rect 32280 65854 33088 65868
rect 33238 65854 33378 65868
rect 33528 65854 34336 65868
rect 34486 65854 34626 65868
rect 34776 65854 35584 65868
rect 35734 65854 35874 65868
rect 36024 65854 36832 65868
rect 36982 65854 37122 65868
rect 37272 65854 38080 65868
rect 38230 65854 38370 65868
rect 38520 65854 39328 65868
rect 39478 65854 39618 65868
rect 39768 65854 40576 65868
rect 40726 65854 40866 65868
rect 41016 65854 41824 65868
rect 41974 65854 42114 65868
rect 42264 65854 43072 65868
rect 43222 65854 43362 65868
rect 43512 65854 44320 65868
rect 44470 65854 44610 65868
rect 44760 65854 45568 65868
rect 45718 65854 45858 65868
rect 46008 65854 46816 65868
rect 46966 65854 47106 65868
rect 47256 65854 48064 65868
rect 48214 65854 48354 65868
rect 48504 65854 49312 65868
rect 49462 65854 49602 65868
rect 49752 65854 50560 65868
rect 50710 65854 50850 65868
rect 51000 65854 51808 65868
rect 51958 65854 52098 65868
rect 52248 65854 53056 65868
rect 53206 65854 53346 65868
rect 53496 65854 54304 65868
rect 54454 65854 54594 65868
rect 54744 65854 55552 65868
rect 55702 65854 55842 65868
rect 55992 65854 56800 65868
rect 56950 65854 57090 65868
rect 57240 65854 58048 65868
rect 58198 65854 58338 65868
rect 58488 65854 58934 65868
rect 16418 65806 58934 65854
rect 16418 65792 16864 65806
rect 17014 65792 17154 65806
rect 17304 65792 18112 65806
rect 18262 65792 18402 65806
rect 18552 65792 19360 65806
rect 19510 65792 19650 65806
rect 19800 65792 20608 65806
rect 20758 65792 20898 65806
rect 21048 65792 21856 65806
rect 22006 65792 22146 65806
rect 22296 65792 23104 65806
rect 23254 65792 23394 65806
rect 23544 65792 24352 65806
rect 24502 65792 24642 65806
rect 24792 65792 25600 65806
rect 25750 65792 25890 65806
rect 26040 65792 26848 65806
rect 26998 65792 27138 65806
rect 27288 65792 28096 65806
rect 28246 65792 28386 65806
rect 28536 65792 29344 65806
rect 29494 65792 29634 65806
rect 29784 65792 30592 65806
rect 30742 65792 30882 65806
rect 31032 65792 31840 65806
rect 31990 65792 32130 65806
rect 32280 65792 33088 65806
rect 33238 65792 33378 65806
rect 33528 65792 34336 65806
rect 34486 65792 34626 65806
rect 34776 65792 35584 65806
rect 35734 65792 35874 65806
rect 36024 65792 36832 65806
rect 36982 65792 37122 65806
rect 37272 65792 38080 65806
rect 38230 65792 38370 65806
rect 38520 65792 39328 65806
rect 39478 65792 39618 65806
rect 39768 65792 40576 65806
rect 40726 65792 40866 65806
rect 41016 65792 41824 65806
rect 41974 65792 42114 65806
rect 42264 65792 43072 65806
rect 43222 65792 43362 65806
rect 43512 65792 44320 65806
rect 44470 65792 44610 65806
rect 44760 65792 45568 65806
rect 45718 65792 45858 65806
rect 46008 65792 46816 65806
rect 46966 65792 47106 65806
rect 47256 65792 48064 65806
rect 48214 65792 48354 65806
rect 48504 65792 49312 65806
rect 49462 65792 49602 65806
rect 49752 65792 50560 65806
rect 50710 65792 50850 65806
rect 51000 65792 51808 65806
rect 51958 65792 52098 65806
rect 52248 65792 53056 65806
rect 53206 65792 53346 65806
rect 53496 65792 54304 65806
rect 54454 65792 54594 65806
rect 54744 65792 55552 65806
rect 55702 65792 55842 65806
rect 55992 65792 56800 65806
rect 56950 65792 57090 65806
rect 57240 65792 58048 65806
rect 58198 65792 58338 65806
rect 58488 65792 58934 65806
rect 16898 65744 16980 65758
rect 17188 65744 17270 65758
rect 18146 65744 18228 65758
rect 18436 65744 18518 65758
rect 19394 65744 19476 65758
rect 19684 65744 19766 65758
rect 20642 65744 20724 65758
rect 20932 65744 21014 65758
rect 21890 65744 21972 65758
rect 22180 65744 22262 65758
rect 23138 65744 23220 65758
rect 23428 65744 23510 65758
rect 24386 65744 24468 65758
rect 24676 65744 24758 65758
rect 25634 65744 25716 65758
rect 25924 65744 26006 65758
rect 26882 65744 26964 65758
rect 27172 65744 27254 65758
rect 28130 65744 28212 65758
rect 28420 65744 28502 65758
rect 29378 65744 29460 65758
rect 29668 65744 29750 65758
rect 30626 65744 30708 65758
rect 30916 65744 30998 65758
rect 31874 65744 31956 65758
rect 32164 65744 32246 65758
rect 33122 65744 33204 65758
rect 33412 65744 33494 65758
rect 34370 65744 34452 65758
rect 34660 65744 34742 65758
rect 35618 65744 35700 65758
rect 35908 65744 35990 65758
rect 36866 65744 36948 65758
rect 37156 65744 37238 65758
rect 38114 65744 38196 65758
rect 38404 65744 38486 65758
rect 39362 65744 39444 65758
rect 39652 65744 39734 65758
rect 40610 65744 40692 65758
rect 40900 65744 40982 65758
rect 41858 65744 41940 65758
rect 42148 65744 42230 65758
rect 43106 65744 43188 65758
rect 43396 65744 43478 65758
rect 44354 65744 44436 65758
rect 44644 65744 44726 65758
rect 45602 65744 45684 65758
rect 45892 65744 45974 65758
rect 46850 65744 46932 65758
rect 47140 65744 47222 65758
rect 48098 65744 48180 65758
rect 48388 65744 48470 65758
rect 49346 65744 49428 65758
rect 49636 65744 49718 65758
rect 50594 65744 50676 65758
rect 50884 65744 50966 65758
rect 51842 65744 51924 65758
rect 52132 65744 52214 65758
rect 53090 65744 53172 65758
rect 53380 65744 53462 65758
rect 54338 65744 54420 65758
rect 54628 65744 54710 65758
rect 55586 65744 55668 65758
rect 55876 65744 55958 65758
rect 56834 65744 56916 65758
rect 57124 65744 57206 65758
rect 58082 65744 58164 65758
rect 58372 65744 58454 65758
rect 16418 65696 58934 65744
rect 16418 65538 58934 65648
rect 16418 65442 58934 65490
rect 16898 65428 16980 65442
rect 17188 65428 17270 65442
rect 18146 65428 18228 65442
rect 18436 65428 18518 65442
rect 19394 65428 19476 65442
rect 19684 65428 19766 65442
rect 20642 65428 20724 65442
rect 20932 65428 21014 65442
rect 21890 65428 21972 65442
rect 22180 65428 22262 65442
rect 23138 65428 23220 65442
rect 23428 65428 23510 65442
rect 24386 65428 24468 65442
rect 24676 65428 24758 65442
rect 25634 65428 25716 65442
rect 25924 65428 26006 65442
rect 26882 65428 26964 65442
rect 27172 65428 27254 65442
rect 28130 65428 28212 65442
rect 28420 65428 28502 65442
rect 29378 65428 29460 65442
rect 29668 65428 29750 65442
rect 30626 65428 30708 65442
rect 30916 65428 30998 65442
rect 31874 65428 31956 65442
rect 32164 65428 32246 65442
rect 33122 65428 33204 65442
rect 33412 65428 33494 65442
rect 34370 65428 34452 65442
rect 34660 65428 34742 65442
rect 35618 65428 35700 65442
rect 35908 65428 35990 65442
rect 36866 65428 36948 65442
rect 37156 65428 37238 65442
rect 38114 65428 38196 65442
rect 38404 65428 38486 65442
rect 39362 65428 39444 65442
rect 39652 65428 39734 65442
rect 40610 65428 40692 65442
rect 40900 65428 40982 65442
rect 41858 65428 41940 65442
rect 42148 65428 42230 65442
rect 43106 65428 43188 65442
rect 43396 65428 43478 65442
rect 44354 65428 44436 65442
rect 44644 65428 44726 65442
rect 45602 65428 45684 65442
rect 45892 65428 45974 65442
rect 46850 65428 46932 65442
rect 47140 65428 47222 65442
rect 48098 65428 48180 65442
rect 48388 65428 48470 65442
rect 49346 65428 49428 65442
rect 49636 65428 49718 65442
rect 50594 65428 50676 65442
rect 50884 65428 50966 65442
rect 51842 65428 51924 65442
rect 52132 65428 52214 65442
rect 53090 65428 53172 65442
rect 53380 65428 53462 65442
rect 54338 65428 54420 65442
rect 54628 65428 54710 65442
rect 55586 65428 55668 65442
rect 55876 65428 55958 65442
rect 56834 65428 56916 65442
rect 57124 65428 57206 65442
rect 58082 65428 58164 65442
rect 58372 65428 58454 65442
rect 16418 65380 16864 65394
rect 17014 65380 17154 65394
rect 17304 65380 18112 65394
rect 18262 65380 18402 65394
rect 18552 65380 19360 65394
rect 19510 65380 19650 65394
rect 19800 65380 20608 65394
rect 20758 65380 20898 65394
rect 21048 65380 21856 65394
rect 22006 65380 22146 65394
rect 22296 65380 23104 65394
rect 23254 65380 23394 65394
rect 23544 65380 24352 65394
rect 24502 65380 24642 65394
rect 24792 65380 25600 65394
rect 25750 65380 25890 65394
rect 26040 65380 26848 65394
rect 26998 65380 27138 65394
rect 27288 65380 28096 65394
rect 28246 65380 28386 65394
rect 28536 65380 29344 65394
rect 29494 65380 29634 65394
rect 29784 65380 30592 65394
rect 30742 65380 30882 65394
rect 31032 65380 31840 65394
rect 31990 65380 32130 65394
rect 32280 65380 33088 65394
rect 33238 65380 33378 65394
rect 33528 65380 34336 65394
rect 34486 65380 34626 65394
rect 34776 65380 35584 65394
rect 35734 65380 35874 65394
rect 36024 65380 36832 65394
rect 36982 65380 37122 65394
rect 37272 65380 38080 65394
rect 38230 65380 38370 65394
rect 38520 65380 39328 65394
rect 39478 65380 39618 65394
rect 39768 65380 40576 65394
rect 40726 65380 40866 65394
rect 41016 65380 41824 65394
rect 41974 65380 42114 65394
rect 42264 65380 43072 65394
rect 43222 65380 43362 65394
rect 43512 65380 44320 65394
rect 44470 65380 44610 65394
rect 44760 65380 45568 65394
rect 45718 65380 45858 65394
rect 46008 65380 46816 65394
rect 46966 65380 47106 65394
rect 47256 65380 48064 65394
rect 48214 65380 48354 65394
rect 48504 65380 49312 65394
rect 49462 65380 49602 65394
rect 49752 65380 50560 65394
rect 50710 65380 50850 65394
rect 51000 65380 51808 65394
rect 51958 65380 52098 65394
rect 52248 65380 53056 65394
rect 53206 65380 53346 65394
rect 53496 65380 54304 65394
rect 54454 65380 54594 65394
rect 54744 65380 55552 65394
rect 55702 65380 55842 65394
rect 55992 65380 56800 65394
rect 56950 65380 57090 65394
rect 57240 65380 58048 65394
rect 58198 65380 58338 65394
rect 58488 65380 58934 65394
rect 16418 65332 58934 65380
rect 16418 65318 16864 65332
rect 17014 65318 17154 65332
rect 17304 65318 18112 65332
rect 18262 65318 18402 65332
rect 18552 65318 19360 65332
rect 19510 65318 19650 65332
rect 19800 65318 20608 65332
rect 20758 65318 20898 65332
rect 21048 65318 21856 65332
rect 22006 65318 22146 65332
rect 22296 65318 23104 65332
rect 23254 65318 23394 65332
rect 23544 65318 24352 65332
rect 24502 65318 24642 65332
rect 24792 65318 25600 65332
rect 25750 65318 25890 65332
rect 26040 65318 26848 65332
rect 26998 65318 27138 65332
rect 27288 65318 28096 65332
rect 28246 65318 28386 65332
rect 28536 65318 29344 65332
rect 29494 65318 29634 65332
rect 29784 65318 30592 65332
rect 30742 65318 30882 65332
rect 31032 65318 31840 65332
rect 31990 65318 32130 65332
rect 32280 65318 33088 65332
rect 33238 65318 33378 65332
rect 33528 65318 34336 65332
rect 34486 65318 34626 65332
rect 34776 65318 35584 65332
rect 35734 65318 35874 65332
rect 36024 65318 36832 65332
rect 36982 65318 37122 65332
rect 37272 65318 38080 65332
rect 38230 65318 38370 65332
rect 38520 65318 39328 65332
rect 39478 65318 39618 65332
rect 39768 65318 40576 65332
rect 40726 65318 40866 65332
rect 41016 65318 41824 65332
rect 41974 65318 42114 65332
rect 42264 65318 43072 65332
rect 43222 65318 43362 65332
rect 43512 65318 44320 65332
rect 44470 65318 44610 65332
rect 44760 65318 45568 65332
rect 45718 65318 45858 65332
rect 46008 65318 46816 65332
rect 46966 65318 47106 65332
rect 47256 65318 48064 65332
rect 48214 65318 48354 65332
rect 48504 65318 49312 65332
rect 49462 65318 49602 65332
rect 49752 65318 50560 65332
rect 50710 65318 50850 65332
rect 51000 65318 51808 65332
rect 51958 65318 52098 65332
rect 52248 65318 53056 65332
rect 53206 65318 53346 65332
rect 53496 65318 54304 65332
rect 54454 65318 54594 65332
rect 54744 65318 55552 65332
rect 55702 65318 55842 65332
rect 55992 65318 56800 65332
rect 56950 65318 57090 65332
rect 57240 65318 58048 65332
rect 58198 65318 58338 65332
rect 58488 65318 58934 65332
rect 16898 65270 16980 65284
rect 17188 65270 17270 65284
rect 18146 65270 18228 65284
rect 18436 65270 18518 65284
rect 19394 65270 19476 65284
rect 19684 65270 19766 65284
rect 20642 65270 20724 65284
rect 20932 65270 21014 65284
rect 21890 65270 21972 65284
rect 22180 65270 22262 65284
rect 23138 65270 23220 65284
rect 23428 65270 23510 65284
rect 24386 65270 24468 65284
rect 24676 65270 24758 65284
rect 25634 65270 25716 65284
rect 25924 65270 26006 65284
rect 26882 65270 26964 65284
rect 27172 65270 27254 65284
rect 28130 65270 28212 65284
rect 28420 65270 28502 65284
rect 29378 65270 29460 65284
rect 29668 65270 29750 65284
rect 30626 65270 30708 65284
rect 30916 65270 30998 65284
rect 31874 65270 31956 65284
rect 32164 65270 32246 65284
rect 33122 65270 33204 65284
rect 33412 65270 33494 65284
rect 34370 65270 34452 65284
rect 34660 65270 34742 65284
rect 35618 65270 35700 65284
rect 35908 65270 35990 65284
rect 36866 65270 36948 65284
rect 37156 65270 37238 65284
rect 38114 65270 38196 65284
rect 38404 65270 38486 65284
rect 39362 65270 39444 65284
rect 39652 65270 39734 65284
rect 40610 65270 40692 65284
rect 40900 65270 40982 65284
rect 41858 65270 41940 65284
rect 42148 65270 42230 65284
rect 43106 65270 43188 65284
rect 43396 65270 43478 65284
rect 44354 65270 44436 65284
rect 44644 65270 44726 65284
rect 45602 65270 45684 65284
rect 45892 65270 45974 65284
rect 46850 65270 46932 65284
rect 47140 65270 47222 65284
rect 48098 65270 48180 65284
rect 48388 65270 48470 65284
rect 49346 65270 49428 65284
rect 49636 65270 49718 65284
rect 50594 65270 50676 65284
rect 50884 65270 50966 65284
rect 51842 65270 51924 65284
rect 52132 65270 52214 65284
rect 53090 65270 53172 65284
rect 53380 65270 53462 65284
rect 54338 65270 54420 65284
rect 54628 65270 54710 65284
rect 55586 65270 55668 65284
rect 55876 65270 55958 65284
rect 56834 65270 56916 65284
rect 57124 65270 57206 65284
rect 58082 65270 58164 65284
rect 58372 65270 58454 65284
rect 16418 65222 58934 65270
rect 16418 65126 58934 65174
rect 16898 65112 16980 65126
rect 17188 65112 17270 65126
rect 18146 65112 18228 65126
rect 18436 65112 18518 65126
rect 19394 65112 19476 65126
rect 19684 65112 19766 65126
rect 20642 65112 20724 65126
rect 20932 65112 21014 65126
rect 21890 65112 21972 65126
rect 22180 65112 22262 65126
rect 23138 65112 23220 65126
rect 23428 65112 23510 65126
rect 24386 65112 24468 65126
rect 24676 65112 24758 65126
rect 25634 65112 25716 65126
rect 25924 65112 26006 65126
rect 26882 65112 26964 65126
rect 27172 65112 27254 65126
rect 28130 65112 28212 65126
rect 28420 65112 28502 65126
rect 29378 65112 29460 65126
rect 29668 65112 29750 65126
rect 30626 65112 30708 65126
rect 30916 65112 30998 65126
rect 31874 65112 31956 65126
rect 32164 65112 32246 65126
rect 33122 65112 33204 65126
rect 33412 65112 33494 65126
rect 34370 65112 34452 65126
rect 34660 65112 34742 65126
rect 35618 65112 35700 65126
rect 35908 65112 35990 65126
rect 36866 65112 36948 65126
rect 37156 65112 37238 65126
rect 38114 65112 38196 65126
rect 38404 65112 38486 65126
rect 39362 65112 39444 65126
rect 39652 65112 39734 65126
rect 40610 65112 40692 65126
rect 40900 65112 40982 65126
rect 41858 65112 41940 65126
rect 42148 65112 42230 65126
rect 43106 65112 43188 65126
rect 43396 65112 43478 65126
rect 44354 65112 44436 65126
rect 44644 65112 44726 65126
rect 45602 65112 45684 65126
rect 45892 65112 45974 65126
rect 46850 65112 46932 65126
rect 47140 65112 47222 65126
rect 48098 65112 48180 65126
rect 48388 65112 48470 65126
rect 49346 65112 49428 65126
rect 49636 65112 49718 65126
rect 50594 65112 50676 65126
rect 50884 65112 50966 65126
rect 51842 65112 51924 65126
rect 52132 65112 52214 65126
rect 53090 65112 53172 65126
rect 53380 65112 53462 65126
rect 54338 65112 54420 65126
rect 54628 65112 54710 65126
rect 55586 65112 55668 65126
rect 55876 65112 55958 65126
rect 56834 65112 56916 65126
rect 57124 65112 57206 65126
rect 58082 65112 58164 65126
rect 58372 65112 58454 65126
rect 16418 65064 16864 65078
rect 17014 65064 17154 65078
rect 17304 65064 18112 65078
rect 18262 65064 18402 65078
rect 18552 65064 19360 65078
rect 19510 65064 19650 65078
rect 19800 65064 20608 65078
rect 20758 65064 20898 65078
rect 21048 65064 21856 65078
rect 22006 65064 22146 65078
rect 22296 65064 23104 65078
rect 23254 65064 23394 65078
rect 23544 65064 24352 65078
rect 24502 65064 24642 65078
rect 24792 65064 25600 65078
rect 25750 65064 25890 65078
rect 26040 65064 26848 65078
rect 26998 65064 27138 65078
rect 27288 65064 28096 65078
rect 28246 65064 28386 65078
rect 28536 65064 29344 65078
rect 29494 65064 29634 65078
rect 29784 65064 30592 65078
rect 30742 65064 30882 65078
rect 31032 65064 31840 65078
rect 31990 65064 32130 65078
rect 32280 65064 33088 65078
rect 33238 65064 33378 65078
rect 33528 65064 34336 65078
rect 34486 65064 34626 65078
rect 34776 65064 35584 65078
rect 35734 65064 35874 65078
rect 36024 65064 36832 65078
rect 36982 65064 37122 65078
rect 37272 65064 38080 65078
rect 38230 65064 38370 65078
rect 38520 65064 39328 65078
rect 39478 65064 39618 65078
rect 39768 65064 40576 65078
rect 40726 65064 40866 65078
rect 41016 65064 41824 65078
rect 41974 65064 42114 65078
rect 42264 65064 43072 65078
rect 43222 65064 43362 65078
rect 43512 65064 44320 65078
rect 44470 65064 44610 65078
rect 44760 65064 45568 65078
rect 45718 65064 45858 65078
rect 46008 65064 46816 65078
rect 46966 65064 47106 65078
rect 47256 65064 48064 65078
rect 48214 65064 48354 65078
rect 48504 65064 49312 65078
rect 49462 65064 49602 65078
rect 49752 65064 50560 65078
rect 50710 65064 50850 65078
rect 51000 65064 51808 65078
rect 51958 65064 52098 65078
rect 52248 65064 53056 65078
rect 53206 65064 53346 65078
rect 53496 65064 54304 65078
rect 54454 65064 54594 65078
rect 54744 65064 55552 65078
rect 55702 65064 55842 65078
rect 55992 65064 56800 65078
rect 56950 65064 57090 65078
rect 57240 65064 58048 65078
rect 58198 65064 58338 65078
rect 58488 65064 58934 65078
rect 16418 65016 58934 65064
rect 16418 65002 16864 65016
rect 17014 65002 17154 65016
rect 17304 65002 18112 65016
rect 18262 65002 18402 65016
rect 18552 65002 19360 65016
rect 19510 65002 19650 65016
rect 19800 65002 20608 65016
rect 20758 65002 20898 65016
rect 21048 65002 21856 65016
rect 22006 65002 22146 65016
rect 22296 65002 23104 65016
rect 23254 65002 23394 65016
rect 23544 65002 24352 65016
rect 24502 65002 24642 65016
rect 24792 65002 25600 65016
rect 25750 65002 25890 65016
rect 26040 65002 26848 65016
rect 26998 65002 27138 65016
rect 27288 65002 28096 65016
rect 28246 65002 28386 65016
rect 28536 65002 29344 65016
rect 29494 65002 29634 65016
rect 29784 65002 30592 65016
rect 30742 65002 30882 65016
rect 31032 65002 31840 65016
rect 31990 65002 32130 65016
rect 32280 65002 33088 65016
rect 33238 65002 33378 65016
rect 33528 65002 34336 65016
rect 34486 65002 34626 65016
rect 34776 65002 35584 65016
rect 35734 65002 35874 65016
rect 36024 65002 36832 65016
rect 36982 65002 37122 65016
rect 37272 65002 38080 65016
rect 38230 65002 38370 65016
rect 38520 65002 39328 65016
rect 39478 65002 39618 65016
rect 39768 65002 40576 65016
rect 40726 65002 40866 65016
rect 41016 65002 41824 65016
rect 41974 65002 42114 65016
rect 42264 65002 43072 65016
rect 43222 65002 43362 65016
rect 43512 65002 44320 65016
rect 44470 65002 44610 65016
rect 44760 65002 45568 65016
rect 45718 65002 45858 65016
rect 46008 65002 46816 65016
rect 46966 65002 47106 65016
rect 47256 65002 48064 65016
rect 48214 65002 48354 65016
rect 48504 65002 49312 65016
rect 49462 65002 49602 65016
rect 49752 65002 50560 65016
rect 50710 65002 50850 65016
rect 51000 65002 51808 65016
rect 51958 65002 52098 65016
rect 52248 65002 53056 65016
rect 53206 65002 53346 65016
rect 53496 65002 54304 65016
rect 54454 65002 54594 65016
rect 54744 65002 55552 65016
rect 55702 65002 55842 65016
rect 55992 65002 56800 65016
rect 56950 65002 57090 65016
rect 57240 65002 58048 65016
rect 58198 65002 58338 65016
rect 58488 65002 58934 65016
rect 16898 64954 16980 64968
rect 17188 64954 17270 64968
rect 18146 64954 18228 64968
rect 18436 64954 18518 64968
rect 19394 64954 19476 64968
rect 19684 64954 19766 64968
rect 20642 64954 20724 64968
rect 20932 64954 21014 64968
rect 21890 64954 21972 64968
rect 22180 64954 22262 64968
rect 23138 64954 23220 64968
rect 23428 64954 23510 64968
rect 24386 64954 24468 64968
rect 24676 64954 24758 64968
rect 25634 64954 25716 64968
rect 25924 64954 26006 64968
rect 26882 64954 26964 64968
rect 27172 64954 27254 64968
rect 28130 64954 28212 64968
rect 28420 64954 28502 64968
rect 29378 64954 29460 64968
rect 29668 64954 29750 64968
rect 30626 64954 30708 64968
rect 30916 64954 30998 64968
rect 31874 64954 31956 64968
rect 32164 64954 32246 64968
rect 33122 64954 33204 64968
rect 33412 64954 33494 64968
rect 34370 64954 34452 64968
rect 34660 64954 34742 64968
rect 35618 64954 35700 64968
rect 35908 64954 35990 64968
rect 36866 64954 36948 64968
rect 37156 64954 37238 64968
rect 38114 64954 38196 64968
rect 38404 64954 38486 64968
rect 39362 64954 39444 64968
rect 39652 64954 39734 64968
rect 40610 64954 40692 64968
rect 40900 64954 40982 64968
rect 41858 64954 41940 64968
rect 42148 64954 42230 64968
rect 43106 64954 43188 64968
rect 43396 64954 43478 64968
rect 44354 64954 44436 64968
rect 44644 64954 44726 64968
rect 45602 64954 45684 64968
rect 45892 64954 45974 64968
rect 46850 64954 46932 64968
rect 47140 64954 47222 64968
rect 48098 64954 48180 64968
rect 48388 64954 48470 64968
rect 49346 64954 49428 64968
rect 49636 64954 49718 64968
rect 50594 64954 50676 64968
rect 50884 64954 50966 64968
rect 51842 64954 51924 64968
rect 52132 64954 52214 64968
rect 53090 64954 53172 64968
rect 53380 64954 53462 64968
rect 54338 64954 54420 64968
rect 54628 64954 54710 64968
rect 55586 64954 55668 64968
rect 55876 64954 55958 64968
rect 56834 64954 56916 64968
rect 57124 64954 57206 64968
rect 58082 64954 58164 64968
rect 58372 64954 58454 64968
rect 16418 64906 58934 64954
rect 16418 64748 58934 64858
rect 16418 64652 58934 64700
rect 16898 64638 16980 64652
rect 17188 64638 17270 64652
rect 18146 64638 18228 64652
rect 18436 64638 18518 64652
rect 19394 64638 19476 64652
rect 19684 64638 19766 64652
rect 20642 64638 20724 64652
rect 20932 64638 21014 64652
rect 21890 64638 21972 64652
rect 22180 64638 22262 64652
rect 23138 64638 23220 64652
rect 23428 64638 23510 64652
rect 24386 64638 24468 64652
rect 24676 64638 24758 64652
rect 25634 64638 25716 64652
rect 25924 64638 26006 64652
rect 26882 64638 26964 64652
rect 27172 64638 27254 64652
rect 28130 64638 28212 64652
rect 28420 64638 28502 64652
rect 29378 64638 29460 64652
rect 29668 64638 29750 64652
rect 30626 64638 30708 64652
rect 30916 64638 30998 64652
rect 31874 64638 31956 64652
rect 32164 64638 32246 64652
rect 33122 64638 33204 64652
rect 33412 64638 33494 64652
rect 34370 64638 34452 64652
rect 34660 64638 34742 64652
rect 35618 64638 35700 64652
rect 35908 64638 35990 64652
rect 36866 64638 36948 64652
rect 37156 64638 37238 64652
rect 38114 64638 38196 64652
rect 38404 64638 38486 64652
rect 39362 64638 39444 64652
rect 39652 64638 39734 64652
rect 40610 64638 40692 64652
rect 40900 64638 40982 64652
rect 41858 64638 41940 64652
rect 42148 64638 42230 64652
rect 43106 64638 43188 64652
rect 43396 64638 43478 64652
rect 44354 64638 44436 64652
rect 44644 64638 44726 64652
rect 45602 64638 45684 64652
rect 45892 64638 45974 64652
rect 46850 64638 46932 64652
rect 47140 64638 47222 64652
rect 48098 64638 48180 64652
rect 48388 64638 48470 64652
rect 49346 64638 49428 64652
rect 49636 64638 49718 64652
rect 50594 64638 50676 64652
rect 50884 64638 50966 64652
rect 51842 64638 51924 64652
rect 52132 64638 52214 64652
rect 53090 64638 53172 64652
rect 53380 64638 53462 64652
rect 54338 64638 54420 64652
rect 54628 64638 54710 64652
rect 55586 64638 55668 64652
rect 55876 64638 55958 64652
rect 56834 64638 56916 64652
rect 57124 64638 57206 64652
rect 58082 64638 58164 64652
rect 58372 64638 58454 64652
rect 16418 64590 16864 64604
rect 17014 64590 17154 64604
rect 17304 64590 18112 64604
rect 18262 64590 18402 64604
rect 18552 64590 19360 64604
rect 19510 64590 19650 64604
rect 19800 64590 20608 64604
rect 20758 64590 20898 64604
rect 21048 64590 21856 64604
rect 22006 64590 22146 64604
rect 22296 64590 23104 64604
rect 23254 64590 23394 64604
rect 23544 64590 24352 64604
rect 24502 64590 24642 64604
rect 24792 64590 25600 64604
rect 25750 64590 25890 64604
rect 26040 64590 26848 64604
rect 26998 64590 27138 64604
rect 27288 64590 28096 64604
rect 28246 64590 28386 64604
rect 28536 64590 29344 64604
rect 29494 64590 29634 64604
rect 29784 64590 30592 64604
rect 30742 64590 30882 64604
rect 31032 64590 31840 64604
rect 31990 64590 32130 64604
rect 32280 64590 33088 64604
rect 33238 64590 33378 64604
rect 33528 64590 34336 64604
rect 34486 64590 34626 64604
rect 34776 64590 35584 64604
rect 35734 64590 35874 64604
rect 36024 64590 36832 64604
rect 36982 64590 37122 64604
rect 37272 64590 38080 64604
rect 38230 64590 38370 64604
rect 38520 64590 39328 64604
rect 39478 64590 39618 64604
rect 39768 64590 40576 64604
rect 40726 64590 40866 64604
rect 41016 64590 41824 64604
rect 41974 64590 42114 64604
rect 42264 64590 43072 64604
rect 43222 64590 43362 64604
rect 43512 64590 44320 64604
rect 44470 64590 44610 64604
rect 44760 64590 45568 64604
rect 45718 64590 45858 64604
rect 46008 64590 46816 64604
rect 46966 64590 47106 64604
rect 47256 64590 48064 64604
rect 48214 64590 48354 64604
rect 48504 64590 49312 64604
rect 49462 64590 49602 64604
rect 49752 64590 50560 64604
rect 50710 64590 50850 64604
rect 51000 64590 51808 64604
rect 51958 64590 52098 64604
rect 52248 64590 53056 64604
rect 53206 64590 53346 64604
rect 53496 64590 54304 64604
rect 54454 64590 54594 64604
rect 54744 64590 55552 64604
rect 55702 64590 55842 64604
rect 55992 64590 56800 64604
rect 56950 64590 57090 64604
rect 57240 64590 58048 64604
rect 58198 64590 58338 64604
rect 58488 64590 58934 64604
rect 16418 64542 58934 64590
rect 16418 64528 16864 64542
rect 17014 64528 17154 64542
rect 17304 64528 18112 64542
rect 18262 64528 18402 64542
rect 18552 64528 19360 64542
rect 19510 64528 19650 64542
rect 19800 64528 20608 64542
rect 20758 64528 20898 64542
rect 21048 64528 21856 64542
rect 22006 64528 22146 64542
rect 22296 64528 23104 64542
rect 23254 64528 23394 64542
rect 23544 64528 24352 64542
rect 24502 64528 24642 64542
rect 24792 64528 25600 64542
rect 25750 64528 25890 64542
rect 26040 64528 26848 64542
rect 26998 64528 27138 64542
rect 27288 64528 28096 64542
rect 28246 64528 28386 64542
rect 28536 64528 29344 64542
rect 29494 64528 29634 64542
rect 29784 64528 30592 64542
rect 30742 64528 30882 64542
rect 31032 64528 31840 64542
rect 31990 64528 32130 64542
rect 32280 64528 33088 64542
rect 33238 64528 33378 64542
rect 33528 64528 34336 64542
rect 34486 64528 34626 64542
rect 34776 64528 35584 64542
rect 35734 64528 35874 64542
rect 36024 64528 36832 64542
rect 36982 64528 37122 64542
rect 37272 64528 38080 64542
rect 38230 64528 38370 64542
rect 38520 64528 39328 64542
rect 39478 64528 39618 64542
rect 39768 64528 40576 64542
rect 40726 64528 40866 64542
rect 41016 64528 41824 64542
rect 41974 64528 42114 64542
rect 42264 64528 43072 64542
rect 43222 64528 43362 64542
rect 43512 64528 44320 64542
rect 44470 64528 44610 64542
rect 44760 64528 45568 64542
rect 45718 64528 45858 64542
rect 46008 64528 46816 64542
rect 46966 64528 47106 64542
rect 47256 64528 48064 64542
rect 48214 64528 48354 64542
rect 48504 64528 49312 64542
rect 49462 64528 49602 64542
rect 49752 64528 50560 64542
rect 50710 64528 50850 64542
rect 51000 64528 51808 64542
rect 51958 64528 52098 64542
rect 52248 64528 53056 64542
rect 53206 64528 53346 64542
rect 53496 64528 54304 64542
rect 54454 64528 54594 64542
rect 54744 64528 55552 64542
rect 55702 64528 55842 64542
rect 55992 64528 56800 64542
rect 56950 64528 57090 64542
rect 57240 64528 58048 64542
rect 58198 64528 58338 64542
rect 58488 64528 58934 64542
rect 16898 64480 16980 64494
rect 17188 64480 17270 64494
rect 18146 64480 18228 64494
rect 18436 64480 18518 64494
rect 19394 64480 19476 64494
rect 19684 64480 19766 64494
rect 20642 64480 20724 64494
rect 20932 64480 21014 64494
rect 21890 64480 21972 64494
rect 22180 64480 22262 64494
rect 23138 64480 23220 64494
rect 23428 64480 23510 64494
rect 24386 64480 24468 64494
rect 24676 64480 24758 64494
rect 25634 64480 25716 64494
rect 25924 64480 26006 64494
rect 26882 64480 26964 64494
rect 27172 64480 27254 64494
rect 28130 64480 28212 64494
rect 28420 64480 28502 64494
rect 29378 64480 29460 64494
rect 29668 64480 29750 64494
rect 30626 64480 30708 64494
rect 30916 64480 30998 64494
rect 31874 64480 31956 64494
rect 32164 64480 32246 64494
rect 33122 64480 33204 64494
rect 33412 64480 33494 64494
rect 34370 64480 34452 64494
rect 34660 64480 34742 64494
rect 35618 64480 35700 64494
rect 35908 64480 35990 64494
rect 36866 64480 36948 64494
rect 37156 64480 37238 64494
rect 38114 64480 38196 64494
rect 38404 64480 38486 64494
rect 39362 64480 39444 64494
rect 39652 64480 39734 64494
rect 40610 64480 40692 64494
rect 40900 64480 40982 64494
rect 41858 64480 41940 64494
rect 42148 64480 42230 64494
rect 43106 64480 43188 64494
rect 43396 64480 43478 64494
rect 44354 64480 44436 64494
rect 44644 64480 44726 64494
rect 45602 64480 45684 64494
rect 45892 64480 45974 64494
rect 46850 64480 46932 64494
rect 47140 64480 47222 64494
rect 48098 64480 48180 64494
rect 48388 64480 48470 64494
rect 49346 64480 49428 64494
rect 49636 64480 49718 64494
rect 50594 64480 50676 64494
rect 50884 64480 50966 64494
rect 51842 64480 51924 64494
rect 52132 64480 52214 64494
rect 53090 64480 53172 64494
rect 53380 64480 53462 64494
rect 54338 64480 54420 64494
rect 54628 64480 54710 64494
rect 55586 64480 55668 64494
rect 55876 64480 55958 64494
rect 56834 64480 56916 64494
rect 57124 64480 57206 64494
rect 58082 64480 58164 64494
rect 58372 64480 58454 64494
rect 16418 64432 58934 64480
rect 16418 64336 58934 64384
rect 16898 64322 16980 64336
rect 17188 64322 17270 64336
rect 18146 64322 18228 64336
rect 18436 64322 18518 64336
rect 19394 64322 19476 64336
rect 19684 64322 19766 64336
rect 20642 64322 20724 64336
rect 20932 64322 21014 64336
rect 21890 64322 21972 64336
rect 22180 64322 22262 64336
rect 23138 64322 23220 64336
rect 23428 64322 23510 64336
rect 24386 64322 24468 64336
rect 24676 64322 24758 64336
rect 25634 64322 25716 64336
rect 25924 64322 26006 64336
rect 26882 64322 26964 64336
rect 27172 64322 27254 64336
rect 28130 64322 28212 64336
rect 28420 64322 28502 64336
rect 29378 64322 29460 64336
rect 29668 64322 29750 64336
rect 30626 64322 30708 64336
rect 30916 64322 30998 64336
rect 31874 64322 31956 64336
rect 32164 64322 32246 64336
rect 33122 64322 33204 64336
rect 33412 64322 33494 64336
rect 34370 64322 34452 64336
rect 34660 64322 34742 64336
rect 35618 64322 35700 64336
rect 35908 64322 35990 64336
rect 36866 64322 36948 64336
rect 37156 64322 37238 64336
rect 38114 64322 38196 64336
rect 38404 64322 38486 64336
rect 39362 64322 39444 64336
rect 39652 64322 39734 64336
rect 40610 64322 40692 64336
rect 40900 64322 40982 64336
rect 41858 64322 41940 64336
rect 42148 64322 42230 64336
rect 43106 64322 43188 64336
rect 43396 64322 43478 64336
rect 44354 64322 44436 64336
rect 44644 64322 44726 64336
rect 45602 64322 45684 64336
rect 45892 64322 45974 64336
rect 46850 64322 46932 64336
rect 47140 64322 47222 64336
rect 48098 64322 48180 64336
rect 48388 64322 48470 64336
rect 49346 64322 49428 64336
rect 49636 64322 49718 64336
rect 50594 64322 50676 64336
rect 50884 64322 50966 64336
rect 51842 64322 51924 64336
rect 52132 64322 52214 64336
rect 53090 64322 53172 64336
rect 53380 64322 53462 64336
rect 54338 64322 54420 64336
rect 54628 64322 54710 64336
rect 55586 64322 55668 64336
rect 55876 64322 55958 64336
rect 56834 64322 56916 64336
rect 57124 64322 57206 64336
rect 58082 64322 58164 64336
rect 58372 64322 58454 64336
rect 16418 64274 16864 64288
rect 17014 64274 17154 64288
rect 17304 64274 18112 64288
rect 18262 64274 18402 64288
rect 18552 64274 19360 64288
rect 19510 64274 19650 64288
rect 19800 64274 20608 64288
rect 20758 64274 20898 64288
rect 21048 64274 21856 64288
rect 22006 64274 22146 64288
rect 22296 64274 23104 64288
rect 23254 64274 23394 64288
rect 23544 64274 24352 64288
rect 24502 64274 24642 64288
rect 24792 64274 25600 64288
rect 25750 64274 25890 64288
rect 26040 64274 26848 64288
rect 26998 64274 27138 64288
rect 27288 64274 28096 64288
rect 28246 64274 28386 64288
rect 28536 64274 29344 64288
rect 29494 64274 29634 64288
rect 29784 64274 30592 64288
rect 30742 64274 30882 64288
rect 31032 64274 31840 64288
rect 31990 64274 32130 64288
rect 32280 64274 33088 64288
rect 33238 64274 33378 64288
rect 33528 64274 34336 64288
rect 34486 64274 34626 64288
rect 34776 64274 35584 64288
rect 35734 64274 35874 64288
rect 36024 64274 36832 64288
rect 36982 64274 37122 64288
rect 37272 64274 38080 64288
rect 38230 64274 38370 64288
rect 38520 64274 39328 64288
rect 39478 64274 39618 64288
rect 39768 64274 40576 64288
rect 40726 64274 40866 64288
rect 41016 64274 41824 64288
rect 41974 64274 42114 64288
rect 42264 64274 43072 64288
rect 43222 64274 43362 64288
rect 43512 64274 44320 64288
rect 44470 64274 44610 64288
rect 44760 64274 45568 64288
rect 45718 64274 45858 64288
rect 46008 64274 46816 64288
rect 46966 64274 47106 64288
rect 47256 64274 48064 64288
rect 48214 64274 48354 64288
rect 48504 64274 49312 64288
rect 49462 64274 49602 64288
rect 49752 64274 50560 64288
rect 50710 64274 50850 64288
rect 51000 64274 51808 64288
rect 51958 64274 52098 64288
rect 52248 64274 53056 64288
rect 53206 64274 53346 64288
rect 53496 64274 54304 64288
rect 54454 64274 54594 64288
rect 54744 64274 55552 64288
rect 55702 64274 55842 64288
rect 55992 64274 56800 64288
rect 56950 64274 57090 64288
rect 57240 64274 58048 64288
rect 58198 64274 58338 64288
rect 58488 64274 58934 64288
rect 16418 64226 58934 64274
rect 16418 64212 16864 64226
rect 17014 64212 17154 64226
rect 17304 64212 18112 64226
rect 18262 64212 18402 64226
rect 18552 64212 19360 64226
rect 19510 64212 19650 64226
rect 19800 64212 20608 64226
rect 20758 64212 20898 64226
rect 21048 64212 21856 64226
rect 22006 64212 22146 64226
rect 22296 64212 23104 64226
rect 23254 64212 23394 64226
rect 23544 64212 24352 64226
rect 24502 64212 24642 64226
rect 24792 64212 25600 64226
rect 25750 64212 25890 64226
rect 26040 64212 26848 64226
rect 26998 64212 27138 64226
rect 27288 64212 28096 64226
rect 28246 64212 28386 64226
rect 28536 64212 29344 64226
rect 29494 64212 29634 64226
rect 29784 64212 30592 64226
rect 30742 64212 30882 64226
rect 31032 64212 31840 64226
rect 31990 64212 32130 64226
rect 32280 64212 33088 64226
rect 33238 64212 33378 64226
rect 33528 64212 34336 64226
rect 34486 64212 34626 64226
rect 34776 64212 35584 64226
rect 35734 64212 35874 64226
rect 36024 64212 36832 64226
rect 36982 64212 37122 64226
rect 37272 64212 38080 64226
rect 38230 64212 38370 64226
rect 38520 64212 39328 64226
rect 39478 64212 39618 64226
rect 39768 64212 40576 64226
rect 40726 64212 40866 64226
rect 41016 64212 41824 64226
rect 41974 64212 42114 64226
rect 42264 64212 43072 64226
rect 43222 64212 43362 64226
rect 43512 64212 44320 64226
rect 44470 64212 44610 64226
rect 44760 64212 45568 64226
rect 45718 64212 45858 64226
rect 46008 64212 46816 64226
rect 46966 64212 47106 64226
rect 47256 64212 48064 64226
rect 48214 64212 48354 64226
rect 48504 64212 49312 64226
rect 49462 64212 49602 64226
rect 49752 64212 50560 64226
rect 50710 64212 50850 64226
rect 51000 64212 51808 64226
rect 51958 64212 52098 64226
rect 52248 64212 53056 64226
rect 53206 64212 53346 64226
rect 53496 64212 54304 64226
rect 54454 64212 54594 64226
rect 54744 64212 55552 64226
rect 55702 64212 55842 64226
rect 55992 64212 56800 64226
rect 56950 64212 57090 64226
rect 57240 64212 58048 64226
rect 58198 64212 58338 64226
rect 58488 64212 58934 64226
rect 16898 64164 16980 64178
rect 17188 64164 17270 64178
rect 18146 64164 18228 64178
rect 18436 64164 18518 64178
rect 19394 64164 19476 64178
rect 19684 64164 19766 64178
rect 20642 64164 20724 64178
rect 20932 64164 21014 64178
rect 21890 64164 21972 64178
rect 22180 64164 22262 64178
rect 23138 64164 23220 64178
rect 23428 64164 23510 64178
rect 24386 64164 24468 64178
rect 24676 64164 24758 64178
rect 25634 64164 25716 64178
rect 25924 64164 26006 64178
rect 26882 64164 26964 64178
rect 27172 64164 27254 64178
rect 28130 64164 28212 64178
rect 28420 64164 28502 64178
rect 29378 64164 29460 64178
rect 29668 64164 29750 64178
rect 30626 64164 30708 64178
rect 30916 64164 30998 64178
rect 31874 64164 31956 64178
rect 32164 64164 32246 64178
rect 33122 64164 33204 64178
rect 33412 64164 33494 64178
rect 34370 64164 34452 64178
rect 34660 64164 34742 64178
rect 35618 64164 35700 64178
rect 35908 64164 35990 64178
rect 36866 64164 36948 64178
rect 37156 64164 37238 64178
rect 38114 64164 38196 64178
rect 38404 64164 38486 64178
rect 39362 64164 39444 64178
rect 39652 64164 39734 64178
rect 40610 64164 40692 64178
rect 40900 64164 40982 64178
rect 41858 64164 41940 64178
rect 42148 64164 42230 64178
rect 43106 64164 43188 64178
rect 43396 64164 43478 64178
rect 44354 64164 44436 64178
rect 44644 64164 44726 64178
rect 45602 64164 45684 64178
rect 45892 64164 45974 64178
rect 46850 64164 46932 64178
rect 47140 64164 47222 64178
rect 48098 64164 48180 64178
rect 48388 64164 48470 64178
rect 49346 64164 49428 64178
rect 49636 64164 49718 64178
rect 50594 64164 50676 64178
rect 50884 64164 50966 64178
rect 51842 64164 51924 64178
rect 52132 64164 52214 64178
rect 53090 64164 53172 64178
rect 53380 64164 53462 64178
rect 54338 64164 54420 64178
rect 54628 64164 54710 64178
rect 55586 64164 55668 64178
rect 55876 64164 55958 64178
rect 56834 64164 56916 64178
rect 57124 64164 57206 64178
rect 58082 64164 58164 64178
rect 58372 64164 58454 64178
rect 16418 64116 58934 64164
rect 16418 63958 58934 64068
rect 16418 63862 58934 63910
rect 16898 63848 16980 63862
rect 17188 63848 17270 63862
rect 18146 63848 18228 63862
rect 18436 63848 18518 63862
rect 19394 63848 19476 63862
rect 19684 63848 19766 63862
rect 20642 63848 20724 63862
rect 20932 63848 21014 63862
rect 21890 63848 21972 63862
rect 22180 63848 22262 63862
rect 23138 63848 23220 63862
rect 23428 63848 23510 63862
rect 24386 63848 24468 63862
rect 24676 63848 24758 63862
rect 25634 63848 25716 63862
rect 25924 63848 26006 63862
rect 26882 63848 26964 63862
rect 27172 63848 27254 63862
rect 28130 63848 28212 63862
rect 28420 63848 28502 63862
rect 29378 63848 29460 63862
rect 29668 63848 29750 63862
rect 30626 63848 30708 63862
rect 30916 63848 30998 63862
rect 31874 63848 31956 63862
rect 32164 63848 32246 63862
rect 33122 63848 33204 63862
rect 33412 63848 33494 63862
rect 34370 63848 34452 63862
rect 34660 63848 34742 63862
rect 35618 63848 35700 63862
rect 35908 63848 35990 63862
rect 36866 63848 36948 63862
rect 37156 63848 37238 63862
rect 38114 63848 38196 63862
rect 38404 63848 38486 63862
rect 39362 63848 39444 63862
rect 39652 63848 39734 63862
rect 40610 63848 40692 63862
rect 40900 63848 40982 63862
rect 41858 63848 41940 63862
rect 42148 63848 42230 63862
rect 43106 63848 43188 63862
rect 43396 63848 43478 63862
rect 44354 63848 44436 63862
rect 44644 63848 44726 63862
rect 45602 63848 45684 63862
rect 45892 63848 45974 63862
rect 46850 63848 46932 63862
rect 47140 63848 47222 63862
rect 48098 63848 48180 63862
rect 48388 63848 48470 63862
rect 49346 63848 49428 63862
rect 49636 63848 49718 63862
rect 50594 63848 50676 63862
rect 50884 63848 50966 63862
rect 51842 63848 51924 63862
rect 52132 63848 52214 63862
rect 53090 63848 53172 63862
rect 53380 63848 53462 63862
rect 54338 63848 54420 63862
rect 54628 63848 54710 63862
rect 55586 63848 55668 63862
rect 55876 63848 55958 63862
rect 56834 63848 56916 63862
rect 57124 63848 57206 63862
rect 58082 63848 58164 63862
rect 58372 63848 58454 63862
rect 16418 63800 16864 63814
rect 17014 63800 17154 63814
rect 17304 63800 18112 63814
rect 18262 63800 18402 63814
rect 18552 63800 19360 63814
rect 19510 63800 19650 63814
rect 19800 63800 20608 63814
rect 20758 63800 20898 63814
rect 21048 63800 21856 63814
rect 22006 63800 22146 63814
rect 22296 63800 23104 63814
rect 23254 63800 23394 63814
rect 23544 63800 24352 63814
rect 24502 63800 24642 63814
rect 24792 63800 25600 63814
rect 25750 63800 25890 63814
rect 26040 63800 26848 63814
rect 26998 63800 27138 63814
rect 27288 63800 28096 63814
rect 28246 63800 28386 63814
rect 28536 63800 29344 63814
rect 29494 63800 29634 63814
rect 29784 63800 30592 63814
rect 30742 63800 30882 63814
rect 31032 63800 31840 63814
rect 31990 63800 32130 63814
rect 32280 63800 33088 63814
rect 33238 63800 33378 63814
rect 33528 63800 34336 63814
rect 34486 63800 34626 63814
rect 34776 63800 35584 63814
rect 35734 63800 35874 63814
rect 36024 63800 36832 63814
rect 36982 63800 37122 63814
rect 37272 63800 38080 63814
rect 38230 63800 38370 63814
rect 38520 63800 39328 63814
rect 39478 63800 39618 63814
rect 39768 63800 40576 63814
rect 40726 63800 40866 63814
rect 41016 63800 41824 63814
rect 41974 63800 42114 63814
rect 42264 63800 43072 63814
rect 43222 63800 43362 63814
rect 43512 63800 44320 63814
rect 44470 63800 44610 63814
rect 44760 63800 45568 63814
rect 45718 63800 45858 63814
rect 46008 63800 46816 63814
rect 46966 63800 47106 63814
rect 47256 63800 48064 63814
rect 48214 63800 48354 63814
rect 48504 63800 49312 63814
rect 49462 63800 49602 63814
rect 49752 63800 50560 63814
rect 50710 63800 50850 63814
rect 51000 63800 51808 63814
rect 51958 63800 52098 63814
rect 52248 63800 53056 63814
rect 53206 63800 53346 63814
rect 53496 63800 54304 63814
rect 54454 63800 54594 63814
rect 54744 63800 55552 63814
rect 55702 63800 55842 63814
rect 55992 63800 56800 63814
rect 56950 63800 57090 63814
rect 57240 63800 58048 63814
rect 58198 63800 58338 63814
rect 58488 63800 58934 63814
rect 16418 63752 58934 63800
rect 16418 63738 16864 63752
rect 17014 63738 17154 63752
rect 17304 63738 18112 63752
rect 18262 63738 18402 63752
rect 18552 63738 19360 63752
rect 19510 63738 19650 63752
rect 19800 63738 20608 63752
rect 20758 63738 20898 63752
rect 21048 63738 21856 63752
rect 22006 63738 22146 63752
rect 22296 63738 23104 63752
rect 23254 63738 23394 63752
rect 23544 63738 24352 63752
rect 24502 63738 24642 63752
rect 24792 63738 25600 63752
rect 25750 63738 25890 63752
rect 26040 63738 26848 63752
rect 26998 63738 27138 63752
rect 27288 63738 28096 63752
rect 28246 63738 28386 63752
rect 28536 63738 29344 63752
rect 29494 63738 29634 63752
rect 29784 63738 30592 63752
rect 30742 63738 30882 63752
rect 31032 63738 31840 63752
rect 31990 63738 32130 63752
rect 32280 63738 33088 63752
rect 33238 63738 33378 63752
rect 33528 63738 34336 63752
rect 34486 63738 34626 63752
rect 34776 63738 35584 63752
rect 35734 63738 35874 63752
rect 36024 63738 36832 63752
rect 36982 63738 37122 63752
rect 37272 63738 38080 63752
rect 38230 63738 38370 63752
rect 38520 63738 39328 63752
rect 39478 63738 39618 63752
rect 39768 63738 40576 63752
rect 40726 63738 40866 63752
rect 41016 63738 41824 63752
rect 41974 63738 42114 63752
rect 42264 63738 43072 63752
rect 43222 63738 43362 63752
rect 43512 63738 44320 63752
rect 44470 63738 44610 63752
rect 44760 63738 45568 63752
rect 45718 63738 45858 63752
rect 46008 63738 46816 63752
rect 46966 63738 47106 63752
rect 47256 63738 48064 63752
rect 48214 63738 48354 63752
rect 48504 63738 49312 63752
rect 49462 63738 49602 63752
rect 49752 63738 50560 63752
rect 50710 63738 50850 63752
rect 51000 63738 51808 63752
rect 51958 63738 52098 63752
rect 52248 63738 53056 63752
rect 53206 63738 53346 63752
rect 53496 63738 54304 63752
rect 54454 63738 54594 63752
rect 54744 63738 55552 63752
rect 55702 63738 55842 63752
rect 55992 63738 56800 63752
rect 56950 63738 57090 63752
rect 57240 63738 58048 63752
rect 58198 63738 58338 63752
rect 58488 63738 58934 63752
rect 16898 63690 16980 63704
rect 17188 63690 17270 63704
rect 18146 63690 18228 63704
rect 18436 63690 18518 63704
rect 19394 63690 19476 63704
rect 19684 63690 19766 63704
rect 20642 63690 20724 63704
rect 20932 63690 21014 63704
rect 21890 63690 21972 63704
rect 22180 63690 22262 63704
rect 23138 63690 23220 63704
rect 23428 63690 23510 63704
rect 24386 63690 24468 63704
rect 24676 63690 24758 63704
rect 25634 63690 25716 63704
rect 25924 63690 26006 63704
rect 26882 63690 26964 63704
rect 27172 63690 27254 63704
rect 28130 63690 28212 63704
rect 28420 63690 28502 63704
rect 29378 63690 29460 63704
rect 29668 63690 29750 63704
rect 30626 63690 30708 63704
rect 30916 63690 30998 63704
rect 31874 63690 31956 63704
rect 32164 63690 32246 63704
rect 33122 63690 33204 63704
rect 33412 63690 33494 63704
rect 34370 63690 34452 63704
rect 34660 63690 34742 63704
rect 35618 63690 35700 63704
rect 35908 63690 35990 63704
rect 36866 63690 36948 63704
rect 37156 63690 37238 63704
rect 38114 63690 38196 63704
rect 38404 63690 38486 63704
rect 39362 63690 39444 63704
rect 39652 63690 39734 63704
rect 40610 63690 40692 63704
rect 40900 63690 40982 63704
rect 41858 63690 41940 63704
rect 42148 63690 42230 63704
rect 43106 63690 43188 63704
rect 43396 63690 43478 63704
rect 44354 63690 44436 63704
rect 44644 63690 44726 63704
rect 45602 63690 45684 63704
rect 45892 63690 45974 63704
rect 46850 63690 46932 63704
rect 47140 63690 47222 63704
rect 48098 63690 48180 63704
rect 48388 63690 48470 63704
rect 49346 63690 49428 63704
rect 49636 63690 49718 63704
rect 50594 63690 50676 63704
rect 50884 63690 50966 63704
rect 51842 63690 51924 63704
rect 52132 63690 52214 63704
rect 53090 63690 53172 63704
rect 53380 63690 53462 63704
rect 54338 63690 54420 63704
rect 54628 63690 54710 63704
rect 55586 63690 55668 63704
rect 55876 63690 55958 63704
rect 56834 63690 56916 63704
rect 57124 63690 57206 63704
rect 58082 63690 58164 63704
rect 58372 63690 58454 63704
rect 16418 63642 58934 63690
rect 16418 63546 58934 63594
rect 16898 63532 16980 63546
rect 17188 63532 17270 63546
rect 18146 63532 18228 63546
rect 18436 63532 18518 63546
rect 19394 63532 19476 63546
rect 19684 63532 19766 63546
rect 20642 63532 20724 63546
rect 20932 63532 21014 63546
rect 21890 63532 21972 63546
rect 22180 63532 22262 63546
rect 23138 63532 23220 63546
rect 23428 63532 23510 63546
rect 24386 63532 24468 63546
rect 24676 63532 24758 63546
rect 25634 63532 25716 63546
rect 25924 63532 26006 63546
rect 26882 63532 26964 63546
rect 27172 63532 27254 63546
rect 28130 63532 28212 63546
rect 28420 63532 28502 63546
rect 29378 63532 29460 63546
rect 29668 63532 29750 63546
rect 30626 63532 30708 63546
rect 30916 63532 30998 63546
rect 31874 63532 31956 63546
rect 32164 63532 32246 63546
rect 33122 63532 33204 63546
rect 33412 63532 33494 63546
rect 34370 63532 34452 63546
rect 34660 63532 34742 63546
rect 35618 63532 35700 63546
rect 35908 63532 35990 63546
rect 36866 63532 36948 63546
rect 37156 63532 37238 63546
rect 38114 63532 38196 63546
rect 38404 63532 38486 63546
rect 39362 63532 39444 63546
rect 39652 63532 39734 63546
rect 40610 63532 40692 63546
rect 40900 63532 40982 63546
rect 41858 63532 41940 63546
rect 42148 63532 42230 63546
rect 43106 63532 43188 63546
rect 43396 63532 43478 63546
rect 44354 63532 44436 63546
rect 44644 63532 44726 63546
rect 45602 63532 45684 63546
rect 45892 63532 45974 63546
rect 46850 63532 46932 63546
rect 47140 63532 47222 63546
rect 48098 63532 48180 63546
rect 48388 63532 48470 63546
rect 49346 63532 49428 63546
rect 49636 63532 49718 63546
rect 50594 63532 50676 63546
rect 50884 63532 50966 63546
rect 51842 63532 51924 63546
rect 52132 63532 52214 63546
rect 53090 63532 53172 63546
rect 53380 63532 53462 63546
rect 54338 63532 54420 63546
rect 54628 63532 54710 63546
rect 55586 63532 55668 63546
rect 55876 63532 55958 63546
rect 56834 63532 56916 63546
rect 57124 63532 57206 63546
rect 58082 63532 58164 63546
rect 58372 63532 58454 63546
rect 16418 63484 16864 63498
rect 17014 63484 17154 63498
rect 17304 63484 18112 63498
rect 18262 63484 18402 63498
rect 18552 63484 19360 63498
rect 19510 63484 19650 63498
rect 19800 63484 20608 63498
rect 20758 63484 20898 63498
rect 21048 63484 21856 63498
rect 22006 63484 22146 63498
rect 22296 63484 23104 63498
rect 23254 63484 23394 63498
rect 23544 63484 24352 63498
rect 24502 63484 24642 63498
rect 24792 63484 25600 63498
rect 25750 63484 25890 63498
rect 26040 63484 26848 63498
rect 26998 63484 27138 63498
rect 27288 63484 28096 63498
rect 28246 63484 28386 63498
rect 28536 63484 29344 63498
rect 29494 63484 29634 63498
rect 29784 63484 30592 63498
rect 30742 63484 30882 63498
rect 31032 63484 31840 63498
rect 31990 63484 32130 63498
rect 32280 63484 33088 63498
rect 33238 63484 33378 63498
rect 33528 63484 34336 63498
rect 34486 63484 34626 63498
rect 34776 63484 35584 63498
rect 35734 63484 35874 63498
rect 36024 63484 36832 63498
rect 36982 63484 37122 63498
rect 37272 63484 38080 63498
rect 38230 63484 38370 63498
rect 38520 63484 39328 63498
rect 39478 63484 39618 63498
rect 39768 63484 40576 63498
rect 40726 63484 40866 63498
rect 41016 63484 41824 63498
rect 41974 63484 42114 63498
rect 42264 63484 43072 63498
rect 43222 63484 43362 63498
rect 43512 63484 44320 63498
rect 44470 63484 44610 63498
rect 44760 63484 45568 63498
rect 45718 63484 45858 63498
rect 46008 63484 46816 63498
rect 46966 63484 47106 63498
rect 47256 63484 48064 63498
rect 48214 63484 48354 63498
rect 48504 63484 49312 63498
rect 49462 63484 49602 63498
rect 49752 63484 50560 63498
rect 50710 63484 50850 63498
rect 51000 63484 51808 63498
rect 51958 63484 52098 63498
rect 52248 63484 53056 63498
rect 53206 63484 53346 63498
rect 53496 63484 54304 63498
rect 54454 63484 54594 63498
rect 54744 63484 55552 63498
rect 55702 63484 55842 63498
rect 55992 63484 56800 63498
rect 56950 63484 57090 63498
rect 57240 63484 58048 63498
rect 58198 63484 58338 63498
rect 58488 63484 58934 63498
rect 16418 63436 58934 63484
rect 16418 63422 16864 63436
rect 17014 63422 17154 63436
rect 17304 63422 18112 63436
rect 18262 63422 18402 63436
rect 18552 63422 19360 63436
rect 19510 63422 19650 63436
rect 19800 63422 20608 63436
rect 20758 63422 20898 63436
rect 21048 63422 21856 63436
rect 22006 63422 22146 63436
rect 22296 63422 23104 63436
rect 23254 63422 23394 63436
rect 23544 63422 24352 63436
rect 24502 63422 24642 63436
rect 24792 63422 25600 63436
rect 25750 63422 25890 63436
rect 26040 63422 26848 63436
rect 26998 63422 27138 63436
rect 27288 63422 28096 63436
rect 28246 63422 28386 63436
rect 28536 63422 29344 63436
rect 29494 63422 29634 63436
rect 29784 63422 30592 63436
rect 30742 63422 30882 63436
rect 31032 63422 31840 63436
rect 31990 63422 32130 63436
rect 32280 63422 33088 63436
rect 33238 63422 33378 63436
rect 33528 63422 34336 63436
rect 34486 63422 34626 63436
rect 34776 63422 35584 63436
rect 35734 63422 35874 63436
rect 36024 63422 36832 63436
rect 36982 63422 37122 63436
rect 37272 63422 38080 63436
rect 38230 63422 38370 63436
rect 38520 63422 39328 63436
rect 39478 63422 39618 63436
rect 39768 63422 40576 63436
rect 40726 63422 40866 63436
rect 41016 63422 41824 63436
rect 41974 63422 42114 63436
rect 42264 63422 43072 63436
rect 43222 63422 43362 63436
rect 43512 63422 44320 63436
rect 44470 63422 44610 63436
rect 44760 63422 45568 63436
rect 45718 63422 45858 63436
rect 46008 63422 46816 63436
rect 46966 63422 47106 63436
rect 47256 63422 48064 63436
rect 48214 63422 48354 63436
rect 48504 63422 49312 63436
rect 49462 63422 49602 63436
rect 49752 63422 50560 63436
rect 50710 63422 50850 63436
rect 51000 63422 51808 63436
rect 51958 63422 52098 63436
rect 52248 63422 53056 63436
rect 53206 63422 53346 63436
rect 53496 63422 54304 63436
rect 54454 63422 54594 63436
rect 54744 63422 55552 63436
rect 55702 63422 55842 63436
rect 55992 63422 56800 63436
rect 56950 63422 57090 63436
rect 57240 63422 58048 63436
rect 58198 63422 58338 63436
rect 58488 63422 58934 63436
rect 16898 63374 16980 63388
rect 17188 63374 17270 63388
rect 18146 63374 18228 63388
rect 18436 63374 18518 63388
rect 19394 63374 19476 63388
rect 19684 63374 19766 63388
rect 20642 63374 20724 63388
rect 20932 63374 21014 63388
rect 21890 63374 21972 63388
rect 22180 63374 22262 63388
rect 23138 63374 23220 63388
rect 23428 63374 23510 63388
rect 24386 63374 24468 63388
rect 24676 63374 24758 63388
rect 25634 63374 25716 63388
rect 25924 63374 26006 63388
rect 26882 63374 26964 63388
rect 27172 63374 27254 63388
rect 28130 63374 28212 63388
rect 28420 63374 28502 63388
rect 29378 63374 29460 63388
rect 29668 63374 29750 63388
rect 30626 63374 30708 63388
rect 30916 63374 30998 63388
rect 31874 63374 31956 63388
rect 32164 63374 32246 63388
rect 33122 63374 33204 63388
rect 33412 63374 33494 63388
rect 34370 63374 34452 63388
rect 34660 63374 34742 63388
rect 35618 63374 35700 63388
rect 35908 63374 35990 63388
rect 36866 63374 36948 63388
rect 37156 63374 37238 63388
rect 38114 63374 38196 63388
rect 38404 63374 38486 63388
rect 39362 63374 39444 63388
rect 39652 63374 39734 63388
rect 40610 63374 40692 63388
rect 40900 63374 40982 63388
rect 41858 63374 41940 63388
rect 42148 63374 42230 63388
rect 43106 63374 43188 63388
rect 43396 63374 43478 63388
rect 44354 63374 44436 63388
rect 44644 63374 44726 63388
rect 45602 63374 45684 63388
rect 45892 63374 45974 63388
rect 46850 63374 46932 63388
rect 47140 63374 47222 63388
rect 48098 63374 48180 63388
rect 48388 63374 48470 63388
rect 49346 63374 49428 63388
rect 49636 63374 49718 63388
rect 50594 63374 50676 63388
rect 50884 63374 50966 63388
rect 51842 63374 51924 63388
rect 52132 63374 52214 63388
rect 53090 63374 53172 63388
rect 53380 63374 53462 63388
rect 54338 63374 54420 63388
rect 54628 63374 54710 63388
rect 55586 63374 55668 63388
rect 55876 63374 55958 63388
rect 56834 63374 56916 63388
rect 57124 63374 57206 63388
rect 58082 63374 58164 63388
rect 58372 63374 58454 63388
rect 16418 63326 58934 63374
rect 16418 63168 58934 63278
rect 16418 63072 58934 63120
rect 16898 63058 16980 63072
rect 17188 63058 17270 63072
rect 18146 63058 18228 63072
rect 18436 63058 18518 63072
rect 19394 63058 19476 63072
rect 19684 63058 19766 63072
rect 20642 63058 20724 63072
rect 20932 63058 21014 63072
rect 21890 63058 21972 63072
rect 22180 63058 22262 63072
rect 23138 63058 23220 63072
rect 23428 63058 23510 63072
rect 24386 63058 24468 63072
rect 24676 63058 24758 63072
rect 25634 63058 25716 63072
rect 25924 63058 26006 63072
rect 26882 63058 26964 63072
rect 27172 63058 27254 63072
rect 28130 63058 28212 63072
rect 28420 63058 28502 63072
rect 29378 63058 29460 63072
rect 29668 63058 29750 63072
rect 30626 63058 30708 63072
rect 30916 63058 30998 63072
rect 31874 63058 31956 63072
rect 32164 63058 32246 63072
rect 33122 63058 33204 63072
rect 33412 63058 33494 63072
rect 34370 63058 34452 63072
rect 34660 63058 34742 63072
rect 35618 63058 35700 63072
rect 35908 63058 35990 63072
rect 36866 63058 36948 63072
rect 37156 63058 37238 63072
rect 38114 63058 38196 63072
rect 38404 63058 38486 63072
rect 39362 63058 39444 63072
rect 39652 63058 39734 63072
rect 40610 63058 40692 63072
rect 40900 63058 40982 63072
rect 41858 63058 41940 63072
rect 42148 63058 42230 63072
rect 43106 63058 43188 63072
rect 43396 63058 43478 63072
rect 44354 63058 44436 63072
rect 44644 63058 44726 63072
rect 45602 63058 45684 63072
rect 45892 63058 45974 63072
rect 46850 63058 46932 63072
rect 47140 63058 47222 63072
rect 48098 63058 48180 63072
rect 48388 63058 48470 63072
rect 49346 63058 49428 63072
rect 49636 63058 49718 63072
rect 50594 63058 50676 63072
rect 50884 63058 50966 63072
rect 51842 63058 51924 63072
rect 52132 63058 52214 63072
rect 53090 63058 53172 63072
rect 53380 63058 53462 63072
rect 54338 63058 54420 63072
rect 54628 63058 54710 63072
rect 55586 63058 55668 63072
rect 55876 63058 55958 63072
rect 56834 63058 56916 63072
rect 57124 63058 57206 63072
rect 58082 63058 58164 63072
rect 58372 63058 58454 63072
rect 16418 63010 16864 63024
rect 17014 63010 17154 63024
rect 17304 63010 18112 63024
rect 18262 63010 18402 63024
rect 18552 63010 19360 63024
rect 19510 63010 19650 63024
rect 19800 63010 20608 63024
rect 20758 63010 20898 63024
rect 21048 63010 21856 63024
rect 22006 63010 22146 63024
rect 22296 63010 23104 63024
rect 23254 63010 23394 63024
rect 23544 63010 24352 63024
rect 24502 63010 24642 63024
rect 24792 63010 25600 63024
rect 25750 63010 25890 63024
rect 26040 63010 26848 63024
rect 26998 63010 27138 63024
rect 27288 63010 28096 63024
rect 28246 63010 28386 63024
rect 28536 63010 29344 63024
rect 29494 63010 29634 63024
rect 29784 63010 30592 63024
rect 30742 63010 30882 63024
rect 31032 63010 31840 63024
rect 31990 63010 32130 63024
rect 32280 63010 33088 63024
rect 33238 63010 33378 63024
rect 33528 63010 34336 63024
rect 34486 63010 34626 63024
rect 34776 63010 35584 63024
rect 35734 63010 35874 63024
rect 36024 63010 36832 63024
rect 36982 63010 37122 63024
rect 37272 63010 38080 63024
rect 38230 63010 38370 63024
rect 38520 63010 39328 63024
rect 39478 63010 39618 63024
rect 39768 63010 40576 63024
rect 40726 63010 40866 63024
rect 41016 63010 41824 63024
rect 41974 63010 42114 63024
rect 42264 63010 43072 63024
rect 43222 63010 43362 63024
rect 43512 63010 44320 63024
rect 44470 63010 44610 63024
rect 44760 63010 45568 63024
rect 45718 63010 45858 63024
rect 46008 63010 46816 63024
rect 46966 63010 47106 63024
rect 47256 63010 48064 63024
rect 48214 63010 48354 63024
rect 48504 63010 49312 63024
rect 49462 63010 49602 63024
rect 49752 63010 50560 63024
rect 50710 63010 50850 63024
rect 51000 63010 51808 63024
rect 51958 63010 52098 63024
rect 52248 63010 53056 63024
rect 53206 63010 53346 63024
rect 53496 63010 54304 63024
rect 54454 63010 54594 63024
rect 54744 63010 55552 63024
rect 55702 63010 55842 63024
rect 55992 63010 56800 63024
rect 56950 63010 57090 63024
rect 57240 63010 58048 63024
rect 58198 63010 58338 63024
rect 58488 63010 58934 63024
rect 16418 62962 58934 63010
rect 16418 62948 16864 62962
rect 17014 62948 17154 62962
rect 17304 62948 18112 62962
rect 18262 62948 18402 62962
rect 18552 62948 19360 62962
rect 19510 62948 19650 62962
rect 19800 62948 20608 62962
rect 20758 62948 20898 62962
rect 21048 62948 21856 62962
rect 22006 62948 22146 62962
rect 22296 62948 23104 62962
rect 23254 62948 23394 62962
rect 23544 62948 24352 62962
rect 24502 62948 24642 62962
rect 24792 62948 25600 62962
rect 25750 62948 25890 62962
rect 26040 62948 26848 62962
rect 26998 62948 27138 62962
rect 27288 62948 28096 62962
rect 28246 62948 28386 62962
rect 28536 62948 29344 62962
rect 29494 62948 29634 62962
rect 29784 62948 30592 62962
rect 30742 62948 30882 62962
rect 31032 62948 31840 62962
rect 31990 62948 32130 62962
rect 32280 62948 33088 62962
rect 33238 62948 33378 62962
rect 33528 62948 34336 62962
rect 34486 62948 34626 62962
rect 34776 62948 35584 62962
rect 35734 62948 35874 62962
rect 36024 62948 36832 62962
rect 36982 62948 37122 62962
rect 37272 62948 38080 62962
rect 38230 62948 38370 62962
rect 38520 62948 39328 62962
rect 39478 62948 39618 62962
rect 39768 62948 40576 62962
rect 40726 62948 40866 62962
rect 41016 62948 41824 62962
rect 41974 62948 42114 62962
rect 42264 62948 43072 62962
rect 43222 62948 43362 62962
rect 43512 62948 44320 62962
rect 44470 62948 44610 62962
rect 44760 62948 45568 62962
rect 45718 62948 45858 62962
rect 46008 62948 46816 62962
rect 46966 62948 47106 62962
rect 47256 62948 48064 62962
rect 48214 62948 48354 62962
rect 48504 62948 49312 62962
rect 49462 62948 49602 62962
rect 49752 62948 50560 62962
rect 50710 62948 50850 62962
rect 51000 62948 51808 62962
rect 51958 62948 52098 62962
rect 52248 62948 53056 62962
rect 53206 62948 53346 62962
rect 53496 62948 54304 62962
rect 54454 62948 54594 62962
rect 54744 62948 55552 62962
rect 55702 62948 55842 62962
rect 55992 62948 56800 62962
rect 56950 62948 57090 62962
rect 57240 62948 58048 62962
rect 58198 62948 58338 62962
rect 58488 62948 58934 62962
rect 16898 62900 16980 62914
rect 17188 62900 17270 62914
rect 18146 62900 18228 62914
rect 18436 62900 18518 62914
rect 19394 62900 19476 62914
rect 19684 62900 19766 62914
rect 20642 62900 20724 62914
rect 20932 62900 21014 62914
rect 21890 62900 21972 62914
rect 22180 62900 22262 62914
rect 23138 62900 23220 62914
rect 23428 62900 23510 62914
rect 24386 62900 24468 62914
rect 24676 62900 24758 62914
rect 25634 62900 25716 62914
rect 25924 62900 26006 62914
rect 26882 62900 26964 62914
rect 27172 62900 27254 62914
rect 28130 62900 28212 62914
rect 28420 62900 28502 62914
rect 29378 62900 29460 62914
rect 29668 62900 29750 62914
rect 30626 62900 30708 62914
rect 30916 62900 30998 62914
rect 31874 62900 31956 62914
rect 32164 62900 32246 62914
rect 33122 62900 33204 62914
rect 33412 62900 33494 62914
rect 34370 62900 34452 62914
rect 34660 62900 34742 62914
rect 35618 62900 35700 62914
rect 35908 62900 35990 62914
rect 36866 62900 36948 62914
rect 37156 62900 37238 62914
rect 38114 62900 38196 62914
rect 38404 62900 38486 62914
rect 39362 62900 39444 62914
rect 39652 62900 39734 62914
rect 40610 62900 40692 62914
rect 40900 62900 40982 62914
rect 41858 62900 41940 62914
rect 42148 62900 42230 62914
rect 43106 62900 43188 62914
rect 43396 62900 43478 62914
rect 44354 62900 44436 62914
rect 44644 62900 44726 62914
rect 45602 62900 45684 62914
rect 45892 62900 45974 62914
rect 46850 62900 46932 62914
rect 47140 62900 47222 62914
rect 48098 62900 48180 62914
rect 48388 62900 48470 62914
rect 49346 62900 49428 62914
rect 49636 62900 49718 62914
rect 50594 62900 50676 62914
rect 50884 62900 50966 62914
rect 51842 62900 51924 62914
rect 52132 62900 52214 62914
rect 53090 62900 53172 62914
rect 53380 62900 53462 62914
rect 54338 62900 54420 62914
rect 54628 62900 54710 62914
rect 55586 62900 55668 62914
rect 55876 62900 55958 62914
rect 56834 62900 56916 62914
rect 57124 62900 57206 62914
rect 58082 62900 58164 62914
rect 58372 62900 58454 62914
rect 16418 62852 58934 62900
rect 16418 62756 58934 62804
rect 16898 62742 16980 62756
rect 17188 62742 17270 62756
rect 18146 62742 18228 62756
rect 18436 62742 18518 62756
rect 19394 62742 19476 62756
rect 19684 62742 19766 62756
rect 20642 62742 20724 62756
rect 20932 62742 21014 62756
rect 21890 62742 21972 62756
rect 22180 62742 22262 62756
rect 23138 62742 23220 62756
rect 23428 62742 23510 62756
rect 24386 62742 24468 62756
rect 24676 62742 24758 62756
rect 25634 62742 25716 62756
rect 25924 62742 26006 62756
rect 26882 62742 26964 62756
rect 27172 62742 27254 62756
rect 28130 62742 28212 62756
rect 28420 62742 28502 62756
rect 29378 62742 29460 62756
rect 29668 62742 29750 62756
rect 30626 62742 30708 62756
rect 30916 62742 30998 62756
rect 31874 62742 31956 62756
rect 32164 62742 32246 62756
rect 33122 62742 33204 62756
rect 33412 62742 33494 62756
rect 34370 62742 34452 62756
rect 34660 62742 34742 62756
rect 35618 62742 35700 62756
rect 35908 62742 35990 62756
rect 36866 62742 36948 62756
rect 37156 62742 37238 62756
rect 38114 62742 38196 62756
rect 38404 62742 38486 62756
rect 39362 62742 39444 62756
rect 39652 62742 39734 62756
rect 40610 62742 40692 62756
rect 40900 62742 40982 62756
rect 41858 62742 41940 62756
rect 42148 62742 42230 62756
rect 43106 62742 43188 62756
rect 43396 62742 43478 62756
rect 44354 62742 44436 62756
rect 44644 62742 44726 62756
rect 45602 62742 45684 62756
rect 45892 62742 45974 62756
rect 46850 62742 46932 62756
rect 47140 62742 47222 62756
rect 48098 62742 48180 62756
rect 48388 62742 48470 62756
rect 49346 62742 49428 62756
rect 49636 62742 49718 62756
rect 50594 62742 50676 62756
rect 50884 62742 50966 62756
rect 51842 62742 51924 62756
rect 52132 62742 52214 62756
rect 53090 62742 53172 62756
rect 53380 62742 53462 62756
rect 54338 62742 54420 62756
rect 54628 62742 54710 62756
rect 55586 62742 55668 62756
rect 55876 62742 55958 62756
rect 56834 62742 56916 62756
rect 57124 62742 57206 62756
rect 58082 62742 58164 62756
rect 58372 62742 58454 62756
rect 16418 62694 16864 62708
rect 17014 62694 17154 62708
rect 17304 62694 18112 62708
rect 18262 62694 18402 62708
rect 18552 62694 19360 62708
rect 19510 62694 19650 62708
rect 19800 62694 20608 62708
rect 20758 62694 20898 62708
rect 21048 62694 21856 62708
rect 22006 62694 22146 62708
rect 22296 62694 23104 62708
rect 23254 62694 23394 62708
rect 23544 62694 24352 62708
rect 24502 62694 24642 62708
rect 24792 62694 25600 62708
rect 25750 62694 25890 62708
rect 26040 62694 26848 62708
rect 26998 62694 27138 62708
rect 27288 62694 28096 62708
rect 28246 62694 28386 62708
rect 28536 62694 29344 62708
rect 29494 62694 29634 62708
rect 29784 62694 30592 62708
rect 30742 62694 30882 62708
rect 31032 62694 31840 62708
rect 31990 62694 32130 62708
rect 32280 62694 33088 62708
rect 33238 62694 33378 62708
rect 33528 62694 34336 62708
rect 34486 62694 34626 62708
rect 34776 62694 35584 62708
rect 35734 62694 35874 62708
rect 36024 62694 36832 62708
rect 36982 62694 37122 62708
rect 37272 62694 38080 62708
rect 38230 62694 38370 62708
rect 38520 62694 39328 62708
rect 39478 62694 39618 62708
rect 39768 62694 40576 62708
rect 40726 62694 40866 62708
rect 41016 62694 41824 62708
rect 41974 62694 42114 62708
rect 42264 62694 43072 62708
rect 43222 62694 43362 62708
rect 43512 62694 44320 62708
rect 44470 62694 44610 62708
rect 44760 62694 45568 62708
rect 45718 62694 45858 62708
rect 46008 62694 46816 62708
rect 46966 62694 47106 62708
rect 47256 62694 48064 62708
rect 48214 62694 48354 62708
rect 48504 62694 49312 62708
rect 49462 62694 49602 62708
rect 49752 62694 50560 62708
rect 50710 62694 50850 62708
rect 51000 62694 51808 62708
rect 51958 62694 52098 62708
rect 52248 62694 53056 62708
rect 53206 62694 53346 62708
rect 53496 62694 54304 62708
rect 54454 62694 54594 62708
rect 54744 62694 55552 62708
rect 55702 62694 55842 62708
rect 55992 62694 56800 62708
rect 56950 62694 57090 62708
rect 57240 62694 58048 62708
rect 58198 62694 58338 62708
rect 58488 62694 58934 62708
rect 16418 62646 58934 62694
rect 16418 62632 16864 62646
rect 17014 62632 17154 62646
rect 17304 62632 18112 62646
rect 18262 62632 18402 62646
rect 18552 62632 19360 62646
rect 19510 62632 19650 62646
rect 19800 62632 20608 62646
rect 20758 62632 20898 62646
rect 21048 62632 21856 62646
rect 22006 62632 22146 62646
rect 22296 62632 23104 62646
rect 23254 62632 23394 62646
rect 23544 62632 24352 62646
rect 24502 62632 24642 62646
rect 24792 62632 25600 62646
rect 25750 62632 25890 62646
rect 26040 62632 26848 62646
rect 26998 62632 27138 62646
rect 27288 62632 28096 62646
rect 28246 62632 28386 62646
rect 28536 62632 29344 62646
rect 29494 62632 29634 62646
rect 29784 62632 30592 62646
rect 30742 62632 30882 62646
rect 31032 62632 31840 62646
rect 31990 62632 32130 62646
rect 32280 62632 33088 62646
rect 33238 62632 33378 62646
rect 33528 62632 34336 62646
rect 34486 62632 34626 62646
rect 34776 62632 35584 62646
rect 35734 62632 35874 62646
rect 36024 62632 36832 62646
rect 36982 62632 37122 62646
rect 37272 62632 38080 62646
rect 38230 62632 38370 62646
rect 38520 62632 39328 62646
rect 39478 62632 39618 62646
rect 39768 62632 40576 62646
rect 40726 62632 40866 62646
rect 41016 62632 41824 62646
rect 41974 62632 42114 62646
rect 42264 62632 43072 62646
rect 43222 62632 43362 62646
rect 43512 62632 44320 62646
rect 44470 62632 44610 62646
rect 44760 62632 45568 62646
rect 45718 62632 45858 62646
rect 46008 62632 46816 62646
rect 46966 62632 47106 62646
rect 47256 62632 48064 62646
rect 48214 62632 48354 62646
rect 48504 62632 49312 62646
rect 49462 62632 49602 62646
rect 49752 62632 50560 62646
rect 50710 62632 50850 62646
rect 51000 62632 51808 62646
rect 51958 62632 52098 62646
rect 52248 62632 53056 62646
rect 53206 62632 53346 62646
rect 53496 62632 54304 62646
rect 54454 62632 54594 62646
rect 54744 62632 55552 62646
rect 55702 62632 55842 62646
rect 55992 62632 56800 62646
rect 56950 62632 57090 62646
rect 57240 62632 58048 62646
rect 58198 62632 58338 62646
rect 58488 62632 58934 62646
rect 16898 62584 16980 62598
rect 17188 62584 17270 62598
rect 18146 62584 18228 62598
rect 18436 62584 18518 62598
rect 19394 62584 19476 62598
rect 19684 62584 19766 62598
rect 20642 62584 20724 62598
rect 20932 62584 21014 62598
rect 21890 62584 21972 62598
rect 22180 62584 22262 62598
rect 23138 62584 23220 62598
rect 23428 62584 23510 62598
rect 24386 62584 24468 62598
rect 24676 62584 24758 62598
rect 25634 62584 25716 62598
rect 25924 62584 26006 62598
rect 26882 62584 26964 62598
rect 27172 62584 27254 62598
rect 28130 62584 28212 62598
rect 28420 62584 28502 62598
rect 29378 62584 29460 62598
rect 29668 62584 29750 62598
rect 30626 62584 30708 62598
rect 30916 62584 30998 62598
rect 31874 62584 31956 62598
rect 32164 62584 32246 62598
rect 33122 62584 33204 62598
rect 33412 62584 33494 62598
rect 34370 62584 34452 62598
rect 34660 62584 34742 62598
rect 35618 62584 35700 62598
rect 35908 62584 35990 62598
rect 36866 62584 36948 62598
rect 37156 62584 37238 62598
rect 38114 62584 38196 62598
rect 38404 62584 38486 62598
rect 39362 62584 39444 62598
rect 39652 62584 39734 62598
rect 40610 62584 40692 62598
rect 40900 62584 40982 62598
rect 41858 62584 41940 62598
rect 42148 62584 42230 62598
rect 43106 62584 43188 62598
rect 43396 62584 43478 62598
rect 44354 62584 44436 62598
rect 44644 62584 44726 62598
rect 45602 62584 45684 62598
rect 45892 62584 45974 62598
rect 46850 62584 46932 62598
rect 47140 62584 47222 62598
rect 48098 62584 48180 62598
rect 48388 62584 48470 62598
rect 49346 62584 49428 62598
rect 49636 62584 49718 62598
rect 50594 62584 50676 62598
rect 50884 62584 50966 62598
rect 51842 62584 51924 62598
rect 52132 62584 52214 62598
rect 53090 62584 53172 62598
rect 53380 62584 53462 62598
rect 54338 62584 54420 62598
rect 54628 62584 54710 62598
rect 55586 62584 55668 62598
rect 55876 62584 55958 62598
rect 56834 62584 56916 62598
rect 57124 62584 57206 62598
rect 58082 62584 58164 62598
rect 58372 62584 58454 62598
rect 16418 62536 58934 62584
rect 16418 62378 58934 62488
rect 16418 62282 58934 62330
rect 16898 62268 16980 62282
rect 17188 62268 17270 62282
rect 18146 62268 18228 62282
rect 18436 62268 18518 62282
rect 19394 62268 19476 62282
rect 19684 62268 19766 62282
rect 20642 62268 20724 62282
rect 20932 62268 21014 62282
rect 21890 62268 21972 62282
rect 22180 62268 22262 62282
rect 23138 62268 23220 62282
rect 23428 62268 23510 62282
rect 24386 62268 24468 62282
rect 24676 62268 24758 62282
rect 25634 62268 25716 62282
rect 25924 62268 26006 62282
rect 26882 62268 26964 62282
rect 27172 62268 27254 62282
rect 28130 62268 28212 62282
rect 28420 62268 28502 62282
rect 29378 62268 29460 62282
rect 29668 62268 29750 62282
rect 30626 62268 30708 62282
rect 30916 62268 30998 62282
rect 31874 62268 31956 62282
rect 32164 62268 32246 62282
rect 33122 62268 33204 62282
rect 33412 62268 33494 62282
rect 34370 62268 34452 62282
rect 34660 62268 34742 62282
rect 35618 62268 35700 62282
rect 35908 62268 35990 62282
rect 36866 62268 36948 62282
rect 37156 62268 37238 62282
rect 38114 62268 38196 62282
rect 38404 62268 38486 62282
rect 39362 62268 39444 62282
rect 39652 62268 39734 62282
rect 40610 62268 40692 62282
rect 40900 62268 40982 62282
rect 41858 62268 41940 62282
rect 42148 62268 42230 62282
rect 43106 62268 43188 62282
rect 43396 62268 43478 62282
rect 44354 62268 44436 62282
rect 44644 62268 44726 62282
rect 45602 62268 45684 62282
rect 45892 62268 45974 62282
rect 46850 62268 46932 62282
rect 47140 62268 47222 62282
rect 48098 62268 48180 62282
rect 48388 62268 48470 62282
rect 49346 62268 49428 62282
rect 49636 62268 49718 62282
rect 50594 62268 50676 62282
rect 50884 62268 50966 62282
rect 51842 62268 51924 62282
rect 52132 62268 52214 62282
rect 53090 62268 53172 62282
rect 53380 62268 53462 62282
rect 54338 62268 54420 62282
rect 54628 62268 54710 62282
rect 55586 62268 55668 62282
rect 55876 62268 55958 62282
rect 56834 62268 56916 62282
rect 57124 62268 57206 62282
rect 58082 62268 58164 62282
rect 58372 62268 58454 62282
rect 16418 62220 16864 62234
rect 17014 62220 17154 62234
rect 17304 62220 18112 62234
rect 18262 62220 18402 62234
rect 18552 62220 19360 62234
rect 19510 62220 19650 62234
rect 19800 62220 20608 62234
rect 20758 62220 20898 62234
rect 21048 62220 21856 62234
rect 22006 62220 22146 62234
rect 22296 62220 23104 62234
rect 23254 62220 23394 62234
rect 23544 62220 24352 62234
rect 24502 62220 24642 62234
rect 24792 62220 25600 62234
rect 25750 62220 25890 62234
rect 26040 62220 26848 62234
rect 26998 62220 27138 62234
rect 27288 62220 28096 62234
rect 28246 62220 28386 62234
rect 28536 62220 29344 62234
rect 29494 62220 29634 62234
rect 29784 62220 30592 62234
rect 30742 62220 30882 62234
rect 31032 62220 31840 62234
rect 31990 62220 32130 62234
rect 32280 62220 33088 62234
rect 33238 62220 33378 62234
rect 33528 62220 34336 62234
rect 34486 62220 34626 62234
rect 34776 62220 35584 62234
rect 35734 62220 35874 62234
rect 36024 62220 36832 62234
rect 36982 62220 37122 62234
rect 37272 62220 38080 62234
rect 38230 62220 38370 62234
rect 38520 62220 39328 62234
rect 39478 62220 39618 62234
rect 39768 62220 40576 62234
rect 40726 62220 40866 62234
rect 41016 62220 41824 62234
rect 41974 62220 42114 62234
rect 42264 62220 43072 62234
rect 43222 62220 43362 62234
rect 43512 62220 44320 62234
rect 44470 62220 44610 62234
rect 44760 62220 45568 62234
rect 45718 62220 45858 62234
rect 46008 62220 46816 62234
rect 46966 62220 47106 62234
rect 47256 62220 48064 62234
rect 48214 62220 48354 62234
rect 48504 62220 49312 62234
rect 49462 62220 49602 62234
rect 49752 62220 50560 62234
rect 50710 62220 50850 62234
rect 51000 62220 51808 62234
rect 51958 62220 52098 62234
rect 52248 62220 53056 62234
rect 53206 62220 53346 62234
rect 53496 62220 54304 62234
rect 54454 62220 54594 62234
rect 54744 62220 55552 62234
rect 55702 62220 55842 62234
rect 55992 62220 56800 62234
rect 56950 62220 57090 62234
rect 57240 62220 58048 62234
rect 58198 62220 58338 62234
rect 58488 62220 58934 62234
rect 16418 62172 58934 62220
rect 16418 62158 16864 62172
rect 17014 62158 17154 62172
rect 17304 62158 18112 62172
rect 18262 62158 18402 62172
rect 18552 62158 19360 62172
rect 19510 62158 19650 62172
rect 19800 62158 20608 62172
rect 20758 62158 20898 62172
rect 21048 62158 21856 62172
rect 22006 62158 22146 62172
rect 22296 62158 23104 62172
rect 23254 62158 23394 62172
rect 23544 62158 24352 62172
rect 24502 62158 24642 62172
rect 24792 62158 25600 62172
rect 25750 62158 25890 62172
rect 26040 62158 26848 62172
rect 26998 62158 27138 62172
rect 27288 62158 28096 62172
rect 28246 62158 28386 62172
rect 28536 62158 29344 62172
rect 29494 62158 29634 62172
rect 29784 62158 30592 62172
rect 30742 62158 30882 62172
rect 31032 62158 31840 62172
rect 31990 62158 32130 62172
rect 32280 62158 33088 62172
rect 33238 62158 33378 62172
rect 33528 62158 34336 62172
rect 34486 62158 34626 62172
rect 34776 62158 35584 62172
rect 35734 62158 35874 62172
rect 36024 62158 36832 62172
rect 36982 62158 37122 62172
rect 37272 62158 38080 62172
rect 38230 62158 38370 62172
rect 38520 62158 39328 62172
rect 39478 62158 39618 62172
rect 39768 62158 40576 62172
rect 40726 62158 40866 62172
rect 41016 62158 41824 62172
rect 41974 62158 42114 62172
rect 42264 62158 43072 62172
rect 43222 62158 43362 62172
rect 43512 62158 44320 62172
rect 44470 62158 44610 62172
rect 44760 62158 45568 62172
rect 45718 62158 45858 62172
rect 46008 62158 46816 62172
rect 46966 62158 47106 62172
rect 47256 62158 48064 62172
rect 48214 62158 48354 62172
rect 48504 62158 49312 62172
rect 49462 62158 49602 62172
rect 49752 62158 50560 62172
rect 50710 62158 50850 62172
rect 51000 62158 51808 62172
rect 51958 62158 52098 62172
rect 52248 62158 53056 62172
rect 53206 62158 53346 62172
rect 53496 62158 54304 62172
rect 54454 62158 54594 62172
rect 54744 62158 55552 62172
rect 55702 62158 55842 62172
rect 55992 62158 56800 62172
rect 56950 62158 57090 62172
rect 57240 62158 58048 62172
rect 58198 62158 58338 62172
rect 58488 62158 58934 62172
rect 16898 62110 16980 62124
rect 17188 62110 17270 62124
rect 18146 62110 18228 62124
rect 18436 62110 18518 62124
rect 19394 62110 19476 62124
rect 19684 62110 19766 62124
rect 20642 62110 20724 62124
rect 20932 62110 21014 62124
rect 21890 62110 21972 62124
rect 22180 62110 22262 62124
rect 23138 62110 23220 62124
rect 23428 62110 23510 62124
rect 24386 62110 24468 62124
rect 24676 62110 24758 62124
rect 25634 62110 25716 62124
rect 25924 62110 26006 62124
rect 26882 62110 26964 62124
rect 27172 62110 27254 62124
rect 28130 62110 28212 62124
rect 28420 62110 28502 62124
rect 29378 62110 29460 62124
rect 29668 62110 29750 62124
rect 30626 62110 30708 62124
rect 30916 62110 30998 62124
rect 31874 62110 31956 62124
rect 32164 62110 32246 62124
rect 33122 62110 33204 62124
rect 33412 62110 33494 62124
rect 34370 62110 34452 62124
rect 34660 62110 34742 62124
rect 35618 62110 35700 62124
rect 35908 62110 35990 62124
rect 36866 62110 36948 62124
rect 37156 62110 37238 62124
rect 38114 62110 38196 62124
rect 38404 62110 38486 62124
rect 39362 62110 39444 62124
rect 39652 62110 39734 62124
rect 40610 62110 40692 62124
rect 40900 62110 40982 62124
rect 41858 62110 41940 62124
rect 42148 62110 42230 62124
rect 43106 62110 43188 62124
rect 43396 62110 43478 62124
rect 44354 62110 44436 62124
rect 44644 62110 44726 62124
rect 45602 62110 45684 62124
rect 45892 62110 45974 62124
rect 46850 62110 46932 62124
rect 47140 62110 47222 62124
rect 48098 62110 48180 62124
rect 48388 62110 48470 62124
rect 49346 62110 49428 62124
rect 49636 62110 49718 62124
rect 50594 62110 50676 62124
rect 50884 62110 50966 62124
rect 51842 62110 51924 62124
rect 52132 62110 52214 62124
rect 53090 62110 53172 62124
rect 53380 62110 53462 62124
rect 54338 62110 54420 62124
rect 54628 62110 54710 62124
rect 55586 62110 55668 62124
rect 55876 62110 55958 62124
rect 56834 62110 56916 62124
rect 57124 62110 57206 62124
rect 58082 62110 58164 62124
rect 58372 62110 58454 62124
rect 16418 62062 58934 62110
rect 16418 61966 58934 62014
rect 16898 61952 16980 61966
rect 17188 61952 17270 61966
rect 18146 61952 18228 61966
rect 18436 61952 18518 61966
rect 19394 61952 19476 61966
rect 19684 61952 19766 61966
rect 20642 61952 20724 61966
rect 20932 61952 21014 61966
rect 21890 61952 21972 61966
rect 22180 61952 22262 61966
rect 23138 61952 23220 61966
rect 23428 61952 23510 61966
rect 24386 61952 24468 61966
rect 24676 61952 24758 61966
rect 25634 61952 25716 61966
rect 25924 61952 26006 61966
rect 26882 61952 26964 61966
rect 27172 61952 27254 61966
rect 28130 61952 28212 61966
rect 28420 61952 28502 61966
rect 29378 61952 29460 61966
rect 29668 61952 29750 61966
rect 30626 61952 30708 61966
rect 30916 61952 30998 61966
rect 31874 61952 31956 61966
rect 32164 61952 32246 61966
rect 33122 61952 33204 61966
rect 33412 61952 33494 61966
rect 34370 61952 34452 61966
rect 34660 61952 34742 61966
rect 35618 61952 35700 61966
rect 35908 61952 35990 61966
rect 36866 61952 36948 61966
rect 37156 61952 37238 61966
rect 38114 61952 38196 61966
rect 38404 61952 38486 61966
rect 39362 61952 39444 61966
rect 39652 61952 39734 61966
rect 40610 61952 40692 61966
rect 40900 61952 40982 61966
rect 41858 61952 41940 61966
rect 42148 61952 42230 61966
rect 43106 61952 43188 61966
rect 43396 61952 43478 61966
rect 44354 61952 44436 61966
rect 44644 61952 44726 61966
rect 45602 61952 45684 61966
rect 45892 61952 45974 61966
rect 46850 61952 46932 61966
rect 47140 61952 47222 61966
rect 48098 61952 48180 61966
rect 48388 61952 48470 61966
rect 49346 61952 49428 61966
rect 49636 61952 49718 61966
rect 50594 61952 50676 61966
rect 50884 61952 50966 61966
rect 51842 61952 51924 61966
rect 52132 61952 52214 61966
rect 53090 61952 53172 61966
rect 53380 61952 53462 61966
rect 54338 61952 54420 61966
rect 54628 61952 54710 61966
rect 55586 61952 55668 61966
rect 55876 61952 55958 61966
rect 56834 61952 56916 61966
rect 57124 61952 57206 61966
rect 58082 61952 58164 61966
rect 58372 61952 58454 61966
rect 16418 61904 16864 61918
rect 17014 61904 17154 61918
rect 17304 61904 18112 61918
rect 18262 61904 18402 61918
rect 18552 61904 19360 61918
rect 19510 61904 19650 61918
rect 19800 61904 20608 61918
rect 20758 61904 20898 61918
rect 21048 61904 21856 61918
rect 22006 61904 22146 61918
rect 22296 61904 23104 61918
rect 23254 61904 23394 61918
rect 23544 61904 24352 61918
rect 24502 61904 24642 61918
rect 24792 61904 25600 61918
rect 25750 61904 25890 61918
rect 26040 61904 26848 61918
rect 26998 61904 27138 61918
rect 27288 61904 28096 61918
rect 28246 61904 28386 61918
rect 28536 61904 29344 61918
rect 29494 61904 29634 61918
rect 29784 61904 30592 61918
rect 30742 61904 30882 61918
rect 31032 61904 31840 61918
rect 31990 61904 32130 61918
rect 32280 61904 33088 61918
rect 33238 61904 33378 61918
rect 33528 61904 34336 61918
rect 34486 61904 34626 61918
rect 34776 61904 35584 61918
rect 35734 61904 35874 61918
rect 36024 61904 36832 61918
rect 36982 61904 37122 61918
rect 37272 61904 38080 61918
rect 38230 61904 38370 61918
rect 38520 61904 39328 61918
rect 39478 61904 39618 61918
rect 39768 61904 40576 61918
rect 40726 61904 40866 61918
rect 41016 61904 41824 61918
rect 41974 61904 42114 61918
rect 42264 61904 43072 61918
rect 43222 61904 43362 61918
rect 43512 61904 44320 61918
rect 44470 61904 44610 61918
rect 44760 61904 45568 61918
rect 45718 61904 45858 61918
rect 46008 61904 46816 61918
rect 46966 61904 47106 61918
rect 47256 61904 48064 61918
rect 48214 61904 48354 61918
rect 48504 61904 49312 61918
rect 49462 61904 49602 61918
rect 49752 61904 50560 61918
rect 50710 61904 50850 61918
rect 51000 61904 51808 61918
rect 51958 61904 52098 61918
rect 52248 61904 53056 61918
rect 53206 61904 53346 61918
rect 53496 61904 54304 61918
rect 54454 61904 54594 61918
rect 54744 61904 55552 61918
rect 55702 61904 55842 61918
rect 55992 61904 56800 61918
rect 56950 61904 57090 61918
rect 57240 61904 58048 61918
rect 58198 61904 58338 61918
rect 58488 61904 58934 61918
rect 16418 61856 58934 61904
rect 16418 61842 16864 61856
rect 17014 61842 17154 61856
rect 17304 61842 18112 61856
rect 18262 61842 18402 61856
rect 18552 61842 19360 61856
rect 19510 61842 19650 61856
rect 19800 61842 20608 61856
rect 20758 61842 20898 61856
rect 21048 61842 21856 61856
rect 22006 61842 22146 61856
rect 22296 61842 23104 61856
rect 23254 61842 23394 61856
rect 23544 61842 24352 61856
rect 24502 61842 24642 61856
rect 24792 61842 25600 61856
rect 25750 61842 25890 61856
rect 26040 61842 26848 61856
rect 26998 61842 27138 61856
rect 27288 61842 28096 61856
rect 28246 61842 28386 61856
rect 28536 61842 29344 61856
rect 29494 61842 29634 61856
rect 29784 61842 30592 61856
rect 30742 61842 30882 61856
rect 31032 61842 31840 61856
rect 31990 61842 32130 61856
rect 32280 61842 33088 61856
rect 33238 61842 33378 61856
rect 33528 61842 34336 61856
rect 34486 61842 34626 61856
rect 34776 61842 35584 61856
rect 35734 61842 35874 61856
rect 36024 61842 36832 61856
rect 36982 61842 37122 61856
rect 37272 61842 38080 61856
rect 38230 61842 38370 61856
rect 38520 61842 39328 61856
rect 39478 61842 39618 61856
rect 39768 61842 40576 61856
rect 40726 61842 40866 61856
rect 41016 61842 41824 61856
rect 41974 61842 42114 61856
rect 42264 61842 43072 61856
rect 43222 61842 43362 61856
rect 43512 61842 44320 61856
rect 44470 61842 44610 61856
rect 44760 61842 45568 61856
rect 45718 61842 45858 61856
rect 46008 61842 46816 61856
rect 46966 61842 47106 61856
rect 47256 61842 48064 61856
rect 48214 61842 48354 61856
rect 48504 61842 49312 61856
rect 49462 61842 49602 61856
rect 49752 61842 50560 61856
rect 50710 61842 50850 61856
rect 51000 61842 51808 61856
rect 51958 61842 52098 61856
rect 52248 61842 53056 61856
rect 53206 61842 53346 61856
rect 53496 61842 54304 61856
rect 54454 61842 54594 61856
rect 54744 61842 55552 61856
rect 55702 61842 55842 61856
rect 55992 61842 56800 61856
rect 56950 61842 57090 61856
rect 57240 61842 58048 61856
rect 58198 61842 58338 61856
rect 58488 61842 58934 61856
rect 16898 61794 16980 61808
rect 17188 61794 17270 61808
rect 18146 61794 18228 61808
rect 18436 61794 18518 61808
rect 19394 61794 19476 61808
rect 19684 61794 19766 61808
rect 20642 61794 20724 61808
rect 20932 61794 21014 61808
rect 21890 61794 21972 61808
rect 22180 61794 22262 61808
rect 23138 61794 23220 61808
rect 23428 61794 23510 61808
rect 24386 61794 24468 61808
rect 24676 61794 24758 61808
rect 25634 61794 25716 61808
rect 25924 61794 26006 61808
rect 26882 61794 26964 61808
rect 27172 61794 27254 61808
rect 28130 61794 28212 61808
rect 28420 61794 28502 61808
rect 29378 61794 29460 61808
rect 29668 61794 29750 61808
rect 30626 61794 30708 61808
rect 30916 61794 30998 61808
rect 31874 61794 31956 61808
rect 32164 61794 32246 61808
rect 33122 61794 33204 61808
rect 33412 61794 33494 61808
rect 34370 61794 34452 61808
rect 34660 61794 34742 61808
rect 35618 61794 35700 61808
rect 35908 61794 35990 61808
rect 36866 61794 36948 61808
rect 37156 61794 37238 61808
rect 38114 61794 38196 61808
rect 38404 61794 38486 61808
rect 39362 61794 39444 61808
rect 39652 61794 39734 61808
rect 40610 61794 40692 61808
rect 40900 61794 40982 61808
rect 41858 61794 41940 61808
rect 42148 61794 42230 61808
rect 43106 61794 43188 61808
rect 43396 61794 43478 61808
rect 44354 61794 44436 61808
rect 44644 61794 44726 61808
rect 45602 61794 45684 61808
rect 45892 61794 45974 61808
rect 46850 61794 46932 61808
rect 47140 61794 47222 61808
rect 48098 61794 48180 61808
rect 48388 61794 48470 61808
rect 49346 61794 49428 61808
rect 49636 61794 49718 61808
rect 50594 61794 50676 61808
rect 50884 61794 50966 61808
rect 51842 61794 51924 61808
rect 52132 61794 52214 61808
rect 53090 61794 53172 61808
rect 53380 61794 53462 61808
rect 54338 61794 54420 61808
rect 54628 61794 54710 61808
rect 55586 61794 55668 61808
rect 55876 61794 55958 61808
rect 56834 61794 56916 61808
rect 57124 61794 57206 61808
rect 58082 61794 58164 61808
rect 58372 61794 58454 61808
rect 16418 61746 58934 61794
rect 16418 61588 58934 61698
rect 16418 61492 58934 61540
rect 16898 61478 16980 61492
rect 17188 61478 17270 61492
rect 18146 61478 18228 61492
rect 18436 61478 18518 61492
rect 19394 61478 19476 61492
rect 19684 61478 19766 61492
rect 20642 61478 20724 61492
rect 20932 61478 21014 61492
rect 21890 61478 21972 61492
rect 22180 61478 22262 61492
rect 23138 61478 23220 61492
rect 23428 61478 23510 61492
rect 24386 61478 24468 61492
rect 24676 61478 24758 61492
rect 25634 61478 25716 61492
rect 25924 61478 26006 61492
rect 26882 61478 26964 61492
rect 27172 61478 27254 61492
rect 28130 61478 28212 61492
rect 28420 61478 28502 61492
rect 29378 61478 29460 61492
rect 29668 61478 29750 61492
rect 30626 61478 30708 61492
rect 30916 61478 30998 61492
rect 31874 61478 31956 61492
rect 32164 61478 32246 61492
rect 33122 61478 33204 61492
rect 33412 61478 33494 61492
rect 34370 61478 34452 61492
rect 34660 61478 34742 61492
rect 35618 61478 35700 61492
rect 35908 61478 35990 61492
rect 36866 61478 36948 61492
rect 37156 61478 37238 61492
rect 38114 61478 38196 61492
rect 38404 61478 38486 61492
rect 39362 61478 39444 61492
rect 39652 61478 39734 61492
rect 40610 61478 40692 61492
rect 40900 61478 40982 61492
rect 41858 61478 41940 61492
rect 42148 61478 42230 61492
rect 43106 61478 43188 61492
rect 43396 61478 43478 61492
rect 44354 61478 44436 61492
rect 44644 61478 44726 61492
rect 45602 61478 45684 61492
rect 45892 61478 45974 61492
rect 46850 61478 46932 61492
rect 47140 61478 47222 61492
rect 48098 61478 48180 61492
rect 48388 61478 48470 61492
rect 49346 61478 49428 61492
rect 49636 61478 49718 61492
rect 50594 61478 50676 61492
rect 50884 61478 50966 61492
rect 51842 61478 51924 61492
rect 52132 61478 52214 61492
rect 53090 61478 53172 61492
rect 53380 61478 53462 61492
rect 54338 61478 54420 61492
rect 54628 61478 54710 61492
rect 55586 61478 55668 61492
rect 55876 61478 55958 61492
rect 56834 61478 56916 61492
rect 57124 61478 57206 61492
rect 58082 61478 58164 61492
rect 58372 61478 58454 61492
rect 16418 61430 16864 61444
rect 17014 61430 17154 61444
rect 17304 61430 18112 61444
rect 18262 61430 18402 61444
rect 18552 61430 19360 61444
rect 19510 61430 19650 61444
rect 19800 61430 20608 61444
rect 20758 61430 20898 61444
rect 21048 61430 21856 61444
rect 22006 61430 22146 61444
rect 22296 61430 23104 61444
rect 23254 61430 23394 61444
rect 23544 61430 24352 61444
rect 24502 61430 24642 61444
rect 24792 61430 25600 61444
rect 25750 61430 25890 61444
rect 26040 61430 26848 61444
rect 26998 61430 27138 61444
rect 27288 61430 28096 61444
rect 28246 61430 28386 61444
rect 28536 61430 29344 61444
rect 29494 61430 29634 61444
rect 29784 61430 30592 61444
rect 30742 61430 30882 61444
rect 31032 61430 31840 61444
rect 31990 61430 32130 61444
rect 32280 61430 33088 61444
rect 33238 61430 33378 61444
rect 33528 61430 34336 61444
rect 34486 61430 34626 61444
rect 34776 61430 35584 61444
rect 35734 61430 35874 61444
rect 36024 61430 36832 61444
rect 36982 61430 37122 61444
rect 37272 61430 38080 61444
rect 38230 61430 38370 61444
rect 38520 61430 39328 61444
rect 39478 61430 39618 61444
rect 39768 61430 40576 61444
rect 40726 61430 40866 61444
rect 41016 61430 41824 61444
rect 41974 61430 42114 61444
rect 42264 61430 43072 61444
rect 43222 61430 43362 61444
rect 43512 61430 44320 61444
rect 44470 61430 44610 61444
rect 44760 61430 45568 61444
rect 45718 61430 45858 61444
rect 46008 61430 46816 61444
rect 46966 61430 47106 61444
rect 47256 61430 48064 61444
rect 48214 61430 48354 61444
rect 48504 61430 49312 61444
rect 49462 61430 49602 61444
rect 49752 61430 50560 61444
rect 50710 61430 50850 61444
rect 51000 61430 51808 61444
rect 51958 61430 52098 61444
rect 52248 61430 53056 61444
rect 53206 61430 53346 61444
rect 53496 61430 54304 61444
rect 54454 61430 54594 61444
rect 54744 61430 55552 61444
rect 55702 61430 55842 61444
rect 55992 61430 56800 61444
rect 56950 61430 57090 61444
rect 57240 61430 58048 61444
rect 58198 61430 58338 61444
rect 58488 61430 58934 61444
rect 16418 61382 58934 61430
rect 16418 61368 16864 61382
rect 17014 61368 17154 61382
rect 17304 61368 18112 61382
rect 18262 61368 18402 61382
rect 18552 61368 19360 61382
rect 19510 61368 19650 61382
rect 19800 61368 20608 61382
rect 20758 61368 20898 61382
rect 21048 61368 21856 61382
rect 22006 61368 22146 61382
rect 22296 61368 23104 61382
rect 23254 61368 23394 61382
rect 23544 61368 24352 61382
rect 24502 61368 24642 61382
rect 24792 61368 25600 61382
rect 25750 61368 25890 61382
rect 26040 61368 26848 61382
rect 26998 61368 27138 61382
rect 27288 61368 28096 61382
rect 28246 61368 28386 61382
rect 28536 61368 29344 61382
rect 29494 61368 29634 61382
rect 29784 61368 30592 61382
rect 30742 61368 30882 61382
rect 31032 61368 31840 61382
rect 31990 61368 32130 61382
rect 32280 61368 33088 61382
rect 33238 61368 33378 61382
rect 33528 61368 34336 61382
rect 34486 61368 34626 61382
rect 34776 61368 35584 61382
rect 35734 61368 35874 61382
rect 36024 61368 36832 61382
rect 36982 61368 37122 61382
rect 37272 61368 38080 61382
rect 38230 61368 38370 61382
rect 38520 61368 39328 61382
rect 39478 61368 39618 61382
rect 39768 61368 40576 61382
rect 40726 61368 40866 61382
rect 41016 61368 41824 61382
rect 41974 61368 42114 61382
rect 42264 61368 43072 61382
rect 43222 61368 43362 61382
rect 43512 61368 44320 61382
rect 44470 61368 44610 61382
rect 44760 61368 45568 61382
rect 45718 61368 45858 61382
rect 46008 61368 46816 61382
rect 46966 61368 47106 61382
rect 47256 61368 48064 61382
rect 48214 61368 48354 61382
rect 48504 61368 49312 61382
rect 49462 61368 49602 61382
rect 49752 61368 50560 61382
rect 50710 61368 50850 61382
rect 51000 61368 51808 61382
rect 51958 61368 52098 61382
rect 52248 61368 53056 61382
rect 53206 61368 53346 61382
rect 53496 61368 54304 61382
rect 54454 61368 54594 61382
rect 54744 61368 55552 61382
rect 55702 61368 55842 61382
rect 55992 61368 56800 61382
rect 56950 61368 57090 61382
rect 57240 61368 58048 61382
rect 58198 61368 58338 61382
rect 58488 61368 58934 61382
rect 16898 61320 16980 61334
rect 17188 61320 17270 61334
rect 18146 61320 18228 61334
rect 18436 61320 18518 61334
rect 19394 61320 19476 61334
rect 19684 61320 19766 61334
rect 20642 61320 20724 61334
rect 20932 61320 21014 61334
rect 21890 61320 21972 61334
rect 22180 61320 22262 61334
rect 23138 61320 23220 61334
rect 23428 61320 23510 61334
rect 24386 61320 24468 61334
rect 24676 61320 24758 61334
rect 25634 61320 25716 61334
rect 25924 61320 26006 61334
rect 26882 61320 26964 61334
rect 27172 61320 27254 61334
rect 28130 61320 28212 61334
rect 28420 61320 28502 61334
rect 29378 61320 29460 61334
rect 29668 61320 29750 61334
rect 30626 61320 30708 61334
rect 30916 61320 30998 61334
rect 31874 61320 31956 61334
rect 32164 61320 32246 61334
rect 33122 61320 33204 61334
rect 33412 61320 33494 61334
rect 34370 61320 34452 61334
rect 34660 61320 34742 61334
rect 35618 61320 35700 61334
rect 35908 61320 35990 61334
rect 36866 61320 36948 61334
rect 37156 61320 37238 61334
rect 38114 61320 38196 61334
rect 38404 61320 38486 61334
rect 39362 61320 39444 61334
rect 39652 61320 39734 61334
rect 40610 61320 40692 61334
rect 40900 61320 40982 61334
rect 41858 61320 41940 61334
rect 42148 61320 42230 61334
rect 43106 61320 43188 61334
rect 43396 61320 43478 61334
rect 44354 61320 44436 61334
rect 44644 61320 44726 61334
rect 45602 61320 45684 61334
rect 45892 61320 45974 61334
rect 46850 61320 46932 61334
rect 47140 61320 47222 61334
rect 48098 61320 48180 61334
rect 48388 61320 48470 61334
rect 49346 61320 49428 61334
rect 49636 61320 49718 61334
rect 50594 61320 50676 61334
rect 50884 61320 50966 61334
rect 51842 61320 51924 61334
rect 52132 61320 52214 61334
rect 53090 61320 53172 61334
rect 53380 61320 53462 61334
rect 54338 61320 54420 61334
rect 54628 61320 54710 61334
rect 55586 61320 55668 61334
rect 55876 61320 55958 61334
rect 56834 61320 56916 61334
rect 57124 61320 57206 61334
rect 58082 61320 58164 61334
rect 58372 61320 58454 61334
rect 16418 61272 58934 61320
rect 16418 61176 58934 61224
rect 16898 61162 16980 61176
rect 17188 61162 17270 61176
rect 18146 61162 18228 61176
rect 18436 61162 18518 61176
rect 19394 61162 19476 61176
rect 19684 61162 19766 61176
rect 20642 61162 20724 61176
rect 20932 61162 21014 61176
rect 21890 61162 21972 61176
rect 22180 61162 22262 61176
rect 23138 61162 23220 61176
rect 23428 61162 23510 61176
rect 24386 61162 24468 61176
rect 24676 61162 24758 61176
rect 25634 61162 25716 61176
rect 25924 61162 26006 61176
rect 26882 61162 26964 61176
rect 27172 61162 27254 61176
rect 28130 61162 28212 61176
rect 28420 61162 28502 61176
rect 29378 61162 29460 61176
rect 29668 61162 29750 61176
rect 30626 61162 30708 61176
rect 30916 61162 30998 61176
rect 31874 61162 31956 61176
rect 32164 61162 32246 61176
rect 33122 61162 33204 61176
rect 33412 61162 33494 61176
rect 34370 61162 34452 61176
rect 34660 61162 34742 61176
rect 35618 61162 35700 61176
rect 35908 61162 35990 61176
rect 36866 61162 36948 61176
rect 37156 61162 37238 61176
rect 38114 61162 38196 61176
rect 38404 61162 38486 61176
rect 39362 61162 39444 61176
rect 39652 61162 39734 61176
rect 40610 61162 40692 61176
rect 40900 61162 40982 61176
rect 41858 61162 41940 61176
rect 42148 61162 42230 61176
rect 43106 61162 43188 61176
rect 43396 61162 43478 61176
rect 44354 61162 44436 61176
rect 44644 61162 44726 61176
rect 45602 61162 45684 61176
rect 45892 61162 45974 61176
rect 46850 61162 46932 61176
rect 47140 61162 47222 61176
rect 48098 61162 48180 61176
rect 48388 61162 48470 61176
rect 49346 61162 49428 61176
rect 49636 61162 49718 61176
rect 50594 61162 50676 61176
rect 50884 61162 50966 61176
rect 51842 61162 51924 61176
rect 52132 61162 52214 61176
rect 53090 61162 53172 61176
rect 53380 61162 53462 61176
rect 54338 61162 54420 61176
rect 54628 61162 54710 61176
rect 55586 61162 55668 61176
rect 55876 61162 55958 61176
rect 56834 61162 56916 61176
rect 57124 61162 57206 61176
rect 58082 61162 58164 61176
rect 58372 61162 58454 61176
rect 16418 61114 16864 61128
rect 17014 61114 17154 61128
rect 17304 61114 18112 61128
rect 18262 61114 18402 61128
rect 18552 61114 19360 61128
rect 19510 61114 19650 61128
rect 19800 61114 20608 61128
rect 20758 61114 20898 61128
rect 21048 61114 21856 61128
rect 22006 61114 22146 61128
rect 22296 61114 23104 61128
rect 23254 61114 23394 61128
rect 23544 61114 24352 61128
rect 24502 61114 24642 61128
rect 24792 61114 25600 61128
rect 25750 61114 25890 61128
rect 26040 61114 26848 61128
rect 26998 61114 27138 61128
rect 27288 61114 28096 61128
rect 28246 61114 28386 61128
rect 28536 61114 29344 61128
rect 29494 61114 29634 61128
rect 29784 61114 30592 61128
rect 30742 61114 30882 61128
rect 31032 61114 31840 61128
rect 31990 61114 32130 61128
rect 32280 61114 33088 61128
rect 33238 61114 33378 61128
rect 33528 61114 34336 61128
rect 34486 61114 34626 61128
rect 34776 61114 35584 61128
rect 35734 61114 35874 61128
rect 36024 61114 36832 61128
rect 36982 61114 37122 61128
rect 37272 61114 38080 61128
rect 38230 61114 38370 61128
rect 38520 61114 39328 61128
rect 39478 61114 39618 61128
rect 39768 61114 40576 61128
rect 40726 61114 40866 61128
rect 41016 61114 41824 61128
rect 41974 61114 42114 61128
rect 42264 61114 43072 61128
rect 43222 61114 43362 61128
rect 43512 61114 44320 61128
rect 44470 61114 44610 61128
rect 44760 61114 45568 61128
rect 45718 61114 45858 61128
rect 46008 61114 46816 61128
rect 46966 61114 47106 61128
rect 47256 61114 48064 61128
rect 48214 61114 48354 61128
rect 48504 61114 49312 61128
rect 49462 61114 49602 61128
rect 49752 61114 50560 61128
rect 50710 61114 50850 61128
rect 51000 61114 51808 61128
rect 51958 61114 52098 61128
rect 52248 61114 53056 61128
rect 53206 61114 53346 61128
rect 53496 61114 54304 61128
rect 54454 61114 54594 61128
rect 54744 61114 55552 61128
rect 55702 61114 55842 61128
rect 55992 61114 56800 61128
rect 56950 61114 57090 61128
rect 57240 61114 58048 61128
rect 58198 61114 58338 61128
rect 58488 61114 58934 61128
rect 16418 61066 58934 61114
rect 16418 61052 16864 61066
rect 17014 61052 17154 61066
rect 17304 61052 18112 61066
rect 18262 61052 18402 61066
rect 18552 61052 19360 61066
rect 19510 61052 19650 61066
rect 19800 61052 20608 61066
rect 20758 61052 20898 61066
rect 21048 61052 21856 61066
rect 22006 61052 22146 61066
rect 22296 61052 23104 61066
rect 23254 61052 23394 61066
rect 23544 61052 24352 61066
rect 24502 61052 24642 61066
rect 24792 61052 25600 61066
rect 25750 61052 25890 61066
rect 26040 61052 26848 61066
rect 26998 61052 27138 61066
rect 27288 61052 28096 61066
rect 28246 61052 28386 61066
rect 28536 61052 29344 61066
rect 29494 61052 29634 61066
rect 29784 61052 30592 61066
rect 30742 61052 30882 61066
rect 31032 61052 31840 61066
rect 31990 61052 32130 61066
rect 32280 61052 33088 61066
rect 33238 61052 33378 61066
rect 33528 61052 34336 61066
rect 34486 61052 34626 61066
rect 34776 61052 35584 61066
rect 35734 61052 35874 61066
rect 36024 61052 36832 61066
rect 36982 61052 37122 61066
rect 37272 61052 38080 61066
rect 38230 61052 38370 61066
rect 38520 61052 39328 61066
rect 39478 61052 39618 61066
rect 39768 61052 40576 61066
rect 40726 61052 40866 61066
rect 41016 61052 41824 61066
rect 41974 61052 42114 61066
rect 42264 61052 43072 61066
rect 43222 61052 43362 61066
rect 43512 61052 44320 61066
rect 44470 61052 44610 61066
rect 44760 61052 45568 61066
rect 45718 61052 45858 61066
rect 46008 61052 46816 61066
rect 46966 61052 47106 61066
rect 47256 61052 48064 61066
rect 48214 61052 48354 61066
rect 48504 61052 49312 61066
rect 49462 61052 49602 61066
rect 49752 61052 50560 61066
rect 50710 61052 50850 61066
rect 51000 61052 51808 61066
rect 51958 61052 52098 61066
rect 52248 61052 53056 61066
rect 53206 61052 53346 61066
rect 53496 61052 54304 61066
rect 54454 61052 54594 61066
rect 54744 61052 55552 61066
rect 55702 61052 55842 61066
rect 55992 61052 56800 61066
rect 56950 61052 57090 61066
rect 57240 61052 58048 61066
rect 58198 61052 58338 61066
rect 58488 61052 58934 61066
rect 16898 61004 16980 61018
rect 17188 61004 17270 61018
rect 18146 61004 18228 61018
rect 18436 61004 18518 61018
rect 19394 61004 19476 61018
rect 19684 61004 19766 61018
rect 20642 61004 20724 61018
rect 20932 61004 21014 61018
rect 21890 61004 21972 61018
rect 22180 61004 22262 61018
rect 23138 61004 23220 61018
rect 23428 61004 23510 61018
rect 24386 61004 24468 61018
rect 24676 61004 24758 61018
rect 25634 61004 25716 61018
rect 25924 61004 26006 61018
rect 26882 61004 26964 61018
rect 27172 61004 27254 61018
rect 28130 61004 28212 61018
rect 28420 61004 28502 61018
rect 29378 61004 29460 61018
rect 29668 61004 29750 61018
rect 30626 61004 30708 61018
rect 30916 61004 30998 61018
rect 31874 61004 31956 61018
rect 32164 61004 32246 61018
rect 33122 61004 33204 61018
rect 33412 61004 33494 61018
rect 34370 61004 34452 61018
rect 34660 61004 34742 61018
rect 35618 61004 35700 61018
rect 35908 61004 35990 61018
rect 36866 61004 36948 61018
rect 37156 61004 37238 61018
rect 38114 61004 38196 61018
rect 38404 61004 38486 61018
rect 39362 61004 39444 61018
rect 39652 61004 39734 61018
rect 40610 61004 40692 61018
rect 40900 61004 40982 61018
rect 41858 61004 41940 61018
rect 42148 61004 42230 61018
rect 43106 61004 43188 61018
rect 43396 61004 43478 61018
rect 44354 61004 44436 61018
rect 44644 61004 44726 61018
rect 45602 61004 45684 61018
rect 45892 61004 45974 61018
rect 46850 61004 46932 61018
rect 47140 61004 47222 61018
rect 48098 61004 48180 61018
rect 48388 61004 48470 61018
rect 49346 61004 49428 61018
rect 49636 61004 49718 61018
rect 50594 61004 50676 61018
rect 50884 61004 50966 61018
rect 51842 61004 51924 61018
rect 52132 61004 52214 61018
rect 53090 61004 53172 61018
rect 53380 61004 53462 61018
rect 54338 61004 54420 61018
rect 54628 61004 54710 61018
rect 55586 61004 55668 61018
rect 55876 61004 55958 61018
rect 56834 61004 56916 61018
rect 57124 61004 57206 61018
rect 58082 61004 58164 61018
rect 58372 61004 58454 61018
rect 16418 60956 58934 61004
rect 16418 60798 58934 60908
rect 16418 60702 58934 60750
rect 16898 60688 16980 60702
rect 17188 60688 17270 60702
rect 18146 60688 18228 60702
rect 18436 60688 18518 60702
rect 19394 60688 19476 60702
rect 19684 60688 19766 60702
rect 20642 60688 20724 60702
rect 20932 60688 21014 60702
rect 21890 60688 21972 60702
rect 22180 60688 22262 60702
rect 23138 60688 23220 60702
rect 23428 60688 23510 60702
rect 24386 60688 24468 60702
rect 24676 60688 24758 60702
rect 25634 60688 25716 60702
rect 25924 60688 26006 60702
rect 26882 60688 26964 60702
rect 27172 60688 27254 60702
rect 28130 60688 28212 60702
rect 28420 60688 28502 60702
rect 29378 60688 29460 60702
rect 29668 60688 29750 60702
rect 30626 60688 30708 60702
rect 30916 60688 30998 60702
rect 31874 60688 31956 60702
rect 32164 60688 32246 60702
rect 33122 60688 33204 60702
rect 33412 60688 33494 60702
rect 34370 60688 34452 60702
rect 34660 60688 34742 60702
rect 35618 60688 35700 60702
rect 35908 60688 35990 60702
rect 36866 60688 36948 60702
rect 37156 60688 37238 60702
rect 38114 60688 38196 60702
rect 38404 60688 38486 60702
rect 39362 60688 39444 60702
rect 39652 60688 39734 60702
rect 40610 60688 40692 60702
rect 40900 60688 40982 60702
rect 41858 60688 41940 60702
rect 42148 60688 42230 60702
rect 43106 60688 43188 60702
rect 43396 60688 43478 60702
rect 44354 60688 44436 60702
rect 44644 60688 44726 60702
rect 45602 60688 45684 60702
rect 45892 60688 45974 60702
rect 46850 60688 46932 60702
rect 47140 60688 47222 60702
rect 48098 60688 48180 60702
rect 48388 60688 48470 60702
rect 49346 60688 49428 60702
rect 49636 60688 49718 60702
rect 50594 60688 50676 60702
rect 50884 60688 50966 60702
rect 51842 60688 51924 60702
rect 52132 60688 52214 60702
rect 53090 60688 53172 60702
rect 53380 60688 53462 60702
rect 54338 60688 54420 60702
rect 54628 60688 54710 60702
rect 55586 60688 55668 60702
rect 55876 60688 55958 60702
rect 56834 60688 56916 60702
rect 57124 60688 57206 60702
rect 58082 60688 58164 60702
rect 58372 60688 58454 60702
rect 16418 60640 16864 60654
rect 17014 60640 17154 60654
rect 17304 60640 18112 60654
rect 18262 60640 18402 60654
rect 18552 60640 19360 60654
rect 19510 60640 19650 60654
rect 19800 60640 20608 60654
rect 20758 60640 20898 60654
rect 21048 60640 21856 60654
rect 22006 60640 22146 60654
rect 22296 60640 23104 60654
rect 23254 60640 23394 60654
rect 23544 60640 24352 60654
rect 24502 60640 24642 60654
rect 24792 60640 25600 60654
rect 25750 60640 25890 60654
rect 26040 60640 26848 60654
rect 26998 60640 27138 60654
rect 27288 60640 28096 60654
rect 28246 60640 28386 60654
rect 28536 60640 29344 60654
rect 29494 60640 29634 60654
rect 29784 60640 30592 60654
rect 30742 60640 30882 60654
rect 31032 60640 31840 60654
rect 31990 60640 32130 60654
rect 32280 60640 33088 60654
rect 33238 60640 33378 60654
rect 33528 60640 34336 60654
rect 34486 60640 34626 60654
rect 34776 60640 35584 60654
rect 35734 60640 35874 60654
rect 36024 60640 36832 60654
rect 36982 60640 37122 60654
rect 37272 60640 38080 60654
rect 38230 60640 38370 60654
rect 38520 60640 39328 60654
rect 39478 60640 39618 60654
rect 39768 60640 40576 60654
rect 40726 60640 40866 60654
rect 41016 60640 41824 60654
rect 41974 60640 42114 60654
rect 42264 60640 43072 60654
rect 43222 60640 43362 60654
rect 43512 60640 44320 60654
rect 44470 60640 44610 60654
rect 44760 60640 45568 60654
rect 45718 60640 45858 60654
rect 46008 60640 46816 60654
rect 46966 60640 47106 60654
rect 47256 60640 48064 60654
rect 48214 60640 48354 60654
rect 48504 60640 49312 60654
rect 49462 60640 49602 60654
rect 49752 60640 50560 60654
rect 50710 60640 50850 60654
rect 51000 60640 51808 60654
rect 51958 60640 52098 60654
rect 52248 60640 53056 60654
rect 53206 60640 53346 60654
rect 53496 60640 54304 60654
rect 54454 60640 54594 60654
rect 54744 60640 55552 60654
rect 55702 60640 55842 60654
rect 55992 60640 56800 60654
rect 56950 60640 57090 60654
rect 57240 60640 58048 60654
rect 58198 60640 58338 60654
rect 58488 60640 58934 60654
rect 16418 60592 58934 60640
rect 16418 60578 16864 60592
rect 17014 60578 17154 60592
rect 17304 60578 18112 60592
rect 18262 60578 18402 60592
rect 18552 60578 19360 60592
rect 19510 60578 19650 60592
rect 19800 60578 20608 60592
rect 20758 60578 20898 60592
rect 21048 60578 21856 60592
rect 22006 60578 22146 60592
rect 22296 60578 23104 60592
rect 23254 60578 23394 60592
rect 23544 60578 24352 60592
rect 24502 60578 24642 60592
rect 24792 60578 25600 60592
rect 25750 60578 25890 60592
rect 26040 60578 26848 60592
rect 26998 60578 27138 60592
rect 27288 60578 28096 60592
rect 28246 60578 28386 60592
rect 28536 60578 29344 60592
rect 29494 60578 29634 60592
rect 29784 60578 30592 60592
rect 30742 60578 30882 60592
rect 31032 60578 31840 60592
rect 31990 60578 32130 60592
rect 32280 60578 33088 60592
rect 33238 60578 33378 60592
rect 33528 60578 34336 60592
rect 34486 60578 34626 60592
rect 34776 60578 35584 60592
rect 35734 60578 35874 60592
rect 36024 60578 36832 60592
rect 36982 60578 37122 60592
rect 37272 60578 38080 60592
rect 38230 60578 38370 60592
rect 38520 60578 39328 60592
rect 39478 60578 39618 60592
rect 39768 60578 40576 60592
rect 40726 60578 40866 60592
rect 41016 60578 41824 60592
rect 41974 60578 42114 60592
rect 42264 60578 43072 60592
rect 43222 60578 43362 60592
rect 43512 60578 44320 60592
rect 44470 60578 44610 60592
rect 44760 60578 45568 60592
rect 45718 60578 45858 60592
rect 46008 60578 46816 60592
rect 46966 60578 47106 60592
rect 47256 60578 48064 60592
rect 48214 60578 48354 60592
rect 48504 60578 49312 60592
rect 49462 60578 49602 60592
rect 49752 60578 50560 60592
rect 50710 60578 50850 60592
rect 51000 60578 51808 60592
rect 51958 60578 52098 60592
rect 52248 60578 53056 60592
rect 53206 60578 53346 60592
rect 53496 60578 54304 60592
rect 54454 60578 54594 60592
rect 54744 60578 55552 60592
rect 55702 60578 55842 60592
rect 55992 60578 56800 60592
rect 56950 60578 57090 60592
rect 57240 60578 58048 60592
rect 58198 60578 58338 60592
rect 58488 60578 58934 60592
rect 16898 60530 16980 60544
rect 17188 60530 17270 60544
rect 18146 60530 18228 60544
rect 18436 60530 18518 60544
rect 19394 60530 19476 60544
rect 19684 60530 19766 60544
rect 20642 60530 20724 60544
rect 20932 60530 21014 60544
rect 21890 60530 21972 60544
rect 22180 60530 22262 60544
rect 23138 60530 23220 60544
rect 23428 60530 23510 60544
rect 24386 60530 24468 60544
rect 24676 60530 24758 60544
rect 25634 60530 25716 60544
rect 25924 60530 26006 60544
rect 26882 60530 26964 60544
rect 27172 60530 27254 60544
rect 28130 60530 28212 60544
rect 28420 60530 28502 60544
rect 29378 60530 29460 60544
rect 29668 60530 29750 60544
rect 30626 60530 30708 60544
rect 30916 60530 30998 60544
rect 31874 60530 31956 60544
rect 32164 60530 32246 60544
rect 33122 60530 33204 60544
rect 33412 60530 33494 60544
rect 34370 60530 34452 60544
rect 34660 60530 34742 60544
rect 35618 60530 35700 60544
rect 35908 60530 35990 60544
rect 36866 60530 36948 60544
rect 37156 60530 37238 60544
rect 38114 60530 38196 60544
rect 38404 60530 38486 60544
rect 39362 60530 39444 60544
rect 39652 60530 39734 60544
rect 40610 60530 40692 60544
rect 40900 60530 40982 60544
rect 41858 60530 41940 60544
rect 42148 60530 42230 60544
rect 43106 60530 43188 60544
rect 43396 60530 43478 60544
rect 44354 60530 44436 60544
rect 44644 60530 44726 60544
rect 45602 60530 45684 60544
rect 45892 60530 45974 60544
rect 46850 60530 46932 60544
rect 47140 60530 47222 60544
rect 48098 60530 48180 60544
rect 48388 60530 48470 60544
rect 49346 60530 49428 60544
rect 49636 60530 49718 60544
rect 50594 60530 50676 60544
rect 50884 60530 50966 60544
rect 51842 60530 51924 60544
rect 52132 60530 52214 60544
rect 53090 60530 53172 60544
rect 53380 60530 53462 60544
rect 54338 60530 54420 60544
rect 54628 60530 54710 60544
rect 55586 60530 55668 60544
rect 55876 60530 55958 60544
rect 56834 60530 56916 60544
rect 57124 60530 57206 60544
rect 58082 60530 58164 60544
rect 58372 60530 58454 60544
rect 16418 60482 58934 60530
rect 16418 60386 58934 60434
rect 16898 60372 16980 60386
rect 17188 60372 17270 60386
rect 18146 60372 18228 60386
rect 18436 60372 18518 60386
rect 19394 60372 19476 60386
rect 19684 60372 19766 60386
rect 20642 60372 20724 60386
rect 20932 60372 21014 60386
rect 21890 60372 21972 60386
rect 22180 60372 22262 60386
rect 23138 60372 23220 60386
rect 23428 60372 23510 60386
rect 24386 60372 24468 60386
rect 24676 60372 24758 60386
rect 25634 60372 25716 60386
rect 25924 60372 26006 60386
rect 26882 60372 26964 60386
rect 27172 60372 27254 60386
rect 28130 60372 28212 60386
rect 28420 60372 28502 60386
rect 29378 60372 29460 60386
rect 29668 60372 29750 60386
rect 30626 60372 30708 60386
rect 30916 60372 30998 60386
rect 31874 60372 31956 60386
rect 32164 60372 32246 60386
rect 33122 60372 33204 60386
rect 33412 60372 33494 60386
rect 34370 60372 34452 60386
rect 34660 60372 34742 60386
rect 35618 60372 35700 60386
rect 35908 60372 35990 60386
rect 36866 60372 36948 60386
rect 37156 60372 37238 60386
rect 38114 60372 38196 60386
rect 38404 60372 38486 60386
rect 39362 60372 39444 60386
rect 39652 60372 39734 60386
rect 40610 60372 40692 60386
rect 40900 60372 40982 60386
rect 41858 60372 41940 60386
rect 42148 60372 42230 60386
rect 43106 60372 43188 60386
rect 43396 60372 43478 60386
rect 44354 60372 44436 60386
rect 44644 60372 44726 60386
rect 45602 60372 45684 60386
rect 45892 60372 45974 60386
rect 46850 60372 46932 60386
rect 47140 60372 47222 60386
rect 48098 60372 48180 60386
rect 48388 60372 48470 60386
rect 49346 60372 49428 60386
rect 49636 60372 49718 60386
rect 50594 60372 50676 60386
rect 50884 60372 50966 60386
rect 51842 60372 51924 60386
rect 52132 60372 52214 60386
rect 53090 60372 53172 60386
rect 53380 60372 53462 60386
rect 54338 60372 54420 60386
rect 54628 60372 54710 60386
rect 55586 60372 55668 60386
rect 55876 60372 55958 60386
rect 56834 60372 56916 60386
rect 57124 60372 57206 60386
rect 58082 60372 58164 60386
rect 58372 60372 58454 60386
rect 16418 60324 16864 60338
rect 17014 60324 17154 60338
rect 17304 60324 18112 60338
rect 18262 60324 18402 60338
rect 18552 60324 19360 60338
rect 19510 60324 19650 60338
rect 19800 60324 20608 60338
rect 20758 60324 20898 60338
rect 21048 60324 21856 60338
rect 22006 60324 22146 60338
rect 22296 60324 23104 60338
rect 23254 60324 23394 60338
rect 23544 60324 24352 60338
rect 24502 60324 24642 60338
rect 24792 60324 25600 60338
rect 25750 60324 25890 60338
rect 26040 60324 26848 60338
rect 26998 60324 27138 60338
rect 27288 60324 28096 60338
rect 28246 60324 28386 60338
rect 28536 60324 29344 60338
rect 29494 60324 29634 60338
rect 29784 60324 30592 60338
rect 30742 60324 30882 60338
rect 31032 60324 31840 60338
rect 31990 60324 32130 60338
rect 32280 60324 33088 60338
rect 33238 60324 33378 60338
rect 33528 60324 34336 60338
rect 34486 60324 34626 60338
rect 34776 60324 35584 60338
rect 35734 60324 35874 60338
rect 36024 60324 36832 60338
rect 36982 60324 37122 60338
rect 37272 60324 38080 60338
rect 38230 60324 38370 60338
rect 38520 60324 39328 60338
rect 39478 60324 39618 60338
rect 39768 60324 40576 60338
rect 40726 60324 40866 60338
rect 41016 60324 41824 60338
rect 41974 60324 42114 60338
rect 42264 60324 43072 60338
rect 43222 60324 43362 60338
rect 43512 60324 44320 60338
rect 44470 60324 44610 60338
rect 44760 60324 45568 60338
rect 45718 60324 45858 60338
rect 46008 60324 46816 60338
rect 46966 60324 47106 60338
rect 47256 60324 48064 60338
rect 48214 60324 48354 60338
rect 48504 60324 49312 60338
rect 49462 60324 49602 60338
rect 49752 60324 50560 60338
rect 50710 60324 50850 60338
rect 51000 60324 51808 60338
rect 51958 60324 52098 60338
rect 52248 60324 53056 60338
rect 53206 60324 53346 60338
rect 53496 60324 54304 60338
rect 54454 60324 54594 60338
rect 54744 60324 55552 60338
rect 55702 60324 55842 60338
rect 55992 60324 56800 60338
rect 56950 60324 57090 60338
rect 57240 60324 58048 60338
rect 58198 60324 58338 60338
rect 58488 60324 58934 60338
rect 16418 60276 58934 60324
rect 16418 60262 16864 60276
rect 17014 60262 17154 60276
rect 17304 60262 18112 60276
rect 18262 60262 18402 60276
rect 18552 60262 19360 60276
rect 19510 60262 19650 60276
rect 19800 60262 20608 60276
rect 20758 60262 20898 60276
rect 21048 60262 21856 60276
rect 22006 60262 22146 60276
rect 22296 60262 23104 60276
rect 23254 60262 23394 60276
rect 23544 60262 24352 60276
rect 24502 60262 24642 60276
rect 24792 60262 25600 60276
rect 25750 60262 25890 60276
rect 26040 60262 26848 60276
rect 26998 60262 27138 60276
rect 27288 60262 28096 60276
rect 28246 60262 28386 60276
rect 28536 60262 29344 60276
rect 29494 60262 29634 60276
rect 29784 60262 30592 60276
rect 30742 60262 30882 60276
rect 31032 60262 31840 60276
rect 31990 60262 32130 60276
rect 32280 60262 33088 60276
rect 33238 60262 33378 60276
rect 33528 60262 34336 60276
rect 34486 60262 34626 60276
rect 34776 60262 35584 60276
rect 35734 60262 35874 60276
rect 36024 60262 36832 60276
rect 36982 60262 37122 60276
rect 37272 60262 38080 60276
rect 38230 60262 38370 60276
rect 38520 60262 39328 60276
rect 39478 60262 39618 60276
rect 39768 60262 40576 60276
rect 40726 60262 40866 60276
rect 41016 60262 41824 60276
rect 41974 60262 42114 60276
rect 42264 60262 43072 60276
rect 43222 60262 43362 60276
rect 43512 60262 44320 60276
rect 44470 60262 44610 60276
rect 44760 60262 45568 60276
rect 45718 60262 45858 60276
rect 46008 60262 46816 60276
rect 46966 60262 47106 60276
rect 47256 60262 48064 60276
rect 48214 60262 48354 60276
rect 48504 60262 49312 60276
rect 49462 60262 49602 60276
rect 49752 60262 50560 60276
rect 50710 60262 50850 60276
rect 51000 60262 51808 60276
rect 51958 60262 52098 60276
rect 52248 60262 53056 60276
rect 53206 60262 53346 60276
rect 53496 60262 54304 60276
rect 54454 60262 54594 60276
rect 54744 60262 55552 60276
rect 55702 60262 55842 60276
rect 55992 60262 56800 60276
rect 56950 60262 57090 60276
rect 57240 60262 58048 60276
rect 58198 60262 58338 60276
rect 58488 60262 58934 60276
rect 16898 60214 16980 60228
rect 17188 60214 17270 60228
rect 18146 60214 18228 60228
rect 18436 60214 18518 60228
rect 19394 60214 19476 60228
rect 19684 60214 19766 60228
rect 20642 60214 20724 60228
rect 20932 60214 21014 60228
rect 21890 60214 21972 60228
rect 22180 60214 22262 60228
rect 23138 60214 23220 60228
rect 23428 60214 23510 60228
rect 24386 60214 24468 60228
rect 24676 60214 24758 60228
rect 25634 60214 25716 60228
rect 25924 60214 26006 60228
rect 26882 60214 26964 60228
rect 27172 60214 27254 60228
rect 28130 60214 28212 60228
rect 28420 60214 28502 60228
rect 29378 60214 29460 60228
rect 29668 60214 29750 60228
rect 30626 60214 30708 60228
rect 30916 60214 30998 60228
rect 31874 60214 31956 60228
rect 32164 60214 32246 60228
rect 33122 60214 33204 60228
rect 33412 60214 33494 60228
rect 34370 60214 34452 60228
rect 34660 60214 34742 60228
rect 35618 60214 35700 60228
rect 35908 60214 35990 60228
rect 36866 60214 36948 60228
rect 37156 60214 37238 60228
rect 38114 60214 38196 60228
rect 38404 60214 38486 60228
rect 39362 60214 39444 60228
rect 39652 60214 39734 60228
rect 40610 60214 40692 60228
rect 40900 60214 40982 60228
rect 41858 60214 41940 60228
rect 42148 60214 42230 60228
rect 43106 60214 43188 60228
rect 43396 60214 43478 60228
rect 44354 60214 44436 60228
rect 44644 60214 44726 60228
rect 45602 60214 45684 60228
rect 45892 60214 45974 60228
rect 46850 60214 46932 60228
rect 47140 60214 47222 60228
rect 48098 60214 48180 60228
rect 48388 60214 48470 60228
rect 49346 60214 49428 60228
rect 49636 60214 49718 60228
rect 50594 60214 50676 60228
rect 50884 60214 50966 60228
rect 51842 60214 51924 60228
rect 52132 60214 52214 60228
rect 53090 60214 53172 60228
rect 53380 60214 53462 60228
rect 54338 60214 54420 60228
rect 54628 60214 54710 60228
rect 55586 60214 55668 60228
rect 55876 60214 55958 60228
rect 56834 60214 56916 60228
rect 57124 60214 57206 60228
rect 58082 60214 58164 60228
rect 58372 60214 58454 60228
rect 16418 60166 58934 60214
rect 16418 60008 58934 60118
rect 16418 59912 58934 59960
rect 16898 59898 16980 59912
rect 17188 59898 17270 59912
rect 18146 59898 18228 59912
rect 18436 59898 18518 59912
rect 19394 59898 19476 59912
rect 19684 59898 19766 59912
rect 20642 59898 20724 59912
rect 20932 59898 21014 59912
rect 21890 59898 21972 59912
rect 22180 59898 22262 59912
rect 23138 59898 23220 59912
rect 23428 59898 23510 59912
rect 24386 59898 24468 59912
rect 24676 59898 24758 59912
rect 25634 59898 25716 59912
rect 25924 59898 26006 59912
rect 26882 59898 26964 59912
rect 27172 59898 27254 59912
rect 28130 59898 28212 59912
rect 28420 59898 28502 59912
rect 29378 59898 29460 59912
rect 29668 59898 29750 59912
rect 30626 59898 30708 59912
rect 30916 59898 30998 59912
rect 31874 59898 31956 59912
rect 32164 59898 32246 59912
rect 33122 59898 33204 59912
rect 33412 59898 33494 59912
rect 34370 59898 34452 59912
rect 34660 59898 34742 59912
rect 35618 59898 35700 59912
rect 35908 59898 35990 59912
rect 36866 59898 36948 59912
rect 37156 59898 37238 59912
rect 38114 59898 38196 59912
rect 38404 59898 38486 59912
rect 39362 59898 39444 59912
rect 39652 59898 39734 59912
rect 40610 59898 40692 59912
rect 40900 59898 40982 59912
rect 41858 59898 41940 59912
rect 42148 59898 42230 59912
rect 43106 59898 43188 59912
rect 43396 59898 43478 59912
rect 44354 59898 44436 59912
rect 44644 59898 44726 59912
rect 45602 59898 45684 59912
rect 45892 59898 45974 59912
rect 46850 59898 46932 59912
rect 47140 59898 47222 59912
rect 48098 59898 48180 59912
rect 48388 59898 48470 59912
rect 49346 59898 49428 59912
rect 49636 59898 49718 59912
rect 50594 59898 50676 59912
rect 50884 59898 50966 59912
rect 51842 59898 51924 59912
rect 52132 59898 52214 59912
rect 53090 59898 53172 59912
rect 53380 59898 53462 59912
rect 54338 59898 54420 59912
rect 54628 59898 54710 59912
rect 55586 59898 55668 59912
rect 55876 59898 55958 59912
rect 56834 59898 56916 59912
rect 57124 59898 57206 59912
rect 58082 59898 58164 59912
rect 58372 59898 58454 59912
rect 16418 59850 16864 59864
rect 17014 59850 17154 59864
rect 17304 59850 18112 59864
rect 18262 59850 18402 59864
rect 18552 59850 19360 59864
rect 19510 59850 19650 59864
rect 19800 59850 20608 59864
rect 20758 59850 20898 59864
rect 21048 59850 21856 59864
rect 22006 59850 22146 59864
rect 22296 59850 23104 59864
rect 23254 59850 23394 59864
rect 23544 59850 24352 59864
rect 24502 59850 24642 59864
rect 24792 59850 25600 59864
rect 25750 59850 25890 59864
rect 26040 59850 26848 59864
rect 26998 59850 27138 59864
rect 27288 59850 28096 59864
rect 28246 59850 28386 59864
rect 28536 59850 29344 59864
rect 29494 59850 29634 59864
rect 29784 59850 30592 59864
rect 30742 59850 30882 59864
rect 31032 59850 31840 59864
rect 31990 59850 32130 59864
rect 32280 59850 33088 59864
rect 33238 59850 33378 59864
rect 33528 59850 34336 59864
rect 34486 59850 34626 59864
rect 34776 59850 35584 59864
rect 35734 59850 35874 59864
rect 36024 59850 36832 59864
rect 36982 59850 37122 59864
rect 37272 59850 38080 59864
rect 38230 59850 38370 59864
rect 38520 59850 39328 59864
rect 39478 59850 39618 59864
rect 39768 59850 40576 59864
rect 40726 59850 40866 59864
rect 41016 59850 41824 59864
rect 41974 59850 42114 59864
rect 42264 59850 43072 59864
rect 43222 59850 43362 59864
rect 43512 59850 44320 59864
rect 44470 59850 44610 59864
rect 44760 59850 45568 59864
rect 45718 59850 45858 59864
rect 46008 59850 46816 59864
rect 46966 59850 47106 59864
rect 47256 59850 48064 59864
rect 48214 59850 48354 59864
rect 48504 59850 49312 59864
rect 49462 59850 49602 59864
rect 49752 59850 50560 59864
rect 50710 59850 50850 59864
rect 51000 59850 51808 59864
rect 51958 59850 52098 59864
rect 52248 59850 53056 59864
rect 53206 59850 53346 59864
rect 53496 59850 54304 59864
rect 54454 59850 54594 59864
rect 54744 59850 55552 59864
rect 55702 59850 55842 59864
rect 55992 59850 56800 59864
rect 56950 59850 57090 59864
rect 57240 59850 58048 59864
rect 58198 59850 58338 59864
rect 58488 59850 58934 59864
rect 16418 59802 58934 59850
rect 16418 59788 16864 59802
rect 17014 59788 17154 59802
rect 17304 59788 18112 59802
rect 18262 59788 18402 59802
rect 18552 59788 19360 59802
rect 19510 59788 19650 59802
rect 19800 59788 20608 59802
rect 20758 59788 20898 59802
rect 21048 59788 21856 59802
rect 22006 59788 22146 59802
rect 22296 59788 23104 59802
rect 23254 59788 23394 59802
rect 23544 59788 24352 59802
rect 24502 59788 24642 59802
rect 24792 59788 25600 59802
rect 25750 59788 25890 59802
rect 26040 59788 26848 59802
rect 26998 59788 27138 59802
rect 27288 59788 28096 59802
rect 28246 59788 28386 59802
rect 28536 59788 29344 59802
rect 29494 59788 29634 59802
rect 29784 59788 30592 59802
rect 30742 59788 30882 59802
rect 31032 59788 31840 59802
rect 31990 59788 32130 59802
rect 32280 59788 33088 59802
rect 33238 59788 33378 59802
rect 33528 59788 34336 59802
rect 34486 59788 34626 59802
rect 34776 59788 35584 59802
rect 35734 59788 35874 59802
rect 36024 59788 36832 59802
rect 36982 59788 37122 59802
rect 37272 59788 38080 59802
rect 38230 59788 38370 59802
rect 38520 59788 39328 59802
rect 39478 59788 39618 59802
rect 39768 59788 40576 59802
rect 40726 59788 40866 59802
rect 41016 59788 41824 59802
rect 41974 59788 42114 59802
rect 42264 59788 43072 59802
rect 43222 59788 43362 59802
rect 43512 59788 44320 59802
rect 44470 59788 44610 59802
rect 44760 59788 45568 59802
rect 45718 59788 45858 59802
rect 46008 59788 46816 59802
rect 46966 59788 47106 59802
rect 47256 59788 48064 59802
rect 48214 59788 48354 59802
rect 48504 59788 49312 59802
rect 49462 59788 49602 59802
rect 49752 59788 50560 59802
rect 50710 59788 50850 59802
rect 51000 59788 51808 59802
rect 51958 59788 52098 59802
rect 52248 59788 53056 59802
rect 53206 59788 53346 59802
rect 53496 59788 54304 59802
rect 54454 59788 54594 59802
rect 54744 59788 55552 59802
rect 55702 59788 55842 59802
rect 55992 59788 56800 59802
rect 56950 59788 57090 59802
rect 57240 59788 58048 59802
rect 58198 59788 58338 59802
rect 58488 59788 58934 59802
rect 16898 59740 16980 59754
rect 17188 59740 17270 59754
rect 18146 59740 18228 59754
rect 18436 59740 18518 59754
rect 19394 59740 19476 59754
rect 19684 59740 19766 59754
rect 20642 59740 20724 59754
rect 20932 59740 21014 59754
rect 21890 59740 21972 59754
rect 22180 59740 22262 59754
rect 23138 59740 23220 59754
rect 23428 59740 23510 59754
rect 24386 59740 24468 59754
rect 24676 59740 24758 59754
rect 25634 59740 25716 59754
rect 25924 59740 26006 59754
rect 26882 59740 26964 59754
rect 27172 59740 27254 59754
rect 28130 59740 28212 59754
rect 28420 59740 28502 59754
rect 29378 59740 29460 59754
rect 29668 59740 29750 59754
rect 30626 59740 30708 59754
rect 30916 59740 30998 59754
rect 31874 59740 31956 59754
rect 32164 59740 32246 59754
rect 33122 59740 33204 59754
rect 33412 59740 33494 59754
rect 34370 59740 34452 59754
rect 34660 59740 34742 59754
rect 35618 59740 35700 59754
rect 35908 59740 35990 59754
rect 36866 59740 36948 59754
rect 37156 59740 37238 59754
rect 38114 59740 38196 59754
rect 38404 59740 38486 59754
rect 39362 59740 39444 59754
rect 39652 59740 39734 59754
rect 40610 59740 40692 59754
rect 40900 59740 40982 59754
rect 41858 59740 41940 59754
rect 42148 59740 42230 59754
rect 43106 59740 43188 59754
rect 43396 59740 43478 59754
rect 44354 59740 44436 59754
rect 44644 59740 44726 59754
rect 45602 59740 45684 59754
rect 45892 59740 45974 59754
rect 46850 59740 46932 59754
rect 47140 59740 47222 59754
rect 48098 59740 48180 59754
rect 48388 59740 48470 59754
rect 49346 59740 49428 59754
rect 49636 59740 49718 59754
rect 50594 59740 50676 59754
rect 50884 59740 50966 59754
rect 51842 59740 51924 59754
rect 52132 59740 52214 59754
rect 53090 59740 53172 59754
rect 53380 59740 53462 59754
rect 54338 59740 54420 59754
rect 54628 59740 54710 59754
rect 55586 59740 55668 59754
rect 55876 59740 55958 59754
rect 56834 59740 56916 59754
rect 57124 59740 57206 59754
rect 58082 59740 58164 59754
rect 58372 59740 58454 59754
rect 16418 59692 58934 59740
rect 16418 59596 58934 59644
rect 16898 59582 16980 59596
rect 17188 59582 17270 59596
rect 18146 59582 18228 59596
rect 18436 59582 18518 59596
rect 19394 59582 19476 59596
rect 19684 59582 19766 59596
rect 20642 59582 20724 59596
rect 20932 59582 21014 59596
rect 21890 59582 21972 59596
rect 22180 59582 22262 59596
rect 23138 59582 23220 59596
rect 23428 59582 23510 59596
rect 24386 59582 24468 59596
rect 24676 59582 24758 59596
rect 25634 59582 25716 59596
rect 25924 59582 26006 59596
rect 26882 59582 26964 59596
rect 27172 59582 27254 59596
rect 28130 59582 28212 59596
rect 28420 59582 28502 59596
rect 29378 59582 29460 59596
rect 29668 59582 29750 59596
rect 30626 59582 30708 59596
rect 30916 59582 30998 59596
rect 31874 59582 31956 59596
rect 32164 59582 32246 59596
rect 33122 59582 33204 59596
rect 33412 59582 33494 59596
rect 34370 59582 34452 59596
rect 34660 59582 34742 59596
rect 35618 59582 35700 59596
rect 35908 59582 35990 59596
rect 36866 59582 36948 59596
rect 37156 59582 37238 59596
rect 38114 59582 38196 59596
rect 38404 59582 38486 59596
rect 39362 59582 39444 59596
rect 39652 59582 39734 59596
rect 40610 59582 40692 59596
rect 40900 59582 40982 59596
rect 41858 59582 41940 59596
rect 42148 59582 42230 59596
rect 43106 59582 43188 59596
rect 43396 59582 43478 59596
rect 44354 59582 44436 59596
rect 44644 59582 44726 59596
rect 45602 59582 45684 59596
rect 45892 59582 45974 59596
rect 46850 59582 46932 59596
rect 47140 59582 47222 59596
rect 48098 59582 48180 59596
rect 48388 59582 48470 59596
rect 49346 59582 49428 59596
rect 49636 59582 49718 59596
rect 50594 59582 50676 59596
rect 50884 59582 50966 59596
rect 51842 59582 51924 59596
rect 52132 59582 52214 59596
rect 53090 59582 53172 59596
rect 53380 59582 53462 59596
rect 54338 59582 54420 59596
rect 54628 59582 54710 59596
rect 55586 59582 55668 59596
rect 55876 59582 55958 59596
rect 56834 59582 56916 59596
rect 57124 59582 57206 59596
rect 58082 59582 58164 59596
rect 58372 59582 58454 59596
rect 16418 59534 16864 59548
rect 17014 59534 17154 59548
rect 17304 59534 18112 59548
rect 18262 59534 18402 59548
rect 18552 59534 19360 59548
rect 19510 59534 19650 59548
rect 19800 59534 20608 59548
rect 20758 59534 20898 59548
rect 21048 59534 21856 59548
rect 22006 59534 22146 59548
rect 22296 59534 23104 59548
rect 23254 59534 23394 59548
rect 23544 59534 24352 59548
rect 24502 59534 24642 59548
rect 24792 59534 25600 59548
rect 25750 59534 25890 59548
rect 26040 59534 26848 59548
rect 26998 59534 27138 59548
rect 27288 59534 28096 59548
rect 28246 59534 28386 59548
rect 28536 59534 29344 59548
rect 29494 59534 29634 59548
rect 29784 59534 30592 59548
rect 30742 59534 30882 59548
rect 31032 59534 31840 59548
rect 31990 59534 32130 59548
rect 32280 59534 33088 59548
rect 33238 59534 33378 59548
rect 33528 59534 34336 59548
rect 34486 59534 34626 59548
rect 34776 59534 35584 59548
rect 35734 59534 35874 59548
rect 36024 59534 36832 59548
rect 36982 59534 37122 59548
rect 37272 59534 38080 59548
rect 38230 59534 38370 59548
rect 38520 59534 39328 59548
rect 39478 59534 39618 59548
rect 39768 59534 40576 59548
rect 40726 59534 40866 59548
rect 41016 59534 41824 59548
rect 41974 59534 42114 59548
rect 42264 59534 43072 59548
rect 43222 59534 43362 59548
rect 43512 59534 44320 59548
rect 44470 59534 44610 59548
rect 44760 59534 45568 59548
rect 45718 59534 45858 59548
rect 46008 59534 46816 59548
rect 46966 59534 47106 59548
rect 47256 59534 48064 59548
rect 48214 59534 48354 59548
rect 48504 59534 49312 59548
rect 49462 59534 49602 59548
rect 49752 59534 50560 59548
rect 50710 59534 50850 59548
rect 51000 59534 51808 59548
rect 51958 59534 52098 59548
rect 52248 59534 53056 59548
rect 53206 59534 53346 59548
rect 53496 59534 54304 59548
rect 54454 59534 54594 59548
rect 54744 59534 55552 59548
rect 55702 59534 55842 59548
rect 55992 59534 56800 59548
rect 56950 59534 57090 59548
rect 57240 59534 58048 59548
rect 58198 59534 58338 59548
rect 58488 59534 58934 59548
rect 16418 59486 58934 59534
rect 16418 59472 16864 59486
rect 17014 59472 17154 59486
rect 17304 59472 18112 59486
rect 18262 59472 18402 59486
rect 18552 59472 19360 59486
rect 19510 59472 19650 59486
rect 19800 59472 20608 59486
rect 20758 59472 20898 59486
rect 21048 59472 21856 59486
rect 22006 59472 22146 59486
rect 22296 59472 23104 59486
rect 23254 59472 23394 59486
rect 23544 59472 24352 59486
rect 24502 59472 24642 59486
rect 24792 59472 25600 59486
rect 25750 59472 25890 59486
rect 26040 59472 26848 59486
rect 26998 59472 27138 59486
rect 27288 59472 28096 59486
rect 28246 59472 28386 59486
rect 28536 59472 29344 59486
rect 29494 59472 29634 59486
rect 29784 59472 30592 59486
rect 30742 59472 30882 59486
rect 31032 59472 31840 59486
rect 31990 59472 32130 59486
rect 32280 59472 33088 59486
rect 33238 59472 33378 59486
rect 33528 59472 34336 59486
rect 34486 59472 34626 59486
rect 34776 59472 35584 59486
rect 35734 59472 35874 59486
rect 36024 59472 36832 59486
rect 36982 59472 37122 59486
rect 37272 59472 38080 59486
rect 38230 59472 38370 59486
rect 38520 59472 39328 59486
rect 39478 59472 39618 59486
rect 39768 59472 40576 59486
rect 40726 59472 40866 59486
rect 41016 59472 41824 59486
rect 41974 59472 42114 59486
rect 42264 59472 43072 59486
rect 43222 59472 43362 59486
rect 43512 59472 44320 59486
rect 44470 59472 44610 59486
rect 44760 59472 45568 59486
rect 45718 59472 45858 59486
rect 46008 59472 46816 59486
rect 46966 59472 47106 59486
rect 47256 59472 48064 59486
rect 48214 59472 48354 59486
rect 48504 59472 49312 59486
rect 49462 59472 49602 59486
rect 49752 59472 50560 59486
rect 50710 59472 50850 59486
rect 51000 59472 51808 59486
rect 51958 59472 52098 59486
rect 52248 59472 53056 59486
rect 53206 59472 53346 59486
rect 53496 59472 54304 59486
rect 54454 59472 54594 59486
rect 54744 59472 55552 59486
rect 55702 59472 55842 59486
rect 55992 59472 56800 59486
rect 56950 59472 57090 59486
rect 57240 59472 58048 59486
rect 58198 59472 58338 59486
rect 58488 59472 58934 59486
rect 16898 59424 16980 59438
rect 17188 59424 17270 59438
rect 18146 59424 18228 59438
rect 18436 59424 18518 59438
rect 19394 59424 19476 59438
rect 19684 59424 19766 59438
rect 20642 59424 20724 59438
rect 20932 59424 21014 59438
rect 21890 59424 21972 59438
rect 22180 59424 22262 59438
rect 23138 59424 23220 59438
rect 23428 59424 23510 59438
rect 24386 59424 24468 59438
rect 24676 59424 24758 59438
rect 25634 59424 25716 59438
rect 25924 59424 26006 59438
rect 26882 59424 26964 59438
rect 27172 59424 27254 59438
rect 28130 59424 28212 59438
rect 28420 59424 28502 59438
rect 29378 59424 29460 59438
rect 29668 59424 29750 59438
rect 30626 59424 30708 59438
rect 30916 59424 30998 59438
rect 31874 59424 31956 59438
rect 32164 59424 32246 59438
rect 33122 59424 33204 59438
rect 33412 59424 33494 59438
rect 34370 59424 34452 59438
rect 34660 59424 34742 59438
rect 35618 59424 35700 59438
rect 35908 59424 35990 59438
rect 36866 59424 36948 59438
rect 37156 59424 37238 59438
rect 38114 59424 38196 59438
rect 38404 59424 38486 59438
rect 39362 59424 39444 59438
rect 39652 59424 39734 59438
rect 40610 59424 40692 59438
rect 40900 59424 40982 59438
rect 41858 59424 41940 59438
rect 42148 59424 42230 59438
rect 43106 59424 43188 59438
rect 43396 59424 43478 59438
rect 44354 59424 44436 59438
rect 44644 59424 44726 59438
rect 45602 59424 45684 59438
rect 45892 59424 45974 59438
rect 46850 59424 46932 59438
rect 47140 59424 47222 59438
rect 48098 59424 48180 59438
rect 48388 59424 48470 59438
rect 49346 59424 49428 59438
rect 49636 59424 49718 59438
rect 50594 59424 50676 59438
rect 50884 59424 50966 59438
rect 51842 59424 51924 59438
rect 52132 59424 52214 59438
rect 53090 59424 53172 59438
rect 53380 59424 53462 59438
rect 54338 59424 54420 59438
rect 54628 59424 54710 59438
rect 55586 59424 55668 59438
rect 55876 59424 55958 59438
rect 56834 59424 56916 59438
rect 57124 59424 57206 59438
rect 58082 59424 58164 59438
rect 58372 59424 58454 59438
rect 16418 59376 58934 59424
rect 16418 59218 58934 59328
rect 16418 59122 58934 59170
rect 16898 59108 16980 59122
rect 17188 59108 17270 59122
rect 18146 59108 18228 59122
rect 18436 59108 18518 59122
rect 19394 59108 19476 59122
rect 19684 59108 19766 59122
rect 20642 59108 20724 59122
rect 20932 59108 21014 59122
rect 21890 59108 21972 59122
rect 22180 59108 22262 59122
rect 23138 59108 23220 59122
rect 23428 59108 23510 59122
rect 24386 59108 24468 59122
rect 24676 59108 24758 59122
rect 25634 59108 25716 59122
rect 25924 59108 26006 59122
rect 26882 59108 26964 59122
rect 27172 59108 27254 59122
rect 28130 59108 28212 59122
rect 28420 59108 28502 59122
rect 29378 59108 29460 59122
rect 29668 59108 29750 59122
rect 30626 59108 30708 59122
rect 30916 59108 30998 59122
rect 31874 59108 31956 59122
rect 32164 59108 32246 59122
rect 33122 59108 33204 59122
rect 33412 59108 33494 59122
rect 34370 59108 34452 59122
rect 34660 59108 34742 59122
rect 35618 59108 35700 59122
rect 35908 59108 35990 59122
rect 36866 59108 36948 59122
rect 37156 59108 37238 59122
rect 38114 59108 38196 59122
rect 38404 59108 38486 59122
rect 39362 59108 39444 59122
rect 39652 59108 39734 59122
rect 40610 59108 40692 59122
rect 40900 59108 40982 59122
rect 41858 59108 41940 59122
rect 42148 59108 42230 59122
rect 43106 59108 43188 59122
rect 43396 59108 43478 59122
rect 44354 59108 44436 59122
rect 44644 59108 44726 59122
rect 45602 59108 45684 59122
rect 45892 59108 45974 59122
rect 46850 59108 46932 59122
rect 47140 59108 47222 59122
rect 48098 59108 48180 59122
rect 48388 59108 48470 59122
rect 49346 59108 49428 59122
rect 49636 59108 49718 59122
rect 50594 59108 50676 59122
rect 50884 59108 50966 59122
rect 51842 59108 51924 59122
rect 52132 59108 52214 59122
rect 53090 59108 53172 59122
rect 53380 59108 53462 59122
rect 54338 59108 54420 59122
rect 54628 59108 54710 59122
rect 55586 59108 55668 59122
rect 55876 59108 55958 59122
rect 56834 59108 56916 59122
rect 57124 59108 57206 59122
rect 58082 59108 58164 59122
rect 58372 59108 58454 59122
rect 16418 59060 16864 59074
rect 17014 59060 17154 59074
rect 17304 59060 18112 59074
rect 18262 59060 18402 59074
rect 18552 59060 19360 59074
rect 19510 59060 19650 59074
rect 19800 59060 20608 59074
rect 20758 59060 20898 59074
rect 21048 59060 21856 59074
rect 22006 59060 22146 59074
rect 22296 59060 23104 59074
rect 23254 59060 23394 59074
rect 23544 59060 24352 59074
rect 24502 59060 24642 59074
rect 24792 59060 25600 59074
rect 25750 59060 25890 59074
rect 26040 59060 26848 59074
rect 26998 59060 27138 59074
rect 27288 59060 28096 59074
rect 28246 59060 28386 59074
rect 28536 59060 29344 59074
rect 29494 59060 29634 59074
rect 29784 59060 30592 59074
rect 30742 59060 30882 59074
rect 31032 59060 31840 59074
rect 31990 59060 32130 59074
rect 32280 59060 33088 59074
rect 33238 59060 33378 59074
rect 33528 59060 34336 59074
rect 34486 59060 34626 59074
rect 34776 59060 35584 59074
rect 35734 59060 35874 59074
rect 36024 59060 36832 59074
rect 36982 59060 37122 59074
rect 37272 59060 38080 59074
rect 38230 59060 38370 59074
rect 38520 59060 39328 59074
rect 39478 59060 39618 59074
rect 39768 59060 40576 59074
rect 40726 59060 40866 59074
rect 41016 59060 41824 59074
rect 41974 59060 42114 59074
rect 42264 59060 43072 59074
rect 43222 59060 43362 59074
rect 43512 59060 44320 59074
rect 44470 59060 44610 59074
rect 44760 59060 45568 59074
rect 45718 59060 45858 59074
rect 46008 59060 46816 59074
rect 46966 59060 47106 59074
rect 47256 59060 48064 59074
rect 48214 59060 48354 59074
rect 48504 59060 49312 59074
rect 49462 59060 49602 59074
rect 49752 59060 50560 59074
rect 50710 59060 50850 59074
rect 51000 59060 51808 59074
rect 51958 59060 52098 59074
rect 52248 59060 53056 59074
rect 53206 59060 53346 59074
rect 53496 59060 54304 59074
rect 54454 59060 54594 59074
rect 54744 59060 55552 59074
rect 55702 59060 55842 59074
rect 55992 59060 56800 59074
rect 56950 59060 57090 59074
rect 57240 59060 58048 59074
rect 58198 59060 58338 59074
rect 58488 59060 58934 59074
rect 16418 59012 58934 59060
rect 16418 58998 16864 59012
rect 17014 58998 17154 59012
rect 17304 58998 18112 59012
rect 18262 58998 18402 59012
rect 18552 58998 19360 59012
rect 19510 58998 19650 59012
rect 19800 58998 20608 59012
rect 20758 58998 20898 59012
rect 21048 58998 21856 59012
rect 22006 58998 22146 59012
rect 22296 58998 23104 59012
rect 23254 58998 23394 59012
rect 23544 58998 24352 59012
rect 24502 58998 24642 59012
rect 24792 58998 25600 59012
rect 25750 58998 25890 59012
rect 26040 58998 26848 59012
rect 26998 58998 27138 59012
rect 27288 58998 28096 59012
rect 28246 58998 28386 59012
rect 28536 58998 29344 59012
rect 29494 58998 29634 59012
rect 29784 58998 30592 59012
rect 30742 58998 30882 59012
rect 31032 58998 31840 59012
rect 31990 58998 32130 59012
rect 32280 58998 33088 59012
rect 33238 58998 33378 59012
rect 33528 58998 34336 59012
rect 34486 58998 34626 59012
rect 34776 58998 35584 59012
rect 35734 58998 35874 59012
rect 36024 58998 36832 59012
rect 36982 58998 37122 59012
rect 37272 58998 38080 59012
rect 38230 58998 38370 59012
rect 38520 58998 39328 59012
rect 39478 58998 39618 59012
rect 39768 58998 40576 59012
rect 40726 58998 40866 59012
rect 41016 58998 41824 59012
rect 41974 58998 42114 59012
rect 42264 58998 43072 59012
rect 43222 58998 43362 59012
rect 43512 58998 44320 59012
rect 44470 58998 44610 59012
rect 44760 58998 45568 59012
rect 45718 58998 45858 59012
rect 46008 58998 46816 59012
rect 46966 58998 47106 59012
rect 47256 58998 48064 59012
rect 48214 58998 48354 59012
rect 48504 58998 49312 59012
rect 49462 58998 49602 59012
rect 49752 58998 50560 59012
rect 50710 58998 50850 59012
rect 51000 58998 51808 59012
rect 51958 58998 52098 59012
rect 52248 58998 53056 59012
rect 53206 58998 53346 59012
rect 53496 58998 54304 59012
rect 54454 58998 54594 59012
rect 54744 58998 55552 59012
rect 55702 58998 55842 59012
rect 55992 58998 56800 59012
rect 56950 58998 57090 59012
rect 57240 58998 58048 59012
rect 58198 58998 58338 59012
rect 58488 58998 58934 59012
rect 16898 58950 16980 58964
rect 17188 58950 17270 58964
rect 18146 58950 18228 58964
rect 18436 58950 18518 58964
rect 19394 58950 19476 58964
rect 19684 58950 19766 58964
rect 20642 58950 20724 58964
rect 20932 58950 21014 58964
rect 21890 58950 21972 58964
rect 22180 58950 22262 58964
rect 23138 58950 23220 58964
rect 23428 58950 23510 58964
rect 24386 58950 24468 58964
rect 24676 58950 24758 58964
rect 25634 58950 25716 58964
rect 25924 58950 26006 58964
rect 26882 58950 26964 58964
rect 27172 58950 27254 58964
rect 28130 58950 28212 58964
rect 28420 58950 28502 58964
rect 29378 58950 29460 58964
rect 29668 58950 29750 58964
rect 30626 58950 30708 58964
rect 30916 58950 30998 58964
rect 31874 58950 31956 58964
rect 32164 58950 32246 58964
rect 33122 58950 33204 58964
rect 33412 58950 33494 58964
rect 34370 58950 34452 58964
rect 34660 58950 34742 58964
rect 35618 58950 35700 58964
rect 35908 58950 35990 58964
rect 36866 58950 36948 58964
rect 37156 58950 37238 58964
rect 38114 58950 38196 58964
rect 38404 58950 38486 58964
rect 39362 58950 39444 58964
rect 39652 58950 39734 58964
rect 40610 58950 40692 58964
rect 40900 58950 40982 58964
rect 41858 58950 41940 58964
rect 42148 58950 42230 58964
rect 43106 58950 43188 58964
rect 43396 58950 43478 58964
rect 44354 58950 44436 58964
rect 44644 58950 44726 58964
rect 45602 58950 45684 58964
rect 45892 58950 45974 58964
rect 46850 58950 46932 58964
rect 47140 58950 47222 58964
rect 48098 58950 48180 58964
rect 48388 58950 48470 58964
rect 49346 58950 49428 58964
rect 49636 58950 49718 58964
rect 50594 58950 50676 58964
rect 50884 58950 50966 58964
rect 51842 58950 51924 58964
rect 52132 58950 52214 58964
rect 53090 58950 53172 58964
rect 53380 58950 53462 58964
rect 54338 58950 54420 58964
rect 54628 58950 54710 58964
rect 55586 58950 55668 58964
rect 55876 58950 55958 58964
rect 56834 58950 56916 58964
rect 57124 58950 57206 58964
rect 58082 58950 58164 58964
rect 58372 58950 58454 58964
rect 16418 58902 58934 58950
rect 16418 58806 58934 58854
rect 16898 58792 16980 58806
rect 17188 58792 17270 58806
rect 18146 58792 18228 58806
rect 18436 58792 18518 58806
rect 19394 58792 19476 58806
rect 19684 58792 19766 58806
rect 20642 58792 20724 58806
rect 20932 58792 21014 58806
rect 21890 58792 21972 58806
rect 22180 58792 22262 58806
rect 23138 58792 23220 58806
rect 23428 58792 23510 58806
rect 24386 58792 24468 58806
rect 24676 58792 24758 58806
rect 25634 58792 25716 58806
rect 25924 58792 26006 58806
rect 26882 58792 26964 58806
rect 27172 58792 27254 58806
rect 28130 58792 28212 58806
rect 28420 58792 28502 58806
rect 29378 58792 29460 58806
rect 29668 58792 29750 58806
rect 30626 58792 30708 58806
rect 30916 58792 30998 58806
rect 31874 58792 31956 58806
rect 32164 58792 32246 58806
rect 33122 58792 33204 58806
rect 33412 58792 33494 58806
rect 34370 58792 34452 58806
rect 34660 58792 34742 58806
rect 35618 58792 35700 58806
rect 35908 58792 35990 58806
rect 36866 58792 36948 58806
rect 37156 58792 37238 58806
rect 38114 58792 38196 58806
rect 38404 58792 38486 58806
rect 39362 58792 39444 58806
rect 39652 58792 39734 58806
rect 40610 58792 40692 58806
rect 40900 58792 40982 58806
rect 41858 58792 41940 58806
rect 42148 58792 42230 58806
rect 43106 58792 43188 58806
rect 43396 58792 43478 58806
rect 44354 58792 44436 58806
rect 44644 58792 44726 58806
rect 45602 58792 45684 58806
rect 45892 58792 45974 58806
rect 46850 58792 46932 58806
rect 47140 58792 47222 58806
rect 48098 58792 48180 58806
rect 48388 58792 48470 58806
rect 49346 58792 49428 58806
rect 49636 58792 49718 58806
rect 50594 58792 50676 58806
rect 50884 58792 50966 58806
rect 51842 58792 51924 58806
rect 52132 58792 52214 58806
rect 53090 58792 53172 58806
rect 53380 58792 53462 58806
rect 54338 58792 54420 58806
rect 54628 58792 54710 58806
rect 55586 58792 55668 58806
rect 55876 58792 55958 58806
rect 56834 58792 56916 58806
rect 57124 58792 57206 58806
rect 58082 58792 58164 58806
rect 58372 58792 58454 58806
rect 16418 58744 16864 58758
rect 17014 58744 17154 58758
rect 17304 58744 18112 58758
rect 18262 58744 18402 58758
rect 18552 58744 19360 58758
rect 19510 58744 19650 58758
rect 19800 58744 20608 58758
rect 20758 58744 20898 58758
rect 21048 58744 21856 58758
rect 22006 58744 22146 58758
rect 22296 58744 23104 58758
rect 23254 58744 23394 58758
rect 23544 58744 24352 58758
rect 24502 58744 24642 58758
rect 24792 58744 25600 58758
rect 25750 58744 25890 58758
rect 26040 58744 26848 58758
rect 26998 58744 27138 58758
rect 27288 58744 28096 58758
rect 28246 58744 28386 58758
rect 28536 58744 29344 58758
rect 29494 58744 29634 58758
rect 29784 58744 30592 58758
rect 30742 58744 30882 58758
rect 31032 58744 31840 58758
rect 31990 58744 32130 58758
rect 32280 58744 33088 58758
rect 33238 58744 33378 58758
rect 33528 58744 34336 58758
rect 34486 58744 34626 58758
rect 34776 58744 35584 58758
rect 35734 58744 35874 58758
rect 36024 58744 36832 58758
rect 36982 58744 37122 58758
rect 37272 58744 38080 58758
rect 38230 58744 38370 58758
rect 38520 58744 39328 58758
rect 39478 58744 39618 58758
rect 39768 58744 40576 58758
rect 40726 58744 40866 58758
rect 41016 58744 41824 58758
rect 41974 58744 42114 58758
rect 42264 58744 43072 58758
rect 43222 58744 43362 58758
rect 43512 58744 44320 58758
rect 44470 58744 44610 58758
rect 44760 58744 45568 58758
rect 45718 58744 45858 58758
rect 46008 58744 46816 58758
rect 46966 58744 47106 58758
rect 47256 58744 48064 58758
rect 48214 58744 48354 58758
rect 48504 58744 49312 58758
rect 49462 58744 49602 58758
rect 49752 58744 50560 58758
rect 50710 58744 50850 58758
rect 51000 58744 51808 58758
rect 51958 58744 52098 58758
rect 52248 58744 53056 58758
rect 53206 58744 53346 58758
rect 53496 58744 54304 58758
rect 54454 58744 54594 58758
rect 54744 58744 55552 58758
rect 55702 58744 55842 58758
rect 55992 58744 56800 58758
rect 56950 58744 57090 58758
rect 57240 58744 58048 58758
rect 58198 58744 58338 58758
rect 58488 58744 58934 58758
rect 16418 58696 58934 58744
rect 16418 58682 16864 58696
rect 17014 58682 17154 58696
rect 17304 58682 18112 58696
rect 18262 58682 18402 58696
rect 18552 58682 19360 58696
rect 19510 58682 19650 58696
rect 19800 58682 20608 58696
rect 20758 58682 20898 58696
rect 21048 58682 21856 58696
rect 22006 58682 22146 58696
rect 22296 58682 23104 58696
rect 23254 58682 23394 58696
rect 23544 58682 24352 58696
rect 24502 58682 24642 58696
rect 24792 58682 25600 58696
rect 25750 58682 25890 58696
rect 26040 58682 26848 58696
rect 26998 58682 27138 58696
rect 27288 58682 28096 58696
rect 28246 58682 28386 58696
rect 28536 58682 29344 58696
rect 29494 58682 29634 58696
rect 29784 58682 30592 58696
rect 30742 58682 30882 58696
rect 31032 58682 31840 58696
rect 31990 58682 32130 58696
rect 32280 58682 33088 58696
rect 33238 58682 33378 58696
rect 33528 58682 34336 58696
rect 34486 58682 34626 58696
rect 34776 58682 35584 58696
rect 35734 58682 35874 58696
rect 36024 58682 36832 58696
rect 36982 58682 37122 58696
rect 37272 58682 38080 58696
rect 38230 58682 38370 58696
rect 38520 58682 39328 58696
rect 39478 58682 39618 58696
rect 39768 58682 40576 58696
rect 40726 58682 40866 58696
rect 41016 58682 41824 58696
rect 41974 58682 42114 58696
rect 42264 58682 43072 58696
rect 43222 58682 43362 58696
rect 43512 58682 44320 58696
rect 44470 58682 44610 58696
rect 44760 58682 45568 58696
rect 45718 58682 45858 58696
rect 46008 58682 46816 58696
rect 46966 58682 47106 58696
rect 47256 58682 48064 58696
rect 48214 58682 48354 58696
rect 48504 58682 49312 58696
rect 49462 58682 49602 58696
rect 49752 58682 50560 58696
rect 50710 58682 50850 58696
rect 51000 58682 51808 58696
rect 51958 58682 52098 58696
rect 52248 58682 53056 58696
rect 53206 58682 53346 58696
rect 53496 58682 54304 58696
rect 54454 58682 54594 58696
rect 54744 58682 55552 58696
rect 55702 58682 55842 58696
rect 55992 58682 56800 58696
rect 56950 58682 57090 58696
rect 57240 58682 58048 58696
rect 58198 58682 58338 58696
rect 58488 58682 58934 58696
rect 16898 58634 16980 58648
rect 17188 58634 17270 58648
rect 18146 58634 18228 58648
rect 18436 58634 18518 58648
rect 19394 58634 19476 58648
rect 19684 58634 19766 58648
rect 20642 58634 20724 58648
rect 20932 58634 21014 58648
rect 21890 58634 21972 58648
rect 22180 58634 22262 58648
rect 23138 58634 23220 58648
rect 23428 58634 23510 58648
rect 24386 58634 24468 58648
rect 24676 58634 24758 58648
rect 25634 58634 25716 58648
rect 25924 58634 26006 58648
rect 26882 58634 26964 58648
rect 27172 58634 27254 58648
rect 28130 58634 28212 58648
rect 28420 58634 28502 58648
rect 29378 58634 29460 58648
rect 29668 58634 29750 58648
rect 30626 58634 30708 58648
rect 30916 58634 30998 58648
rect 31874 58634 31956 58648
rect 32164 58634 32246 58648
rect 33122 58634 33204 58648
rect 33412 58634 33494 58648
rect 34370 58634 34452 58648
rect 34660 58634 34742 58648
rect 35618 58634 35700 58648
rect 35908 58634 35990 58648
rect 36866 58634 36948 58648
rect 37156 58634 37238 58648
rect 38114 58634 38196 58648
rect 38404 58634 38486 58648
rect 39362 58634 39444 58648
rect 39652 58634 39734 58648
rect 40610 58634 40692 58648
rect 40900 58634 40982 58648
rect 41858 58634 41940 58648
rect 42148 58634 42230 58648
rect 43106 58634 43188 58648
rect 43396 58634 43478 58648
rect 44354 58634 44436 58648
rect 44644 58634 44726 58648
rect 45602 58634 45684 58648
rect 45892 58634 45974 58648
rect 46850 58634 46932 58648
rect 47140 58634 47222 58648
rect 48098 58634 48180 58648
rect 48388 58634 48470 58648
rect 49346 58634 49428 58648
rect 49636 58634 49718 58648
rect 50594 58634 50676 58648
rect 50884 58634 50966 58648
rect 51842 58634 51924 58648
rect 52132 58634 52214 58648
rect 53090 58634 53172 58648
rect 53380 58634 53462 58648
rect 54338 58634 54420 58648
rect 54628 58634 54710 58648
rect 55586 58634 55668 58648
rect 55876 58634 55958 58648
rect 56834 58634 56916 58648
rect 57124 58634 57206 58648
rect 58082 58634 58164 58648
rect 58372 58634 58454 58648
rect 16418 58586 58934 58634
rect 16418 58428 58934 58538
rect 16418 58332 58934 58380
rect 16898 58318 16980 58332
rect 17188 58318 17270 58332
rect 18146 58318 18228 58332
rect 18436 58318 18518 58332
rect 19394 58318 19476 58332
rect 19684 58318 19766 58332
rect 20642 58318 20724 58332
rect 20932 58318 21014 58332
rect 21890 58318 21972 58332
rect 22180 58318 22262 58332
rect 23138 58318 23220 58332
rect 23428 58318 23510 58332
rect 24386 58318 24468 58332
rect 24676 58318 24758 58332
rect 25634 58318 25716 58332
rect 25924 58318 26006 58332
rect 26882 58318 26964 58332
rect 27172 58318 27254 58332
rect 28130 58318 28212 58332
rect 28420 58318 28502 58332
rect 29378 58318 29460 58332
rect 29668 58318 29750 58332
rect 30626 58318 30708 58332
rect 30916 58318 30998 58332
rect 31874 58318 31956 58332
rect 32164 58318 32246 58332
rect 33122 58318 33204 58332
rect 33412 58318 33494 58332
rect 34370 58318 34452 58332
rect 34660 58318 34742 58332
rect 35618 58318 35700 58332
rect 35908 58318 35990 58332
rect 36866 58318 36948 58332
rect 37156 58318 37238 58332
rect 38114 58318 38196 58332
rect 38404 58318 38486 58332
rect 39362 58318 39444 58332
rect 39652 58318 39734 58332
rect 40610 58318 40692 58332
rect 40900 58318 40982 58332
rect 41858 58318 41940 58332
rect 42148 58318 42230 58332
rect 43106 58318 43188 58332
rect 43396 58318 43478 58332
rect 44354 58318 44436 58332
rect 44644 58318 44726 58332
rect 45602 58318 45684 58332
rect 45892 58318 45974 58332
rect 46850 58318 46932 58332
rect 47140 58318 47222 58332
rect 48098 58318 48180 58332
rect 48388 58318 48470 58332
rect 49346 58318 49428 58332
rect 49636 58318 49718 58332
rect 50594 58318 50676 58332
rect 50884 58318 50966 58332
rect 51842 58318 51924 58332
rect 52132 58318 52214 58332
rect 53090 58318 53172 58332
rect 53380 58318 53462 58332
rect 54338 58318 54420 58332
rect 54628 58318 54710 58332
rect 55586 58318 55668 58332
rect 55876 58318 55958 58332
rect 56834 58318 56916 58332
rect 57124 58318 57206 58332
rect 58082 58318 58164 58332
rect 58372 58318 58454 58332
rect 16418 58270 16864 58284
rect 17014 58270 17154 58284
rect 17304 58270 18112 58284
rect 18262 58270 18402 58284
rect 18552 58270 19360 58284
rect 19510 58270 19650 58284
rect 19800 58270 20608 58284
rect 20758 58270 20898 58284
rect 21048 58270 21856 58284
rect 22006 58270 22146 58284
rect 22296 58270 23104 58284
rect 23254 58270 23394 58284
rect 23544 58270 24352 58284
rect 24502 58270 24642 58284
rect 24792 58270 25600 58284
rect 25750 58270 25890 58284
rect 26040 58270 26848 58284
rect 26998 58270 27138 58284
rect 27288 58270 28096 58284
rect 28246 58270 28386 58284
rect 28536 58270 29344 58284
rect 29494 58270 29634 58284
rect 29784 58270 30592 58284
rect 30742 58270 30882 58284
rect 31032 58270 31840 58284
rect 31990 58270 32130 58284
rect 32280 58270 33088 58284
rect 33238 58270 33378 58284
rect 33528 58270 34336 58284
rect 34486 58270 34626 58284
rect 34776 58270 35584 58284
rect 35734 58270 35874 58284
rect 36024 58270 36832 58284
rect 36982 58270 37122 58284
rect 37272 58270 38080 58284
rect 38230 58270 38370 58284
rect 38520 58270 39328 58284
rect 39478 58270 39618 58284
rect 39768 58270 40576 58284
rect 40726 58270 40866 58284
rect 41016 58270 41824 58284
rect 41974 58270 42114 58284
rect 42264 58270 43072 58284
rect 43222 58270 43362 58284
rect 43512 58270 44320 58284
rect 44470 58270 44610 58284
rect 44760 58270 45568 58284
rect 45718 58270 45858 58284
rect 46008 58270 46816 58284
rect 46966 58270 47106 58284
rect 47256 58270 48064 58284
rect 48214 58270 48354 58284
rect 48504 58270 49312 58284
rect 49462 58270 49602 58284
rect 49752 58270 50560 58284
rect 50710 58270 50850 58284
rect 51000 58270 51808 58284
rect 51958 58270 52098 58284
rect 52248 58270 53056 58284
rect 53206 58270 53346 58284
rect 53496 58270 54304 58284
rect 54454 58270 54594 58284
rect 54744 58270 55552 58284
rect 55702 58270 55842 58284
rect 55992 58270 56800 58284
rect 56950 58270 57090 58284
rect 57240 58270 58048 58284
rect 58198 58270 58338 58284
rect 58488 58270 58934 58284
rect 16418 58222 58934 58270
rect 16418 58208 16864 58222
rect 17014 58208 17154 58222
rect 17304 58208 18112 58222
rect 18262 58208 18402 58222
rect 18552 58208 19360 58222
rect 19510 58208 19650 58222
rect 19800 58208 20608 58222
rect 20758 58208 20898 58222
rect 21048 58208 21856 58222
rect 22006 58208 22146 58222
rect 22296 58208 23104 58222
rect 23254 58208 23394 58222
rect 23544 58208 24352 58222
rect 24502 58208 24642 58222
rect 24792 58208 25600 58222
rect 25750 58208 25890 58222
rect 26040 58208 26848 58222
rect 26998 58208 27138 58222
rect 27288 58208 28096 58222
rect 28246 58208 28386 58222
rect 28536 58208 29344 58222
rect 29494 58208 29634 58222
rect 29784 58208 30592 58222
rect 30742 58208 30882 58222
rect 31032 58208 31840 58222
rect 31990 58208 32130 58222
rect 32280 58208 33088 58222
rect 33238 58208 33378 58222
rect 33528 58208 34336 58222
rect 34486 58208 34626 58222
rect 34776 58208 35584 58222
rect 35734 58208 35874 58222
rect 36024 58208 36832 58222
rect 36982 58208 37122 58222
rect 37272 58208 38080 58222
rect 38230 58208 38370 58222
rect 38520 58208 39328 58222
rect 39478 58208 39618 58222
rect 39768 58208 40576 58222
rect 40726 58208 40866 58222
rect 41016 58208 41824 58222
rect 41974 58208 42114 58222
rect 42264 58208 43072 58222
rect 43222 58208 43362 58222
rect 43512 58208 44320 58222
rect 44470 58208 44610 58222
rect 44760 58208 45568 58222
rect 45718 58208 45858 58222
rect 46008 58208 46816 58222
rect 46966 58208 47106 58222
rect 47256 58208 48064 58222
rect 48214 58208 48354 58222
rect 48504 58208 49312 58222
rect 49462 58208 49602 58222
rect 49752 58208 50560 58222
rect 50710 58208 50850 58222
rect 51000 58208 51808 58222
rect 51958 58208 52098 58222
rect 52248 58208 53056 58222
rect 53206 58208 53346 58222
rect 53496 58208 54304 58222
rect 54454 58208 54594 58222
rect 54744 58208 55552 58222
rect 55702 58208 55842 58222
rect 55992 58208 56800 58222
rect 56950 58208 57090 58222
rect 57240 58208 58048 58222
rect 58198 58208 58338 58222
rect 58488 58208 58934 58222
rect 16898 58160 16980 58174
rect 17188 58160 17270 58174
rect 18146 58160 18228 58174
rect 18436 58160 18518 58174
rect 19394 58160 19476 58174
rect 19684 58160 19766 58174
rect 20642 58160 20724 58174
rect 20932 58160 21014 58174
rect 21890 58160 21972 58174
rect 22180 58160 22262 58174
rect 23138 58160 23220 58174
rect 23428 58160 23510 58174
rect 24386 58160 24468 58174
rect 24676 58160 24758 58174
rect 25634 58160 25716 58174
rect 25924 58160 26006 58174
rect 26882 58160 26964 58174
rect 27172 58160 27254 58174
rect 28130 58160 28212 58174
rect 28420 58160 28502 58174
rect 29378 58160 29460 58174
rect 29668 58160 29750 58174
rect 30626 58160 30708 58174
rect 30916 58160 30998 58174
rect 31874 58160 31956 58174
rect 32164 58160 32246 58174
rect 33122 58160 33204 58174
rect 33412 58160 33494 58174
rect 34370 58160 34452 58174
rect 34660 58160 34742 58174
rect 35618 58160 35700 58174
rect 35908 58160 35990 58174
rect 36866 58160 36948 58174
rect 37156 58160 37238 58174
rect 38114 58160 38196 58174
rect 38404 58160 38486 58174
rect 39362 58160 39444 58174
rect 39652 58160 39734 58174
rect 40610 58160 40692 58174
rect 40900 58160 40982 58174
rect 41858 58160 41940 58174
rect 42148 58160 42230 58174
rect 43106 58160 43188 58174
rect 43396 58160 43478 58174
rect 44354 58160 44436 58174
rect 44644 58160 44726 58174
rect 45602 58160 45684 58174
rect 45892 58160 45974 58174
rect 46850 58160 46932 58174
rect 47140 58160 47222 58174
rect 48098 58160 48180 58174
rect 48388 58160 48470 58174
rect 49346 58160 49428 58174
rect 49636 58160 49718 58174
rect 50594 58160 50676 58174
rect 50884 58160 50966 58174
rect 51842 58160 51924 58174
rect 52132 58160 52214 58174
rect 53090 58160 53172 58174
rect 53380 58160 53462 58174
rect 54338 58160 54420 58174
rect 54628 58160 54710 58174
rect 55586 58160 55668 58174
rect 55876 58160 55958 58174
rect 56834 58160 56916 58174
rect 57124 58160 57206 58174
rect 58082 58160 58164 58174
rect 58372 58160 58454 58174
rect 16418 58112 58934 58160
rect 16418 58016 58934 58064
rect 16898 58002 16980 58016
rect 17188 58002 17270 58016
rect 18146 58002 18228 58016
rect 18436 58002 18518 58016
rect 19394 58002 19476 58016
rect 19684 58002 19766 58016
rect 20642 58002 20724 58016
rect 20932 58002 21014 58016
rect 21890 58002 21972 58016
rect 22180 58002 22262 58016
rect 23138 58002 23220 58016
rect 23428 58002 23510 58016
rect 24386 58002 24468 58016
rect 24676 58002 24758 58016
rect 25634 58002 25716 58016
rect 25924 58002 26006 58016
rect 26882 58002 26964 58016
rect 27172 58002 27254 58016
rect 28130 58002 28212 58016
rect 28420 58002 28502 58016
rect 29378 58002 29460 58016
rect 29668 58002 29750 58016
rect 30626 58002 30708 58016
rect 30916 58002 30998 58016
rect 31874 58002 31956 58016
rect 32164 58002 32246 58016
rect 33122 58002 33204 58016
rect 33412 58002 33494 58016
rect 34370 58002 34452 58016
rect 34660 58002 34742 58016
rect 35618 58002 35700 58016
rect 35908 58002 35990 58016
rect 36866 58002 36948 58016
rect 37156 58002 37238 58016
rect 38114 58002 38196 58016
rect 38404 58002 38486 58016
rect 39362 58002 39444 58016
rect 39652 58002 39734 58016
rect 40610 58002 40692 58016
rect 40900 58002 40982 58016
rect 41858 58002 41940 58016
rect 42148 58002 42230 58016
rect 43106 58002 43188 58016
rect 43396 58002 43478 58016
rect 44354 58002 44436 58016
rect 44644 58002 44726 58016
rect 45602 58002 45684 58016
rect 45892 58002 45974 58016
rect 46850 58002 46932 58016
rect 47140 58002 47222 58016
rect 48098 58002 48180 58016
rect 48388 58002 48470 58016
rect 49346 58002 49428 58016
rect 49636 58002 49718 58016
rect 50594 58002 50676 58016
rect 50884 58002 50966 58016
rect 51842 58002 51924 58016
rect 52132 58002 52214 58016
rect 53090 58002 53172 58016
rect 53380 58002 53462 58016
rect 54338 58002 54420 58016
rect 54628 58002 54710 58016
rect 55586 58002 55668 58016
rect 55876 58002 55958 58016
rect 56834 58002 56916 58016
rect 57124 58002 57206 58016
rect 58082 58002 58164 58016
rect 58372 58002 58454 58016
rect 16418 57954 16864 57968
rect 17014 57954 17154 57968
rect 17304 57954 18112 57968
rect 18262 57954 18402 57968
rect 18552 57954 19360 57968
rect 19510 57954 19650 57968
rect 19800 57954 20608 57968
rect 20758 57954 20898 57968
rect 21048 57954 21856 57968
rect 22006 57954 22146 57968
rect 22296 57954 23104 57968
rect 23254 57954 23394 57968
rect 23544 57954 24352 57968
rect 24502 57954 24642 57968
rect 24792 57954 25600 57968
rect 25750 57954 25890 57968
rect 26040 57954 26848 57968
rect 26998 57954 27138 57968
rect 27288 57954 28096 57968
rect 28246 57954 28386 57968
rect 28536 57954 29344 57968
rect 29494 57954 29634 57968
rect 29784 57954 30592 57968
rect 30742 57954 30882 57968
rect 31032 57954 31840 57968
rect 31990 57954 32130 57968
rect 32280 57954 33088 57968
rect 33238 57954 33378 57968
rect 33528 57954 34336 57968
rect 34486 57954 34626 57968
rect 34776 57954 35584 57968
rect 35734 57954 35874 57968
rect 36024 57954 36832 57968
rect 36982 57954 37122 57968
rect 37272 57954 38080 57968
rect 38230 57954 38370 57968
rect 38520 57954 39328 57968
rect 39478 57954 39618 57968
rect 39768 57954 40576 57968
rect 40726 57954 40866 57968
rect 41016 57954 41824 57968
rect 41974 57954 42114 57968
rect 42264 57954 43072 57968
rect 43222 57954 43362 57968
rect 43512 57954 44320 57968
rect 44470 57954 44610 57968
rect 44760 57954 45568 57968
rect 45718 57954 45858 57968
rect 46008 57954 46816 57968
rect 46966 57954 47106 57968
rect 47256 57954 48064 57968
rect 48214 57954 48354 57968
rect 48504 57954 49312 57968
rect 49462 57954 49602 57968
rect 49752 57954 50560 57968
rect 50710 57954 50850 57968
rect 51000 57954 51808 57968
rect 51958 57954 52098 57968
rect 52248 57954 53056 57968
rect 53206 57954 53346 57968
rect 53496 57954 54304 57968
rect 54454 57954 54594 57968
rect 54744 57954 55552 57968
rect 55702 57954 55842 57968
rect 55992 57954 56800 57968
rect 56950 57954 57090 57968
rect 57240 57954 58048 57968
rect 58198 57954 58338 57968
rect 58488 57954 58934 57968
rect 16418 57906 58934 57954
rect 16418 57892 16864 57906
rect 17014 57892 17154 57906
rect 17304 57892 18112 57906
rect 18262 57892 18402 57906
rect 18552 57892 19360 57906
rect 19510 57892 19650 57906
rect 19800 57892 20608 57906
rect 20758 57892 20898 57906
rect 21048 57892 21856 57906
rect 22006 57892 22146 57906
rect 22296 57892 23104 57906
rect 23254 57892 23394 57906
rect 23544 57892 24352 57906
rect 24502 57892 24642 57906
rect 24792 57892 25600 57906
rect 25750 57892 25890 57906
rect 26040 57892 26848 57906
rect 26998 57892 27138 57906
rect 27288 57892 28096 57906
rect 28246 57892 28386 57906
rect 28536 57892 29344 57906
rect 29494 57892 29634 57906
rect 29784 57892 30592 57906
rect 30742 57892 30882 57906
rect 31032 57892 31840 57906
rect 31990 57892 32130 57906
rect 32280 57892 33088 57906
rect 33238 57892 33378 57906
rect 33528 57892 34336 57906
rect 34486 57892 34626 57906
rect 34776 57892 35584 57906
rect 35734 57892 35874 57906
rect 36024 57892 36832 57906
rect 36982 57892 37122 57906
rect 37272 57892 38080 57906
rect 38230 57892 38370 57906
rect 38520 57892 39328 57906
rect 39478 57892 39618 57906
rect 39768 57892 40576 57906
rect 40726 57892 40866 57906
rect 41016 57892 41824 57906
rect 41974 57892 42114 57906
rect 42264 57892 43072 57906
rect 43222 57892 43362 57906
rect 43512 57892 44320 57906
rect 44470 57892 44610 57906
rect 44760 57892 45568 57906
rect 45718 57892 45858 57906
rect 46008 57892 46816 57906
rect 46966 57892 47106 57906
rect 47256 57892 48064 57906
rect 48214 57892 48354 57906
rect 48504 57892 49312 57906
rect 49462 57892 49602 57906
rect 49752 57892 50560 57906
rect 50710 57892 50850 57906
rect 51000 57892 51808 57906
rect 51958 57892 52098 57906
rect 52248 57892 53056 57906
rect 53206 57892 53346 57906
rect 53496 57892 54304 57906
rect 54454 57892 54594 57906
rect 54744 57892 55552 57906
rect 55702 57892 55842 57906
rect 55992 57892 56800 57906
rect 56950 57892 57090 57906
rect 57240 57892 58048 57906
rect 58198 57892 58338 57906
rect 58488 57892 58934 57906
rect 16898 57844 16980 57858
rect 17188 57844 17270 57858
rect 18146 57844 18228 57858
rect 18436 57844 18518 57858
rect 19394 57844 19476 57858
rect 19684 57844 19766 57858
rect 20642 57844 20724 57858
rect 20932 57844 21014 57858
rect 21890 57844 21972 57858
rect 22180 57844 22262 57858
rect 23138 57844 23220 57858
rect 23428 57844 23510 57858
rect 24386 57844 24468 57858
rect 24676 57844 24758 57858
rect 25634 57844 25716 57858
rect 25924 57844 26006 57858
rect 26882 57844 26964 57858
rect 27172 57844 27254 57858
rect 28130 57844 28212 57858
rect 28420 57844 28502 57858
rect 29378 57844 29460 57858
rect 29668 57844 29750 57858
rect 30626 57844 30708 57858
rect 30916 57844 30998 57858
rect 31874 57844 31956 57858
rect 32164 57844 32246 57858
rect 33122 57844 33204 57858
rect 33412 57844 33494 57858
rect 34370 57844 34452 57858
rect 34660 57844 34742 57858
rect 35618 57844 35700 57858
rect 35908 57844 35990 57858
rect 36866 57844 36948 57858
rect 37156 57844 37238 57858
rect 38114 57844 38196 57858
rect 38404 57844 38486 57858
rect 39362 57844 39444 57858
rect 39652 57844 39734 57858
rect 40610 57844 40692 57858
rect 40900 57844 40982 57858
rect 41858 57844 41940 57858
rect 42148 57844 42230 57858
rect 43106 57844 43188 57858
rect 43396 57844 43478 57858
rect 44354 57844 44436 57858
rect 44644 57844 44726 57858
rect 45602 57844 45684 57858
rect 45892 57844 45974 57858
rect 46850 57844 46932 57858
rect 47140 57844 47222 57858
rect 48098 57844 48180 57858
rect 48388 57844 48470 57858
rect 49346 57844 49428 57858
rect 49636 57844 49718 57858
rect 50594 57844 50676 57858
rect 50884 57844 50966 57858
rect 51842 57844 51924 57858
rect 52132 57844 52214 57858
rect 53090 57844 53172 57858
rect 53380 57844 53462 57858
rect 54338 57844 54420 57858
rect 54628 57844 54710 57858
rect 55586 57844 55668 57858
rect 55876 57844 55958 57858
rect 56834 57844 56916 57858
rect 57124 57844 57206 57858
rect 58082 57844 58164 57858
rect 58372 57844 58454 57858
rect 16418 57796 58934 57844
rect 16418 57638 58934 57748
rect 16418 57542 58934 57590
rect 16898 57528 16980 57542
rect 17188 57528 17270 57542
rect 18146 57528 18228 57542
rect 18436 57528 18518 57542
rect 19394 57528 19476 57542
rect 19684 57528 19766 57542
rect 20642 57528 20724 57542
rect 20932 57528 21014 57542
rect 21890 57528 21972 57542
rect 22180 57528 22262 57542
rect 23138 57528 23220 57542
rect 23428 57528 23510 57542
rect 24386 57528 24468 57542
rect 24676 57528 24758 57542
rect 25634 57528 25716 57542
rect 25924 57528 26006 57542
rect 26882 57528 26964 57542
rect 27172 57528 27254 57542
rect 28130 57528 28212 57542
rect 28420 57528 28502 57542
rect 29378 57528 29460 57542
rect 29668 57528 29750 57542
rect 30626 57528 30708 57542
rect 30916 57528 30998 57542
rect 31874 57528 31956 57542
rect 32164 57528 32246 57542
rect 33122 57528 33204 57542
rect 33412 57528 33494 57542
rect 34370 57528 34452 57542
rect 34660 57528 34742 57542
rect 35618 57528 35700 57542
rect 35908 57528 35990 57542
rect 36866 57528 36948 57542
rect 37156 57528 37238 57542
rect 38114 57528 38196 57542
rect 38404 57528 38486 57542
rect 39362 57528 39444 57542
rect 39652 57528 39734 57542
rect 40610 57528 40692 57542
rect 40900 57528 40982 57542
rect 41858 57528 41940 57542
rect 42148 57528 42230 57542
rect 43106 57528 43188 57542
rect 43396 57528 43478 57542
rect 44354 57528 44436 57542
rect 44644 57528 44726 57542
rect 45602 57528 45684 57542
rect 45892 57528 45974 57542
rect 46850 57528 46932 57542
rect 47140 57528 47222 57542
rect 48098 57528 48180 57542
rect 48388 57528 48470 57542
rect 49346 57528 49428 57542
rect 49636 57528 49718 57542
rect 50594 57528 50676 57542
rect 50884 57528 50966 57542
rect 51842 57528 51924 57542
rect 52132 57528 52214 57542
rect 53090 57528 53172 57542
rect 53380 57528 53462 57542
rect 54338 57528 54420 57542
rect 54628 57528 54710 57542
rect 55586 57528 55668 57542
rect 55876 57528 55958 57542
rect 56834 57528 56916 57542
rect 57124 57528 57206 57542
rect 58082 57528 58164 57542
rect 58372 57528 58454 57542
rect 16418 57480 16864 57494
rect 17014 57480 17154 57494
rect 17304 57480 18112 57494
rect 18262 57480 18402 57494
rect 18552 57480 19360 57494
rect 19510 57480 19650 57494
rect 19800 57480 20608 57494
rect 20758 57480 20898 57494
rect 21048 57480 21856 57494
rect 22006 57480 22146 57494
rect 22296 57480 23104 57494
rect 23254 57480 23394 57494
rect 23544 57480 24352 57494
rect 24502 57480 24642 57494
rect 24792 57480 25600 57494
rect 25750 57480 25890 57494
rect 26040 57480 26848 57494
rect 26998 57480 27138 57494
rect 27288 57480 28096 57494
rect 28246 57480 28386 57494
rect 28536 57480 29344 57494
rect 29494 57480 29634 57494
rect 29784 57480 30592 57494
rect 30742 57480 30882 57494
rect 31032 57480 31840 57494
rect 31990 57480 32130 57494
rect 32280 57480 33088 57494
rect 33238 57480 33378 57494
rect 33528 57480 34336 57494
rect 34486 57480 34626 57494
rect 34776 57480 35584 57494
rect 35734 57480 35874 57494
rect 36024 57480 36832 57494
rect 36982 57480 37122 57494
rect 37272 57480 38080 57494
rect 38230 57480 38370 57494
rect 38520 57480 39328 57494
rect 39478 57480 39618 57494
rect 39768 57480 40576 57494
rect 40726 57480 40866 57494
rect 41016 57480 41824 57494
rect 41974 57480 42114 57494
rect 42264 57480 43072 57494
rect 43222 57480 43362 57494
rect 43512 57480 44320 57494
rect 44470 57480 44610 57494
rect 44760 57480 45568 57494
rect 45718 57480 45858 57494
rect 46008 57480 46816 57494
rect 46966 57480 47106 57494
rect 47256 57480 48064 57494
rect 48214 57480 48354 57494
rect 48504 57480 49312 57494
rect 49462 57480 49602 57494
rect 49752 57480 50560 57494
rect 50710 57480 50850 57494
rect 51000 57480 51808 57494
rect 51958 57480 52098 57494
rect 52248 57480 53056 57494
rect 53206 57480 53346 57494
rect 53496 57480 54304 57494
rect 54454 57480 54594 57494
rect 54744 57480 55552 57494
rect 55702 57480 55842 57494
rect 55992 57480 56800 57494
rect 56950 57480 57090 57494
rect 57240 57480 58048 57494
rect 58198 57480 58338 57494
rect 58488 57480 58934 57494
rect 16418 57432 58934 57480
rect 16418 57418 16864 57432
rect 17014 57418 17154 57432
rect 17304 57418 18112 57432
rect 18262 57418 18402 57432
rect 18552 57418 19360 57432
rect 19510 57418 19650 57432
rect 19800 57418 20608 57432
rect 20758 57418 20898 57432
rect 21048 57418 21856 57432
rect 22006 57418 22146 57432
rect 22296 57418 23104 57432
rect 23254 57418 23394 57432
rect 23544 57418 24352 57432
rect 24502 57418 24642 57432
rect 24792 57418 25600 57432
rect 25750 57418 25890 57432
rect 26040 57418 26848 57432
rect 26998 57418 27138 57432
rect 27288 57418 28096 57432
rect 28246 57418 28386 57432
rect 28536 57418 29344 57432
rect 29494 57418 29634 57432
rect 29784 57418 30592 57432
rect 30742 57418 30882 57432
rect 31032 57418 31840 57432
rect 31990 57418 32130 57432
rect 32280 57418 33088 57432
rect 33238 57418 33378 57432
rect 33528 57418 34336 57432
rect 34486 57418 34626 57432
rect 34776 57418 35584 57432
rect 35734 57418 35874 57432
rect 36024 57418 36832 57432
rect 36982 57418 37122 57432
rect 37272 57418 38080 57432
rect 38230 57418 38370 57432
rect 38520 57418 39328 57432
rect 39478 57418 39618 57432
rect 39768 57418 40576 57432
rect 40726 57418 40866 57432
rect 41016 57418 41824 57432
rect 41974 57418 42114 57432
rect 42264 57418 43072 57432
rect 43222 57418 43362 57432
rect 43512 57418 44320 57432
rect 44470 57418 44610 57432
rect 44760 57418 45568 57432
rect 45718 57418 45858 57432
rect 46008 57418 46816 57432
rect 46966 57418 47106 57432
rect 47256 57418 48064 57432
rect 48214 57418 48354 57432
rect 48504 57418 49312 57432
rect 49462 57418 49602 57432
rect 49752 57418 50560 57432
rect 50710 57418 50850 57432
rect 51000 57418 51808 57432
rect 51958 57418 52098 57432
rect 52248 57418 53056 57432
rect 53206 57418 53346 57432
rect 53496 57418 54304 57432
rect 54454 57418 54594 57432
rect 54744 57418 55552 57432
rect 55702 57418 55842 57432
rect 55992 57418 56800 57432
rect 56950 57418 57090 57432
rect 57240 57418 58048 57432
rect 58198 57418 58338 57432
rect 58488 57418 58934 57432
rect 16898 57370 16980 57384
rect 17188 57370 17270 57384
rect 18146 57370 18228 57384
rect 18436 57370 18518 57384
rect 19394 57370 19476 57384
rect 19684 57370 19766 57384
rect 20642 57370 20724 57384
rect 20932 57370 21014 57384
rect 21890 57370 21972 57384
rect 22180 57370 22262 57384
rect 23138 57370 23220 57384
rect 23428 57370 23510 57384
rect 24386 57370 24468 57384
rect 24676 57370 24758 57384
rect 25634 57370 25716 57384
rect 25924 57370 26006 57384
rect 26882 57370 26964 57384
rect 27172 57370 27254 57384
rect 28130 57370 28212 57384
rect 28420 57370 28502 57384
rect 29378 57370 29460 57384
rect 29668 57370 29750 57384
rect 30626 57370 30708 57384
rect 30916 57370 30998 57384
rect 31874 57370 31956 57384
rect 32164 57370 32246 57384
rect 33122 57370 33204 57384
rect 33412 57370 33494 57384
rect 34370 57370 34452 57384
rect 34660 57370 34742 57384
rect 35618 57370 35700 57384
rect 35908 57370 35990 57384
rect 36866 57370 36948 57384
rect 37156 57370 37238 57384
rect 38114 57370 38196 57384
rect 38404 57370 38486 57384
rect 39362 57370 39444 57384
rect 39652 57370 39734 57384
rect 40610 57370 40692 57384
rect 40900 57370 40982 57384
rect 41858 57370 41940 57384
rect 42148 57370 42230 57384
rect 43106 57370 43188 57384
rect 43396 57370 43478 57384
rect 44354 57370 44436 57384
rect 44644 57370 44726 57384
rect 45602 57370 45684 57384
rect 45892 57370 45974 57384
rect 46850 57370 46932 57384
rect 47140 57370 47222 57384
rect 48098 57370 48180 57384
rect 48388 57370 48470 57384
rect 49346 57370 49428 57384
rect 49636 57370 49718 57384
rect 50594 57370 50676 57384
rect 50884 57370 50966 57384
rect 51842 57370 51924 57384
rect 52132 57370 52214 57384
rect 53090 57370 53172 57384
rect 53380 57370 53462 57384
rect 54338 57370 54420 57384
rect 54628 57370 54710 57384
rect 55586 57370 55668 57384
rect 55876 57370 55958 57384
rect 56834 57370 56916 57384
rect 57124 57370 57206 57384
rect 58082 57370 58164 57384
rect 58372 57370 58454 57384
rect 16418 57322 58934 57370
rect 16418 57226 58934 57274
rect 16898 57212 16980 57226
rect 17188 57212 17270 57226
rect 18146 57212 18228 57226
rect 18436 57212 18518 57226
rect 19394 57212 19476 57226
rect 19684 57212 19766 57226
rect 20642 57212 20724 57226
rect 20932 57212 21014 57226
rect 21890 57212 21972 57226
rect 22180 57212 22262 57226
rect 23138 57212 23220 57226
rect 23428 57212 23510 57226
rect 24386 57212 24468 57226
rect 24676 57212 24758 57226
rect 25634 57212 25716 57226
rect 25924 57212 26006 57226
rect 26882 57212 26964 57226
rect 27172 57212 27254 57226
rect 28130 57212 28212 57226
rect 28420 57212 28502 57226
rect 29378 57212 29460 57226
rect 29668 57212 29750 57226
rect 30626 57212 30708 57226
rect 30916 57212 30998 57226
rect 31874 57212 31956 57226
rect 32164 57212 32246 57226
rect 33122 57212 33204 57226
rect 33412 57212 33494 57226
rect 34370 57212 34452 57226
rect 34660 57212 34742 57226
rect 35618 57212 35700 57226
rect 35908 57212 35990 57226
rect 36866 57212 36948 57226
rect 37156 57212 37238 57226
rect 38114 57212 38196 57226
rect 38404 57212 38486 57226
rect 39362 57212 39444 57226
rect 39652 57212 39734 57226
rect 40610 57212 40692 57226
rect 40900 57212 40982 57226
rect 41858 57212 41940 57226
rect 42148 57212 42230 57226
rect 43106 57212 43188 57226
rect 43396 57212 43478 57226
rect 44354 57212 44436 57226
rect 44644 57212 44726 57226
rect 45602 57212 45684 57226
rect 45892 57212 45974 57226
rect 46850 57212 46932 57226
rect 47140 57212 47222 57226
rect 48098 57212 48180 57226
rect 48388 57212 48470 57226
rect 49346 57212 49428 57226
rect 49636 57212 49718 57226
rect 50594 57212 50676 57226
rect 50884 57212 50966 57226
rect 51842 57212 51924 57226
rect 52132 57212 52214 57226
rect 53090 57212 53172 57226
rect 53380 57212 53462 57226
rect 54338 57212 54420 57226
rect 54628 57212 54710 57226
rect 55586 57212 55668 57226
rect 55876 57212 55958 57226
rect 56834 57212 56916 57226
rect 57124 57212 57206 57226
rect 58082 57212 58164 57226
rect 58372 57212 58454 57226
rect 16418 57164 16864 57178
rect 17014 57164 17154 57178
rect 17304 57164 18112 57178
rect 18262 57164 18402 57178
rect 18552 57164 19360 57178
rect 19510 57164 19650 57178
rect 19800 57164 20608 57178
rect 20758 57164 20898 57178
rect 21048 57164 21856 57178
rect 22006 57164 22146 57178
rect 22296 57164 23104 57178
rect 23254 57164 23394 57178
rect 23544 57164 24352 57178
rect 24502 57164 24642 57178
rect 24792 57164 25600 57178
rect 25750 57164 25890 57178
rect 26040 57164 26848 57178
rect 26998 57164 27138 57178
rect 27288 57164 28096 57178
rect 28246 57164 28386 57178
rect 28536 57164 29344 57178
rect 29494 57164 29634 57178
rect 29784 57164 30592 57178
rect 30742 57164 30882 57178
rect 31032 57164 31840 57178
rect 31990 57164 32130 57178
rect 32280 57164 33088 57178
rect 33238 57164 33378 57178
rect 33528 57164 34336 57178
rect 34486 57164 34626 57178
rect 34776 57164 35584 57178
rect 35734 57164 35874 57178
rect 36024 57164 36832 57178
rect 36982 57164 37122 57178
rect 37272 57164 38080 57178
rect 38230 57164 38370 57178
rect 38520 57164 39328 57178
rect 39478 57164 39618 57178
rect 39768 57164 40576 57178
rect 40726 57164 40866 57178
rect 41016 57164 41824 57178
rect 41974 57164 42114 57178
rect 42264 57164 43072 57178
rect 43222 57164 43362 57178
rect 43512 57164 44320 57178
rect 44470 57164 44610 57178
rect 44760 57164 45568 57178
rect 45718 57164 45858 57178
rect 46008 57164 46816 57178
rect 46966 57164 47106 57178
rect 47256 57164 48064 57178
rect 48214 57164 48354 57178
rect 48504 57164 49312 57178
rect 49462 57164 49602 57178
rect 49752 57164 50560 57178
rect 50710 57164 50850 57178
rect 51000 57164 51808 57178
rect 51958 57164 52098 57178
rect 52248 57164 53056 57178
rect 53206 57164 53346 57178
rect 53496 57164 54304 57178
rect 54454 57164 54594 57178
rect 54744 57164 55552 57178
rect 55702 57164 55842 57178
rect 55992 57164 56800 57178
rect 56950 57164 57090 57178
rect 57240 57164 58048 57178
rect 58198 57164 58338 57178
rect 58488 57164 58934 57178
rect 16418 57116 58934 57164
rect 16418 57102 16864 57116
rect 17014 57102 17154 57116
rect 17304 57102 18112 57116
rect 18262 57102 18402 57116
rect 18552 57102 19360 57116
rect 19510 57102 19650 57116
rect 19800 57102 20608 57116
rect 20758 57102 20898 57116
rect 21048 57102 21856 57116
rect 22006 57102 22146 57116
rect 22296 57102 23104 57116
rect 23254 57102 23394 57116
rect 23544 57102 24352 57116
rect 24502 57102 24642 57116
rect 24792 57102 25600 57116
rect 25750 57102 25890 57116
rect 26040 57102 26848 57116
rect 26998 57102 27138 57116
rect 27288 57102 28096 57116
rect 28246 57102 28386 57116
rect 28536 57102 29344 57116
rect 29494 57102 29634 57116
rect 29784 57102 30592 57116
rect 30742 57102 30882 57116
rect 31032 57102 31840 57116
rect 31990 57102 32130 57116
rect 32280 57102 33088 57116
rect 33238 57102 33378 57116
rect 33528 57102 34336 57116
rect 34486 57102 34626 57116
rect 34776 57102 35584 57116
rect 35734 57102 35874 57116
rect 36024 57102 36832 57116
rect 36982 57102 37122 57116
rect 37272 57102 38080 57116
rect 38230 57102 38370 57116
rect 38520 57102 39328 57116
rect 39478 57102 39618 57116
rect 39768 57102 40576 57116
rect 40726 57102 40866 57116
rect 41016 57102 41824 57116
rect 41974 57102 42114 57116
rect 42264 57102 43072 57116
rect 43222 57102 43362 57116
rect 43512 57102 44320 57116
rect 44470 57102 44610 57116
rect 44760 57102 45568 57116
rect 45718 57102 45858 57116
rect 46008 57102 46816 57116
rect 46966 57102 47106 57116
rect 47256 57102 48064 57116
rect 48214 57102 48354 57116
rect 48504 57102 49312 57116
rect 49462 57102 49602 57116
rect 49752 57102 50560 57116
rect 50710 57102 50850 57116
rect 51000 57102 51808 57116
rect 51958 57102 52098 57116
rect 52248 57102 53056 57116
rect 53206 57102 53346 57116
rect 53496 57102 54304 57116
rect 54454 57102 54594 57116
rect 54744 57102 55552 57116
rect 55702 57102 55842 57116
rect 55992 57102 56800 57116
rect 56950 57102 57090 57116
rect 57240 57102 58048 57116
rect 58198 57102 58338 57116
rect 58488 57102 58934 57116
rect 16898 57054 16980 57068
rect 17188 57054 17270 57068
rect 18146 57054 18228 57068
rect 18436 57054 18518 57068
rect 19394 57054 19476 57068
rect 19684 57054 19766 57068
rect 20642 57054 20724 57068
rect 20932 57054 21014 57068
rect 21890 57054 21972 57068
rect 22180 57054 22262 57068
rect 23138 57054 23220 57068
rect 23428 57054 23510 57068
rect 24386 57054 24468 57068
rect 24676 57054 24758 57068
rect 25634 57054 25716 57068
rect 25924 57054 26006 57068
rect 26882 57054 26964 57068
rect 27172 57054 27254 57068
rect 28130 57054 28212 57068
rect 28420 57054 28502 57068
rect 29378 57054 29460 57068
rect 29668 57054 29750 57068
rect 30626 57054 30708 57068
rect 30916 57054 30998 57068
rect 31874 57054 31956 57068
rect 32164 57054 32246 57068
rect 33122 57054 33204 57068
rect 33412 57054 33494 57068
rect 34370 57054 34452 57068
rect 34660 57054 34742 57068
rect 35618 57054 35700 57068
rect 35908 57054 35990 57068
rect 36866 57054 36948 57068
rect 37156 57054 37238 57068
rect 38114 57054 38196 57068
rect 38404 57054 38486 57068
rect 39362 57054 39444 57068
rect 39652 57054 39734 57068
rect 40610 57054 40692 57068
rect 40900 57054 40982 57068
rect 41858 57054 41940 57068
rect 42148 57054 42230 57068
rect 43106 57054 43188 57068
rect 43396 57054 43478 57068
rect 44354 57054 44436 57068
rect 44644 57054 44726 57068
rect 45602 57054 45684 57068
rect 45892 57054 45974 57068
rect 46850 57054 46932 57068
rect 47140 57054 47222 57068
rect 48098 57054 48180 57068
rect 48388 57054 48470 57068
rect 49346 57054 49428 57068
rect 49636 57054 49718 57068
rect 50594 57054 50676 57068
rect 50884 57054 50966 57068
rect 51842 57054 51924 57068
rect 52132 57054 52214 57068
rect 53090 57054 53172 57068
rect 53380 57054 53462 57068
rect 54338 57054 54420 57068
rect 54628 57054 54710 57068
rect 55586 57054 55668 57068
rect 55876 57054 55958 57068
rect 56834 57054 56916 57068
rect 57124 57054 57206 57068
rect 58082 57054 58164 57068
rect 58372 57054 58454 57068
rect 16418 57006 58934 57054
rect 16418 56848 58934 56958
rect 16418 56752 58934 56800
rect 16898 56738 16980 56752
rect 17188 56738 17270 56752
rect 18146 56738 18228 56752
rect 18436 56738 18518 56752
rect 19394 56738 19476 56752
rect 19684 56738 19766 56752
rect 20642 56738 20724 56752
rect 20932 56738 21014 56752
rect 21890 56738 21972 56752
rect 22180 56738 22262 56752
rect 23138 56738 23220 56752
rect 23428 56738 23510 56752
rect 24386 56738 24468 56752
rect 24676 56738 24758 56752
rect 25634 56738 25716 56752
rect 25924 56738 26006 56752
rect 26882 56738 26964 56752
rect 27172 56738 27254 56752
rect 28130 56738 28212 56752
rect 28420 56738 28502 56752
rect 29378 56738 29460 56752
rect 29668 56738 29750 56752
rect 30626 56738 30708 56752
rect 30916 56738 30998 56752
rect 31874 56738 31956 56752
rect 32164 56738 32246 56752
rect 33122 56738 33204 56752
rect 33412 56738 33494 56752
rect 34370 56738 34452 56752
rect 34660 56738 34742 56752
rect 35618 56738 35700 56752
rect 35908 56738 35990 56752
rect 36866 56738 36948 56752
rect 37156 56738 37238 56752
rect 38114 56738 38196 56752
rect 38404 56738 38486 56752
rect 39362 56738 39444 56752
rect 39652 56738 39734 56752
rect 40610 56738 40692 56752
rect 40900 56738 40982 56752
rect 41858 56738 41940 56752
rect 42148 56738 42230 56752
rect 43106 56738 43188 56752
rect 43396 56738 43478 56752
rect 44354 56738 44436 56752
rect 44644 56738 44726 56752
rect 45602 56738 45684 56752
rect 45892 56738 45974 56752
rect 46850 56738 46932 56752
rect 47140 56738 47222 56752
rect 48098 56738 48180 56752
rect 48388 56738 48470 56752
rect 49346 56738 49428 56752
rect 49636 56738 49718 56752
rect 50594 56738 50676 56752
rect 50884 56738 50966 56752
rect 51842 56738 51924 56752
rect 52132 56738 52214 56752
rect 53090 56738 53172 56752
rect 53380 56738 53462 56752
rect 54338 56738 54420 56752
rect 54628 56738 54710 56752
rect 55586 56738 55668 56752
rect 55876 56738 55958 56752
rect 56834 56738 56916 56752
rect 57124 56738 57206 56752
rect 58082 56738 58164 56752
rect 58372 56738 58454 56752
rect 16418 56690 16864 56704
rect 17014 56690 17154 56704
rect 17304 56690 18112 56704
rect 18262 56690 18402 56704
rect 18552 56690 19360 56704
rect 19510 56690 19650 56704
rect 19800 56690 20608 56704
rect 20758 56690 20898 56704
rect 21048 56690 21856 56704
rect 22006 56690 22146 56704
rect 22296 56690 23104 56704
rect 23254 56690 23394 56704
rect 23544 56690 24352 56704
rect 24502 56690 24642 56704
rect 24792 56690 25600 56704
rect 25750 56690 25890 56704
rect 26040 56690 26848 56704
rect 26998 56690 27138 56704
rect 27288 56690 28096 56704
rect 28246 56690 28386 56704
rect 28536 56690 29344 56704
rect 29494 56690 29634 56704
rect 29784 56690 30592 56704
rect 30742 56690 30882 56704
rect 31032 56690 31840 56704
rect 31990 56690 32130 56704
rect 32280 56690 33088 56704
rect 33238 56690 33378 56704
rect 33528 56690 34336 56704
rect 34486 56690 34626 56704
rect 34776 56690 35584 56704
rect 35734 56690 35874 56704
rect 36024 56690 36832 56704
rect 36982 56690 37122 56704
rect 37272 56690 38080 56704
rect 38230 56690 38370 56704
rect 38520 56690 39328 56704
rect 39478 56690 39618 56704
rect 39768 56690 40576 56704
rect 40726 56690 40866 56704
rect 41016 56690 41824 56704
rect 41974 56690 42114 56704
rect 42264 56690 43072 56704
rect 43222 56690 43362 56704
rect 43512 56690 44320 56704
rect 44470 56690 44610 56704
rect 44760 56690 45568 56704
rect 45718 56690 45858 56704
rect 46008 56690 46816 56704
rect 46966 56690 47106 56704
rect 47256 56690 48064 56704
rect 48214 56690 48354 56704
rect 48504 56690 49312 56704
rect 49462 56690 49602 56704
rect 49752 56690 50560 56704
rect 50710 56690 50850 56704
rect 51000 56690 51808 56704
rect 51958 56690 52098 56704
rect 52248 56690 53056 56704
rect 53206 56690 53346 56704
rect 53496 56690 54304 56704
rect 54454 56690 54594 56704
rect 54744 56690 55552 56704
rect 55702 56690 55842 56704
rect 55992 56690 56800 56704
rect 56950 56690 57090 56704
rect 57240 56690 58048 56704
rect 58198 56690 58338 56704
rect 58488 56690 58934 56704
rect 16418 56642 58934 56690
rect 16418 56628 16864 56642
rect 17014 56628 17154 56642
rect 17304 56628 18112 56642
rect 18262 56628 18402 56642
rect 18552 56628 19360 56642
rect 19510 56628 19650 56642
rect 19800 56628 20608 56642
rect 20758 56628 20898 56642
rect 21048 56628 21856 56642
rect 22006 56628 22146 56642
rect 22296 56628 23104 56642
rect 23254 56628 23394 56642
rect 23544 56628 24352 56642
rect 24502 56628 24642 56642
rect 24792 56628 25600 56642
rect 25750 56628 25890 56642
rect 26040 56628 26848 56642
rect 26998 56628 27138 56642
rect 27288 56628 28096 56642
rect 28246 56628 28386 56642
rect 28536 56628 29344 56642
rect 29494 56628 29634 56642
rect 29784 56628 30592 56642
rect 30742 56628 30882 56642
rect 31032 56628 31840 56642
rect 31990 56628 32130 56642
rect 32280 56628 33088 56642
rect 33238 56628 33378 56642
rect 33528 56628 34336 56642
rect 34486 56628 34626 56642
rect 34776 56628 35584 56642
rect 35734 56628 35874 56642
rect 36024 56628 36832 56642
rect 36982 56628 37122 56642
rect 37272 56628 38080 56642
rect 38230 56628 38370 56642
rect 38520 56628 39328 56642
rect 39478 56628 39618 56642
rect 39768 56628 40576 56642
rect 40726 56628 40866 56642
rect 41016 56628 41824 56642
rect 41974 56628 42114 56642
rect 42264 56628 43072 56642
rect 43222 56628 43362 56642
rect 43512 56628 44320 56642
rect 44470 56628 44610 56642
rect 44760 56628 45568 56642
rect 45718 56628 45858 56642
rect 46008 56628 46816 56642
rect 46966 56628 47106 56642
rect 47256 56628 48064 56642
rect 48214 56628 48354 56642
rect 48504 56628 49312 56642
rect 49462 56628 49602 56642
rect 49752 56628 50560 56642
rect 50710 56628 50850 56642
rect 51000 56628 51808 56642
rect 51958 56628 52098 56642
rect 52248 56628 53056 56642
rect 53206 56628 53346 56642
rect 53496 56628 54304 56642
rect 54454 56628 54594 56642
rect 54744 56628 55552 56642
rect 55702 56628 55842 56642
rect 55992 56628 56800 56642
rect 56950 56628 57090 56642
rect 57240 56628 58048 56642
rect 58198 56628 58338 56642
rect 58488 56628 58934 56642
rect 16898 56580 16980 56594
rect 17188 56580 17270 56594
rect 18146 56580 18228 56594
rect 18436 56580 18518 56594
rect 19394 56580 19476 56594
rect 19684 56580 19766 56594
rect 20642 56580 20724 56594
rect 20932 56580 21014 56594
rect 21890 56580 21972 56594
rect 22180 56580 22262 56594
rect 23138 56580 23220 56594
rect 23428 56580 23510 56594
rect 24386 56580 24468 56594
rect 24676 56580 24758 56594
rect 25634 56580 25716 56594
rect 25924 56580 26006 56594
rect 26882 56580 26964 56594
rect 27172 56580 27254 56594
rect 28130 56580 28212 56594
rect 28420 56580 28502 56594
rect 29378 56580 29460 56594
rect 29668 56580 29750 56594
rect 30626 56580 30708 56594
rect 30916 56580 30998 56594
rect 31874 56580 31956 56594
rect 32164 56580 32246 56594
rect 33122 56580 33204 56594
rect 33412 56580 33494 56594
rect 34370 56580 34452 56594
rect 34660 56580 34742 56594
rect 35618 56580 35700 56594
rect 35908 56580 35990 56594
rect 36866 56580 36948 56594
rect 37156 56580 37238 56594
rect 38114 56580 38196 56594
rect 38404 56580 38486 56594
rect 39362 56580 39444 56594
rect 39652 56580 39734 56594
rect 40610 56580 40692 56594
rect 40900 56580 40982 56594
rect 41858 56580 41940 56594
rect 42148 56580 42230 56594
rect 43106 56580 43188 56594
rect 43396 56580 43478 56594
rect 44354 56580 44436 56594
rect 44644 56580 44726 56594
rect 45602 56580 45684 56594
rect 45892 56580 45974 56594
rect 46850 56580 46932 56594
rect 47140 56580 47222 56594
rect 48098 56580 48180 56594
rect 48388 56580 48470 56594
rect 49346 56580 49428 56594
rect 49636 56580 49718 56594
rect 50594 56580 50676 56594
rect 50884 56580 50966 56594
rect 51842 56580 51924 56594
rect 52132 56580 52214 56594
rect 53090 56580 53172 56594
rect 53380 56580 53462 56594
rect 54338 56580 54420 56594
rect 54628 56580 54710 56594
rect 55586 56580 55668 56594
rect 55876 56580 55958 56594
rect 56834 56580 56916 56594
rect 57124 56580 57206 56594
rect 58082 56580 58164 56594
rect 58372 56580 58454 56594
rect 16418 56532 58934 56580
rect 16418 56436 58934 56484
rect 16898 56422 16980 56436
rect 17188 56422 17270 56436
rect 18146 56422 18228 56436
rect 18436 56422 18518 56436
rect 19394 56422 19476 56436
rect 19684 56422 19766 56436
rect 20642 56422 20724 56436
rect 20932 56422 21014 56436
rect 21890 56422 21972 56436
rect 22180 56422 22262 56436
rect 23138 56422 23220 56436
rect 23428 56422 23510 56436
rect 24386 56422 24468 56436
rect 24676 56422 24758 56436
rect 25634 56422 25716 56436
rect 25924 56422 26006 56436
rect 26882 56422 26964 56436
rect 27172 56422 27254 56436
rect 28130 56422 28212 56436
rect 28420 56422 28502 56436
rect 29378 56422 29460 56436
rect 29668 56422 29750 56436
rect 30626 56422 30708 56436
rect 30916 56422 30998 56436
rect 31874 56422 31956 56436
rect 32164 56422 32246 56436
rect 33122 56422 33204 56436
rect 33412 56422 33494 56436
rect 34370 56422 34452 56436
rect 34660 56422 34742 56436
rect 35618 56422 35700 56436
rect 35908 56422 35990 56436
rect 36866 56422 36948 56436
rect 37156 56422 37238 56436
rect 38114 56422 38196 56436
rect 38404 56422 38486 56436
rect 39362 56422 39444 56436
rect 39652 56422 39734 56436
rect 40610 56422 40692 56436
rect 40900 56422 40982 56436
rect 41858 56422 41940 56436
rect 42148 56422 42230 56436
rect 43106 56422 43188 56436
rect 43396 56422 43478 56436
rect 44354 56422 44436 56436
rect 44644 56422 44726 56436
rect 45602 56422 45684 56436
rect 45892 56422 45974 56436
rect 46850 56422 46932 56436
rect 47140 56422 47222 56436
rect 48098 56422 48180 56436
rect 48388 56422 48470 56436
rect 49346 56422 49428 56436
rect 49636 56422 49718 56436
rect 50594 56422 50676 56436
rect 50884 56422 50966 56436
rect 51842 56422 51924 56436
rect 52132 56422 52214 56436
rect 53090 56422 53172 56436
rect 53380 56422 53462 56436
rect 54338 56422 54420 56436
rect 54628 56422 54710 56436
rect 55586 56422 55668 56436
rect 55876 56422 55958 56436
rect 56834 56422 56916 56436
rect 57124 56422 57206 56436
rect 58082 56422 58164 56436
rect 58372 56422 58454 56436
rect 16418 56374 16864 56388
rect 17014 56374 17154 56388
rect 17304 56374 18112 56388
rect 18262 56374 18402 56388
rect 18552 56374 19360 56388
rect 19510 56374 19650 56388
rect 19800 56374 20608 56388
rect 20758 56374 20898 56388
rect 21048 56374 21856 56388
rect 22006 56374 22146 56388
rect 22296 56374 23104 56388
rect 23254 56374 23394 56388
rect 23544 56374 24352 56388
rect 24502 56374 24642 56388
rect 24792 56374 25600 56388
rect 25750 56374 25890 56388
rect 26040 56374 26848 56388
rect 26998 56374 27138 56388
rect 27288 56374 28096 56388
rect 28246 56374 28386 56388
rect 28536 56374 29344 56388
rect 29494 56374 29634 56388
rect 29784 56374 30592 56388
rect 30742 56374 30882 56388
rect 31032 56374 31840 56388
rect 31990 56374 32130 56388
rect 32280 56374 33088 56388
rect 33238 56374 33378 56388
rect 33528 56374 34336 56388
rect 34486 56374 34626 56388
rect 34776 56374 35584 56388
rect 35734 56374 35874 56388
rect 36024 56374 36832 56388
rect 36982 56374 37122 56388
rect 37272 56374 38080 56388
rect 38230 56374 38370 56388
rect 38520 56374 39328 56388
rect 39478 56374 39618 56388
rect 39768 56374 40576 56388
rect 40726 56374 40866 56388
rect 41016 56374 41824 56388
rect 41974 56374 42114 56388
rect 42264 56374 43072 56388
rect 43222 56374 43362 56388
rect 43512 56374 44320 56388
rect 44470 56374 44610 56388
rect 44760 56374 45568 56388
rect 45718 56374 45858 56388
rect 46008 56374 46816 56388
rect 46966 56374 47106 56388
rect 47256 56374 48064 56388
rect 48214 56374 48354 56388
rect 48504 56374 49312 56388
rect 49462 56374 49602 56388
rect 49752 56374 50560 56388
rect 50710 56374 50850 56388
rect 51000 56374 51808 56388
rect 51958 56374 52098 56388
rect 52248 56374 53056 56388
rect 53206 56374 53346 56388
rect 53496 56374 54304 56388
rect 54454 56374 54594 56388
rect 54744 56374 55552 56388
rect 55702 56374 55842 56388
rect 55992 56374 56800 56388
rect 56950 56374 57090 56388
rect 57240 56374 58048 56388
rect 58198 56374 58338 56388
rect 58488 56374 58934 56388
rect 16418 56326 58934 56374
rect 16418 56312 16864 56326
rect 17014 56312 17154 56326
rect 17304 56312 18112 56326
rect 18262 56312 18402 56326
rect 18552 56312 19360 56326
rect 19510 56312 19650 56326
rect 19800 56312 20608 56326
rect 20758 56312 20898 56326
rect 21048 56312 21856 56326
rect 22006 56312 22146 56326
rect 22296 56312 23104 56326
rect 23254 56312 23394 56326
rect 23544 56312 24352 56326
rect 24502 56312 24642 56326
rect 24792 56312 25600 56326
rect 25750 56312 25890 56326
rect 26040 56312 26848 56326
rect 26998 56312 27138 56326
rect 27288 56312 28096 56326
rect 28246 56312 28386 56326
rect 28536 56312 29344 56326
rect 29494 56312 29634 56326
rect 29784 56312 30592 56326
rect 30742 56312 30882 56326
rect 31032 56312 31840 56326
rect 31990 56312 32130 56326
rect 32280 56312 33088 56326
rect 33238 56312 33378 56326
rect 33528 56312 34336 56326
rect 34486 56312 34626 56326
rect 34776 56312 35584 56326
rect 35734 56312 35874 56326
rect 36024 56312 36832 56326
rect 36982 56312 37122 56326
rect 37272 56312 38080 56326
rect 38230 56312 38370 56326
rect 38520 56312 39328 56326
rect 39478 56312 39618 56326
rect 39768 56312 40576 56326
rect 40726 56312 40866 56326
rect 41016 56312 41824 56326
rect 41974 56312 42114 56326
rect 42264 56312 43072 56326
rect 43222 56312 43362 56326
rect 43512 56312 44320 56326
rect 44470 56312 44610 56326
rect 44760 56312 45568 56326
rect 45718 56312 45858 56326
rect 46008 56312 46816 56326
rect 46966 56312 47106 56326
rect 47256 56312 48064 56326
rect 48214 56312 48354 56326
rect 48504 56312 49312 56326
rect 49462 56312 49602 56326
rect 49752 56312 50560 56326
rect 50710 56312 50850 56326
rect 51000 56312 51808 56326
rect 51958 56312 52098 56326
rect 52248 56312 53056 56326
rect 53206 56312 53346 56326
rect 53496 56312 54304 56326
rect 54454 56312 54594 56326
rect 54744 56312 55552 56326
rect 55702 56312 55842 56326
rect 55992 56312 56800 56326
rect 56950 56312 57090 56326
rect 57240 56312 58048 56326
rect 58198 56312 58338 56326
rect 58488 56312 58934 56326
rect 16898 56264 16980 56278
rect 17188 56264 17270 56278
rect 18146 56264 18228 56278
rect 18436 56264 18518 56278
rect 19394 56264 19476 56278
rect 19684 56264 19766 56278
rect 20642 56264 20724 56278
rect 20932 56264 21014 56278
rect 21890 56264 21972 56278
rect 22180 56264 22262 56278
rect 23138 56264 23220 56278
rect 23428 56264 23510 56278
rect 24386 56264 24468 56278
rect 24676 56264 24758 56278
rect 25634 56264 25716 56278
rect 25924 56264 26006 56278
rect 26882 56264 26964 56278
rect 27172 56264 27254 56278
rect 28130 56264 28212 56278
rect 28420 56264 28502 56278
rect 29378 56264 29460 56278
rect 29668 56264 29750 56278
rect 30626 56264 30708 56278
rect 30916 56264 30998 56278
rect 31874 56264 31956 56278
rect 32164 56264 32246 56278
rect 33122 56264 33204 56278
rect 33412 56264 33494 56278
rect 34370 56264 34452 56278
rect 34660 56264 34742 56278
rect 35618 56264 35700 56278
rect 35908 56264 35990 56278
rect 36866 56264 36948 56278
rect 37156 56264 37238 56278
rect 38114 56264 38196 56278
rect 38404 56264 38486 56278
rect 39362 56264 39444 56278
rect 39652 56264 39734 56278
rect 40610 56264 40692 56278
rect 40900 56264 40982 56278
rect 41858 56264 41940 56278
rect 42148 56264 42230 56278
rect 43106 56264 43188 56278
rect 43396 56264 43478 56278
rect 44354 56264 44436 56278
rect 44644 56264 44726 56278
rect 45602 56264 45684 56278
rect 45892 56264 45974 56278
rect 46850 56264 46932 56278
rect 47140 56264 47222 56278
rect 48098 56264 48180 56278
rect 48388 56264 48470 56278
rect 49346 56264 49428 56278
rect 49636 56264 49718 56278
rect 50594 56264 50676 56278
rect 50884 56264 50966 56278
rect 51842 56264 51924 56278
rect 52132 56264 52214 56278
rect 53090 56264 53172 56278
rect 53380 56264 53462 56278
rect 54338 56264 54420 56278
rect 54628 56264 54710 56278
rect 55586 56264 55668 56278
rect 55876 56264 55958 56278
rect 56834 56264 56916 56278
rect 57124 56264 57206 56278
rect 58082 56264 58164 56278
rect 58372 56264 58454 56278
rect 16418 56216 58934 56264
rect 16418 56058 58934 56168
rect 16418 55962 58934 56010
rect 16898 55948 16980 55962
rect 17188 55948 17270 55962
rect 18146 55948 18228 55962
rect 18436 55948 18518 55962
rect 19394 55948 19476 55962
rect 19684 55948 19766 55962
rect 20642 55948 20724 55962
rect 20932 55948 21014 55962
rect 21890 55948 21972 55962
rect 22180 55948 22262 55962
rect 23138 55948 23220 55962
rect 23428 55948 23510 55962
rect 24386 55948 24468 55962
rect 24676 55948 24758 55962
rect 25634 55948 25716 55962
rect 25924 55948 26006 55962
rect 26882 55948 26964 55962
rect 27172 55948 27254 55962
rect 28130 55948 28212 55962
rect 28420 55948 28502 55962
rect 29378 55948 29460 55962
rect 29668 55948 29750 55962
rect 30626 55948 30708 55962
rect 30916 55948 30998 55962
rect 31874 55948 31956 55962
rect 32164 55948 32246 55962
rect 33122 55948 33204 55962
rect 33412 55948 33494 55962
rect 34370 55948 34452 55962
rect 34660 55948 34742 55962
rect 35618 55948 35700 55962
rect 35908 55948 35990 55962
rect 36866 55948 36948 55962
rect 37156 55948 37238 55962
rect 38114 55948 38196 55962
rect 38404 55948 38486 55962
rect 39362 55948 39444 55962
rect 39652 55948 39734 55962
rect 40610 55948 40692 55962
rect 40900 55948 40982 55962
rect 41858 55948 41940 55962
rect 42148 55948 42230 55962
rect 43106 55948 43188 55962
rect 43396 55948 43478 55962
rect 44354 55948 44436 55962
rect 44644 55948 44726 55962
rect 45602 55948 45684 55962
rect 45892 55948 45974 55962
rect 46850 55948 46932 55962
rect 47140 55948 47222 55962
rect 48098 55948 48180 55962
rect 48388 55948 48470 55962
rect 49346 55948 49428 55962
rect 49636 55948 49718 55962
rect 50594 55948 50676 55962
rect 50884 55948 50966 55962
rect 51842 55948 51924 55962
rect 52132 55948 52214 55962
rect 53090 55948 53172 55962
rect 53380 55948 53462 55962
rect 54338 55948 54420 55962
rect 54628 55948 54710 55962
rect 55586 55948 55668 55962
rect 55876 55948 55958 55962
rect 56834 55948 56916 55962
rect 57124 55948 57206 55962
rect 58082 55948 58164 55962
rect 58372 55948 58454 55962
rect 16418 55900 16864 55914
rect 17014 55900 17154 55914
rect 17304 55900 18112 55914
rect 18262 55900 18402 55914
rect 18552 55900 19360 55914
rect 19510 55900 19650 55914
rect 19800 55900 20608 55914
rect 20758 55900 20898 55914
rect 21048 55900 21856 55914
rect 22006 55900 22146 55914
rect 22296 55900 23104 55914
rect 23254 55900 23394 55914
rect 23544 55900 24352 55914
rect 24502 55900 24642 55914
rect 24792 55900 25600 55914
rect 25750 55900 25890 55914
rect 26040 55900 26848 55914
rect 26998 55900 27138 55914
rect 27288 55900 28096 55914
rect 28246 55900 28386 55914
rect 28536 55900 29344 55914
rect 29494 55900 29634 55914
rect 29784 55900 30592 55914
rect 30742 55900 30882 55914
rect 31032 55900 31840 55914
rect 31990 55900 32130 55914
rect 32280 55900 33088 55914
rect 33238 55900 33378 55914
rect 33528 55900 34336 55914
rect 34486 55900 34626 55914
rect 34776 55900 35584 55914
rect 35734 55900 35874 55914
rect 36024 55900 36832 55914
rect 36982 55900 37122 55914
rect 37272 55900 38080 55914
rect 38230 55900 38370 55914
rect 38520 55900 39328 55914
rect 39478 55900 39618 55914
rect 39768 55900 40576 55914
rect 40726 55900 40866 55914
rect 41016 55900 41824 55914
rect 41974 55900 42114 55914
rect 42264 55900 43072 55914
rect 43222 55900 43362 55914
rect 43512 55900 44320 55914
rect 44470 55900 44610 55914
rect 44760 55900 45568 55914
rect 45718 55900 45858 55914
rect 46008 55900 46816 55914
rect 46966 55900 47106 55914
rect 47256 55900 48064 55914
rect 48214 55900 48354 55914
rect 48504 55900 49312 55914
rect 49462 55900 49602 55914
rect 49752 55900 50560 55914
rect 50710 55900 50850 55914
rect 51000 55900 51808 55914
rect 51958 55900 52098 55914
rect 52248 55900 53056 55914
rect 53206 55900 53346 55914
rect 53496 55900 54304 55914
rect 54454 55900 54594 55914
rect 54744 55900 55552 55914
rect 55702 55900 55842 55914
rect 55992 55900 56800 55914
rect 56950 55900 57090 55914
rect 57240 55900 58048 55914
rect 58198 55900 58338 55914
rect 58488 55900 58934 55914
rect 16418 55852 58934 55900
rect 16418 55838 16864 55852
rect 17014 55838 17154 55852
rect 17304 55838 18112 55852
rect 18262 55838 18402 55852
rect 18552 55838 19360 55852
rect 19510 55838 19650 55852
rect 19800 55838 20608 55852
rect 20758 55838 20898 55852
rect 21048 55838 21856 55852
rect 22006 55838 22146 55852
rect 22296 55838 23104 55852
rect 23254 55838 23394 55852
rect 23544 55838 24352 55852
rect 24502 55838 24642 55852
rect 24792 55838 25600 55852
rect 25750 55838 25890 55852
rect 26040 55838 26848 55852
rect 26998 55838 27138 55852
rect 27288 55838 28096 55852
rect 28246 55838 28386 55852
rect 28536 55838 29344 55852
rect 29494 55838 29634 55852
rect 29784 55838 30592 55852
rect 30742 55838 30882 55852
rect 31032 55838 31840 55852
rect 31990 55838 32130 55852
rect 32280 55838 33088 55852
rect 33238 55838 33378 55852
rect 33528 55838 34336 55852
rect 34486 55838 34626 55852
rect 34776 55838 35584 55852
rect 35734 55838 35874 55852
rect 36024 55838 36832 55852
rect 36982 55838 37122 55852
rect 37272 55838 38080 55852
rect 38230 55838 38370 55852
rect 38520 55838 39328 55852
rect 39478 55838 39618 55852
rect 39768 55838 40576 55852
rect 40726 55838 40866 55852
rect 41016 55838 41824 55852
rect 41974 55838 42114 55852
rect 42264 55838 43072 55852
rect 43222 55838 43362 55852
rect 43512 55838 44320 55852
rect 44470 55838 44610 55852
rect 44760 55838 45568 55852
rect 45718 55838 45858 55852
rect 46008 55838 46816 55852
rect 46966 55838 47106 55852
rect 47256 55838 48064 55852
rect 48214 55838 48354 55852
rect 48504 55838 49312 55852
rect 49462 55838 49602 55852
rect 49752 55838 50560 55852
rect 50710 55838 50850 55852
rect 51000 55838 51808 55852
rect 51958 55838 52098 55852
rect 52248 55838 53056 55852
rect 53206 55838 53346 55852
rect 53496 55838 54304 55852
rect 54454 55838 54594 55852
rect 54744 55838 55552 55852
rect 55702 55838 55842 55852
rect 55992 55838 56800 55852
rect 56950 55838 57090 55852
rect 57240 55838 58048 55852
rect 58198 55838 58338 55852
rect 58488 55838 58934 55852
rect 16898 55790 16980 55804
rect 17188 55790 17270 55804
rect 18146 55790 18228 55804
rect 18436 55790 18518 55804
rect 19394 55790 19476 55804
rect 19684 55790 19766 55804
rect 20642 55790 20724 55804
rect 20932 55790 21014 55804
rect 21890 55790 21972 55804
rect 22180 55790 22262 55804
rect 23138 55790 23220 55804
rect 23428 55790 23510 55804
rect 24386 55790 24468 55804
rect 24676 55790 24758 55804
rect 25634 55790 25716 55804
rect 25924 55790 26006 55804
rect 26882 55790 26964 55804
rect 27172 55790 27254 55804
rect 28130 55790 28212 55804
rect 28420 55790 28502 55804
rect 29378 55790 29460 55804
rect 29668 55790 29750 55804
rect 30626 55790 30708 55804
rect 30916 55790 30998 55804
rect 31874 55790 31956 55804
rect 32164 55790 32246 55804
rect 33122 55790 33204 55804
rect 33412 55790 33494 55804
rect 34370 55790 34452 55804
rect 34660 55790 34742 55804
rect 35618 55790 35700 55804
rect 35908 55790 35990 55804
rect 36866 55790 36948 55804
rect 37156 55790 37238 55804
rect 38114 55790 38196 55804
rect 38404 55790 38486 55804
rect 39362 55790 39444 55804
rect 39652 55790 39734 55804
rect 40610 55790 40692 55804
rect 40900 55790 40982 55804
rect 41858 55790 41940 55804
rect 42148 55790 42230 55804
rect 43106 55790 43188 55804
rect 43396 55790 43478 55804
rect 44354 55790 44436 55804
rect 44644 55790 44726 55804
rect 45602 55790 45684 55804
rect 45892 55790 45974 55804
rect 46850 55790 46932 55804
rect 47140 55790 47222 55804
rect 48098 55790 48180 55804
rect 48388 55790 48470 55804
rect 49346 55790 49428 55804
rect 49636 55790 49718 55804
rect 50594 55790 50676 55804
rect 50884 55790 50966 55804
rect 51842 55790 51924 55804
rect 52132 55790 52214 55804
rect 53090 55790 53172 55804
rect 53380 55790 53462 55804
rect 54338 55790 54420 55804
rect 54628 55790 54710 55804
rect 55586 55790 55668 55804
rect 55876 55790 55958 55804
rect 56834 55790 56916 55804
rect 57124 55790 57206 55804
rect 58082 55790 58164 55804
rect 58372 55790 58454 55804
rect 16418 55742 58934 55790
rect 16418 55646 58934 55694
rect 16898 55632 16980 55646
rect 17188 55632 17270 55646
rect 18146 55632 18228 55646
rect 18436 55632 18518 55646
rect 19394 55632 19476 55646
rect 19684 55632 19766 55646
rect 20642 55632 20724 55646
rect 20932 55632 21014 55646
rect 21890 55632 21972 55646
rect 22180 55632 22262 55646
rect 23138 55632 23220 55646
rect 23428 55632 23510 55646
rect 24386 55632 24468 55646
rect 24676 55632 24758 55646
rect 25634 55632 25716 55646
rect 25924 55632 26006 55646
rect 26882 55632 26964 55646
rect 27172 55632 27254 55646
rect 28130 55632 28212 55646
rect 28420 55632 28502 55646
rect 29378 55632 29460 55646
rect 29668 55632 29750 55646
rect 30626 55632 30708 55646
rect 30916 55632 30998 55646
rect 31874 55632 31956 55646
rect 32164 55632 32246 55646
rect 33122 55632 33204 55646
rect 33412 55632 33494 55646
rect 34370 55632 34452 55646
rect 34660 55632 34742 55646
rect 35618 55632 35700 55646
rect 35908 55632 35990 55646
rect 36866 55632 36948 55646
rect 37156 55632 37238 55646
rect 38114 55632 38196 55646
rect 38404 55632 38486 55646
rect 39362 55632 39444 55646
rect 39652 55632 39734 55646
rect 40610 55632 40692 55646
rect 40900 55632 40982 55646
rect 41858 55632 41940 55646
rect 42148 55632 42230 55646
rect 43106 55632 43188 55646
rect 43396 55632 43478 55646
rect 44354 55632 44436 55646
rect 44644 55632 44726 55646
rect 45602 55632 45684 55646
rect 45892 55632 45974 55646
rect 46850 55632 46932 55646
rect 47140 55632 47222 55646
rect 48098 55632 48180 55646
rect 48388 55632 48470 55646
rect 49346 55632 49428 55646
rect 49636 55632 49718 55646
rect 50594 55632 50676 55646
rect 50884 55632 50966 55646
rect 51842 55632 51924 55646
rect 52132 55632 52214 55646
rect 53090 55632 53172 55646
rect 53380 55632 53462 55646
rect 54338 55632 54420 55646
rect 54628 55632 54710 55646
rect 55586 55632 55668 55646
rect 55876 55632 55958 55646
rect 56834 55632 56916 55646
rect 57124 55632 57206 55646
rect 58082 55632 58164 55646
rect 58372 55632 58454 55646
rect 16418 55584 16864 55598
rect 17014 55584 17154 55598
rect 17304 55584 18112 55598
rect 18262 55584 18402 55598
rect 18552 55584 19360 55598
rect 19510 55584 19650 55598
rect 19800 55584 20608 55598
rect 20758 55584 20898 55598
rect 21048 55584 21856 55598
rect 22006 55584 22146 55598
rect 22296 55584 23104 55598
rect 23254 55584 23394 55598
rect 23544 55584 24352 55598
rect 24502 55584 24642 55598
rect 24792 55584 25600 55598
rect 25750 55584 25890 55598
rect 26040 55584 26848 55598
rect 26998 55584 27138 55598
rect 27288 55584 28096 55598
rect 28246 55584 28386 55598
rect 28536 55584 29344 55598
rect 29494 55584 29634 55598
rect 29784 55584 30592 55598
rect 30742 55584 30882 55598
rect 31032 55584 31840 55598
rect 31990 55584 32130 55598
rect 32280 55584 33088 55598
rect 33238 55584 33378 55598
rect 33528 55584 34336 55598
rect 34486 55584 34626 55598
rect 34776 55584 35584 55598
rect 35734 55584 35874 55598
rect 36024 55584 36832 55598
rect 36982 55584 37122 55598
rect 37272 55584 38080 55598
rect 38230 55584 38370 55598
rect 38520 55584 39328 55598
rect 39478 55584 39618 55598
rect 39768 55584 40576 55598
rect 40726 55584 40866 55598
rect 41016 55584 41824 55598
rect 41974 55584 42114 55598
rect 42264 55584 43072 55598
rect 43222 55584 43362 55598
rect 43512 55584 44320 55598
rect 44470 55584 44610 55598
rect 44760 55584 45568 55598
rect 45718 55584 45858 55598
rect 46008 55584 46816 55598
rect 46966 55584 47106 55598
rect 47256 55584 48064 55598
rect 48214 55584 48354 55598
rect 48504 55584 49312 55598
rect 49462 55584 49602 55598
rect 49752 55584 50560 55598
rect 50710 55584 50850 55598
rect 51000 55584 51808 55598
rect 51958 55584 52098 55598
rect 52248 55584 53056 55598
rect 53206 55584 53346 55598
rect 53496 55584 54304 55598
rect 54454 55584 54594 55598
rect 54744 55584 55552 55598
rect 55702 55584 55842 55598
rect 55992 55584 56800 55598
rect 56950 55584 57090 55598
rect 57240 55584 58048 55598
rect 58198 55584 58338 55598
rect 58488 55584 58934 55598
rect 16418 55536 58934 55584
rect 16418 55522 16864 55536
rect 17014 55522 17154 55536
rect 17304 55522 18112 55536
rect 18262 55522 18402 55536
rect 18552 55522 19360 55536
rect 19510 55522 19650 55536
rect 19800 55522 20608 55536
rect 20758 55522 20898 55536
rect 21048 55522 21856 55536
rect 22006 55522 22146 55536
rect 22296 55522 23104 55536
rect 23254 55522 23394 55536
rect 23544 55522 24352 55536
rect 24502 55522 24642 55536
rect 24792 55522 25600 55536
rect 25750 55522 25890 55536
rect 26040 55522 26848 55536
rect 26998 55522 27138 55536
rect 27288 55522 28096 55536
rect 28246 55522 28386 55536
rect 28536 55522 29344 55536
rect 29494 55522 29634 55536
rect 29784 55522 30592 55536
rect 30742 55522 30882 55536
rect 31032 55522 31840 55536
rect 31990 55522 32130 55536
rect 32280 55522 33088 55536
rect 33238 55522 33378 55536
rect 33528 55522 34336 55536
rect 34486 55522 34626 55536
rect 34776 55522 35584 55536
rect 35734 55522 35874 55536
rect 36024 55522 36832 55536
rect 36982 55522 37122 55536
rect 37272 55522 38080 55536
rect 38230 55522 38370 55536
rect 38520 55522 39328 55536
rect 39478 55522 39618 55536
rect 39768 55522 40576 55536
rect 40726 55522 40866 55536
rect 41016 55522 41824 55536
rect 41974 55522 42114 55536
rect 42264 55522 43072 55536
rect 43222 55522 43362 55536
rect 43512 55522 44320 55536
rect 44470 55522 44610 55536
rect 44760 55522 45568 55536
rect 45718 55522 45858 55536
rect 46008 55522 46816 55536
rect 46966 55522 47106 55536
rect 47256 55522 48064 55536
rect 48214 55522 48354 55536
rect 48504 55522 49312 55536
rect 49462 55522 49602 55536
rect 49752 55522 50560 55536
rect 50710 55522 50850 55536
rect 51000 55522 51808 55536
rect 51958 55522 52098 55536
rect 52248 55522 53056 55536
rect 53206 55522 53346 55536
rect 53496 55522 54304 55536
rect 54454 55522 54594 55536
rect 54744 55522 55552 55536
rect 55702 55522 55842 55536
rect 55992 55522 56800 55536
rect 56950 55522 57090 55536
rect 57240 55522 58048 55536
rect 58198 55522 58338 55536
rect 58488 55522 58934 55536
rect 16898 55474 16980 55488
rect 17188 55474 17270 55488
rect 18146 55474 18228 55488
rect 18436 55474 18518 55488
rect 19394 55474 19476 55488
rect 19684 55474 19766 55488
rect 20642 55474 20724 55488
rect 20932 55474 21014 55488
rect 21890 55474 21972 55488
rect 22180 55474 22262 55488
rect 23138 55474 23220 55488
rect 23428 55474 23510 55488
rect 24386 55474 24468 55488
rect 24676 55474 24758 55488
rect 25634 55474 25716 55488
rect 25924 55474 26006 55488
rect 26882 55474 26964 55488
rect 27172 55474 27254 55488
rect 28130 55474 28212 55488
rect 28420 55474 28502 55488
rect 29378 55474 29460 55488
rect 29668 55474 29750 55488
rect 30626 55474 30708 55488
rect 30916 55474 30998 55488
rect 31874 55474 31956 55488
rect 32164 55474 32246 55488
rect 33122 55474 33204 55488
rect 33412 55474 33494 55488
rect 34370 55474 34452 55488
rect 34660 55474 34742 55488
rect 35618 55474 35700 55488
rect 35908 55474 35990 55488
rect 36866 55474 36948 55488
rect 37156 55474 37238 55488
rect 38114 55474 38196 55488
rect 38404 55474 38486 55488
rect 39362 55474 39444 55488
rect 39652 55474 39734 55488
rect 40610 55474 40692 55488
rect 40900 55474 40982 55488
rect 41858 55474 41940 55488
rect 42148 55474 42230 55488
rect 43106 55474 43188 55488
rect 43396 55474 43478 55488
rect 44354 55474 44436 55488
rect 44644 55474 44726 55488
rect 45602 55474 45684 55488
rect 45892 55474 45974 55488
rect 46850 55474 46932 55488
rect 47140 55474 47222 55488
rect 48098 55474 48180 55488
rect 48388 55474 48470 55488
rect 49346 55474 49428 55488
rect 49636 55474 49718 55488
rect 50594 55474 50676 55488
rect 50884 55474 50966 55488
rect 51842 55474 51924 55488
rect 52132 55474 52214 55488
rect 53090 55474 53172 55488
rect 53380 55474 53462 55488
rect 54338 55474 54420 55488
rect 54628 55474 54710 55488
rect 55586 55474 55668 55488
rect 55876 55474 55958 55488
rect 56834 55474 56916 55488
rect 57124 55474 57206 55488
rect 58082 55474 58164 55488
rect 58372 55474 58454 55488
rect 16418 55426 58934 55474
rect 16418 55268 58934 55378
rect 16418 55172 58934 55220
rect 16898 55158 16980 55172
rect 17188 55158 17270 55172
rect 18146 55158 18228 55172
rect 18436 55158 18518 55172
rect 19394 55158 19476 55172
rect 19684 55158 19766 55172
rect 20642 55158 20724 55172
rect 20932 55158 21014 55172
rect 21890 55158 21972 55172
rect 22180 55158 22262 55172
rect 23138 55158 23220 55172
rect 23428 55158 23510 55172
rect 24386 55158 24468 55172
rect 24676 55158 24758 55172
rect 25634 55158 25716 55172
rect 25924 55158 26006 55172
rect 26882 55158 26964 55172
rect 27172 55158 27254 55172
rect 28130 55158 28212 55172
rect 28420 55158 28502 55172
rect 29378 55158 29460 55172
rect 29668 55158 29750 55172
rect 30626 55158 30708 55172
rect 30916 55158 30998 55172
rect 31874 55158 31956 55172
rect 32164 55158 32246 55172
rect 33122 55158 33204 55172
rect 33412 55158 33494 55172
rect 34370 55158 34452 55172
rect 34660 55158 34742 55172
rect 35618 55158 35700 55172
rect 35908 55158 35990 55172
rect 36866 55158 36948 55172
rect 37156 55158 37238 55172
rect 38114 55158 38196 55172
rect 38404 55158 38486 55172
rect 39362 55158 39444 55172
rect 39652 55158 39734 55172
rect 40610 55158 40692 55172
rect 40900 55158 40982 55172
rect 41858 55158 41940 55172
rect 42148 55158 42230 55172
rect 43106 55158 43188 55172
rect 43396 55158 43478 55172
rect 44354 55158 44436 55172
rect 44644 55158 44726 55172
rect 45602 55158 45684 55172
rect 45892 55158 45974 55172
rect 46850 55158 46932 55172
rect 47140 55158 47222 55172
rect 48098 55158 48180 55172
rect 48388 55158 48470 55172
rect 49346 55158 49428 55172
rect 49636 55158 49718 55172
rect 50594 55158 50676 55172
rect 50884 55158 50966 55172
rect 51842 55158 51924 55172
rect 52132 55158 52214 55172
rect 53090 55158 53172 55172
rect 53380 55158 53462 55172
rect 54338 55158 54420 55172
rect 54628 55158 54710 55172
rect 55586 55158 55668 55172
rect 55876 55158 55958 55172
rect 56834 55158 56916 55172
rect 57124 55158 57206 55172
rect 58082 55158 58164 55172
rect 58372 55158 58454 55172
rect 16418 55110 16864 55124
rect 17014 55110 17154 55124
rect 17304 55110 18112 55124
rect 18262 55110 18402 55124
rect 18552 55110 19360 55124
rect 19510 55110 19650 55124
rect 19800 55110 20608 55124
rect 20758 55110 20898 55124
rect 21048 55110 21856 55124
rect 22006 55110 22146 55124
rect 22296 55110 23104 55124
rect 23254 55110 23394 55124
rect 23544 55110 24352 55124
rect 24502 55110 24642 55124
rect 24792 55110 25600 55124
rect 25750 55110 25890 55124
rect 26040 55110 26848 55124
rect 26998 55110 27138 55124
rect 27288 55110 28096 55124
rect 28246 55110 28386 55124
rect 28536 55110 29344 55124
rect 29494 55110 29634 55124
rect 29784 55110 30592 55124
rect 30742 55110 30882 55124
rect 31032 55110 31840 55124
rect 31990 55110 32130 55124
rect 32280 55110 33088 55124
rect 33238 55110 33378 55124
rect 33528 55110 34336 55124
rect 34486 55110 34626 55124
rect 34776 55110 35584 55124
rect 35734 55110 35874 55124
rect 36024 55110 36832 55124
rect 36982 55110 37122 55124
rect 37272 55110 38080 55124
rect 38230 55110 38370 55124
rect 38520 55110 39328 55124
rect 39478 55110 39618 55124
rect 39768 55110 40576 55124
rect 40726 55110 40866 55124
rect 41016 55110 41824 55124
rect 41974 55110 42114 55124
rect 42264 55110 43072 55124
rect 43222 55110 43362 55124
rect 43512 55110 44320 55124
rect 44470 55110 44610 55124
rect 44760 55110 45568 55124
rect 45718 55110 45858 55124
rect 46008 55110 46816 55124
rect 46966 55110 47106 55124
rect 47256 55110 48064 55124
rect 48214 55110 48354 55124
rect 48504 55110 49312 55124
rect 49462 55110 49602 55124
rect 49752 55110 50560 55124
rect 50710 55110 50850 55124
rect 51000 55110 51808 55124
rect 51958 55110 52098 55124
rect 52248 55110 53056 55124
rect 53206 55110 53346 55124
rect 53496 55110 54304 55124
rect 54454 55110 54594 55124
rect 54744 55110 55552 55124
rect 55702 55110 55842 55124
rect 55992 55110 56800 55124
rect 56950 55110 57090 55124
rect 57240 55110 58048 55124
rect 58198 55110 58338 55124
rect 58488 55110 58934 55124
rect 16418 55062 58934 55110
rect 16418 55048 16864 55062
rect 17014 55048 17154 55062
rect 17304 55048 18112 55062
rect 18262 55048 18402 55062
rect 18552 55048 19360 55062
rect 19510 55048 19650 55062
rect 19800 55048 20608 55062
rect 20758 55048 20898 55062
rect 21048 55048 21856 55062
rect 22006 55048 22146 55062
rect 22296 55048 23104 55062
rect 23254 55048 23394 55062
rect 23544 55048 24352 55062
rect 24502 55048 24642 55062
rect 24792 55048 25600 55062
rect 25750 55048 25890 55062
rect 26040 55048 26848 55062
rect 26998 55048 27138 55062
rect 27288 55048 28096 55062
rect 28246 55048 28386 55062
rect 28536 55048 29344 55062
rect 29494 55048 29634 55062
rect 29784 55048 30592 55062
rect 30742 55048 30882 55062
rect 31032 55048 31840 55062
rect 31990 55048 32130 55062
rect 32280 55048 33088 55062
rect 33238 55048 33378 55062
rect 33528 55048 34336 55062
rect 34486 55048 34626 55062
rect 34776 55048 35584 55062
rect 35734 55048 35874 55062
rect 36024 55048 36832 55062
rect 36982 55048 37122 55062
rect 37272 55048 38080 55062
rect 38230 55048 38370 55062
rect 38520 55048 39328 55062
rect 39478 55048 39618 55062
rect 39768 55048 40576 55062
rect 40726 55048 40866 55062
rect 41016 55048 41824 55062
rect 41974 55048 42114 55062
rect 42264 55048 43072 55062
rect 43222 55048 43362 55062
rect 43512 55048 44320 55062
rect 44470 55048 44610 55062
rect 44760 55048 45568 55062
rect 45718 55048 45858 55062
rect 46008 55048 46816 55062
rect 46966 55048 47106 55062
rect 47256 55048 48064 55062
rect 48214 55048 48354 55062
rect 48504 55048 49312 55062
rect 49462 55048 49602 55062
rect 49752 55048 50560 55062
rect 50710 55048 50850 55062
rect 51000 55048 51808 55062
rect 51958 55048 52098 55062
rect 52248 55048 53056 55062
rect 53206 55048 53346 55062
rect 53496 55048 54304 55062
rect 54454 55048 54594 55062
rect 54744 55048 55552 55062
rect 55702 55048 55842 55062
rect 55992 55048 56800 55062
rect 56950 55048 57090 55062
rect 57240 55048 58048 55062
rect 58198 55048 58338 55062
rect 58488 55048 58934 55062
rect 16898 55000 16980 55014
rect 17188 55000 17270 55014
rect 18146 55000 18228 55014
rect 18436 55000 18518 55014
rect 19394 55000 19476 55014
rect 19684 55000 19766 55014
rect 20642 55000 20724 55014
rect 20932 55000 21014 55014
rect 21890 55000 21972 55014
rect 22180 55000 22262 55014
rect 23138 55000 23220 55014
rect 23428 55000 23510 55014
rect 24386 55000 24468 55014
rect 24676 55000 24758 55014
rect 25634 55000 25716 55014
rect 25924 55000 26006 55014
rect 26882 55000 26964 55014
rect 27172 55000 27254 55014
rect 28130 55000 28212 55014
rect 28420 55000 28502 55014
rect 29378 55000 29460 55014
rect 29668 55000 29750 55014
rect 30626 55000 30708 55014
rect 30916 55000 30998 55014
rect 31874 55000 31956 55014
rect 32164 55000 32246 55014
rect 33122 55000 33204 55014
rect 33412 55000 33494 55014
rect 34370 55000 34452 55014
rect 34660 55000 34742 55014
rect 35618 55000 35700 55014
rect 35908 55000 35990 55014
rect 36866 55000 36948 55014
rect 37156 55000 37238 55014
rect 38114 55000 38196 55014
rect 38404 55000 38486 55014
rect 39362 55000 39444 55014
rect 39652 55000 39734 55014
rect 40610 55000 40692 55014
rect 40900 55000 40982 55014
rect 41858 55000 41940 55014
rect 42148 55000 42230 55014
rect 43106 55000 43188 55014
rect 43396 55000 43478 55014
rect 44354 55000 44436 55014
rect 44644 55000 44726 55014
rect 45602 55000 45684 55014
rect 45892 55000 45974 55014
rect 46850 55000 46932 55014
rect 47140 55000 47222 55014
rect 48098 55000 48180 55014
rect 48388 55000 48470 55014
rect 49346 55000 49428 55014
rect 49636 55000 49718 55014
rect 50594 55000 50676 55014
rect 50884 55000 50966 55014
rect 51842 55000 51924 55014
rect 52132 55000 52214 55014
rect 53090 55000 53172 55014
rect 53380 55000 53462 55014
rect 54338 55000 54420 55014
rect 54628 55000 54710 55014
rect 55586 55000 55668 55014
rect 55876 55000 55958 55014
rect 56834 55000 56916 55014
rect 57124 55000 57206 55014
rect 58082 55000 58164 55014
rect 58372 55000 58454 55014
rect 16418 54952 58934 55000
rect 16418 54856 58934 54904
rect 16898 54842 16980 54856
rect 17188 54842 17270 54856
rect 18146 54842 18228 54856
rect 18436 54842 18518 54856
rect 19394 54842 19476 54856
rect 19684 54842 19766 54856
rect 20642 54842 20724 54856
rect 20932 54842 21014 54856
rect 21890 54842 21972 54856
rect 22180 54842 22262 54856
rect 23138 54842 23220 54856
rect 23428 54842 23510 54856
rect 24386 54842 24468 54856
rect 24676 54842 24758 54856
rect 25634 54842 25716 54856
rect 25924 54842 26006 54856
rect 26882 54842 26964 54856
rect 27172 54842 27254 54856
rect 28130 54842 28212 54856
rect 28420 54842 28502 54856
rect 29378 54842 29460 54856
rect 29668 54842 29750 54856
rect 30626 54842 30708 54856
rect 30916 54842 30998 54856
rect 31874 54842 31956 54856
rect 32164 54842 32246 54856
rect 33122 54842 33204 54856
rect 33412 54842 33494 54856
rect 34370 54842 34452 54856
rect 34660 54842 34742 54856
rect 35618 54842 35700 54856
rect 35908 54842 35990 54856
rect 36866 54842 36948 54856
rect 37156 54842 37238 54856
rect 38114 54842 38196 54856
rect 38404 54842 38486 54856
rect 39362 54842 39444 54856
rect 39652 54842 39734 54856
rect 40610 54842 40692 54856
rect 40900 54842 40982 54856
rect 41858 54842 41940 54856
rect 42148 54842 42230 54856
rect 43106 54842 43188 54856
rect 43396 54842 43478 54856
rect 44354 54842 44436 54856
rect 44644 54842 44726 54856
rect 45602 54842 45684 54856
rect 45892 54842 45974 54856
rect 46850 54842 46932 54856
rect 47140 54842 47222 54856
rect 48098 54842 48180 54856
rect 48388 54842 48470 54856
rect 49346 54842 49428 54856
rect 49636 54842 49718 54856
rect 50594 54842 50676 54856
rect 50884 54842 50966 54856
rect 51842 54842 51924 54856
rect 52132 54842 52214 54856
rect 53090 54842 53172 54856
rect 53380 54842 53462 54856
rect 54338 54842 54420 54856
rect 54628 54842 54710 54856
rect 55586 54842 55668 54856
rect 55876 54842 55958 54856
rect 56834 54842 56916 54856
rect 57124 54842 57206 54856
rect 58082 54842 58164 54856
rect 58372 54842 58454 54856
rect 16418 54794 16864 54808
rect 17014 54794 17154 54808
rect 17304 54794 18112 54808
rect 18262 54794 18402 54808
rect 18552 54794 19360 54808
rect 19510 54794 19650 54808
rect 19800 54794 20608 54808
rect 20758 54794 20898 54808
rect 21048 54794 21856 54808
rect 22006 54794 22146 54808
rect 22296 54794 23104 54808
rect 23254 54794 23394 54808
rect 23544 54794 24352 54808
rect 24502 54794 24642 54808
rect 24792 54794 25600 54808
rect 25750 54794 25890 54808
rect 26040 54794 26848 54808
rect 26998 54794 27138 54808
rect 27288 54794 28096 54808
rect 28246 54794 28386 54808
rect 28536 54794 29344 54808
rect 29494 54794 29634 54808
rect 29784 54794 30592 54808
rect 30742 54794 30882 54808
rect 31032 54794 31840 54808
rect 31990 54794 32130 54808
rect 32280 54794 33088 54808
rect 33238 54794 33378 54808
rect 33528 54794 34336 54808
rect 34486 54794 34626 54808
rect 34776 54794 35584 54808
rect 35734 54794 35874 54808
rect 36024 54794 36832 54808
rect 36982 54794 37122 54808
rect 37272 54794 38080 54808
rect 38230 54794 38370 54808
rect 38520 54794 39328 54808
rect 39478 54794 39618 54808
rect 39768 54794 40576 54808
rect 40726 54794 40866 54808
rect 41016 54794 41824 54808
rect 41974 54794 42114 54808
rect 42264 54794 43072 54808
rect 43222 54794 43362 54808
rect 43512 54794 44320 54808
rect 44470 54794 44610 54808
rect 44760 54794 45568 54808
rect 45718 54794 45858 54808
rect 46008 54794 46816 54808
rect 46966 54794 47106 54808
rect 47256 54794 48064 54808
rect 48214 54794 48354 54808
rect 48504 54794 49312 54808
rect 49462 54794 49602 54808
rect 49752 54794 50560 54808
rect 50710 54794 50850 54808
rect 51000 54794 51808 54808
rect 51958 54794 52098 54808
rect 52248 54794 53056 54808
rect 53206 54794 53346 54808
rect 53496 54794 54304 54808
rect 54454 54794 54594 54808
rect 54744 54794 55552 54808
rect 55702 54794 55842 54808
rect 55992 54794 56800 54808
rect 56950 54794 57090 54808
rect 57240 54794 58048 54808
rect 58198 54794 58338 54808
rect 58488 54794 58934 54808
rect 16418 54746 58934 54794
rect 16418 54732 16864 54746
rect 17014 54732 17154 54746
rect 17304 54732 18112 54746
rect 18262 54732 18402 54746
rect 18552 54732 19360 54746
rect 19510 54732 19650 54746
rect 19800 54732 20608 54746
rect 20758 54732 20898 54746
rect 21048 54732 21856 54746
rect 22006 54732 22146 54746
rect 22296 54732 23104 54746
rect 23254 54732 23394 54746
rect 23544 54732 24352 54746
rect 24502 54732 24642 54746
rect 24792 54732 25600 54746
rect 25750 54732 25890 54746
rect 26040 54732 26848 54746
rect 26998 54732 27138 54746
rect 27288 54732 28096 54746
rect 28246 54732 28386 54746
rect 28536 54732 29344 54746
rect 29494 54732 29634 54746
rect 29784 54732 30592 54746
rect 30742 54732 30882 54746
rect 31032 54732 31840 54746
rect 31990 54732 32130 54746
rect 32280 54732 33088 54746
rect 33238 54732 33378 54746
rect 33528 54732 34336 54746
rect 34486 54732 34626 54746
rect 34776 54732 35584 54746
rect 35734 54732 35874 54746
rect 36024 54732 36832 54746
rect 36982 54732 37122 54746
rect 37272 54732 38080 54746
rect 38230 54732 38370 54746
rect 38520 54732 39328 54746
rect 39478 54732 39618 54746
rect 39768 54732 40576 54746
rect 40726 54732 40866 54746
rect 41016 54732 41824 54746
rect 41974 54732 42114 54746
rect 42264 54732 43072 54746
rect 43222 54732 43362 54746
rect 43512 54732 44320 54746
rect 44470 54732 44610 54746
rect 44760 54732 45568 54746
rect 45718 54732 45858 54746
rect 46008 54732 46816 54746
rect 46966 54732 47106 54746
rect 47256 54732 48064 54746
rect 48214 54732 48354 54746
rect 48504 54732 49312 54746
rect 49462 54732 49602 54746
rect 49752 54732 50560 54746
rect 50710 54732 50850 54746
rect 51000 54732 51808 54746
rect 51958 54732 52098 54746
rect 52248 54732 53056 54746
rect 53206 54732 53346 54746
rect 53496 54732 54304 54746
rect 54454 54732 54594 54746
rect 54744 54732 55552 54746
rect 55702 54732 55842 54746
rect 55992 54732 56800 54746
rect 56950 54732 57090 54746
rect 57240 54732 58048 54746
rect 58198 54732 58338 54746
rect 58488 54732 58934 54746
rect 16898 54684 16980 54698
rect 17188 54684 17270 54698
rect 18146 54684 18228 54698
rect 18436 54684 18518 54698
rect 19394 54684 19476 54698
rect 19684 54684 19766 54698
rect 20642 54684 20724 54698
rect 20932 54684 21014 54698
rect 21890 54684 21972 54698
rect 22180 54684 22262 54698
rect 23138 54684 23220 54698
rect 23428 54684 23510 54698
rect 24386 54684 24468 54698
rect 24676 54684 24758 54698
rect 25634 54684 25716 54698
rect 25924 54684 26006 54698
rect 26882 54684 26964 54698
rect 27172 54684 27254 54698
rect 28130 54684 28212 54698
rect 28420 54684 28502 54698
rect 29378 54684 29460 54698
rect 29668 54684 29750 54698
rect 30626 54684 30708 54698
rect 30916 54684 30998 54698
rect 31874 54684 31956 54698
rect 32164 54684 32246 54698
rect 33122 54684 33204 54698
rect 33412 54684 33494 54698
rect 34370 54684 34452 54698
rect 34660 54684 34742 54698
rect 35618 54684 35700 54698
rect 35908 54684 35990 54698
rect 36866 54684 36948 54698
rect 37156 54684 37238 54698
rect 38114 54684 38196 54698
rect 38404 54684 38486 54698
rect 39362 54684 39444 54698
rect 39652 54684 39734 54698
rect 40610 54684 40692 54698
rect 40900 54684 40982 54698
rect 41858 54684 41940 54698
rect 42148 54684 42230 54698
rect 43106 54684 43188 54698
rect 43396 54684 43478 54698
rect 44354 54684 44436 54698
rect 44644 54684 44726 54698
rect 45602 54684 45684 54698
rect 45892 54684 45974 54698
rect 46850 54684 46932 54698
rect 47140 54684 47222 54698
rect 48098 54684 48180 54698
rect 48388 54684 48470 54698
rect 49346 54684 49428 54698
rect 49636 54684 49718 54698
rect 50594 54684 50676 54698
rect 50884 54684 50966 54698
rect 51842 54684 51924 54698
rect 52132 54684 52214 54698
rect 53090 54684 53172 54698
rect 53380 54684 53462 54698
rect 54338 54684 54420 54698
rect 54628 54684 54710 54698
rect 55586 54684 55668 54698
rect 55876 54684 55958 54698
rect 56834 54684 56916 54698
rect 57124 54684 57206 54698
rect 58082 54684 58164 54698
rect 58372 54684 58454 54698
rect 16418 54636 58934 54684
rect 16418 54478 58934 54588
rect 16418 54382 58934 54430
rect 16898 54368 16980 54382
rect 17188 54368 17270 54382
rect 18146 54368 18228 54382
rect 18436 54368 18518 54382
rect 19394 54368 19476 54382
rect 19684 54368 19766 54382
rect 20642 54368 20724 54382
rect 20932 54368 21014 54382
rect 21890 54368 21972 54382
rect 22180 54368 22262 54382
rect 23138 54368 23220 54382
rect 23428 54368 23510 54382
rect 24386 54368 24468 54382
rect 24676 54368 24758 54382
rect 25634 54368 25716 54382
rect 25924 54368 26006 54382
rect 26882 54368 26964 54382
rect 27172 54368 27254 54382
rect 28130 54368 28212 54382
rect 28420 54368 28502 54382
rect 29378 54368 29460 54382
rect 29668 54368 29750 54382
rect 30626 54368 30708 54382
rect 30916 54368 30998 54382
rect 31874 54368 31956 54382
rect 32164 54368 32246 54382
rect 33122 54368 33204 54382
rect 33412 54368 33494 54382
rect 34370 54368 34452 54382
rect 34660 54368 34742 54382
rect 35618 54368 35700 54382
rect 35908 54368 35990 54382
rect 36866 54368 36948 54382
rect 37156 54368 37238 54382
rect 38114 54368 38196 54382
rect 38404 54368 38486 54382
rect 39362 54368 39444 54382
rect 39652 54368 39734 54382
rect 40610 54368 40692 54382
rect 40900 54368 40982 54382
rect 41858 54368 41940 54382
rect 42148 54368 42230 54382
rect 43106 54368 43188 54382
rect 43396 54368 43478 54382
rect 44354 54368 44436 54382
rect 44644 54368 44726 54382
rect 45602 54368 45684 54382
rect 45892 54368 45974 54382
rect 46850 54368 46932 54382
rect 47140 54368 47222 54382
rect 48098 54368 48180 54382
rect 48388 54368 48470 54382
rect 49346 54368 49428 54382
rect 49636 54368 49718 54382
rect 50594 54368 50676 54382
rect 50884 54368 50966 54382
rect 51842 54368 51924 54382
rect 52132 54368 52214 54382
rect 53090 54368 53172 54382
rect 53380 54368 53462 54382
rect 54338 54368 54420 54382
rect 54628 54368 54710 54382
rect 55586 54368 55668 54382
rect 55876 54368 55958 54382
rect 56834 54368 56916 54382
rect 57124 54368 57206 54382
rect 58082 54368 58164 54382
rect 58372 54368 58454 54382
rect 16418 54320 16864 54334
rect 17014 54320 17154 54334
rect 17304 54320 18112 54334
rect 18262 54320 18402 54334
rect 18552 54320 19360 54334
rect 19510 54320 19650 54334
rect 19800 54320 20608 54334
rect 20758 54320 20898 54334
rect 21048 54320 21856 54334
rect 22006 54320 22146 54334
rect 22296 54320 23104 54334
rect 23254 54320 23394 54334
rect 23544 54320 24352 54334
rect 24502 54320 24642 54334
rect 24792 54320 25600 54334
rect 25750 54320 25890 54334
rect 26040 54320 26848 54334
rect 26998 54320 27138 54334
rect 27288 54320 28096 54334
rect 28246 54320 28386 54334
rect 28536 54320 29344 54334
rect 29494 54320 29634 54334
rect 29784 54320 30592 54334
rect 30742 54320 30882 54334
rect 31032 54320 31840 54334
rect 31990 54320 32130 54334
rect 32280 54320 33088 54334
rect 33238 54320 33378 54334
rect 33528 54320 34336 54334
rect 34486 54320 34626 54334
rect 34776 54320 35584 54334
rect 35734 54320 35874 54334
rect 36024 54320 36832 54334
rect 36982 54320 37122 54334
rect 37272 54320 38080 54334
rect 38230 54320 38370 54334
rect 38520 54320 39328 54334
rect 39478 54320 39618 54334
rect 39768 54320 40576 54334
rect 40726 54320 40866 54334
rect 41016 54320 41824 54334
rect 41974 54320 42114 54334
rect 42264 54320 43072 54334
rect 43222 54320 43362 54334
rect 43512 54320 44320 54334
rect 44470 54320 44610 54334
rect 44760 54320 45568 54334
rect 45718 54320 45858 54334
rect 46008 54320 46816 54334
rect 46966 54320 47106 54334
rect 47256 54320 48064 54334
rect 48214 54320 48354 54334
rect 48504 54320 49312 54334
rect 49462 54320 49602 54334
rect 49752 54320 50560 54334
rect 50710 54320 50850 54334
rect 51000 54320 51808 54334
rect 51958 54320 52098 54334
rect 52248 54320 53056 54334
rect 53206 54320 53346 54334
rect 53496 54320 54304 54334
rect 54454 54320 54594 54334
rect 54744 54320 55552 54334
rect 55702 54320 55842 54334
rect 55992 54320 56800 54334
rect 56950 54320 57090 54334
rect 57240 54320 58048 54334
rect 58198 54320 58338 54334
rect 58488 54320 58934 54334
rect 16418 54272 58934 54320
rect 16418 54258 16864 54272
rect 17014 54258 17154 54272
rect 17304 54258 18112 54272
rect 18262 54258 18402 54272
rect 18552 54258 19360 54272
rect 19510 54258 19650 54272
rect 19800 54258 20608 54272
rect 20758 54258 20898 54272
rect 21048 54258 21856 54272
rect 22006 54258 22146 54272
rect 22296 54258 23104 54272
rect 23254 54258 23394 54272
rect 23544 54258 24352 54272
rect 24502 54258 24642 54272
rect 24792 54258 25600 54272
rect 25750 54258 25890 54272
rect 26040 54258 26848 54272
rect 26998 54258 27138 54272
rect 27288 54258 28096 54272
rect 28246 54258 28386 54272
rect 28536 54258 29344 54272
rect 29494 54258 29634 54272
rect 29784 54258 30592 54272
rect 30742 54258 30882 54272
rect 31032 54258 31840 54272
rect 31990 54258 32130 54272
rect 32280 54258 33088 54272
rect 33238 54258 33378 54272
rect 33528 54258 34336 54272
rect 34486 54258 34626 54272
rect 34776 54258 35584 54272
rect 35734 54258 35874 54272
rect 36024 54258 36832 54272
rect 36982 54258 37122 54272
rect 37272 54258 38080 54272
rect 38230 54258 38370 54272
rect 38520 54258 39328 54272
rect 39478 54258 39618 54272
rect 39768 54258 40576 54272
rect 40726 54258 40866 54272
rect 41016 54258 41824 54272
rect 41974 54258 42114 54272
rect 42264 54258 43072 54272
rect 43222 54258 43362 54272
rect 43512 54258 44320 54272
rect 44470 54258 44610 54272
rect 44760 54258 45568 54272
rect 45718 54258 45858 54272
rect 46008 54258 46816 54272
rect 46966 54258 47106 54272
rect 47256 54258 48064 54272
rect 48214 54258 48354 54272
rect 48504 54258 49312 54272
rect 49462 54258 49602 54272
rect 49752 54258 50560 54272
rect 50710 54258 50850 54272
rect 51000 54258 51808 54272
rect 51958 54258 52098 54272
rect 52248 54258 53056 54272
rect 53206 54258 53346 54272
rect 53496 54258 54304 54272
rect 54454 54258 54594 54272
rect 54744 54258 55552 54272
rect 55702 54258 55842 54272
rect 55992 54258 56800 54272
rect 56950 54258 57090 54272
rect 57240 54258 58048 54272
rect 58198 54258 58338 54272
rect 58488 54258 58934 54272
rect 16898 54210 16980 54224
rect 17188 54210 17270 54224
rect 18146 54210 18228 54224
rect 18436 54210 18518 54224
rect 19394 54210 19476 54224
rect 19684 54210 19766 54224
rect 20642 54210 20724 54224
rect 20932 54210 21014 54224
rect 21890 54210 21972 54224
rect 22180 54210 22262 54224
rect 23138 54210 23220 54224
rect 23428 54210 23510 54224
rect 24386 54210 24468 54224
rect 24676 54210 24758 54224
rect 25634 54210 25716 54224
rect 25924 54210 26006 54224
rect 26882 54210 26964 54224
rect 27172 54210 27254 54224
rect 28130 54210 28212 54224
rect 28420 54210 28502 54224
rect 29378 54210 29460 54224
rect 29668 54210 29750 54224
rect 30626 54210 30708 54224
rect 30916 54210 30998 54224
rect 31874 54210 31956 54224
rect 32164 54210 32246 54224
rect 33122 54210 33204 54224
rect 33412 54210 33494 54224
rect 34370 54210 34452 54224
rect 34660 54210 34742 54224
rect 35618 54210 35700 54224
rect 35908 54210 35990 54224
rect 36866 54210 36948 54224
rect 37156 54210 37238 54224
rect 38114 54210 38196 54224
rect 38404 54210 38486 54224
rect 39362 54210 39444 54224
rect 39652 54210 39734 54224
rect 40610 54210 40692 54224
rect 40900 54210 40982 54224
rect 41858 54210 41940 54224
rect 42148 54210 42230 54224
rect 43106 54210 43188 54224
rect 43396 54210 43478 54224
rect 44354 54210 44436 54224
rect 44644 54210 44726 54224
rect 45602 54210 45684 54224
rect 45892 54210 45974 54224
rect 46850 54210 46932 54224
rect 47140 54210 47222 54224
rect 48098 54210 48180 54224
rect 48388 54210 48470 54224
rect 49346 54210 49428 54224
rect 49636 54210 49718 54224
rect 50594 54210 50676 54224
rect 50884 54210 50966 54224
rect 51842 54210 51924 54224
rect 52132 54210 52214 54224
rect 53090 54210 53172 54224
rect 53380 54210 53462 54224
rect 54338 54210 54420 54224
rect 54628 54210 54710 54224
rect 55586 54210 55668 54224
rect 55876 54210 55958 54224
rect 56834 54210 56916 54224
rect 57124 54210 57206 54224
rect 58082 54210 58164 54224
rect 58372 54210 58454 54224
rect 16418 54162 58934 54210
rect 16418 54066 58934 54114
rect 16898 54052 16980 54066
rect 17188 54052 17270 54066
rect 18146 54052 18228 54066
rect 18436 54052 18518 54066
rect 19394 54052 19476 54066
rect 19684 54052 19766 54066
rect 20642 54052 20724 54066
rect 20932 54052 21014 54066
rect 21890 54052 21972 54066
rect 22180 54052 22262 54066
rect 23138 54052 23220 54066
rect 23428 54052 23510 54066
rect 24386 54052 24468 54066
rect 24676 54052 24758 54066
rect 25634 54052 25716 54066
rect 25924 54052 26006 54066
rect 26882 54052 26964 54066
rect 27172 54052 27254 54066
rect 28130 54052 28212 54066
rect 28420 54052 28502 54066
rect 29378 54052 29460 54066
rect 29668 54052 29750 54066
rect 30626 54052 30708 54066
rect 30916 54052 30998 54066
rect 31874 54052 31956 54066
rect 32164 54052 32246 54066
rect 33122 54052 33204 54066
rect 33412 54052 33494 54066
rect 34370 54052 34452 54066
rect 34660 54052 34742 54066
rect 35618 54052 35700 54066
rect 35908 54052 35990 54066
rect 36866 54052 36948 54066
rect 37156 54052 37238 54066
rect 38114 54052 38196 54066
rect 38404 54052 38486 54066
rect 39362 54052 39444 54066
rect 39652 54052 39734 54066
rect 40610 54052 40692 54066
rect 40900 54052 40982 54066
rect 41858 54052 41940 54066
rect 42148 54052 42230 54066
rect 43106 54052 43188 54066
rect 43396 54052 43478 54066
rect 44354 54052 44436 54066
rect 44644 54052 44726 54066
rect 45602 54052 45684 54066
rect 45892 54052 45974 54066
rect 46850 54052 46932 54066
rect 47140 54052 47222 54066
rect 48098 54052 48180 54066
rect 48388 54052 48470 54066
rect 49346 54052 49428 54066
rect 49636 54052 49718 54066
rect 50594 54052 50676 54066
rect 50884 54052 50966 54066
rect 51842 54052 51924 54066
rect 52132 54052 52214 54066
rect 53090 54052 53172 54066
rect 53380 54052 53462 54066
rect 54338 54052 54420 54066
rect 54628 54052 54710 54066
rect 55586 54052 55668 54066
rect 55876 54052 55958 54066
rect 56834 54052 56916 54066
rect 57124 54052 57206 54066
rect 58082 54052 58164 54066
rect 58372 54052 58454 54066
rect 16418 54004 16864 54018
rect 17014 54004 17154 54018
rect 17304 54004 18112 54018
rect 18262 54004 18402 54018
rect 18552 54004 19360 54018
rect 19510 54004 19650 54018
rect 19800 54004 20608 54018
rect 20758 54004 20898 54018
rect 21048 54004 21856 54018
rect 22006 54004 22146 54018
rect 22296 54004 23104 54018
rect 23254 54004 23394 54018
rect 23544 54004 24352 54018
rect 24502 54004 24642 54018
rect 24792 54004 25600 54018
rect 25750 54004 25890 54018
rect 26040 54004 26848 54018
rect 26998 54004 27138 54018
rect 27288 54004 28096 54018
rect 28246 54004 28386 54018
rect 28536 54004 29344 54018
rect 29494 54004 29634 54018
rect 29784 54004 30592 54018
rect 30742 54004 30882 54018
rect 31032 54004 31840 54018
rect 31990 54004 32130 54018
rect 32280 54004 33088 54018
rect 33238 54004 33378 54018
rect 33528 54004 34336 54018
rect 34486 54004 34626 54018
rect 34776 54004 35584 54018
rect 35734 54004 35874 54018
rect 36024 54004 36832 54018
rect 36982 54004 37122 54018
rect 37272 54004 38080 54018
rect 38230 54004 38370 54018
rect 38520 54004 39328 54018
rect 39478 54004 39618 54018
rect 39768 54004 40576 54018
rect 40726 54004 40866 54018
rect 41016 54004 41824 54018
rect 41974 54004 42114 54018
rect 42264 54004 43072 54018
rect 43222 54004 43362 54018
rect 43512 54004 44320 54018
rect 44470 54004 44610 54018
rect 44760 54004 45568 54018
rect 45718 54004 45858 54018
rect 46008 54004 46816 54018
rect 46966 54004 47106 54018
rect 47256 54004 48064 54018
rect 48214 54004 48354 54018
rect 48504 54004 49312 54018
rect 49462 54004 49602 54018
rect 49752 54004 50560 54018
rect 50710 54004 50850 54018
rect 51000 54004 51808 54018
rect 51958 54004 52098 54018
rect 52248 54004 53056 54018
rect 53206 54004 53346 54018
rect 53496 54004 54304 54018
rect 54454 54004 54594 54018
rect 54744 54004 55552 54018
rect 55702 54004 55842 54018
rect 55992 54004 56800 54018
rect 56950 54004 57090 54018
rect 57240 54004 58048 54018
rect 58198 54004 58338 54018
rect 58488 54004 58934 54018
rect 16418 53956 58934 54004
rect 16418 53942 16864 53956
rect 17014 53942 17154 53956
rect 17304 53942 18112 53956
rect 18262 53942 18402 53956
rect 18552 53942 19360 53956
rect 19510 53942 19650 53956
rect 19800 53942 20608 53956
rect 20758 53942 20898 53956
rect 21048 53942 21856 53956
rect 22006 53942 22146 53956
rect 22296 53942 23104 53956
rect 23254 53942 23394 53956
rect 23544 53942 24352 53956
rect 24502 53942 24642 53956
rect 24792 53942 25600 53956
rect 25750 53942 25890 53956
rect 26040 53942 26848 53956
rect 26998 53942 27138 53956
rect 27288 53942 28096 53956
rect 28246 53942 28386 53956
rect 28536 53942 29344 53956
rect 29494 53942 29634 53956
rect 29784 53942 30592 53956
rect 30742 53942 30882 53956
rect 31032 53942 31840 53956
rect 31990 53942 32130 53956
rect 32280 53942 33088 53956
rect 33238 53942 33378 53956
rect 33528 53942 34336 53956
rect 34486 53942 34626 53956
rect 34776 53942 35584 53956
rect 35734 53942 35874 53956
rect 36024 53942 36832 53956
rect 36982 53942 37122 53956
rect 37272 53942 38080 53956
rect 38230 53942 38370 53956
rect 38520 53942 39328 53956
rect 39478 53942 39618 53956
rect 39768 53942 40576 53956
rect 40726 53942 40866 53956
rect 41016 53942 41824 53956
rect 41974 53942 42114 53956
rect 42264 53942 43072 53956
rect 43222 53942 43362 53956
rect 43512 53942 44320 53956
rect 44470 53942 44610 53956
rect 44760 53942 45568 53956
rect 45718 53942 45858 53956
rect 46008 53942 46816 53956
rect 46966 53942 47106 53956
rect 47256 53942 48064 53956
rect 48214 53942 48354 53956
rect 48504 53942 49312 53956
rect 49462 53942 49602 53956
rect 49752 53942 50560 53956
rect 50710 53942 50850 53956
rect 51000 53942 51808 53956
rect 51958 53942 52098 53956
rect 52248 53942 53056 53956
rect 53206 53942 53346 53956
rect 53496 53942 54304 53956
rect 54454 53942 54594 53956
rect 54744 53942 55552 53956
rect 55702 53942 55842 53956
rect 55992 53942 56800 53956
rect 56950 53942 57090 53956
rect 57240 53942 58048 53956
rect 58198 53942 58338 53956
rect 58488 53942 58934 53956
rect 16898 53894 16980 53908
rect 17188 53894 17270 53908
rect 18146 53894 18228 53908
rect 18436 53894 18518 53908
rect 19394 53894 19476 53908
rect 19684 53894 19766 53908
rect 20642 53894 20724 53908
rect 20932 53894 21014 53908
rect 21890 53894 21972 53908
rect 22180 53894 22262 53908
rect 23138 53894 23220 53908
rect 23428 53894 23510 53908
rect 24386 53894 24468 53908
rect 24676 53894 24758 53908
rect 25634 53894 25716 53908
rect 25924 53894 26006 53908
rect 26882 53894 26964 53908
rect 27172 53894 27254 53908
rect 28130 53894 28212 53908
rect 28420 53894 28502 53908
rect 29378 53894 29460 53908
rect 29668 53894 29750 53908
rect 30626 53894 30708 53908
rect 30916 53894 30998 53908
rect 31874 53894 31956 53908
rect 32164 53894 32246 53908
rect 33122 53894 33204 53908
rect 33412 53894 33494 53908
rect 34370 53894 34452 53908
rect 34660 53894 34742 53908
rect 35618 53894 35700 53908
rect 35908 53894 35990 53908
rect 36866 53894 36948 53908
rect 37156 53894 37238 53908
rect 38114 53894 38196 53908
rect 38404 53894 38486 53908
rect 39362 53894 39444 53908
rect 39652 53894 39734 53908
rect 40610 53894 40692 53908
rect 40900 53894 40982 53908
rect 41858 53894 41940 53908
rect 42148 53894 42230 53908
rect 43106 53894 43188 53908
rect 43396 53894 43478 53908
rect 44354 53894 44436 53908
rect 44644 53894 44726 53908
rect 45602 53894 45684 53908
rect 45892 53894 45974 53908
rect 46850 53894 46932 53908
rect 47140 53894 47222 53908
rect 48098 53894 48180 53908
rect 48388 53894 48470 53908
rect 49346 53894 49428 53908
rect 49636 53894 49718 53908
rect 50594 53894 50676 53908
rect 50884 53894 50966 53908
rect 51842 53894 51924 53908
rect 52132 53894 52214 53908
rect 53090 53894 53172 53908
rect 53380 53894 53462 53908
rect 54338 53894 54420 53908
rect 54628 53894 54710 53908
rect 55586 53894 55668 53908
rect 55876 53894 55958 53908
rect 56834 53894 56916 53908
rect 57124 53894 57206 53908
rect 58082 53894 58164 53908
rect 58372 53894 58454 53908
rect 16418 53846 58934 53894
rect 16418 53688 58934 53798
rect 16418 53592 58934 53640
rect 16898 53578 16980 53592
rect 17188 53578 17270 53592
rect 18146 53578 18228 53592
rect 18436 53578 18518 53592
rect 19394 53578 19476 53592
rect 19684 53578 19766 53592
rect 20642 53578 20724 53592
rect 20932 53578 21014 53592
rect 21890 53578 21972 53592
rect 22180 53578 22262 53592
rect 23138 53578 23220 53592
rect 23428 53578 23510 53592
rect 24386 53578 24468 53592
rect 24676 53578 24758 53592
rect 25634 53578 25716 53592
rect 25924 53578 26006 53592
rect 26882 53578 26964 53592
rect 27172 53578 27254 53592
rect 28130 53578 28212 53592
rect 28420 53578 28502 53592
rect 29378 53578 29460 53592
rect 29668 53578 29750 53592
rect 30626 53578 30708 53592
rect 30916 53578 30998 53592
rect 31874 53578 31956 53592
rect 32164 53578 32246 53592
rect 33122 53578 33204 53592
rect 33412 53578 33494 53592
rect 34370 53578 34452 53592
rect 34660 53578 34742 53592
rect 35618 53578 35700 53592
rect 35908 53578 35990 53592
rect 36866 53578 36948 53592
rect 37156 53578 37238 53592
rect 38114 53578 38196 53592
rect 38404 53578 38486 53592
rect 39362 53578 39444 53592
rect 39652 53578 39734 53592
rect 40610 53578 40692 53592
rect 40900 53578 40982 53592
rect 41858 53578 41940 53592
rect 42148 53578 42230 53592
rect 43106 53578 43188 53592
rect 43396 53578 43478 53592
rect 44354 53578 44436 53592
rect 44644 53578 44726 53592
rect 45602 53578 45684 53592
rect 45892 53578 45974 53592
rect 46850 53578 46932 53592
rect 47140 53578 47222 53592
rect 48098 53578 48180 53592
rect 48388 53578 48470 53592
rect 49346 53578 49428 53592
rect 49636 53578 49718 53592
rect 50594 53578 50676 53592
rect 50884 53578 50966 53592
rect 51842 53578 51924 53592
rect 52132 53578 52214 53592
rect 53090 53578 53172 53592
rect 53380 53578 53462 53592
rect 54338 53578 54420 53592
rect 54628 53578 54710 53592
rect 55586 53578 55668 53592
rect 55876 53578 55958 53592
rect 56834 53578 56916 53592
rect 57124 53578 57206 53592
rect 58082 53578 58164 53592
rect 58372 53578 58454 53592
rect 16418 53530 16864 53544
rect 17014 53530 17154 53544
rect 17304 53530 18112 53544
rect 18262 53530 18402 53544
rect 18552 53530 19360 53544
rect 19510 53530 19650 53544
rect 19800 53530 20608 53544
rect 20758 53530 20898 53544
rect 21048 53530 21856 53544
rect 22006 53530 22146 53544
rect 22296 53530 23104 53544
rect 23254 53530 23394 53544
rect 23544 53530 24352 53544
rect 24502 53530 24642 53544
rect 24792 53530 25600 53544
rect 25750 53530 25890 53544
rect 26040 53530 26848 53544
rect 26998 53530 27138 53544
rect 27288 53530 28096 53544
rect 28246 53530 28386 53544
rect 28536 53530 29344 53544
rect 29494 53530 29634 53544
rect 29784 53530 30592 53544
rect 30742 53530 30882 53544
rect 31032 53530 31840 53544
rect 31990 53530 32130 53544
rect 32280 53530 33088 53544
rect 33238 53530 33378 53544
rect 33528 53530 34336 53544
rect 34486 53530 34626 53544
rect 34776 53530 35584 53544
rect 35734 53530 35874 53544
rect 36024 53530 36832 53544
rect 36982 53530 37122 53544
rect 37272 53530 38080 53544
rect 38230 53530 38370 53544
rect 38520 53530 39328 53544
rect 39478 53530 39618 53544
rect 39768 53530 40576 53544
rect 40726 53530 40866 53544
rect 41016 53530 41824 53544
rect 41974 53530 42114 53544
rect 42264 53530 43072 53544
rect 43222 53530 43362 53544
rect 43512 53530 44320 53544
rect 44470 53530 44610 53544
rect 44760 53530 45568 53544
rect 45718 53530 45858 53544
rect 46008 53530 46816 53544
rect 46966 53530 47106 53544
rect 47256 53530 48064 53544
rect 48214 53530 48354 53544
rect 48504 53530 49312 53544
rect 49462 53530 49602 53544
rect 49752 53530 50560 53544
rect 50710 53530 50850 53544
rect 51000 53530 51808 53544
rect 51958 53530 52098 53544
rect 52248 53530 53056 53544
rect 53206 53530 53346 53544
rect 53496 53530 54304 53544
rect 54454 53530 54594 53544
rect 54744 53530 55552 53544
rect 55702 53530 55842 53544
rect 55992 53530 56800 53544
rect 56950 53530 57090 53544
rect 57240 53530 58048 53544
rect 58198 53530 58338 53544
rect 58488 53530 58934 53544
rect 16418 53482 58934 53530
rect 16418 53468 16864 53482
rect 17014 53468 17154 53482
rect 17304 53468 18112 53482
rect 18262 53468 18402 53482
rect 18552 53468 19360 53482
rect 19510 53468 19650 53482
rect 19800 53468 20608 53482
rect 20758 53468 20898 53482
rect 21048 53468 21856 53482
rect 22006 53468 22146 53482
rect 22296 53468 23104 53482
rect 23254 53468 23394 53482
rect 23544 53468 24352 53482
rect 24502 53468 24642 53482
rect 24792 53468 25600 53482
rect 25750 53468 25890 53482
rect 26040 53468 26848 53482
rect 26998 53468 27138 53482
rect 27288 53468 28096 53482
rect 28246 53468 28386 53482
rect 28536 53468 29344 53482
rect 29494 53468 29634 53482
rect 29784 53468 30592 53482
rect 30742 53468 30882 53482
rect 31032 53468 31840 53482
rect 31990 53468 32130 53482
rect 32280 53468 33088 53482
rect 33238 53468 33378 53482
rect 33528 53468 34336 53482
rect 34486 53468 34626 53482
rect 34776 53468 35584 53482
rect 35734 53468 35874 53482
rect 36024 53468 36832 53482
rect 36982 53468 37122 53482
rect 37272 53468 38080 53482
rect 38230 53468 38370 53482
rect 38520 53468 39328 53482
rect 39478 53468 39618 53482
rect 39768 53468 40576 53482
rect 40726 53468 40866 53482
rect 41016 53468 41824 53482
rect 41974 53468 42114 53482
rect 42264 53468 43072 53482
rect 43222 53468 43362 53482
rect 43512 53468 44320 53482
rect 44470 53468 44610 53482
rect 44760 53468 45568 53482
rect 45718 53468 45858 53482
rect 46008 53468 46816 53482
rect 46966 53468 47106 53482
rect 47256 53468 48064 53482
rect 48214 53468 48354 53482
rect 48504 53468 49312 53482
rect 49462 53468 49602 53482
rect 49752 53468 50560 53482
rect 50710 53468 50850 53482
rect 51000 53468 51808 53482
rect 51958 53468 52098 53482
rect 52248 53468 53056 53482
rect 53206 53468 53346 53482
rect 53496 53468 54304 53482
rect 54454 53468 54594 53482
rect 54744 53468 55552 53482
rect 55702 53468 55842 53482
rect 55992 53468 56800 53482
rect 56950 53468 57090 53482
rect 57240 53468 58048 53482
rect 58198 53468 58338 53482
rect 58488 53468 58934 53482
rect 16898 53420 16980 53434
rect 17188 53420 17270 53434
rect 18146 53420 18228 53434
rect 18436 53420 18518 53434
rect 19394 53420 19476 53434
rect 19684 53420 19766 53434
rect 20642 53420 20724 53434
rect 20932 53420 21014 53434
rect 21890 53420 21972 53434
rect 22180 53420 22262 53434
rect 23138 53420 23220 53434
rect 23428 53420 23510 53434
rect 24386 53420 24468 53434
rect 24676 53420 24758 53434
rect 25634 53420 25716 53434
rect 25924 53420 26006 53434
rect 26882 53420 26964 53434
rect 27172 53420 27254 53434
rect 28130 53420 28212 53434
rect 28420 53420 28502 53434
rect 29378 53420 29460 53434
rect 29668 53420 29750 53434
rect 30626 53420 30708 53434
rect 30916 53420 30998 53434
rect 31874 53420 31956 53434
rect 32164 53420 32246 53434
rect 33122 53420 33204 53434
rect 33412 53420 33494 53434
rect 34370 53420 34452 53434
rect 34660 53420 34742 53434
rect 35618 53420 35700 53434
rect 35908 53420 35990 53434
rect 36866 53420 36948 53434
rect 37156 53420 37238 53434
rect 38114 53420 38196 53434
rect 38404 53420 38486 53434
rect 39362 53420 39444 53434
rect 39652 53420 39734 53434
rect 40610 53420 40692 53434
rect 40900 53420 40982 53434
rect 41858 53420 41940 53434
rect 42148 53420 42230 53434
rect 43106 53420 43188 53434
rect 43396 53420 43478 53434
rect 44354 53420 44436 53434
rect 44644 53420 44726 53434
rect 45602 53420 45684 53434
rect 45892 53420 45974 53434
rect 46850 53420 46932 53434
rect 47140 53420 47222 53434
rect 48098 53420 48180 53434
rect 48388 53420 48470 53434
rect 49346 53420 49428 53434
rect 49636 53420 49718 53434
rect 50594 53420 50676 53434
rect 50884 53420 50966 53434
rect 51842 53420 51924 53434
rect 52132 53420 52214 53434
rect 53090 53420 53172 53434
rect 53380 53420 53462 53434
rect 54338 53420 54420 53434
rect 54628 53420 54710 53434
rect 55586 53420 55668 53434
rect 55876 53420 55958 53434
rect 56834 53420 56916 53434
rect 57124 53420 57206 53434
rect 58082 53420 58164 53434
rect 58372 53420 58454 53434
rect 16418 53372 58934 53420
rect 16418 53276 58934 53324
rect 16898 53262 16980 53276
rect 17188 53262 17270 53276
rect 18146 53262 18228 53276
rect 18436 53262 18518 53276
rect 19394 53262 19476 53276
rect 19684 53262 19766 53276
rect 20642 53262 20724 53276
rect 20932 53262 21014 53276
rect 21890 53262 21972 53276
rect 22180 53262 22262 53276
rect 23138 53262 23220 53276
rect 23428 53262 23510 53276
rect 24386 53262 24468 53276
rect 24676 53262 24758 53276
rect 25634 53262 25716 53276
rect 25924 53262 26006 53276
rect 26882 53262 26964 53276
rect 27172 53262 27254 53276
rect 28130 53262 28212 53276
rect 28420 53262 28502 53276
rect 29378 53262 29460 53276
rect 29668 53262 29750 53276
rect 30626 53262 30708 53276
rect 30916 53262 30998 53276
rect 31874 53262 31956 53276
rect 32164 53262 32246 53276
rect 33122 53262 33204 53276
rect 33412 53262 33494 53276
rect 34370 53262 34452 53276
rect 34660 53262 34742 53276
rect 35618 53262 35700 53276
rect 35908 53262 35990 53276
rect 36866 53262 36948 53276
rect 37156 53262 37238 53276
rect 38114 53262 38196 53276
rect 38404 53262 38486 53276
rect 39362 53262 39444 53276
rect 39652 53262 39734 53276
rect 40610 53262 40692 53276
rect 40900 53262 40982 53276
rect 41858 53262 41940 53276
rect 42148 53262 42230 53276
rect 43106 53262 43188 53276
rect 43396 53262 43478 53276
rect 44354 53262 44436 53276
rect 44644 53262 44726 53276
rect 45602 53262 45684 53276
rect 45892 53262 45974 53276
rect 46850 53262 46932 53276
rect 47140 53262 47222 53276
rect 48098 53262 48180 53276
rect 48388 53262 48470 53276
rect 49346 53262 49428 53276
rect 49636 53262 49718 53276
rect 50594 53262 50676 53276
rect 50884 53262 50966 53276
rect 51842 53262 51924 53276
rect 52132 53262 52214 53276
rect 53090 53262 53172 53276
rect 53380 53262 53462 53276
rect 54338 53262 54420 53276
rect 54628 53262 54710 53276
rect 55586 53262 55668 53276
rect 55876 53262 55958 53276
rect 56834 53262 56916 53276
rect 57124 53262 57206 53276
rect 58082 53262 58164 53276
rect 58372 53262 58454 53276
rect 16418 53214 16864 53228
rect 17014 53214 17154 53228
rect 17304 53214 18112 53228
rect 18262 53214 18402 53228
rect 18552 53214 19360 53228
rect 19510 53214 19650 53228
rect 19800 53214 20608 53228
rect 20758 53214 20898 53228
rect 21048 53214 21856 53228
rect 22006 53214 22146 53228
rect 22296 53214 23104 53228
rect 23254 53214 23394 53228
rect 23544 53214 24352 53228
rect 24502 53214 24642 53228
rect 24792 53214 25600 53228
rect 25750 53214 25890 53228
rect 26040 53214 26848 53228
rect 26998 53214 27138 53228
rect 27288 53214 28096 53228
rect 28246 53214 28386 53228
rect 28536 53214 29344 53228
rect 29494 53214 29634 53228
rect 29784 53214 30592 53228
rect 30742 53214 30882 53228
rect 31032 53214 31840 53228
rect 31990 53214 32130 53228
rect 32280 53214 33088 53228
rect 33238 53214 33378 53228
rect 33528 53214 34336 53228
rect 34486 53214 34626 53228
rect 34776 53214 35584 53228
rect 35734 53214 35874 53228
rect 36024 53214 36832 53228
rect 36982 53214 37122 53228
rect 37272 53214 38080 53228
rect 38230 53214 38370 53228
rect 38520 53214 39328 53228
rect 39478 53214 39618 53228
rect 39768 53214 40576 53228
rect 40726 53214 40866 53228
rect 41016 53214 41824 53228
rect 41974 53214 42114 53228
rect 42264 53214 43072 53228
rect 43222 53214 43362 53228
rect 43512 53214 44320 53228
rect 44470 53214 44610 53228
rect 44760 53214 45568 53228
rect 45718 53214 45858 53228
rect 46008 53214 46816 53228
rect 46966 53214 47106 53228
rect 47256 53214 48064 53228
rect 48214 53214 48354 53228
rect 48504 53214 49312 53228
rect 49462 53214 49602 53228
rect 49752 53214 50560 53228
rect 50710 53214 50850 53228
rect 51000 53214 51808 53228
rect 51958 53214 52098 53228
rect 52248 53214 53056 53228
rect 53206 53214 53346 53228
rect 53496 53214 54304 53228
rect 54454 53214 54594 53228
rect 54744 53214 55552 53228
rect 55702 53214 55842 53228
rect 55992 53214 56800 53228
rect 56950 53214 57090 53228
rect 57240 53214 58048 53228
rect 58198 53214 58338 53228
rect 58488 53214 58934 53228
rect 16418 53166 58934 53214
rect 16418 53152 16864 53166
rect 17014 53152 17154 53166
rect 17304 53152 18112 53166
rect 18262 53152 18402 53166
rect 18552 53152 19360 53166
rect 19510 53152 19650 53166
rect 19800 53152 20608 53166
rect 20758 53152 20898 53166
rect 21048 53152 21856 53166
rect 22006 53152 22146 53166
rect 22296 53152 23104 53166
rect 23254 53152 23394 53166
rect 23544 53152 24352 53166
rect 24502 53152 24642 53166
rect 24792 53152 25600 53166
rect 25750 53152 25890 53166
rect 26040 53152 26848 53166
rect 26998 53152 27138 53166
rect 27288 53152 28096 53166
rect 28246 53152 28386 53166
rect 28536 53152 29344 53166
rect 29494 53152 29634 53166
rect 29784 53152 30592 53166
rect 30742 53152 30882 53166
rect 31032 53152 31840 53166
rect 31990 53152 32130 53166
rect 32280 53152 33088 53166
rect 33238 53152 33378 53166
rect 33528 53152 34336 53166
rect 34486 53152 34626 53166
rect 34776 53152 35584 53166
rect 35734 53152 35874 53166
rect 36024 53152 36832 53166
rect 36982 53152 37122 53166
rect 37272 53152 38080 53166
rect 38230 53152 38370 53166
rect 38520 53152 39328 53166
rect 39478 53152 39618 53166
rect 39768 53152 40576 53166
rect 40726 53152 40866 53166
rect 41016 53152 41824 53166
rect 41974 53152 42114 53166
rect 42264 53152 43072 53166
rect 43222 53152 43362 53166
rect 43512 53152 44320 53166
rect 44470 53152 44610 53166
rect 44760 53152 45568 53166
rect 45718 53152 45858 53166
rect 46008 53152 46816 53166
rect 46966 53152 47106 53166
rect 47256 53152 48064 53166
rect 48214 53152 48354 53166
rect 48504 53152 49312 53166
rect 49462 53152 49602 53166
rect 49752 53152 50560 53166
rect 50710 53152 50850 53166
rect 51000 53152 51808 53166
rect 51958 53152 52098 53166
rect 52248 53152 53056 53166
rect 53206 53152 53346 53166
rect 53496 53152 54304 53166
rect 54454 53152 54594 53166
rect 54744 53152 55552 53166
rect 55702 53152 55842 53166
rect 55992 53152 56800 53166
rect 56950 53152 57090 53166
rect 57240 53152 58048 53166
rect 58198 53152 58338 53166
rect 58488 53152 58934 53166
rect 16898 53104 16980 53118
rect 17188 53104 17270 53118
rect 18146 53104 18228 53118
rect 18436 53104 18518 53118
rect 19394 53104 19476 53118
rect 19684 53104 19766 53118
rect 20642 53104 20724 53118
rect 20932 53104 21014 53118
rect 21890 53104 21972 53118
rect 22180 53104 22262 53118
rect 23138 53104 23220 53118
rect 23428 53104 23510 53118
rect 24386 53104 24468 53118
rect 24676 53104 24758 53118
rect 25634 53104 25716 53118
rect 25924 53104 26006 53118
rect 26882 53104 26964 53118
rect 27172 53104 27254 53118
rect 28130 53104 28212 53118
rect 28420 53104 28502 53118
rect 29378 53104 29460 53118
rect 29668 53104 29750 53118
rect 30626 53104 30708 53118
rect 30916 53104 30998 53118
rect 31874 53104 31956 53118
rect 32164 53104 32246 53118
rect 33122 53104 33204 53118
rect 33412 53104 33494 53118
rect 34370 53104 34452 53118
rect 34660 53104 34742 53118
rect 35618 53104 35700 53118
rect 35908 53104 35990 53118
rect 36866 53104 36948 53118
rect 37156 53104 37238 53118
rect 38114 53104 38196 53118
rect 38404 53104 38486 53118
rect 39362 53104 39444 53118
rect 39652 53104 39734 53118
rect 40610 53104 40692 53118
rect 40900 53104 40982 53118
rect 41858 53104 41940 53118
rect 42148 53104 42230 53118
rect 43106 53104 43188 53118
rect 43396 53104 43478 53118
rect 44354 53104 44436 53118
rect 44644 53104 44726 53118
rect 45602 53104 45684 53118
rect 45892 53104 45974 53118
rect 46850 53104 46932 53118
rect 47140 53104 47222 53118
rect 48098 53104 48180 53118
rect 48388 53104 48470 53118
rect 49346 53104 49428 53118
rect 49636 53104 49718 53118
rect 50594 53104 50676 53118
rect 50884 53104 50966 53118
rect 51842 53104 51924 53118
rect 52132 53104 52214 53118
rect 53090 53104 53172 53118
rect 53380 53104 53462 53118
rect 54338 53104 54420 53118
rect 54628 53104 54710 53118
rect 55586 53104 55668 53118
rect 55876 53104 55958 53118
rect 56834 53104 56916 53118
rect 57124 53104 57206 53118
rect 58082 53104 58164 53118
rect 58372 53104 58454 53118
rect 16418 53056 58934 53104
rect 16418 52898 58934 53008
rect 16418 52802 58934 52850
rect 16898 52788 16980 52802
rect 17188 52788 17270 52802
rect 18146 52788 18228 52802
rect 18436 52788 18518 52802
rect 19394 52788 19476 52802
rect 19684 52788 19766 52802
rect 20642 52788 20724 52802
rect 20932 52788 21014 52802
rect 21890 52788 21972 52802
rect 22180 52788 22262 52802
rect 23138 52788 23220 52802
rect 23428 52788 23510 52802
rect 24386 52788 24468 52802
rect 24676 52788 24758 52802
rect 25634 52788 25716 52802
rect 25924 52788 26006 52802
rect 26882 52788 26964 52802
rect 27172 52788 27254 52802
rect 28130 52788 28212 52802
rect 28420 52788 28502 52802
rect 29378 52788 29460 52802
rect 29668 52788 29750 52802
rect 30626 52788 30708 52802
rect 30916 52788 30998 52802
rect 31874 52788 31956 52802
rect 32164 52788 32246 52802
rect 33122 52788 33204 52802
rect 33412 52788 33494 52802
rect 34370 52788 34452 52802
rect 34660 52788 34742 52802
rect 35618 52788 35700 52802
rect 35908 52788 35990 52802
rect 36866 52788 36948 52802
rect 37156 52788 37238 52802
rect 38114 52788 38196 52802
rect 38404 52788 38486 52802
rect 39362 52788 39444 52802
rect 39652 52788 39734 52802
rect 40610 52788 40692 52802
rect 40900 52788 40982 52802
rect 41858 52788 41940 52802
rect 42148 52788 42230 52802
rect 43106 52788 43188 52802
rect 43396 52788 43478 52802
rect 44354 52788 44436 52802
rect 44644 52788 44726 52802
rect 45602 52788 45684 52802
rect 45892 52788 45974 52802
rect 46850 52788 46932 52802
rect 47140 52788 47222 52802
rect 48098 52788 48180 52802
rect 48388 52788 48470 52802
rect 49346 52788 49428 52802
rect 49636 52788 49718 52802
rect 50594 52788 50676 52802
rect 50884 52788 50966 52802
rect 51842 52788 51924 52802
rect 52132 52788 52214 52802
rect 53090 52788 53172 52802
rect 53380 52788 53462 52802
rect 54338 52788 54420 52802
rect 54628 52788 54710 52802
rect 55586 52788 55668 52802
rect 55876 52788 55958 52802
rect 56834 52788 56916 52802
rect 57124 52788 57206 52802
rect 58082 52788 58164 52802
rect 58372 52788 58454 52802
rect 16418 52740 16864 52754
rect 17014 52740 17154 52754
rect 17304 52740 18112 52754
rect 18262 52740 18402 52754
rect 18552 52740 19360 52754
rect 19510 52740 19650 52754
rect 19800 52740 20608 52754
rect 20758 52740 20898 52754
rect 21048 52740 21856 52754
rect 22006 52740 22146 52754
rect 22296 52740 23104 52754
rect 23254 52740 23394 52754
rect 23544 52740 24352 52754
rect 24502 52740 24642 52754
rect 24792 52740 25600 52754
rect 25750 52740 25890 52754
rect 26040 52740 26848 52754
rect 26998 52740 27138 52754
rect 27288 52740 28096 52754
rect 28246 52740 28386 52754
rect 28536 52740 29344 52754
rect 29494 52740 29634 52754
rect 29784 52740 30592 52754
rect 30742 52740 30882 52754
rect 31032 52740 31840 52754
rect 31990 52740 32130 52754
rect 32280 52740 33088 52754
rect 33238 52740 33378 52754
rect 33528 52740 34336 52754
rect 34486 52740 34626 52754
rect 34776 52740 35584 52754
rect 35734 52740 35874 52754
rect 36024 52740 36832 52754
rect 36982 52740 37122 52754
rect 37272 52740 38080 52754
rect 38230 52740 38370 52754
rect 38520 52740 39328 52754
rect 39478 52740 39618 52754
rect 39768 52740 40576 52754
rect 40726 52740 40866 52754
rect 41016 52740 41824 52754
rect 41974 52740 42114 52754
rect 42264 52740 43072 52754
rect 43222 52740 43362 52754
rect 43512 52740 44320 52754
rect 44470 52740 44610 52754
rect 44760 52740 45568 52754
rect 45718 52740 45858 52754
rect 46008 52740 46816 52754
rect 46966 52740 47106 52754
rect 47256 52740 48064 52754
rect 48214 52740 48354 52754
rect 48504 52740 49312 52754
rect 49462 52740 49602 52754
rect 49752 52740 50560 52754
rect 50710 52740 50850 52754
rect 51000 52740 51808 52754
rect 51958 52740 52098 52754
rect 52248 52740 53056 52754
rect 53206 52740 53346 52754
rect 53496 52740 54304 52754
rect 54454 52740 54594 52754
rect 54744 52740 55552 52754
rect 55702 52740 55842 52754
rect 55992 52740 56800 52754
rect 56950 52740 57090 52754
rect 57240 52740 58048 52754
rect 58198 52740 58338 52754
rect 58488 52740 58934 52754
rect 16418 52692 58934 52740
rect 16418 52678 16864 52692
rect 17014 52678 17154 52692
rect 17304 52678 18112 52692
rect 18262 52678 18402 52692
rect 18552 52678 19360 52692
rect 19510 52678 19650 52692
rect 19800 52678 20608 52692
rect 20758 52678 20898 52692
rect 21048 52678 21856 52692
rect 22006 52678 22146 52692
rect 22296 52678 23104 52692
rect 23254 52678 23394 52692
rect 23544 52678 24352 52692
rect 24502 52678 24642 52692
rect 24792 52678 25600 52692
rect 25750 52678 25890 52692
rect 26040 52678 26848 52692
rect 26998 52678 27138 52692
rect 27288 52678 28096 52692
rect 28246 52678 28386 52692
rect 28536 52678 29344 52692
rect 29494 52678 29634 52692
rect 29784 52678 30592 52692
rect 30742 52678 30882 52692
rect 31032 52678 31840 52692
rect 31990 52678 32130 52692
rect 32280 52678 33088 52692
rect 33238 52678 33378 52692
rect 33528 52678 34336 52692
rect 34486 52678 34626 52692
rect 34776 52678 35584 52692
rect 35734 52678 35874 52692
rect 36024 52678 36832 52692
rect 36982 52678 37122 52692
rect 37272 52678 38080 52692
rect 38230 52678 38370 52692
rect 38520 52678 39328 52692
rect 39478 52678 39618 52692
rect 39768 52678 40576 52692
rect 40726 52678 40866 52692
rect 41016 52678 41824 52692
rect 41974 52678 42114 52692
rect 42264 52678 43072 52692
rect 43222 52678 43362 52692
rect 43512 52678 44320 52692
rect 44470 52678 44610 52692
rect 44760 52678 45568 52692
rect 45718 52678 45858 52692
rect 46008 52678 46816 52692
rect 46966 52678 47106 52692
rect 47256 52678 48064 52692
rect 48214 52678 48354 52692
rect 48504 52678 49312 52692
rect 49462 52678 49602 52692
rect 49752 52678 50560 52692
rect 50710 52678 50850 52692
rect 51000 52678 51808 52692
rect 51958 52678 52098 52692
rect 52248 52678 53056 52692
rect 53206 52678 53346 52692
rect 53496 52678 54304 52692
rect 54454 52678 54594 52692
rect 54744 52678 55552 52692
rect 55702 52678 55842 52692
rect 55992 52678 56800 52692
rect 56950 52678 57090 52692
rect 57240 52678 58048 52692
rect 58198 52678 58338 52692
rect 58488 52678 58934 52692
rect 16898 52630 16980 52644
rect 17188 52630 17270 52644
rect 18146 52630 18228 52644
rect 18436 52630 18518 52644
rect 19394 52630 19476 52644
rect 19684 52630 19766 52644
rect 20642 52630 20724 52644
rect 20932 52630 21014 52644
rect 21890 52630 21972 52644
rect 22180 52630 22262 52644
rect 23138 52630 23220 52644
rect 23428 52630 23510 52644
rect 24386 52630 24468 52644
rect 24676 52630 24758 52644
rect 25634 52630 25716 52644
rect 25924 52630 26006 52644
rect 26882 52630 26964 52644
rect 27172 52630 27254 52644
rect 28130 52630 28212 52644
rect 28420 52630 28502 52644
rect 29378 52630 29460 52644
rect 29668 52630 29750 52644
rect 30626 52630 30708 52644
rect 30916 52630 30998 52644
rect 31874 52630 31956 52644
rect 32164 52630 32246 52644
rect 33122 52630 33204 52644
rect 33412 52630 33494 52644
rect 34370 52630 34452 52644
rect 34660 52630 34742 52644
rect 35618 52630 35700 52644
rect 35908 52630 35990 52644
rect 36866 52630 36948 52644
rect 37156 52630 37238 52644
rect 38114 52630 38196 52644
rect 38404 52630 38486 52644
rect 39362 52630 39444 52644
rect 39652 52630 39734 52644
rect 40610 52630 40692 52644
rect 40900 52630 40982 52644
rect 41858 52630 41940 52644
rect 42148 52630 42230 52644
rect 43106 52630 43188 52644
rect 43396 52630 43478 52644
rect 44354 52630 44436 52644
rect 44644 52630 44726 52644
rect 45602 52630 45684 52644
rect 45892 52630 45974 52644
rect 46850 52630 46932 52644
rect 47140 52630 47222 52644
rect 48098 52630 48180 52644
rect 48388 52630 48470 52644
rect 49346 52630 49428 52644
rect 49636 52630 49718 52644
rect 50594 52630 50676 52644
rect 50884 52630 50966 52644
rect 51842 52630 51924 52644
rect 52132 52630 52214 52644
rect 53090 52630 53172 52644
rect 53380 52630 53462 52644
rect 54338 52630 54420 52644
rect 54628 52630 54710 52644
rect 55586 52630 55668 52644
rect 55876 52630 55958 52644
rect 56834 52630 56916 52644
rect 57124 52630 57206 52644
rect 58082 52630 58164 52644
rect 58372 52630 58454 52644
rect 16418 52582 58934 52630
rect 16418 52486 58934 52534
rect 16898 52472 16980 52486
rect 17188 52472 17270 52486
rect 18146 52472 18228 52486
rect 18436 52472 18518 52486
rect 19394 52472 19476 52486
rect 19684 52472 19766 52486
rect 20642 52472 20724 52486
rect 20932 52472 21014 52486
rect 21890 52472 21972 52486
rect 22180 52472 22262 52486
rect 23138 52472 23220 52486
rect 23428 52472 23510 52486
rect 24386 52472 24468 52486
rect 24676 52472 24758 52486
rect 25634 52472 25716 52486
rect 25924 52472 26006 52486
rect 26882 52472 26964 52486
rect 27172 52472 27254 52486
rect 28130 52472 28212 52486
rect 28420 52472 28502 52486
rect 29378 52472 29460 52486
rect 29668 52472 29750 52486
rect 30626 52472 30708 52486
rect 30916 52472 30998 52486
rect 31874 52472 31956 52486
rect 32164 52472 32246 52486
rect 33122 52472 33204 52486
rect 33412 52472 33494 52486
rect 34370 52472 34452 52486
rect 34660 52472 34742 52486
rect 35618 52472 35700 52486
rect 35908 52472 35990 52486
rect 36866 52472 36948 52486
rect 37156 52472 37238 52486
rect 38114 52472 38196 52486
rect 38404 52472 38486 52486
rect 39362 52472 39444 52486
rect 39652 52472 39734 52486
rect 40610 52472 40692 52486
rect 40900 52472 40982 52486
rect 41858 52472 41940 52486
rect 42148 52472 42230 52486
rect 43106 52472 43188 52486
rect 43396 52472 43478 52486
rect 44354 52472 44436 52486
rect 44644 52472 44726 52486
rect 45602 52472 45684 52486
rect 45892 52472 45974 52486
rect 46850 52472 46932 52486
rect 47140 52472 47222 52486
rect 48098 52472 48180 52486
rect 48388 52472 48470 52486
rect 49346 52472 49428 52486
rect 49636 52472 49718 52486
rect 50594 52472 50676 52486
rect 50884 52472 50966 52486
rect 51842 52472 51924 52486
rect 52132 52472 52214 52486
rect 53090 52472 53172 52486
rect 53380 52472 53462 52486
rect 54338 52472 54420 52486
rect 54628 52472 54710 52486
rect 55586 52472 55668 52486
rect 55876 52472 55958 52486
rect 56834 52472 56916 52486
rect 57124 52472 57206 52486
rect 58082 52472 58164 52486
rect 58372 52472 58454 52486
rect 16418 52424 16864 52438
rect 17014 52424 17154 52438
rect 17304 52424 18112 52438
rect 18262 52424 18402 52438
rect 18552 52424 19360 52438
rect 19510 52424 19650 52438
rect 19800 52424 20608 52438
rect 20758 52424 20898 52438
rect 21048 52424 21856 52438
rect 22006 52424 22146 52438
rect 22296 52424 23104 52438
rect 23254 52424 23394 52438
rect 23544 52424 24352 52438
rect 24502 52424 24642 52438
rect 24792 52424 25600 52438
rect 25750 52424 25890 52438
rect 26040 52424 26848 52438
rect 26998 52424 27138 52438
rect 27288 52424 28096 52438
rect 28246 52424 28386 52438
rect 28536 52424 29344 52438
rect 29494 52424 29634 52438
rect 29784 52424 30592 52438
rect 30742 52424 30882 52438
rect 31032 52424 31840 52438
rect 31990 52424 32130 52438
rect 32280 52424 33088 52438
rect 33238 52424 33378 52438
rect 33528 52424 34336 52438
rect 34486 52424 34626 52438
rect 34776 52424 35584 52438
rect 35734 52424 35874 52438
rect 36024 52424 36832 52438
rect 36982 52424 37122 52438
rect 37272 52424 38080 52438
rect 38230 52424 38370 52438
rect 38520 52424 39328 52438
rect 39478 52424 39618 52438
rect 39768 52424 40576 52438
rect 40726 52424 40866 52438
rect 41016 52424 41824 52438
rect 41974 52424 42114 52438
rect 42264 52424 43072 52438
rect 43222 52424 43362 52438
rect 43512 52424 44320 52438
rect 44470 52424 44610 52438
rect 44760 52424 45568 52438
rect 45718 52424 45858 52438
rect 46008 52424 46816 52438
rect 46966 52424 47106 52438
rect 47256 52424 48064 52438
rect 48214 52424 48354 52438
rect 48504 52424 49312 52438
rect 49462 52424 49602 52438
rect 49752 52424 50560 52438
rect 50710 52424 50850 52438
rect 51000 52424 51808 52438
rect 51958 52424 52098 52438
rect 52248 52424 53056 52438
rect 53206 52424 53346 52438
rect 53496 52424 54304 52438
rect 54454 52424 54594 52438
rect 54744 52424 55552 52438
rect 55702 52424 55842 52438
rect 55992 52424 56800 52438
rect 56950 52424 57090 52438
rect 57240 52424 58048 52438
rect 58198 52424 58338 52438
rect 58488 52424 58934 52438
rect 16418 52376 58934 52424
rect 16418 52362 16864 52376
rect 17014 52362 17154 52376
rect 17304 52362 18112 52376
rect 18262 52362 18402 52376
rect 18552 52362 19360 52376
rect 19510 52362 19650 52376
rect 19800 52362 20608 52376
rect 20758 52362 20898 52376
rect 21048 52362 21856 52376
rect 22006 52362 22146 52376
rect 22296 52362 23104 52376
rect 23254 52362 23394 52376
rect 23544 52362 24352 52376
rect 24502 52362 24642 52376
rect 24792 52362 25600 52376
rect 25750 52362 25890 52376
rect 26040 52362 26848 52376
rect 26998 52362 27138 52376
rect 27288 52362 28096 52376
rect 28246 52362 28386 52376
rect 28536 52362 29344 52376
rect 29494 52362 29634 52376
rect 29784 52362 30592 52376
rect 30742 52362 30882 52376
rect 31032 52362 31840 52376
rect 31990 52362 32130 52376
rect 32280 52362 33088 52376
rect 33238 52362 33378 52376
rect 33528 52362 34336 52376
rect 34486 52362 34626 52376
rect 34776 52362 35584 52376
rect 35734 52362 35874 52376
rect 36024 52362 36832 52376
rect 36982 52362 37122 52376
rect 37272 52362 38080 52376
rect 38230 52362 38370 52376
rect 38520 52362 39328 52376
rect 39478 52362 39618 52376
rect 39768 52362 40576 52376
rect 40726 52362 40866 52376
rect 41016 52362 41824 52376
rect 41974 52362 42114 52376
rect 42264 52362 43072 52376
rect 43222 52362 43362 52376
rect 43512 52362 44320 52376
rect 44470 52362 44610 52376
rect 44760 52362 45568 52376
rect 45718 52362 45858 52376
rect 46008 52362 46816 52376
rect 46966 52362 47106 52376
rect 47256 52362 48064 52376
rect 48214 52362 48354 52376
rect 48504 52362 49312 52376
rect 49462 52362 49602 52376
rect 49752 52362 50560 52376
rect 50710 52362 50850 52376
rect 51000 52362 51808 52376
rect 51958 52362 52098 52376
rect 52248 52362 53056 52376
rect 53206 52362 53346 52376
rect 53496 52362 54304 52376
rect 54454 52362 54594 52376
rect 54744 52362 55552 52376
rect 55702 52362 55842 52376
rect 55992 52362 56800 52376
rect 56950 52362 57090 52376
rect 57240 52362 58048 52376
rect 58198 52362 58338 52376
rect 58488 52362 58934 52376
rect 16898 52314 16980 52328
rect 17188 52314 17270 52328
rect 18146 52314 18228 52328
rect 18436 52314 18518 52328
rect 19394 52314 19476 52328
rect 19684 52314 19766 52328
rect 20642 52314 20724 52328
rect 20932 52314 21014 52328
rect 21890 52314 21972 52328
rect 22180 52314 22262 52328
rect 23138 52314 23220 52328
rect 23428 52314 23510 52328
rect 24386 52314 24468 52328
rect 24676 52314 24758 52328
rect 25634 52314 25716 52328
rect 25924 52314 26006 52328
rect 26882 52314 26964 52328
rect 27172 52314 27254 52328
rect 28130 52314 28212 52328
rect 28420 52314 28502 52328
rect 29378 52314 29460 52328
rect 29668 52314 29750 52328
rect 30626 52314 30708 52328
rect 30916 52314 30998 52328
rect 31874 52314 31956 52328
rect 32164 52314 32246 52328
rect 33122 52314 33204 52328
rect 33412 52314 33494 52328
rect 34370 52314 34452 52328
rect 34660 52314 34742 52328
rect 35618 52314 35700 52328
rect 35908 52314 35990 52328
rect 36866 52314 36948 52328
rect 37156 52314 37238 52328
rect 38114 52314 38196 52328
rect 38404 52314 38486 52328
rect 39362 52314 39444 52328
rect 39652 52314 39734 52328
rect 40610 52314 40692 52328
rect 40900 52314 40982 52328
rect 41858 52314 41940 52328
rect 42148 52314 42230 52328
rect 43106 52314 43188 52328
rect 43396 52314 43478 52328
rect 44354 52314 44436 52328
rect 44644 52314 44726 52328
rect 45602 52314 45684 52328
rect 45892 52314 45974 52328
rect 46850 52314 46932 52328
rect 47140 52314 47222 52328
rect 48098 52314 48180 52328
rect 48388 52314 48470 52328
rect 49346 52314 49428 52328
rect 49636 52314 49718 52328
rect 50594 52314 50676 52328
rect 50884 52314 50966 52328
rect 51842 52314 51924 52328
rect 52132 52314 52214 52328
rect 53090 52314 53172 52328
rect 53380 52314 53462 52328
rect 54338 52314 54420 52328
rect 54628 52314 54710 52328
rect 55586 52314 55668 52328
rect 55876 52314 55958 52328
rect 56834 52314 56916 52328
rect 57124 52314 57206 52328
rect 58082 52314 58164 52328
rect 58372 52314 58454 52328
rect 16418 52266 58934 52314
rect 16418 52108 58934 52218
rect 16418 52012 58934 52060
rect 16898 51998 16980 52012
rect 17188 51998 17270 52012
rect 18146 51998 18228 52012
rect 18436 51998 18518 52012
rect 19394 51998 19476 52012
rect 19684 51998 19766 52012
rect 20642 51998 20724 52012
rect 20932 51998 21014 52012
rect 21890 51998 21972 52012
rect 22180 51998 22262 52012
rect 23138 51998 23220 52012
rect 23428 51998 23510 52012
rect 24386 51998 24468 52012
rect 24676 51998 24758 52012
rect 25634 51998 25716 52012
rect 25924 51998 26006 52012
rect 26882 51998 26964 52012
rect 27172 51998 27254 52012
rect 28130 51998 28212 52012
rect 28420 51998 28502 52012
rect 29378 51998 29460 52012
rect 29668 51998 29750 52012
rect 30626 51998 30708 52012
rect 30916 51998 30998 52012
rect 31874 51998 31956 52012
rect 32164 51998 32246 52012
rect 33122 51998 33204 52012
rect 33412 51998 33494 52012
rect 34370 51998 34452 52012
rect 34660 51998 34742 52012
rect 35618 51998 35700 52012
rect 35908 51998 35990 52012
rect 36866 51998 36948 52012
rect 37156 51998 37238 52012
rect 38114 51998 38196 52012
rect 38404 51998 38486 52012
rect 39362 51998 39444 52012
rect 39652 51998 39734 52012
rect 40610 51998 40692 52012
rect 40900 51998 40982 52012
rect 41858 51998 41940 52012
rect 42148 51998 42230 52012
rect 43106 51998 43188 52012
rect 43396 51998 43478 52012
rect 44354 51998 44436 52012
rect 44644 51998 44726 52012
rect 45602 51998 45684 52012
rect 45892 51998 45974 52012
rect 46850 51998 46932 52012
rect 47140 51998 47222 52012
rect 48098 51998 48180 52012
rect 48388 51998 48470 52012
rect 49346 51998 49428 52012
rect 49636 51998 49718 52012
rect 50594 51998 50676 52012
rect 50884 51998 50966 52012
rect 51842 51998 51924 52012
rect 52132 51998 52214 52012
rect 53090 51998 53172 52012
rect 53380 51998 53462 52012
rect 54338 51998 54420 52012
rect 54628 51998 54710 52012
rect 55586 51998 55668 52012
rect 55876 51998 55958 52012
rect 56834 51998 56916 52012
rect 57124 51998 57206 52012
rect 58082 51998 58164 52012
rect 58372 51998 58454 52012
rect 16418 51950 16864 51964
rect 17014 51950 17154 51964
rect 17304 51950 18112 51964
rect 18262 51950 18402 51964
rect 18552 51950 19360 51964
rect 19510 51950 19650 51964
rect 19800 51950 20608 51964
rect 20758 51950 20898 51964
rect 21048 51950 21856 51964
rect 22006 51950 22146 51964
rect 22296 51950 23104 51964
rect 23254 51950 23394 51964
rect 23544 51950 24352 51964
rect 24502 51950 24642 51964
rect 24792 51950 25600 51964
rect 25750 51950 25890 51964
rect 26040 51950 26848 51964
rect 26998 51950 27138 51964
rect 27288 51950 28096 51964
rect 28246 51950 28386 51964
rect 28536 51950 29344 51964
rect 29494 51950 29634 51964
rect 29784 51950 30592 51964
rect 30742 51950 30882 51964
rect 31032 51950 31840 51964
rect 31990 51950 32130 51964
rect 32280 51950 33088 51964
rect 33238 51950 33378 51964
rect 33528 51950 34336 51964
rect 34486 51950 34626 51964
rect 34776 51950 35584 51964
rect 35734 51950 35874 51964
rect 36024 51950 36832 51964
rect 36982 51950 37122 51964
rect 37272 51950 38080 51964
rect 38230 51950 38370 51964
rect 38520 51950 39328 51964
rect 39478 51950 39618 51964
rect 39768 51950 40576 51964
rect 40726 51950 40866 51964
rect 41016 51950 41824 51964
rect 41974 51950 42114 51964
rect 42264 51950 43072 51964
rect 43222 51950 43362 51964
rect 43512 51950 44320 51964
rect 44470 51950 44610 51964
rect 44760 51950 45568 51964
rect 45718 51950 45858 51964
rect 46008 51950 46816 51964
rect 46966 51950 47106 51964
rect 47256 51950 48064 51964
rect 48214 51950 48354 51964
rect 48504 51950 49312 51964
rect 49462 51950 49602 51964
rect 49752 51950 50560 51964
rect 50710 51950 50850 51964
rect 51000 51950 51808 51964
rect 51958 51950 52098 51964
rect 52248 51950 53056 51964
rect 53206 51950 53346 51964
rect 53496 51950 54304 51964
rect 54454 51950 54594 51964
rect 54744 51950 55552 51964
rect 55702 51950 55842 51964
rect 55992 51950 56800 51964
rect 56950 51950 57090 51964
rect 57240 51950 58048 51964
rect 58198 51950 58338 51964
rect 58488 51950 58934 51964
rect 16418 51902 58934 51950
rect 16418 51888 16864 51902
rect 17014 51888 17154 51902
rect 17304 51888 18112 51902
rect 18262 51888 18402 51902
rect 18552 51888 19360 51902
rect 19510 51888 19650 51902
rect 19800 51888 20608 51902
rect 20758 51888 20898 51902
rect 21048 51888 21856 51902
rect 22006 51888 22146 51902
rect 22296 51888 23104 51902
rect 23254 51888 23394 51902
rect 23544 51888 24352 51902
rect 24502 51888 24642 51902
rect 24792 51888 25600 51902
rect 25750 51888 25890 51902
rect 26040 51888 26848 51902
rect 26998 51888 27138 51902
rect 27288 51888 28096 51902
rect 28246 51888 28386 51902
rect 28536 51888 29344 51902
rect 29494 51888 29634 51902
rect 29784 51888 30592 51902
rect 30742 51888 30882 51902
rect 31032 51888 31840 51902
rect 31990 51888 32130 51902
rect 32280 51888 33088 51902
rect 33238 51888 33378 51902
rect 33528 51888 34336 51902
rect 34486 51888 34626 51902
rect 34776 51888 35584 51902
rect 35734 51888 35874 51902
rect 36024 51888 36832 51902
rect 36982 51888 37122 51902
rect 37272 51888 38080 51902
rect 38230 51888 38370 51902
rect 38520 51888 39328 51902
rect 39478 51888 39618 51902
rect 39768 51888 40576 51902
rect 40726 51888 40866 51902
rect 41016 51888 41824 51902
rect 41974 51888 42114 51902
rect 42264 51888 43072 51902
rect 43222 51888 43362 51902
rect 43512 51888 44320 51902
rect 44470 51888 44610 51902
rect 44760 51888 45568 51902
rect 45718 51888 45858 51902
rect 46008 51888 46816 51902
rect 46966 51888 47106 51902
rect 47256 51888 48064 51902
rect 48214 51888 48354 51902
rect 48504 51888 49312 51902
rect 49462 51888 49602 51902
rect 49752 51888 50560 51902
rect 50710 51888 50850 51902
rect 51000 51888 51808 51902
rect 51958 51888 52098 51902
rect 52248 51888 53056 51902
rect 53206 51888 53346 51902
rect 53496 51888 54304 51902
rect 54454 51888 54594 51902
rect 54744 51888 55552 51902
rect 55702 51888 55842 51902
rect 55992 51888 56800 51902
rect 56950 51888 57090 51902
rect 57240 51888 58048 51902
rect 58198 51888 58338 51902
rect 58488 51888 58934 51902
rect 16898 51840 16980 51854
rect 17188 51840 17270 51854
rect 18146 51840 18228 51854
rect 18436 51840 18518 51854
rect 19394 51840 19476 51854
rect 19684 51840 19766 51854
rect 20642 51840 20724 51854
rect 20932 51840 21014 51854
rect 21890 51840 21972 51854
rect 22180 51840 22262 51854
rect 23138 51840 23220 51854
rect 23428 51840 23510 51854
rect 24386 51840 24468 51854
rect 24676 51840 24758 51854
rect 25634 51840 25716 51854
rect 25924 51840 26006 51854
rect 26882 51840 26964 51854
rect 27172 51840 27254 51854
rect 28130 51840 28212 51854
rect 28420 51840 28502 51854
rect 29378 51840 29460 51854
rect 29668 51840 29750 51854
rect 30626 51840 30708 51854
rect 30916 51840 30998 51854
rect 31874 51840 31956 51854
rect 32164 51840 32246 51854
rect 33122 51840 33204 51854
rect 33412 51840 33494 51854
rect 34370 51840 34452 51854
rect 34660 51840 34742 51854
rect 35618 51840 35700 51854
rect 35908 51840 35990 51854
rect 36866 51840 36948 51854
rect 37156 51840 37238 51854
rect 38114 51840 38196 51854
rect 38404 51840 38486 51854
rect 39362 51840 39444 51854
rect 39652 51840 39734 51854
rect 40610 51840 40692 51854
rect 40900 51840 40982 51854
rect 41858 51840 41940 51854
rect 42148 51840 42230 51854
rect 43106 51840 43188 51854
rect 43396 51840 43478 51854
rect 44354 51840 44436 51854
rect 44644 51840 44726 51854
rect 45602 51840 45684 51854
rect 45892 51840 45974 51854
rect 46850 51840 46932 51854
rect 47140 51840 47222 51854
rect 48098 51840 48180 51854
rect 48388 51840 48470 51854
rect 49346 51840 49428 51854
rect 49636 51840 49718 51854
rect 50594 51840 50676 51854
rect 50884 51840 50966 51854
rect 51842 51840 51924 51854
rect 52132 51840 52214 51854
rect 53090 51840 53172 51854
rect 53380 51840 53462 51854
rect 54338 51840 54420 51854
rect 54628 51840 54710 51854
rect 55586 51840 55668 51854
rect 55876 51840 55958 51854
rect 56834 51840 56916 51854
rect 57124 51840 57206 51854
rect 58082 51840 58164 51854
rect 58372 51840 58454 51854
rect 16418 51792 58934 51840
rect 16418 51696 58934 51744
rect 16898 51682 16980 51696
rect 17188 51682 17270 51696
rect 18146 51682 18228 51696
rect 18436 51682 18518 51696
rect 19394 51682 19476 51696
rect 19684 51682 19766 51696
rect 20642 51682 20724 51696
rect 20932 51682 21014 51696
rect 21890 51682 21972 51696
rect 22180 51682 22262 51696
rect 23138 51682 23220 51696
rect 23428 51682 23510 51696
rect 24386 51682 24468 51696
rect 24676 51682 24758 51696
rect 25634 51682 25716 51696
rect 25924 51682 26006 51696
rect 26882 51682 26964 51696
rect 27172 51682 27254 51696
rect 28130 51682 28212 51696
rect 28420 51682 28502 51696
rect 29378 51682 29460 51696
rect 29668 51682 29750 51696
rect 30626 51682 30708 51696
rect 30916 51682 30998 51696
rect 31874 51682 31956 51696
rect 32164 51682 32246 51696
rect 33122 51682 33204 51696
rect 33412 51682 33494 51696
rect 34370 51682 34452 51696
rect 34660 51682 34742 51696
rect 35618 51682 35700 51696
rect 35908 51682 35990 51696
rect 36866 51682 36948 51696
rect 37156 51682 37238 51696
rect 38114 51682 38196 51696
rect 38404 51682 38486 51696
rect 39362 51682 39444 51696
rect 39652 51682 39734 51696
rect 40610 51682 40692 51696
rect 40900 51682 40982 51696
rect 41858 51682 41940 51696
rect 42148 51682 42230 51696
rect 43106 51682 43188 51696
rect 43396 51682 43478 51696
rect 44354 51682 44436 51696
rect 44644 51682 44726 51696
rect 45602 51682 45684 51696
rect 45892 51682 45974 51696
rect 46850 51682 46932 51696
rect 47140 51682 47222 51696
rect 48098 51682 48180 51696
rect 48388 51682 48470 51696
rect 49346 51682 49428 51696
rect 49636 51682 49718 51696
rect 50594 51682 50676 51696
rect 50884 51682 50966 51696
rect 51842 51682 51924 51696
rect 52132 51682 52214 51696
rect 53090 51682 53172 51696
rect 53380 51682 53462 51696
rect 54338 51682 54420 51696
rect 54628 51682 54710 51696
rect 55586 51682 55668 51696
rect 55876 51682 55958 51696
rect 56834 51682 56916 51696
rect 57124 51682 57206 51696
rect 58082 51682 58164 51696
rect 58372 51682 58454 51696
rect 16418 51634 16864 51648
rect 17014 51634 17154 51648
rect 17304 51634 18112 51648
rect 18262 51634 18402 51648
rect 18552 51634 19360 51648
rect 19510 51634 19650 51648
rect 19800 51634 20608 51648
rect 20758 51634 20898 51648
rect 21048 51634 21856 51648
rect 22006 51634 22146 51648
rect 22296 51634 23104 51648
rect 23254 51634 23394 51648
rect 23544 51634 24352 51648
rect 24502 51634 24642 51648
rect 24792 51634 25600 51648
rect 25750 51634 25890 51648
rect 26040 51634 26848 51648
rect 26998 51634 27138 51648
rect 27288 51634 28096 51648
rect 28246 51634 28386 51648
rect 28536 51634 29344 51648
rect 29494 51634 29634 51648
rect 29784 51634 30592 51648
rect 30742 51634 30882 51648
rect 31032 51634 31840 51648
rect 31990 51634 32130 51648
rect 32280 51634 33088 51648
rect 33238 51634 33378 51648
rect 33528 51634 34336 51648
rect 34486 51634 34626 51648
rect 34776 51634 35584 51648
rect 35734 51634 35874 51648
rect 36024 51634 36832 51648
rect 36982 51634 37122 51648
rect 37272 51634 38080 51648
rect 38230 51634 38370 51648
rect 38520 51634 39328 51648
rect 39478 51634 39618 51648
rect 39768 51634 40576 51648
rect 40726 51634 40866 51648
rect 41016 51634 41824 51648
rect 41974 51634 42114 51648
rect 42264 51634 43072 51648
rect 43222 51634 43362 51648
rect 43512 51634 44320 51648
rect 44470 51634 44610 51648
rect 44760 51634 45568 51648
rect 45718 51634 45858 51648
rect 46008 51634 46816 51648
rect 46966 51634 47106 51648
rect 47256 51634 48064 51648
rect 48214 51634 48354 51648
rect 48504 51634 49312 51648
rect 49462 51634 49602 51648
rect 49752 51634 50560 51648
rect 50710 51634 50850 51648
rect 51000 51634 51808 51648
rect 51958 51634 52098 51648
rect 52248 51634 53056 51648
rect 53206 51634 53346 51648
rect 53496 51634 54304 51648
rect 54454 51634 54594 51648
rect 54744 51634 55552 51648
rect 55702 51634 55842 51648
rect 55992 51634 56800 51648
rect 56950 51634 57090 51648
rect 57240 51634 58048 51648
rect 58198 51634 58338 51648
rect 58488 51634 58934 51648
rect 16418 51586 58934 51634
rect 16418 51572 16864 51586
rect 17014 51572 17154 51586
rect 17304 51572 18112 51586
rect 18262 51572 18402 51586
rect 18552 51572 19360 51586
rect 19510 51572 19650 51586
rect 19800 51572 20608 51586
rect 20758 51572 20898 51586
rect 21048 51572 21856 51586
rect 22006 51572 22146 51586
rect 22296 51572 23104 51586
rect 23254 51572 23394 51586
rect 23544 51572 24352 51586
rect 24502 51572 24642 51586
rect 24792 51572 25600 51586
rect 25750 51572 25890 51586
rect 26040 51572 26848 51586
rect 26998 51572 27138 51586
rect 27288 51572 28096 51586
rect 28246 51572 28386 51586
rect 28536 51572 29344 51586
rect 29494 51572 29634 51586
rect 29784 51572 30592 51586
rect 30742 51572 30882 51586
rect 31032 51572 31840 51586
rect 31990 51572 32130 51586
rect 32280 51572 33088 51586
rect 33238 51572 33378 51586
rect 33528 51572 34336 51586
rect 34486 51572 34626 51586
rect 34776 51572 35584 51586
rect 35734 51572 35874 51586
rect 36024 51572 36832 51586
rect 36982 51572 37122 51586
rect 37272 51572 38080 51586
rect 38230 51572 38370 51586
rect 38520 51572 39328 51586
rect 39478 51572 39618 51586
rect 39768 51572 40576 51586
rect 40726 51572 40866 51586
rect 41016 51572 41824 51586
rect 41974 51572 42114 51586
rect 42264 51572 43072 51586
rect 43222 51572 43362 51586
rect 43512 51572 44320 51586
rect 44470 51572 44610 51586
rect 44760 51572 45568 51586
rect 45718 51572 45858 51586
rect 46008 51572 46816 51586
rect 46966 51572 47106 51586
rect 47256 51572 48064 51586
rect 48214 51572 48354 51586
rect 48504 51572 49312 51586
rect 49462 51572 49602 51586
rect 49752 51572 50560 51586
rect 50710 51572 50850 51586
rect 51000 51572 51808 51586
rect 51958 51572 52098 51586
rect 52248 51572 53056 51586
rect 53206 51572 53346 51586
rect 53496 51572 54304 51586
rect 54454 51572 54594 51586
rect 54744 51572 55552 51586
rect 55702 51572 55842 51586
rect 55992 51572 56800 51586
rect 56950 51572 57090 51586
rect 57240 51572 58048 51586
rect 58198 51572 58338 51586
rect 58488 51572 58934 51586
rect 16898 51524 16980 51538
rect 17188 51524 17270 51538
rect 18146 51524 18228 51538
rect 18436 51524 18518 51538
rect 19394 51524 19476 51538
rect 19684 51524 19766 51538
rect 20642 51524 20724 51538
rect 20932 51524 21014 51538
rect 21890 51524 21972 51538
rect 22180 51524 22262 51538
rect 23138 51524 23220 51538
rect 23428 51524 23510 51538
rect 24386 51524 24468 51538
rect 24676 51524 24758 51538
rect 25634 51524 25716 51538
rect 25924 51524 26006 51538
rect 26882 51524 26964 51538
rect 27172 51524 27254 51538
rect 28130 51524 28212 51538
rect 28420 51524 28502 51538
rect 29378 51524 29460 51538
rect 29668 51524 29750 51538
rect 30626 51524 30708 51538
rect 30916 51524 30998 51538
rect 31874 51524 31956 51538
rect 32164 51524 32246 51538
rect 33122 51524 33204 51538
rect 33412 51524 33494 51538
rect 34370 51524 34452 51538
rect 34660 51524 34742 51538
rect 35618 51524 35700 51538
rect 35908 51524 35990 51538
rect 36866 51524 36948 51538
rect 37156 51524 37238 51538
rect 38114 51524 38196 51538
rect 38404 51524 38486 51538
rect 39362 51524 39444 51538
rect 39652 51524 39734 51538
rect 40610 51524 40692 51538
rect 40900 51524 40982 51538
rect 41858 51524 41940 51538
rect 42148 51524 42230 51538
rect 43106 51524 43188 51538
rect 43396 51524 43478 51538
rect 44354 51524 44436 51538
rect 44644 51524 44726 51538
rect 45602 51524 45684 51538
rect 45892 51524 45974 51538
rect 46850 51524 46932 51538
rect 47140 51524 47222 51538
rect 48098 51524 48180 51538
rect 48388 51524 48470 51538
rect 49346 51524 49428 51538
rect 49636 51524 49718 51538
rect 50594 51524 50676 51538
rect 50884 51524 50966 51538
rect 51842 51524 51924 51538
rect 52132 51524 52214 51538
rect 53090 51524 53172 51538
rect 53380 51524 53462 51538
rect 54338 51524 54420 51538
rect 54628 51524 54710 51538
rect 55586 51524 55668 51538
rect 55876 51524 55958 51538
rect 56834 51524 56916 51538
rect 57124 51524 57206 51538
rect 58082 51524 58164 51538
rect 58372 51524 58454 51538
rect 16418 51476 58934 51524
rect 16418 51318 58934 51428
rect 16418 51222 58934 51270
rect 16898 51208 16980 51222
rect 17188 51208 17270 51222
rect 18146 51208 18228 51222
rect 18436 51208 18518 51222
rect 19394 51208 19476 51222
rect 19684 51208 19766 51222
rect 20642 51208 20724 51222
rect 20932 51208 21014 51222
rect 21890 51208 21972 51222
rect 22180 51208 22262 51222
rect 23138 51208 23220 51222
rect 23428 51208 23510 51222
rect 24386 51208 24468 51222
rect 24676 51208 24758 51222
rect 25634 51208 25716 51222
rect 25924 51208 26006 51222
rect 26882 51208 26964 51222
rect 27172 51208 27254 51222
rect 28130 51208 28212 51222
rect 28420 51208 28502 51222
rect 29378 51208 29460 51222
rect 29668 51208 29750 51222
rect 30626 51208 30708 51222
rect 30916 51208 30998 51222
rect 31874 51208 31956 51222
rect 32164 51208 32246 51222
rect 33122 51208 33204 51222
rect 33412 51208 33494 51222
rect 34370 51208 34452 51222
rect 34660 51208 34742 51222
rect 35618 51208 35700 51222
rect 35908 51208 35990 51222
rect 36866 51208 36948 51222
rect 37156 51208 37238 51222
rect 38114 51208 38196 51222
rect 38404 51208 38486 51222
rect 39362 51208 39444 51222
rect 39652 51208 39734 51222
rect 40610 51208 40692 51222
rect 40900 51208 40982 51222
rect 41858 51208 41940 51222
rect 42148 51208 42230 51222
rect 43106 51208 43188 51222
rect 43396 51208 43478 51222
rect 44354 51208 44436 51222
rect 44644 51208 44726 51222
rect 45602 51208 45684 51222
rect 45892 51208 45974 51222
rect 46850 51208 46932 51222
rect 47140 51208 47222 51222
rect 48098 51208 48180 51222
rect 48388 51208 48470 51222
rect 49346 51208 49428 51222
rect 49636 51208 49718 51222
rect 50594 51208 50676 51222
rect 50884 51208 50966 51222
rect 51842 51208 51924 51222
rect 52132 51208 52214 51222
rect 53090 51208 53172 51222
rect 53380 51208 53462 51222
rect 54338 51208 54420 51222
rect 54628 51208 54710 51222
rect 55586 51208 55668 51222
rect 55876 51208 55958 51222
rect 56834 51208 56916 51222
rect 57124 51208 57206 51222
rect 58082 51208 58164 51222
rect 58372 51208 58454 51222
rect 16418 51160 16864 51174
rect 17014 51160 17154 51174
rect 17304 51160 18112 51174
rect 18262 51160 18402 51174
rect 18552 51160 19360 51174
rect 19510 51160 19650 51174
rect 19800 51160 20608 51174
rect 20758 51160 20898 51174
rect 21048 51160 21856 51174
rect 22006 51160 22146 51174
rect 22296 51160 23104 51174
rect 23254 51160 23394 51174
rect 23544 51160 24352 51174
rect 24502 51160 24642 51174
rect 24792 51160 25600 51174
rect 25750 51160 25890 51174
rect 26040 51160 26848 51174
rect 26998 51160 27138 51174
rect 27288 51160 28096 51174
rect 28246 51160 28386 51174
rect 28536 51160 29344 51174
rect 29494 51160 29634 51174
rect 29784 51160 30592 51174
rect 30742 51160 30882 51174
rect 31032 51160 31840 51174
rect 31990 51160 32130 51174
rect 32280 51160 33088 51174
rect 33238 51160 33378 51174
rect 33528 51160 34336 51174
rect 34486 51160 34626 51174
rect 34776 51160 35584 51174
rect 35734 51160 35874 51174
rect 36024 51160 36832 51174
rect 36982 51160 37122 51174
rect 37272 51160 38080 51174
rect 38230 51160 38370 51174
rect 38520 51160 39328 51174
rect 39478 51160 39618 51174
rect 39768 51160 40576 51174
rect 40726 51160 40866 51174
rect 41016 51160 41824 51174
rect 41974 51160 42114 51174
rect 42264 51160 43072 51174
rect 43222 51160 43362 51174
rect 43512 51160 44320 51174
rect 44470 51160 44610 51174
rect 44760 51160 45568 51174
rect 45718 51160 45858 51174
rect 46008 51160 46816 51174
rect 46966 51160 47106 51174
rect 47256 51160 48064 51174
rect 48214 51160 48354 51174
rect 48504 51160 49312 51174
rect 49462 51160 49602 51174
rect 49752 51160 50560 51174
rect 50710 51160 50850 51174
rect 51000 51160 51808 51174
rect 51958 51160 52098 51174
rect 52248 51160 53056 51174
rect 53206 51160 53346 51174
rect 53496 51160 54304 51174
rect 54454 51160 54594 51174
rect 54744 51160 55552 51174
rect 55702 51160 55842 51174
rect 55992 51160 56800 51174
rect 56950 51160 57090 51174
rect 57240 51160 58048 51174
rect 58198 51160 58338 51174
rect 58488 51160 58934 51174
rect 16418 51112 58934 51160
rect 16418 51098 16864 51112
rect 17014 51098 17154 51112
rect 17304 51098 18112 51112
rect 18262 51098 18402 51112
rect 18552 51098 19360 51112
rect 19510 51098 19650 51112
rect 19800 51098 20608 51112
rect 20758 51098 20898 51112
rect 21048 51098 21856 51112
rect 22006 51098 22146 51112
rect 22296 51098 23104 51112
rect 23254 51098 23394 51112
rect 23544 51098 24352 51112
rect 24502 51098 24642 51112
rect 24792 51098 25600 51112
rect 25750 51098 25890 51112
rect 26040 51098 26848 51112
rect 26998 51098 27138 51112
rect 27288 51098 28096 51112
rect 28246 51098 28386 51112
rect 28536 51098 29344 51112
rect 29494 51098 29634 51112
rect 29784 51098 30592 51112
rect 30742 51098 30882 51112
rect 31032 51098 31840 51112
rect 31990 51098 32130 51112
rect 32280 51098 33088 51112
rect 33238 51098 33378 51112
rect 33528 51098 34336 51112
rect 34486 51098 34626 51112
rect 34776 51098 35584 51112
rect 35734 51098 35874 51112
rect 36024 51098 36832 51112
rect 36982 51098 37122 51112
rect 37272 51098 38080 51112
rect 38230 51098 38370 51112
rect 38520 51098 39328 51112
rect 39478 51098 39618 51112
rect 39768 51098 40576 51112
rect 40726 51098 40866 51112
rect 41016 51098 41824 51112
rect 41974 51098 42114 51112
rect 42264 51098 43072 51112
rect 43222 51098 43362 51112
rect 43512 51098 44320 51112
rect 44470 51098 44610 51112
rect 44760 51098 45568 51112
rect 45718 51098 45858 51112
rect 46008 51098 46816 51112
rect 46966 51098 47106 51112
rect 47256 51098 48064 51112
rect 48214 51098 48354 51112
rect 48504 51098 49312 51112
rect 49462 51098 49602 51112
rect 49752 51098 50560 51112
rect 50710 51098 50850 51112
rect 51000 51098 51808 51112
rect 51958 51098 52098 51112
rect 52248 51098 53056 51112
rect 53206 51098 53346 51112
rect 53496 51098 54304 51112
rect 54454 51098 54594 51112
rect 54744 51098 55552 51112
rect 55702 51098 55842 51112
rect 55992 51098 56800 51112
rect 56950 51098 57090 51112
rect 57240 51098 58048 51112
rect 58198 51098 58338 51112
rect 58488 51098 58934 51112
rect 16898 51050 16980 51064
rect 17188 51050 17270 51064
rect 18146 51050 18228 51064
rect 18436 51050 18518 51064
rect 19394 51050 19476 51064
rect 19684 51050 19766 51064
rect 20642 51050 20724 51064
rect 20932 51050 21014 51064
rect 21890 51050 21972 51064
rect 22180 51050 22262 51064
rect 23138 51050 23220 51064
rect 23428 51050 23510 51064
rect 24386 51050 24468 51064
rect 24676 51050 24758 51064
rect 25634 51050 25716 51064
rect 25924 51050 26006 51064
rect 26882 51050 26964 51064
rect 27172 51050 27254 51064
rect 28130 51050 28212 51064
rect 28420 51050 28502 51064
rect 29378 51050 29460 51064
rect 29668 51050 29750 51064
rect 30626 51050 30708 51064
rect 30916 51050 30998 51064
rect 31874 51050 31956 51064
rect 32164 51050 32246 51064
rect 33122 51050 33204 51064
rect 33412 51050 33494 51064
rect 34370 51050 34452 51064
rect 34660 51050 34742 51064
rect 35618 51050 35700 51064
rect 35908 51050 35990 51064
rect 36866 51050 36948 51064
rect 37156 51050 37238 51064
rect 38114 51050 38196 51064
rect 38404 51050 38486 51064
rect 39362 51050 39444 51064
rect 39652 51050 39734 51064
rect 40610 51050 40692 51064
rect 40900 51050 40982 51064
rect 41858 51050 41940 51064
rect 42148 51050 42230 51064
rect 43106 51050 43188 51064
rect 43396 51050 43478 51064
rect 44354 51050 44436 51064
rect 44644 51050 44726 51064
rect 45602 51050 45684 51064
rect 45892 51050 45974 51064
rect 46850 51050 46932 51064
rect 47140 51050 47222 51064
rect 48098 51050 48180 51064
rect 48388 51050 48470 51064
rect 49346 51050 49428 51064
rect 49636 51050 49718 51064
rect 50594 51050 50676 51064
rect 50884 51050 50966 51064
rect 51842 51050 51924 51064
rect 52132 51050 52214 51064
rect 53090 51050 53172 51064
rect 53380 51050 53462 51064
rect 54338 51050 54420 51064
rect 54628 51050 54710 51064
rect 55586 51050 55668 51064
rect 55876 51050 55958 51064
rect 56834 51050 56916 51064
rect 57124 51050 57206 51064
rect 58082 51050 58164 51064
rect 58372 51050 58454 51064
rect 16418 51002 58934 51050
rect 16418 50906 58934 50954
rect 16898 50892 16980 50906
rect 17188 50892 17270 50906
rect 18146 50892 18228 50906
rect 18436 50892 18518 50906
rect 19394 50892 19476 50906
rect 19684 50892 19766 50906
rect 20642 50892 20724 50906
rect 20932 50892 21014 50906
rect 21890 50892 21972 50906
rect 22180 50892 22262 50906
rect 23138 50892 23220 50906
rect 23428 50892 23510 50906
rect 24386 50892 24468 50906
rect 24676 50892 24758 50906
rect 25634 50892 25716 50906
rect 25924 50892 26006 50906
rect 26882 50892 26964 50906
rect 27172 50892 27254 50906
rect 28130 50892 28212 50906
rect 28420 50892 28502 50906
rect 29378 50892 29460 50906
rect 29668 50892 29750 50906
rect 30626 50892 30708 50906
rect 30916 50892 30998 50906
rect 31874 50892 31956 50906
rect 32164 50892 32246 50906
rect 33122 50892 33204 50906
rect 33412 50892 33494 50906
rect 34370 50892 34452 50906
rect 34660 50892 34742 50906
rect 35618 50892 35700 50906
rect 35908 50892 35990 50906
rect 36866 50892 36948 50906
rect 37156 50892 37238 50906
rect 38114 50892 38196 50906
rect 38404 50892 38486 50906
rect 39362 50892 39444 50906
rect 39652 50892 39734 50906
rect 40610 50892 40692 50906
rect 40900 50892 40982 50906
rect 41858 50892 41940 50906
rect 42148 50892 42230 50906
rect 43106 50892 43188 50906
rect 43396 50892 43478 50906
rect 44354 50892 44436 50906
rect 44644 50892 44726 50906
rect 45602 50892 45684 50906
rect 45892 50892 45974 50906
rect 46850 50892 46932 50906
rect 47140 50892 47222 50906
rect 48098 50892 48180 50906
rect 48388 50892 48470 50906
rect 49346 50892 49428 50906
rect 49636 50892 49718 50906
rect 50594 50892 50676 50906
rect 50884 50892 50966 50906
rect 51842 50892 51924 50906
rect 52132 50892 52214 50906
rect 53090 50892 53172 50906
rect 53380 50892 53462 50906
rect 54338 50892 54420 50906
rect 54628 50892 54710 50906
rect 55586 50892 55668 50906
rect 55876 50892 55958 50906
rect 56834 50892 56916 50906
rect 57124 50892 57206 50906
rect 58082 50892 58164 50906
rect 58372 50892 58454 50906
rect 16418 50844 16864 50858
rect 17014 50844 17154 50858
rect 17304 50844 18112 50858
rect 18262 50844 18402 50858
rect 18552 50844 19360 50858
rect 19510 50844 19650 50858
rect 19800 50844 20608 50858
rect 20758 50844 20898 50858
rect 21048 50844 21856 50858
rect 22006 50844 22146 50858
rect 22296 50844 23104 50858
rect 23254 50844 23394 50858
rect 23544 50844 24352 50858
rect 24502 50844 24642 50858
rect 24792 50844 25600 50858
rect 25750 50844 25890 50858
rect 26040 50844 26848 50858
rect 26998 50844 27138 50858
rect 27288 50844 28096 50858
rect 28246 50844 28386 50858
rect 28536 50844 29344 50858
rect 29494 50844 29634 50858
rect 29784 50844 30592 50858
rect 30742 50844 30882 50858
rect 31032 50844 31840 50858
rect 31990 50844 32130 50858
rect 32280 50844 33088 50858
rect 33238 50844 33378 50858
rect 33528 50844 34336 50858
rect 34486 50844 34626 50858
rect 34776 50844 35584 50858
rect 35734 50844 35874 50858
rect 36024 50844 36832 50858
rect 36982 50844 37122 50858
rect 37272 50844 38080 50858
rect 38230 50844 38370 50858
rect 38520 50844 39328 50858
rect 39478 50844 39618 50858
rect 39768 50844 40576 50858
rect 40726 50844 40866 50858
rect 41016 50844 41824 50858
rect 41974 50844 42114 50858
rect 42264 50844 43072 50858
rect 43222 50844 43362 50858
rect 43512 50844 44320 50858
rect 44470 50844 44610 50858
rect 44760 50844 45568 50858
rect 45718 50844 45858 50858
rect 46008 50844 46816 50858
rect 46966 50844 47106 50858
rect 47256 50844 48064 50858
rect 48214 50844 48354 50858
rect 48504 50844 49312 50858
rect 49462 50844 49602 50858
rect 49752 50844 50560 50858
rect 50710 50844 50850 50858
rect 51000 50844 51808 50858
rect 51958 50844 52098 50858
rect 52248 50844 53056 50858
rect 53206 50844 53346 50858
rect 53496 50844 54304 50858
rect 54454 50844 54594 50858
rect 54744 50844 55552 50858
rect 55702 50844 55842 50858
rect 55992 50844 56800 50858
rect 56950 50844 57090 50858
rect 57240 50844 58048 50858
rect 58198 50844 58338 50858
rect 58488 50844 58934 50858
rect 16418 50796 58934 50844
rect 16418 50782 16864 50796
rect 17014 50782 17154 50796
rect 17304 50782 18112 50796
rect 18262 50782 18402 50796
rect 18552 50782 19360 50796
rect 19510 50782 19650 50796
rect 19800 50782 20608 50796
rect 20758 50782 20898 50796
rect 21048 50782 21856 50796
rect 22006 50782 22146 50796
rect 22296 50782 23104 50796
rect 23254 50782 23394 50796
rect 23544 50782 24352 50796
rect 24502 50782 24642 50796
rect 24792 50782 25600 50796
rect 25750 50782 25890 50796
rect 26040 50782 26848 50796
rect 26998 50782 27138 50796
rect 27288 50782 28096 50796
rect 28246 50782 28386 50796
rect 28536 50782 29344 50796
rect 29494 50782 29634 50796
rect 29784 50782 30592 50796
rect 30742 50782 30882 50796
rect 31032 50782 31840 50796
rect 31990 50782 32130 50796
rect 32280 50782 33088 50796
rect 33238 50782 33378 50796
rect 33528 50782 34336 50796
rect 34486 50782 34626 50796
rect 34776 50782 35584 50796
rect 35734 50782 35874 50796
rect 36024 50782 36832 50796
rect 36982 50782 37122 50796
rect 37272 50782 38080 50796
rect 38230 50782 38370 50796
rect 38520 50782 39328 50796
rect 39478 50782 39618 50796
rect 39768 50782 40576 50796
rect 40726 50782 40866 50796
rect 41016 50782 41824 50796
rect 41974 50782 42114 50796
rect 42264 50782 43072 50796
rect 43222 50782 43362 50796
rect 43512 50782 44320 50796
rect 44470 50782 44610 50796
rect 44760 50782 45568 50796
rect 45718 50782 45858 50796
rect 46008 50782 46816 50796
rect 46966 50782 47106 50796
rect 47256 50782 48064 50796
rect 48214 50782 48354 50796
rect 48504 50782 49312 50796
rect 49462 50782 49602 50796
rect 49752 50782 50560 50796
rect 50710 50782 50850 50796
rect 51000 50782 51808 50796
rect 51958 50782 52098 50796
rect 52248 50782 53056 50796
rect 53206 50782 53346 50796
rect 53496 50782 54304 50796
rect 54454 50782 54594 50796
rect 54744 50782 55552 50796
rect 55702 50782 55842 50796
rect 55992 50782 56800 50796
rect 56950 50782 57090 50796
rect 57240 50782 58048 50796
rect 58198 50782 58338 50796
rect 58488 50782 58934 50796
rect 16898 50734 16980 50748
rect 17188 50734 17270 50748
rect 18146 50734 18228 50748
rect 18436 50734 18518 50748
rect 19394 50734 19476 50748
rect 19684 50734 19766 50748
rect 20642 50734 20724 50748
rect 20932 50734 21014 50748
rect 21890 50734 21972 50748
rect 22180 50734 22262 50748
rect 23138 50734 23220 50748
rect 23428 50734 23510 50748
rect 24386 50734 24468 50748
rect 24676 50734 24758 50748
rect 25634 50734 25716 50748
rect 25924 50734 26006 50748
rect 26882 50734 26964 50748
rect 27172 50734 27254 50748
rect 28130 50734 28212 50748
rect 28420 50734 28502 50748
rect 29378 50734 29460 50748
rect 29668 50734 29750 50748
rect 30626 50734 30708 50748
rect 30916 50734 30998 50748
rect 31874 50734 31956 50748
rect 32164 50734 32246 50748
rect 33122 50734 33204 50748
rect 33412 50734 33494 50748
rect 34370 50734 34452 50748
rect 34660 50734 34742 50748
rect 35618 50734 35700 50748
rect 35908 50734 35990 50748
rect 36866 50734 36948 50748
rect 37156 50734 37238 50748
rect 38114 50734 38196 50748
rect 38404 50734 38486 50748
rect 39362 50734 39444 50748
rect 39652 50734 39734 50748
rect 40610 50734 40692 50748
rect 40900 50734 40982 50748
rect 41858 50734 41940 50748
rect 42148 50734 42230 50748
rect 43106 50734 43188 50748
rect 43396 50734 43478 50748
rect 44354 50734 44436 50748
rect 44644 50734 44726 50748
rect 45602 50734 45684 50748
rect 45892 50734 45974 50748
rect 46850 50734 46932 50748
rect 47140 50734 47222 50748
rect 48098 50734 48180 50748
rect 48388 50734 48470 50748
rect 49346 50734 49428 50748
rect 49636 50734 49718 50748
rect 50594 50734 50676 50748
rect 50884 50734 50966 50748
rect 51842 50734 51924 50748
rect 52132 50734 52214 50748
rect 53090 50734 53172 50748
rect 53380 50734 53462 50748
rect 54338 50734 54420 50748
rect 54628 50734 54710 50748
rect 55586 50734 55668 50748
rect 55876 50734 55958 50748
rect 56834 50734 56916 50748
rect 57124 50734 57206 50748
rect 58082 50734 58164 50748
rect 58372 50734 58454 50748
rect 16418 50686 58934 50734
rect 16418 50528 58934 50638
rect 16418 50432 58934 50480
rect 16898 50418 16980 50432
rect 17188 50418 17270 50432
rect 18146 50418 18228 50432
rect 18436 50418 18518 50432
rect 19394 50418 19476 50432
rect 19684 50418 19766 50432
rect 20642 50418 20724 50432
rect 20932 50418 21014 50432
rect 21890 50418 21972 50432
rect 22180 50418 22262 50432
rect 23138 50418 23220 50432
rect 23428 50418 23510 50432
rect 24386 50418 24468 50432
rect 24676 50418 24758 50432
rect 25634 50418 25716 50432
rect 25924 50418 26006 50432
rect 26882 50418 26964 50432
rect 27172 50418 27254 50432
rect 28130 50418 28212 50432
rect 28420 50418 28502 50432
rect 29378 50418 29460 50432
rect 29668 50418 29750 50432
rect 30626 50418 30708 50432
rect 30916 50418 30998 50432
rect 31874 50418 31956 50432
rect 32164 50418 32246 50432
rect 33122 50418 33204 50432
rect 33412 50418 33494 50432
rect 34370 50418 34452 50432
rect 34660 50418 34742 50432
rect 35618 50418 35700 50432
rect 35908 50418 35990 50432
rect 36866 50418 36948 50432
rect 37156 50418 37238 50432
rect 38114 50418 38196 50432
rect 38404 50418 38486 50432
rect 39362 50418 39444 50432
rect 39652 50418 39734 50432
rect 40610 50418 40692 50432
rect 40900 50418 40982 50432
rect 41858 50418 41940 50432
rect 42148 50418 42230 50432
rect 43106 50418 43188 50432
rect 43396 50418 43478 50432
rect 44354 50418 44436 50432
rect 44644 50418 44726 50432
rect 45602 50418 45684 50432
rect 45892 50418 45974 50432
rect 46850 50418 46932 50432
rect 47140 50418 47222 50432
rect 48098 50418 48180 50432
rect 48388 50418 48470 50432
rect 49346 50418 49428 50432
rect 49636 50418 49718 50432
rect 50594 50418 50676 50432
rect 50884 50418 50966 50432
rect 51842 50418 51924 50432
rect 52132 50418 52214 50432
rect 53090 50418 53172 50432
rect 53380 50418 53462 50432
rect 54338 50418 54420 50432
rect 54628 50418 54710 50432
rect 55586 50418 55668 50432
rect 55876 50418 55958 50432
rect 56834 50418 56916 50432
rect 57124 50418 57206 50432
rect 58082 50418 58164 50432
rect 58372 50418 58454 50432
rect 16418 50370 16864 50384
rect 17014 50370 17154 50384
rect 17304 50370 18112 50384
rect 18262 50370 18402 50384
rect 18552 50370 19360 50384
rect 19510 50370 19650 50384
rect 19800 50370 20608 50384
rect 20758 50370 20898 50384
rect 21048 50370 21856 50384
rect 22006 50370 22146 50384
rect 22296 50370 23104 50384
rect 23254 50370 23394 50384
rect 23544 50370 24352 50384
rect 24502 50370 24642 50384
rect 24792 50370 25600 50384
rect 25750 50370 25890 50384
rect 26040 50370 26848 50384
rect 26998 50370 27138 50384
rect 27288 50370 28096 50384
rect 28246 50370 28386 50384
rect 28536 50370 29344 50384
rect 29494 50370 29634 50384
rect 29784 50370 30592 50384
rect 30742 50370 30882 50384
rect 31032 50370 31840 50384
rect 31990 50370 32130 50384
rect 32280 50370 33088 50384
rect 33238 50370 33378 50384
rect 33528 50370 34336 50384
rect 34486 50370 34626 50384
rect 34776 50370 35584 50384
rect 35734 50370 35874 50384
rect 36024 50370 36832 50384
rect 36982 50370 37122 50384
rect 37272 50370 38080 50384
rect 38230 50370 38370 50384
rect 38520 50370 39328 50384
rect 39478 50370 39618 50384
rect 39768 50370 40576 50384
rect 40726 50370 40866 50384
rect 41016 50370 41824 50384
rect 41974 50370 42114 50384
rect 42264 50370 43072 50384
rect 43222 50370 43362 50384
rect 43512 50370 44320 50384
rect 44470 50370 44610 50384
rect 44760 50370 45568 50384
rect 45718 50370 45858 50384
rect 46008 50370 46816 50384
rect 46966 50370 47106 50384
rect 47256 50370 48064 50384
rect 48214 50370 48354 50384
rect 48504 50370 49312 50384
rect 49462 50370 49602 50384
rect 49752 50370 50560 50384
rect 50710 50370 50850 50384
rect 51000 50370 51808 50384
rect 51958 50370 52098 50384
rect 52248 50370 53056 50384
rect 53206 50370 53346 50384
rect 53496 50370 54304 50384
rect 54454 50370 54594 50384
rect 54744 50370 55552 50384
rect 55702 50370 55842 50384
rect 55992 50370 56800 50384
rect 56950 50370 57090 50384
rect 57240 50370 58048 50384
rect 58198 50370 58338 50384
rect 58488 50370 58934 50384
rect 16418 50322 58934 50370
rect 16418 50308 16864 50322
rect 17014 50308 17154 50322
rect 17304 50308 18112 50322
rect 18262 50308 18402 50322
rect 18552 50308 19360 50322
rect 19510 50308 19650 50322
rect 19800 50308 20608 50322
rect 20758 50308 20898 50322
rect 21048 50308 21856 50322
rect 22006 50308 22146 50322
rect 22296 50308 23104 50322
rect 23254 50308 23394 50322
rect 23544 50308 24352 50322
rect 24502 50308 24642 50322
rect 24792 50308 25600 50322
rect 25750 50308 25890 50322
rect 26040 50308 26848 50322
rect 26998 50308 27138 50322
rect 27288 50308 28096 50322
rect 28246 50308 28386 50322
rect 28536 50308 29344 50322
rect 29494 50308 29634 50322
rect 29784 50308 30592 50322
rect 30742 50308 30882 50322
rect 31032 50308 31840 50322
rect 31990 50308 32130 50322
rect 32280 50308 33088 50322
rect 33238 50308 33378 50322
rect 33528 50308 34336 50322
rect 34486 50308 34626 50322
rect 34776 50308 35584 50322
rect 35734 50308 35874 50322
rect 36024 50308 36832 50322
rect 36982 50308 37122 50322
rect 37272 50308 38080 50322
rect 38230 50308 38370 50322
rect 38520 50308 39328 50322
rect 39478 50308 39618 50322
rect 39768 50308 40576 50322
rect 40726 50308 40866 50322
rect 41016 50308 41824 50322
rect 41974 50308 42114 50322
rect 42264 50308 43072 50322
rect 43222 50308 43362 50322
rect 43512 50308 44320 50322
rect 44470 50308 44610 50322
rect 44760 50308 45568 50322
rect 45718 50308 45858 50322
rect 46008 50308 46816 50322
rect 46966 50308 47106 50322
rect 47256 50308 48064 50322
rect 48214 50308 48354 50322
rect 48504 50308 49312 50322
rect 49462 50308 49602 50322
rect 49752 50308 50560 50322
rect 50710 50308 50850 50322
rect 51000 50308 51808 50322
rect 51958 50308 52098 50322
rect 52248 50308 53056 50322
rect 53206 50308 53346 50322
rect 53496 50308 54304 50322
rect 54454 50308 54594 50322
rect 54744 50308 55552 50322
rect 55702 50308 55842 50322
rect 55992 50308 56800 50322
rect 56950 50308 57090 50322
rect 57240 50308 58048 50322
rect 58198 50308 58338 50322
rect 58488 50308 58934 50322
rect 16898 50260 16980 50274
rect 17188 50260 17270 50274
rect 18146 50260 18228 50274
rect 18436 50260 18518 50274
rect 19394 50260 19476 50274
rect 19684 50260 19766 50274
rect 20642 50260 20724 50274
rect 20932 50260 21014 50274
rect 21890 50260 21972 50274
rect 22180 50260 22262 50274
rect 23138 50260 23220 50274
rect 23428 50260 23510 50274
rect 24386 50260 24468 50274
rect 24676 50260 24758 50274
rect 25634 50260 25716 50274
rect 25924 50260 26006 50274
rect 26882 50260 26964 50274
rect 27172 50260 27254 50274
rect 28130 50260 28212 50274
rect 28420 50260 28502 50274
rect 29378 50260 29460 50274
rect 29668 50260 29750 50274
rect 30626 50260 30708 50274
rect 30916 50260 30998 50274
rect 31874 50260 31956 50274
rect 32164 50260 32246 50274
rect 33122 50260 33204 50274
rect 33412 50260 33494 50274
rect 34370 50260 34452 50274
rect 34660 50260 34742 50274
rect 35618 50260 35700 50274
rect 35908 50260 35990 50274
rect 36866 50260 36948 50274
rect 37156 50260 37238 50274
rect 38114 50260 38196 50274
rect 38404 50260 38486 50274
rect 39362 50260 39444 50274
rect 39652 50260 39734 50274
rect 40610 50260 40692 50274
rect 40900 50260 40982 50274
rect 41858 50260 41940 50274
rect 42148 50260 42230 50274
rect 43106 50260 43188 50274
rect 43396 50260 43478 50274
rect 44354 50260 44436 50274
rect 44644 50260 44726 50274
rect 45602 50260 45684 50274
rect 45892 50260 45974 50274
rect 46850 50260 46932 50274
rect 47140 50260 47222 50274
rect 48098 50260 48180 50274
rect 48388 50260 48470 50274
rect 49346 50260 49428 50274
rect 49636 50260 49718 50274
rect 50594 50260 50676 50274
rect 50884 50260 50966 50274
rect 51842 50260 51924 50274
rect 52132 50260 52214 50274
rect 53090 50260 53172 50274
rect 53380 50260 53462 50274
rect 54338 50260 54420 50274
rect 54628 50260 54710 50274
rect 55586 50260 55668 50274
rect 55876 50260 55958 50274
rect 56834 50260 56916 50274
rect 57124 50260 57206 50274
rect 58082 50260 58164 50274
rect 58372 50260 58454 50274
rect 16418 50212 58934 50260
rect 16418 50116 58934 50164
rect 16898 50102 16980 50116
rect 17188 50102 17270 50116
rect 18146 50102 18228 50116
rect 18436 50102 18518 50116
rect 19394 50102 19476 50116
rect 19684 50102 19766 50116
rect 20642 50102 20724 50116
rect 20932 50102 21014 50116
rect 21890 50102 21972 50116
rect 22180 50102 22262 50116
rect 23138 50102 23220 50116
rect 23428 50102 23510 50116
rect 24386 50102 24468 50116
rect 24676 50102 24758 50116
rect 25634 50102 25716 50116
rect 25924 50102 26006 50116
rect 26882 50102 26964 50116
rect 27172 50102 27254 50116
rect 28130 50102 28212 50116
rect 28420 50102 28502 50116
rect 29378 50102 29460 50116
rect 29668 50102 29750 50116
rect 30626 50102 30708 50116
rect 30916 50102 30998 50116
rect 31874 50102 31956 50116
rect 32164 50102 32246 50116
rect 33122 50102 33204 50116
rect 33412 50102 33494 50116
rect 34370 50102 34452 50116
rect 34660 50102 34742 50116
rect 35618 50102 35700 50116
rect 35908 50102 35990 50116
rect 36866 50102 36948 50116
rect 37156 50102 37238 50116
rect 38114 50102 38196 50116
rect 38404 50102 38486 50116
rect 39362 50102 39444 50116
rect 39652 50102 39734 50116
rect 40610 50102 40692 50116
rect 40900 50102 40982 50116
rect 41858 50102 41940 50116
rect 42148 50102 42230 50116
rect 43106 50102 43188 50116
rect 43396 50102 43478 50116
rect 44354 50102 44436 50116
rect 44644 50102 44726 50116
rect 45602 50102 45684 50116
rect 45892 50102 45974 50116
rect 46850 50102 46932 50116
rect 47140 50102 47222 50116
rect 48098 50102 48180 50116
rect 48388 50102 48470 50116
rect 49346 50102 49428 50116
rect 49636 50102 49718 50116
rect 50594 50102 50676 50116
rect 50884 50102 50966 50116
rect 51842 50102 51924 50116
rect 52132 50102 52214 50116
rect 53090 50102 53172 50116
rect 53380 50102 53462 50116
rect 54338 50102 54420 50116
rect 54628 50102 54710 50116
rect 55586 50102 55668 50116
rect 55876 50102 55958 50116
rect 56834 50102 56916 50116
rect 57124 50102 57206 50116
rect 58082 50102 58164 50116
rect 58372 50102 58454 50116
rect 16418 50054 16864 50068
rect 17014 50054 17154 50068
rect 17304 50054 18112 50068
rect 18262 50054 18402 50068
rect 18552 50054 19360 50068
rect 19510 50054 19650 50068
rect 19800 50054 20608 50068
rect 20758 50054 20898 50068
rect 21048 50054 21856 50068
rect 22006 50054 22146 50068
rect 22296 50054 23104 50068
rect 23254 50054 23394 50068
rect 23544 50054 24352 50068
rect 24502 50054 24642 50068
rect 24792 50054 25600 50068
rect 25750 50054 25890 50068
rect 26040 50054 26848 50068
rect 26998 50054 27138 50068
rect 27288 50054 28096 50068
rect 28246 50054 28386 50068
rect 28536 50054 29344 50068
rect 29494 50054 29634 50068
rect 29784 50054 30592 50068
rect 30742 50054 30882 50068
rect 31032 50054 31840 50068
rect 31990 50054 32130 50068
rect 32280 50054 33088 50068
rect 33238 50054 33378 50068
rect 33528 50054 34336 50068
rect 34486 50054 34626 50068
rect 34776 50054 35584 50068
rect 35734 50054 35874 50068
rect 36024 50054 36832 50068
rect 36982 50054 37122 50068
rect 37272 50054 38080 50068
rect 38230 50054 38370 50068
rect 38520 50054 39328 50068
rect 39478 50054 39618 50068
rect 39768 50054 40576 50068
rect 40726 50054 40866 50068
rect 41016 50054 41824 50068
rect 41974 50054 42114 50068
rect 42264 50054 43072 50068
rect 43222 50054 43362 50068
rect 43512 50054 44320 50068
rect 44470 50054 44610 50068
rect 44760 50054 45568 50068
rect 45718 50054 45858 50068
rect 46008 50054 46816 50068
rect 46966 50054 47106 50068
rect 47256 50054 48064 50068
rect 48214 50054 48354 50068
rect 48504 50054 49312 50068
rect 49462 50054 49602 50068
rect 49752 50054 50560 50068
rect 50710 50054 50850 50068
rect 51000 50054 51808 50068
rect 51958 50054 52098 50068
rect 52248 50054 53056 50068
rect 53206 50054 53346 50068
rect 53496 50054 54304 50068
rect 54454 50054 54594 50068
rect 54744 50054 55552 50068
rect 55702 50054 55842 50068
rect 55992 50054 56800 50068
rect 56950 50054 57090 50068
rect 57240 50054 58048 50068
rect 58198 50054 58338 50068
rect 58488 50054 58934 50068
rect 16418 50006 58934 50054
rect 16418 49992 16864 50006
rect 17014 49992 17154 50006
rect 17304 49992 18112 50006
rect 18262 49992 18402 50006
rect 18552 49992 19360 50006
rect 19510 49992 19650 50006
rect 19800 49992 20608 50006
rect 20758 49992 20898 50006
rect 21048 49992 21856 50006
rect 22006 49992 22146 50006
rect 22296 49992 23104 50006
rect 23254 49992 23394 50006
rect 23544 49992 24352 50006
rect 24502 49992 24642 50006
rect 24792 49992 25600 50006
rect 25750 49992 25890 50006
rect 26040 49992 26848 50006
rect 26998 49992 27138 50006
rect 27288 49992 28096 50006
rect 28246 49992 28386 50006
rect 28536 49992 29344 50006
rect 29494 49992 29634 50006
rect 29784 49992 30592 50006
rect 30742 49992 30882 50006
rect 31032 49992 31840 50006
rect 31990 49992 32130 50006
rect 32280 49992 33088 50006
rect 33238 49992 33378 50006
rect 33528 49992 34336 50006
rect 34486 49992 34626 50006
rect 34776 49992 35584 50006
rect 35734 49992 35874 50006
rect 36024 49992 36832 50006
rect 36982 49992 37122 50006
rect 37272 49992 38080 50006
rect 38230 49992 38370 50006
rect 38520 49992 39328 50006
rect 39478 49992 39618 50006
rect 39768 49992 40576 50006
rect 40726 49992 40866 50006
rect 41016 49992 41824 50006
rect 41974 49992 42114 50006
rect 42264 49992 43072 50006
rect 43222 49992 43362 50006
rect 43512 49992 44320 50006
rect 44470 49992 44610 50006
rect 44760 49992 45568 50006
rect 45718 49992 45858 50006
rect 46008 49992 46816 50006
rect 46966 49992 47106 50006
rect 47256 49992 48064 50006
rect 48214 49992 48354 50006
rect 48504 49992 49312 50006
rect 49462 49992 49602 50006
rect 49752 49992 50560 50006
rect 50710 49992 50850 50006
rect 51000 49992 51808 50006
rect 51958 49992 52098 50006
rect 52248 49992 53056 50006
rect 53206 49992 53346 50006
rect 53496 49992 54304 50006
rect 54454 49992 54594 50006
rect 54744 49992 55552 50006
rect 55702 49992 55842 50006
rect 55992 49992 56800 50006
rect 56950 49992 57090 50006
rect 57240 49992 58048 50006
rect 58198 49992 58338 50006
rect 58488 49992 58934 50006
rect 16898 49944 16980 49958
rect 17188 49944 17270 49958
rect 18146 49944 18228 49958
rect 18436 49944 18518 49958
rect 19394 49944 19476 49958
rect 19684 49944 19766 49958
rect 20642 49944 20724 49958
rect 20932 49944 21014 49958
rect 21890 49944 21972 49958
rect 22180 49944 22262 49958
rect 23138 49944 23220 49958
rect 23428 49944 23510 49958
rect 24386 49944 24468 49958
rect 24676 49944 24758 49958
rect 25634 49944 25716 49958
rect 25924 49944 26006 49958
rect 26882 49944 26964 49958
rect 27172 49944 27254 49958
rect 28130 49944 28212 49958
rect 28420 49944 28502 49958
rect 29378 49944 29460 49958
rect 29668 49944 29750 49958
rect 30626 49944 30708 49958
rect 30916 49944 30998 49958
rect 31874 49944 31956 49958
rect 32164 49944 32246 49958
rect 33122 49944 33204 49958
rect 33412 49944 33494 49958
rect 34370 49944 34452 49958
rect 34660 49944 34742 49958
rect 35618 49944 35700 49958
rect 35908 49944 35990 49958
rect 36866 49944 36948 49958
rect 37156 49944 37238 49958
rect 38114 49944 38196 49958
rect 38404 49944 38486 49958
rect 39362 49944 39444 49958
rect 39652 49944 39734 49958
rect 40610 49944 40692 49958
rect 40900 49944 40982 49958
rect 41858 49944 41940 49958
rect 42148 49944 42230 49958
rect 43106 49944 43188 49958
rect 43396 49944 43478 49958
rect 44354 49944 44436 49958
rect 44644 49944 44726 49958
rect 45602 49944 45684 49958
rect 45892 49944 45974 49958
rect 46850 49944 46932 49958
rect 47140 49944 47222 49958
rect 48098 49944 48180 49958
rect 48388 49944 48470 49958
rect 49346 49944 49428 49958
rect 49636 49944 49718 49958
rect 50594 49944 50676 49958
rect 50884 49944 50966 49958
rect 51842 49944 51924 49958
rect 52132 49944 52214 49958
rect 53090 49944 53172 49958
rect 53380 49944 53462 49958
rect 54338 49944 54420 49958
rect 54628 49944 54710 49958
rect 55586 49944 55668 49958
rect 55876 49944 55958 49958
rect 56834 49944 56916 49958
rect 57124 49944 57206 49958
rect 58082 49944 58164 49958
rect 58372 49944 58454 49958
rect 16418 49896 58934 49944
rect 16418 49738 58934 49848
rect 16418 49642 58934 49690
rect 16898 49628 16980 49642
rect 17188 49628 17270 49642
rect 18146 49628 18228 49642
rect 18436 49628 18518 49642
rect 19394 49628 19476 49642
rect 19684 49628 19766 49642
rect 20642 49628 20724 49642
rect 20932 49628 21014 49642
rect 21890 49628 21972 49642
rect 22180 49628 22262 49642
rect 23138 49628 23220 49642
rect 23428 49628 23510 49642
rect 24386 49628 24468 49642
rect 24676 49628 24758 49642
rect 25634 49628 25716 49642
rect 25924 49628 26006 49642
rect 26882 49628 26964 49642
rect 27172 49628 27254 49642
rect 28130 49628 28212 49642
rect 28420 49628 28502 49642
rect 29378 49628 29460 49642
rect 29668 49628 29750 49642
rect 30626 49628 30708 49642
rect 30916 49628 30998 49642
rect 31874 49628 31956 49642
rect 32164 49628 32246 49642
rect 33122 49628 33204 49642
rect 33412 49628 33494 49642
rect 34370 49628 34452 49642
rect 34660 49628 34742 49642
rect 35618 49628 35700 49642
rect 35908 49628 35990 49642
rect 36866 49628 36948 49642
rect 37156 49628 37238 49642
rect 38114 49628 38196 49642
rect 38404 49628 38486 49642
rect 39362 49628 39444 49642
rect 39652 49628 39734 49642
rect 40610 49628 40692 49642
rect 40900 49628 40982 49642
rect 41858 49628 41940 49642
rect 42148 49628 42230 49642
rect 43106 49628 43188 49642
rect 43396 49628 43478 49642
rect 44354 49628 44436 49642
rect 44644 49628 44726 49642
rect 45602 49628 45684 49642
rect 45892 49628 45974 49642
rect 46850 49628 46932 49642
rect 47140 49628 47222 49642
rect 48098 49628 48180 49642
rect 48388 49628 48470 49642
rect 49346 49628 49428 49642
rect 49636 49628 49718 49642
rect 50594 49628 50676 49642
rect 50884 49628 50966 49642
rect 51842 49628 51924 49642
rect 52132 49628 52214 49642
rect 53090 49628 53172 49642
rect 53380 49628 53462 49642
rect 54338 49628 54420 49642
rect 54628 49628 54710 49642
rect 55586 49628 55668 49642
rect 55876 49628 55958 49642
rect 56834 49628 56916 49642
rect 57124 49628 57206 49642
rect 58082 49628 58164 49642
rect 58372 49628 58454 49642
rect 16418 49580 16864 49594
rect 17014 49580 17154 49594
rect 17304 49580 18112 49594
rect 18262 49580 18402 49594
rect 18552 49580 19360 49594
rect 19510 49580 19650 49594
rect 19800 49580 20608 49594
rect 20758 49580 20898 49594
rect 21048 49580 21856 49594
rect 22006 49580 22146 49594
rect 22296 49580 23104 49594
rect 23254 49580 23394 49594
rect 23544 49580 24352 49594
rect 24502 49580 24642 49594
rect 24792 49580 25600 49594
rect 25750 49580 25890 49594
rect 26040 49580 26848 49594
rect 26998 49580 27138 49594
rect 27288 49580 28096 49594
rect 28246 49580 28386 49594
rect 28536 49580 29344 49594
rect 29494 49580 29634 49594
rect 29784 49580 30592 49594
rect 30742 49580 30882 49594
rect 31032 49580 31840 49594
rect 31990 49580 32130 49594
rect 32280 49580 33088 49594
rect 33238 49580 33378 49594
rect 33528 49580 34336 49594
rect 34486 49580 34626 49594
rect 34776 49580 35584 49594
rect 35734 49580 35874 49594
rect 36024 49580 36832 49594
rect 36982 49580 37122 49594
rect 37272 49580 38080 49594
rect 38230 49580 38370 49594
rect 38520 49580 39328 49594
rect 39478 49580 39618 49594
rect 39768 49580 40576 49594
rect 40726 49580 40866 49594
rect 41016 49580 41824 49594
rect 41974 49580 42114 49594
rect 42264 49580 43072 49594
rect 43222 49580 43362 49594
rect 43512 49580 44320 49594
rect 44470 49580 44610 49594
rect 44760 49580 45568 49594
rect 45718 49580 45858 49594
rect 46008 49580 46816 49594
rect 46966 49580 47106 49594
rect 47256 49580 48064 49594
rect 48214 49580 48354 49594
rect 48504 49580 49312 49594
rect 49462 49580 49602 49594
rect 49752 49580 50560 49594
rect 50710 49580 50850 49594
rect 51000 49580 51808 49594
rect 51958 49580 52098 49594
rect 52248 49580 53056 49594
rect 53206 49580 53346 49594
rect 53496 49580 54304 49594
rect 54454 49580 54594 49594
rect 54744 49580 55552 49594
rect 55702 49580 55842 49594
rect 55992 49580 56800 49594
rect 56950 49580 57090 49594
rect 57240 49580 58048 49594
rect 58198 49580 58338 49594
rect 58488 49580 58934 49594
rect 16418 49532 58934 49580
rect 16418 49518 16864 49532
rect 17014 49518 17154 49532
rect 17304 49518 18112 49532
rect 18262 49518 18402 49532
rect 18552 49518 19360 49532
rect 19510 49518 19650 49532
rect 19800 49518 20608 49532
rect 20758 49518 20898 49532
rect 21048 49518 21856 49532
rect 22006 49518 22146 49532
rect 22296 49518 23104 49532
rect 23254 49518 23394 49532
rect 23544 49518 24352 49532
rect 24502 49518 24642 49532
rect 24792 49518 25600 49532
rect 25750 49518 25890 49532
rect 26040 49518 26848 49532
rect 26998 49518 27138 49532
rect 27288 49518 28096 49532
rect 28246 49518 28386 49532
rect 28536 49518 29344 49532
rect 29494 49518 29634 49532
rect 29784 49518 30592 49532
rect 30742 49518 30882 49532
rect 31032 49518 31840 49532
rect 31990 49518 32130 49532
rect 32280 49518 33088 49532
rect 33238 49518 33378 49532
rect 33528 49518 34336 49532
rect 34486 49518 34626 49532
rect 34776 49518 35584 49532
rect 35734 49518 35874 49532
rect 36024 49518 36832 49532
rect 36982 49518 37122 49532
rect 37272 49518 38080 49532
rect 38230 49518 38370 49532
rect 38520 49518 39328 49532
rect 39478 49518 39618 49532
rect 39768 49518 40576 49532
rect 40726 49518 40866 49532
rect 41016 49518 41824 49532
rect 41974 49518 42114 49532
rect 42264 49518 43072 49532
rect 43222 49518 43362 49532
rect 43512 49518 44320 49532
rect 44470 49518 44610 49532
rect 44760 49518 45568 49532
rect 45718 49518 45858 49532
rect 46008 49518 46816 49532
rect 46966 49518 47106 49532
rect 47256 49518 48064 49532
rect 48214 49518 48354 49532
rect 48504 49518 49312 49532
rect 49462 49518 49602 49532
rect 49752 49518 50560 49532
rect 50710 49518 50850 49532
rect 51000 49518 51808 49532
rect 51958 49518 52098 49532
rect 52248 49518 53056 49532
rect 53206 49518 53346 49532
rect 53496 49518 54304 49532
rect 54454 49518 54594 49532
rect 54744 49518 55552 49532
rect 55702 49518 55842 49532
rect 55992 49518 56800 49532
rect 56950 49518 57090 49532
rect 57240 49518 58048 49532
rect 58198 49518 58338 49532
rect 58488 49518 58934 49532
rect 16898 49470 16980 49484
rect 17188 49470 17270 49484
rect 18146 49470 18228 49484
rect 18436 49470 18518 49484
rect 19394 49470 19476 49484
rect 19684 49470 19766 49484
rect 20642 49470 20724 49484
rect 20932 49470 21014 49484
rect 21890 49470 21972 49484
rect 22180 49470 22262 49484
rect 23138 49470 23220 49484
rect 23428 49470 23510 49484
rect 24386 49470 24468 49484
rect 24676 49470 24758 49484
rect 25634 49470 25716 49484
rect 25924 49470 26006 49484
rect 26882 49470 26964 49484
rect 27172 49470 27254 49484
rect 28130 49470 28212 49484
rect 28420 49470 28502 49484
rect 29378 49470 29460 49484
rect 29668 49470 29750 49484
rect 30626 49470 30708 49484
rect 30916 49470 30998 49484
rect 31874 49470 31956 49484
rect 32164 49470 32246 49484
rect 33122 49470 33204 49484
rect 33412 49470 33494 49484
rect 34370 49470 34452 49484
rect 34660 49470 34742 49484
rect 35618 49470 35700 49484
rect 35908 49470 35990 49484
rect 36866 49470 36948 49484
rect 37156 49470 37238 49484
rect 38114 49470 38196 49484
rect 38404 49470 38486 49484
rect 39362 49470 39444 49484
rect 39652 49470 39734 49484
rect 40610 49470 40692 49484
rect 40900 49470 40982 49484
rect 41858 49470 41940 49484
rect 42148 49470 42230 49484
rect 43106 49470 43188 49484
rect 43396 49470 43478 49484
rect 44354 49470 44436 49484
rect 44644 49470 44726 49484
rect 45602 49470 45684 49484
rect 45892 49470 45974 49484
rect 46850 49470 46932 49484
rect 47140 49470 47222 49484
rect 48098 49470 48180 49484
rect 48388 49470 48470 49484
rect 49346 49470 49428 49484
rect 49636 49470 49718 49484
rect 50594 49470 50676 49484
rect 50884 49470 50966 49484
rect 51842 49470 51924 49484
rect 52132 49470 52214 49484
rect 53090 49470 53172 49484
rect 53380 49470 53462 49484
rect 54338 49470 54420 49484
rect 54628 49470 54710 49484
rect 55586 49470 55668 49484
rect 55876 49470 55958 49484
rect 56834 49470 56916 49484
rect 57124 49470 57206 49484
rect 58082 49470 58164 49484
rect 58372 49470 58454 49484
rect 16418 49422 58934 49470
rect 16418 49326 58934 49374
rect 16898 49312 16980 49326
rect 17188 49312 17270 49326
rect 18146 49312 18228 49326
rect 18436 49312 18518 49326
rect 19394 49312 19476 49326
rect 19684 49312 19766 49326
rect 20642 49312 20724 49326
rect 20932 49312 21014 49326
rect 21890 49312 21972 49326
rect 22180 49312 22262 49326
rect 23138 49312 23220 49326
rect 23428 49312 23510 49326
rect 24386 49312 24468 49326
rect 24676 49312 24758 49326
rect 25634 49312 25716 49326
rect 25924 49312 26006 49326
rect 26882 49312 26964 49326
rect 27172 49312 27254 49326
rect 28130 49312 28212 49326
rect 28420 49312 28502 49326
rect 29378 49312 29460 49326
rect 29668 49312 29750 49326
rect 30626 49312 30708 49326
rect 30916 49312 30998 49326
rect 31874 49312 31956 49326
rect 32164 49312 32246 49326
rect 33122 49312 33204 49326
rect 33412 49312 33494 49326
rect 34370 49312 34452 49326
rect 34660 49312 34742 49326
rect 35618 49312 35700 49326
rect 35908 49312 35990 49326
rect 36866 49312 36948 49326
rect 37156 49312 37238 49326
rect 38114 49312 38196 49326
rect 38404 49312 38486 49326
rect 39362 49312 39444 49326
rect 39652 49312 39734 49326
rect 40610 49312 40692 49326
rect 40900 49312 40982 49326
rect 41858 49312 41940 49326
rect 42148 49312 42230 49326
rect 43106 49312 43188 49326
rect 43396 49312 43478 49326
rect 44354 49312 44436 49326
rect 44644 49312 44726 49326
rect 45602 49312 45684 49326
rect 45892 49312 45974 49326
rect 46850 49312 46932 49326
rect 47140 49312 47222 49326
rect 48098 49312 48180 49326
rect 48388 49312 48470 49326
rect 49346 49312 49428 49326
rect 49636 49312 49718 49326
rect 50594 49312 50676 49326
rect 50884 49312 50966 49326
rect 51842 49312 51924 49326
rect 52132 49312 52214 49326
rect 53090 49312 53172 49326
rect 53380 49312 53462 49326
rect 54338 49312 54420 49326
rect 54628 49312 54710 49326
rect 55586 49312 55668 49326
rect 55876 49312 55958 49326
rect 56834 49312 56916 49326
rect 57124 49312 57206 49326
rect 58082 49312 58164 49326
rect 58372 49312 58454 49326
rect 16418 49264 16864 49278
rect 17014 49264 17154 49278
rect 17304 49264 18112 49278
rect 18262 49264 18402 49278
rect 18552 49264 19360 49278
rect 19510 49264 19650 49278
rect 19800 49264 20608 49278
rect 20758 49264 20898 49278
rect 21048 49264 21856 49278
rect 22006 49264 22146 49278
rect 22296 49264 23104 49278
rect 23254 49264 23394 49278
rect 23544 49264 24352 49278
rect 24502 49264 24642 49278
rect 24792 49264 25600 49278
rect 25750 49264 25890 49278
rect 26040 49264 26848 49278
rect 26998 49264 27138 49278
rect 27288 49264 28096 49278
rect 28246 49264 28386 49278
rect 28536 49264 29344 49278
rect 29494 49264 29634 49278
rect 29784 49264 30592 49278
rect 30742 49264 30882 49278
rect 31032 49264 31840 49278
rect 31990 49264 32130 49278
rect 32280 49264 33088 49278
rect 33238 49264 33378 49278
rect 33528 49264 34336 49278
rect 34486 49264 34626 49278
rect 34776 49264 35584 49278
rect 35734 49264 35874 49278
rect 36024 49264 36832 49278
rect 36982 49264 37122 49278
rect 37272 49264 38080 49278
rect 38230 49264 38370 49278
rect 38520 49264 39328 49278
rect 39478 49264 39618 49278
rect 39768 49264 40576 49278
rect 40726 49264 40866 49278
rect 41016 49264 41824 49278
rect 41974 49264 42114 49278
rect 42264 49264 43072 49278
rect 43222 49264 43362 49278
rect 43512 49264 44320 49278
rect 44470 49264 44610 49278
rect 44760 49264 45568 49278
rect 45718 49264 45858 49278
rect 46008 49264 46816 49278
rect 46966 49264 47106 49278
rect 47256 49264 48064 49278
rect 48214 49264 48354 49278
rect 48504 49264 49312 49278
rect 49462 49264 49602 49278
rect 49752 49264 50560 49278
rect 50710 49264 50850 49278
rect 51000 49264 51808 49278
rect 51958 49264 52098 49278
rect 52248 49264 53056 49278
rect 53206 49264 53346 49278
rect 53496 49264 54304 49278
rect 54454 49264 54594 49278
rect 54744 49264 55552 49278
rect 55702 49264 55842 49278
rect 55992 49264 56800 49278
rect 56950 49264 57090 49278
rect 57240 49264 58048 49278
rect 58198 49264 58338 49278
rect 58488 49264 58934 49278
rect 16418 49216 58934 49264
rect 16418 49202 16864 49216
rect 17014 49202 17154 49216
rect 17304 49202 18112 49216
rect 18262 49202 18402 49216
rect 18552 49202 19360 49216
rect 19510 49202 19650 49216
rect 19800 49202 20608 49216
rect 20758 49202 20898 49216
rect 21048 49202 21856 49216
rect 22006 49202 22146 49216
rect 22296 49202 23104 49216
rect 23254 49202 23394 49216
rect 23544 49202 24352 49216
rect 24502 49202 24642 49216
rect 24792 49202 25600 49216
rect 25750 49202 25890 49216
rect 26040 49202 26848 49216
rect 26998 49202 27138 49216
rect 27288 49202 28096 49216
rect 28246 49202 28386 49216
rect 28536 49202 29344 49216
rect 29494 49202 29634 49216
rect 29784 49202 30592 49216
rect 30742 49202 30882 49216
rect 31032 49202 31840 49216
rect 31990 49202 32130 49216
rect 32280 49202 33088 49216
rect 33238 49202 33378 49216
rect 33528 49202 34336 49216
rect 34486 49202 34626 49216
rect 34776 49202 35584 49216
rect 35734 49202 35874 49216
rect 36024 49202 36832 49216
rect 36982 49202 37122 49216
rect 37272 49202 38080 49216
rect 38230 49202 38370 49216
rect 38520 49202 39328 49216
rect 39478 49202 39618 49216
rect 39768 49202 40576 49216
rect 40726 49202 40866 49216
rect 41016 49202 41824 49216
rect 41974 49202 42114 49216
rect 42264 49202 43072 49216
rect 43222 49202 43362 49216
rect 43512 49202 44320 49216
rect 44470 49202 44610 49216
rect 44760 49202 45568 49216
rect 45718 49202 45858 49216
rect 46008 49202 46816 49216
rect 46966 49202 47106 49216
rect 47256 49202 48064 49216
rect 48214 49202 48354 49216
rect 48504 49202 49312 49216
rect 49462 49202 49602 49216
rect 49752 49202 50560 49216
rect 50710 49202 50850 49216
rect 51000 49202 51808 49216
rect 51958 49202 52098 49216
rect 52248 49202 53056 49216
rect 53206 49202 53346 49216
rect 53496 49202 54304 49216
rect 54454 49202 54594 49216
rect 54744 49202 55552 49216
rect 55702 49202 55842 49216
rect 55992 49202 56800 49216
rect 56950 49202 57090 49216
rect 57240 49202 58048 49216
rect 58198 49202 58338 49216
rect 58488 49202 58934 49216
rect 16898 49154 16980 49168
rect 17188 49154 17270 49168
rect 18146 49154 18228 49168
rect 18436 49154 18518 49168
rect 19394 49154 19476 49168
rect 19684 49154 19766 49168
rect 20642 49154 20724 49168
rect 20932 49154 21014 49168
rect 21890 49154 21972 49168
rect 22180 49154 22262 49168
rect 23138 49154 23220 49168
rect 23428 49154 23510 49168
rect 24386 49154 24468 49168
rect 24676 49154 24758 49168
rect 25634 49154 25716 49168
rect 25924 49154 26006 49168
rect 26882 49154 26964 49168
rect 27172 49154 27254 49168
rect 28130 49154 28212 49168
rect 28420 49154 28502 49168
rect 29378 49154 29460 49168
rect 29668 49154 29750 49168
rect 30626 49154 30708 49168
rect 30916 49154 30998 49168
rect 31874 49154 31956 49168
rect 32164 49154 32246 49168
rect 33122 49154 33204 49168
rect 33412 49154 33494 49168
rect 34370 49154 34452 49168
rect 34660 49154 34742 49168
rect 35618 49154 35700 49168
rect 35908 49154 35990 49168
rect 36866 49154 36948 49168
rect 37156 49154 37238 49168
rect 38114 49154 38196 49168
rect 38404 49154 38486 49168
rect 39362 49154 39444 49168
rect 39652 49154 39734 49168
rect 40610 49154 40692 49168
rect 40900 49154 40982 49168
rect 41858 49154 41940 49168
rect 42148 49154 42230 49168
rect 43106 49154 43188 49168
rect 43396 49154 43478 49168
rect 44354 49154 44436 49168
rect 44644 49154 44726 49168
rect 45602 49154 45684 49168
rect 45892 49154 45974 49168
rect 46850 49154 46932 49168
rect 47140 49154 47222 49168
rect 48098 49154 48180 49168
rect 48388 49154 48470 49168
rect 49346 49154 49428 49168
rect 49636 49154 49718 49168
rect 50594 49154 50676 49168
rect 50884 49154 50966 49168
rect 51842 49154 51924 49168
rect 52132 49154 52214 49168
rect 53090 49154 53172 49168
rect 53380 49154 53462 49168
rect 54338 49154 54420 49168
rect 54628 49154 54710 49168
rect 55586 49154 55668 49168
rect 55876 49154 55958 49168
rect 56834 49154 56916 49168
rect 57124 49154 57206 49168
rect 58082 49154 58164 49168
rect 58372 49154 58454 49168
rect 16418 49106 58934 49154
rect 16418 48948 58934 49058
rect 16418 48852 58934 48900
rect 16898 48838 16980 48852
rect 17188 48838 17270 48852
rect 18146 48838 18228 48852
rect 18436 48838 18518 48852
rect 19394 48838 19476 48852
rect 19684 48838 19766 48852
rect 20642 48838 20724 48852
rect 20932 48838 21014 48852
rect 21890 48838 21972 48852
rect 22180 48838 22262 48852
rect 23138 48838 23220 48852
rect 23428 48838 23510 48852
rect 24386 48838 24468 48852
rect 24676 48838 24758 48852
rect 25634 48838 25716 48852
rect 25924 48838 26006 48852
rect 26882 48838 26964 48852
rect 27172 48838 27254 48852
rect 28130 48838 28212 48852
rect 28420 48838 28502 48852
rect 29378 48838 29460 48852
rect 29668 48838 29750 48852
rect 30626 48838 30708 48852
rect 30916 48838 30998 48852
rect 31874 48838 31956 48852
rect 32164 48838 32246 48852
rect 33122 48838 33204 48852
rect 33412 48838 33494 48852
rect 34370 48838 34452 48852
rect 34660 48838 34742 48852
rect 35618 48838 35700 48852
rect 35908 48838 35990 48852
rect 36866 48838 36948 48852
rect 37156 48838 37238 48852
rect 38114 48838 38196 48852
rect 38404 48838 38486 48852
rect 39362 48838 39444 48852
rect 39652 48838 39734 48852
rect 40610 48838 40692 48852
rect 40900 48838 40982 48852
rect 41858 48838 41940 48852
rect 42148 48838 42230 48852
rect 43106 48838 43188 48852
rect 43396 48838 43478 48852
rect 44354 48838 44436 48852
rect 44644 48838 44726 48852
rect 45602 48838 45684 48852
rect 45892 48838 45974 48852
rect 46850 48838 46932 48852
rect 47140 48838 47222 48852
rect 48098 48838 48180 48852
rect 48388 48838 48470 48852
rect 49346 48838 49428 48852
rect 49636 48838 49718 48852
rect 50594 48838 50676 48852
rect 50884 48838 50966 48852
rect 51842 48838 51924 48852
rect 52132 48838 52214 48852
rect 53090 48838 53172 48852
rect 53380 48838 53462 48852
rect 54338 48838 54420 48852
rect 54628 48838 54710 48852
rect 55586 48838 55668 48852
rect 55876 48838 55958 48852
rect 56834 48838 56916 48852
rect 57124 48838 57206 48852
rect 58082 48838 58164 48852
rect 58372 48838 58454 48852
rect 16418 48790 16864 48804
rect 17014 48790 17154 48804
rect 17304 48790 18112 48804
rect 18262 48790 18402 48804
rect 18552 48790 19360 48804
rect 19510 48790 19650 48804
rect 19800 48790 20608 48804
rect 20758 48790 20898 48804
rect 21048 48790 21856 48804
rect 22006 48790 22146 48804
rect 22296 48790 23104 48804
rect 23254 48790 23394 48804
rect 23544 48790 24352 48804
rect 24502 48790 24642 48804
rect 24792 48790 25600 48804
rect 25750 48790 25890 48804
rect 26040 48790 26848 48804
rect 26998 48790 27138 48804
rect 27288 48790 28096 48804
rect 28246 48790 28386 48804
rect 28536 48790 29344 48804
rect 29494 48790 29634 48804
rect 29784 48790 30592 48804
rect 30742 48790 30882 48804
rect 31032 48790 31840 48804
rect 31990 48790 32130 48804
rect 32280 48790 33088 48804
rect 33238 48790 33378 48804
rect 33528 48790 34336 48804
rect 34486 48790 34626 48804
rect 34776 48790 35584 48804
rect 35734 48790 35874 48804
rect 36024 48790 36832 48804
rect 36982 48790 37122 48804
rect 37272 48790 38080 48804
rect 38230 48790 38370 48804
rect 38520 48790 39328 48804
rect 39478 48790 39618 48804
rect 39768 48790 40576 48804
rect 40726 48790 40866 48804
rect 41016 48790 41824 48804
rect 41974 48790 42114 48804
rect 42264 48790 43072 48804
rect 43222 48790 43362 48804
rect 43512 48790 44320 48804
rect 44470 48790 44610 48804
rect 44760 48790 45568 48804
rect 45718 48790 45858 48804
rect 46008 48790 46816 48804
rect 46966 48790 47106 48804
rect 47256 48790 48064 48804
rect 48214 48790 48354 48804
rect 48504 48790 49312 48804
rect 49462 48790 49602 48804
rect 49752 48790 50560 48804
rect 50710 48790 50850 48804
rect 51000 48790 51808 48804
rect 51958 48790 52098 48804
rect 52248 48790 53056 48804
rect 53206 48790 53346 48804
rect 53496 48790 54304 48804
rect 54454 48790 54594 48804
rect 54744 48790 55552 48804
rect 55702 48790 55842 48804
rect 55992 48790 56800 48804
rect 56950 48790 57090 48804
rect 57240 48790 58048 48804
rect 58198 48790 58338 48804
rect 58488 48790 58934 48804
rect 16418 48742 58934 48790
rect 16418 48728 16864 48742
rect 17014 48728 17154 48742
rect 17304 48728 18112 48742
rect 18262 48728 18402 48742
rect 18552 48728 19360 48742
rect 19510 48728 19650 48742
rect 19800 48728 20608 48742
rect 20758 48728 20898 48742
rect 21048 48728 21856 48742
rect 22006 48728 22146 48742
rect 22296 48728 23104 48742
rect 23254 48728 23394 48742
rect 23544 48728 24352 48742
rect 24502 48728 24642 48742
rect 24792 48728 25600 48742
rect 25750 48728 25890 48742
rect 26040 48728 26848 48742
rect 26998 48728 27138 48742
rect 27288 48728 28096 48742
rect 28246 48728 28386 48742
rect 28536 48728 29344 48742
rect 29494 48728 29634 48742
rect 29784 48728 30592 48742
rect 30742 48728 30882 48742
rect 31032 48728 31840 48742
rect 31990 48728 32130 48742
rect 32280 48728 33088 48742
rect 33238 48728 33378 48742
rect 33528 48728 34336 48742
rect 34486 48728 34626 48742
rect 34776 48728 35584 48742
rect 35734 48728 35874 48742
rect 36024 48728 36832 48742
rect 36982 48728 37122 48742
rect 37272 48728 38080 48742
rect 38230 48728 38370 48742
rect 38520 48728 39328 48742
rect 39478 48728 39618 48742
rect 39768 48728 40576 48742
rect 40726 48728 40866 48742
rect 41016 48728 41824 48742
rect 41974 48728 42114 48742
rect 42264 48728 43072 48742
rect 43222 48728 43362 48742
rect 43512 48728 44320 48742
rect 44470 48728 44610 48742
rect 44760 48728 45568 48742
rect 45718 48728 45858 48742
rect 46008 48728 46816 48742
rect 46966 48728 47106 48742
rect 47256 48728 48064 48742
rect 48214 48728 48354 48742
rect 48504 48728 49312 48742
rect 49462 48728 49602 48742
rect 49752 48728 50560 48742
rect 50710 48728 50850 48742
rect 51000 48728 51808 48742
rect 51958 48728 52098 48742
rect 52248 48728 53056 48742
rect 53206 48728 53346 48742
rect 53496 48728 54304 48742
rect 54454 48728 54594 48742
rect 54744 48728 55552 48742
rect 55702 48728 55842 48742
rect 55992 48728 56800 48742
rect 56950 48728 57090 48742
rect 57240 48728 58048 48742
rect 58198 48728 58338 48742
rect 58488 48728 58934 48742
rect 16898 48680 16980 48694
rect 17188 48680 17270 48694
rect 18146 48680 18228 48694
rect 18436 48680 18518 48694
rect 19394 48680 19476 48694
rect 19684 48680 19766 48694
rect 20642 48680 20724 48694
rect 20932 48680 21014 48694
rect 21890 48680 21972 48694
rect 22180 48680 22262 48694
rect 23138 48680 23220 48694
rect 23428 48680 23510 48694
rect 24386 48680 24468 48694
rect 24676 48680 24758 48694
rect 25634 48680 25716 48694
rect 25924 48680 26006 48694
rect 26882 48680 26964 48694
rect 27172 48680 27254 48694
rect 28130 48680 28212 48694
rect 28420 48680 28502 48694
rect 29378 48680 29460 48694
rect 29668 48680 29750 48694
rect 30626 48680 30708 48694
rect 30916 48680 30998 48694
rect 31874 48680 31956 48694
rect 32164 48680 32246 48694
rect 33122 48680 33204 48694
rect 33412 48680 33494 48694
rect 34370 48680 34452 48694
rect 34660 48680 34742 48694
rect 35618 48680 35700 48694
rect 35908 48680 35990 48694
rect 36866 48680 36948 48694
rect 37156 48680 37238 48694
rect 38114 48680 38196 48694
rect 38404 48680 38486 48694
rect 39362 48680 39444 48694
rect 39652 48680 39734 48694
rect 40610 48680 40692 48694
rect 40900 48680 40982 48694
rect 41858 48680 41940 48694
rect 42148 48680 42230 48694
rect 43106 48680 43188 48694
rect 43396 48680 43478 48694
rect 44354 48680 44436 48694
rect 44644 48680 44726 48694
rect 45602 48680 45684 48694
rect 45892 48680 45974 48694
rect 46850 48680 46932 48694
rect 47140 48680 47222 48694
rect 48098 48680 48180 48694
rect 48388 48680 48470 48694
rect 49346 48680 49428 48694
rect 49636 48680 49718 48694
rect 50594 48680 50676 48694
rect 50884 48680 50966 48694
rect 51842 48680 51924 48694
rect 52132 48680 52214 48694
rect 53090 48680 53172 48694
rect 53380 48680 53462 48694
rect 54338 48680 54420 48694
rect 54628 48680 54710 48694
rect 55586 48680 55668 48694
rect 55876 48680 55958 48694
rect 56834 48680 56916 48694
rect 57124 48680 57206 48694
rect 58082 48680 58164 48694
rect 58372 48680 58454 48694
rect 16418 48632 58934 48680
rect 16418 48536 58934 48584
rect 16898 48522 16980 48536
rect 17188 48522 17270 48536
rect 18146 48522 18228 48536
rect 18436 48522 18518 48536
rect 19394 48522 19476 48536
rect 19684 48522 19766 48536
rect 20642 48522 20724 48536
rect 20932 48522 21014 48536
rect 21890 48522 21972 48536
rect 22180 48522 22262 48536
rect 23138 48522 23220 48536
rect 23428 48522 23510 48536
rect 24386 48522 24468 48536
rect 24676 48522 24758 48536
rect 25634 48522 25716 48536
rect 25924 48522 26006 48536
rect 26882 48522 26964 48536
rect 27172 48522 27254 48536
rect 28130 48522 28212 48536
rect 28420 48522 28502 48536
rect 29378 48522 29460 48536
rect 29668 48522 29750 48536
rect 30626 48522 30708 48536
rect 30916 48522 30998 48536
rect 31874 48522 31956 48536
rect 32164 48522 32246 48536
rect 33122 48522 33204 48536
rect 33412 48522 33494 48536
rect 34370 48522 34452 48536
rect 34660 48522 34742 48536
rect 35618 48522 35700 48536
rect 35908 48522 35990 48536
rect 36866 48522 36948 48536
rect 37156 48522 37238 48536
rect 38114 48522 38196 48536
rect 38404 48522 38486 48536
rect 39362 48522 39444 48536
rect 39652 48522 39734 48536
rect 40610 48522 40692 48536
rect 40900 48522 40982 48536
rect 41858 48522 41940 48536
rect 42148 48522 42230 48536
rect 43106 48522 43188 48536
rect 43396 48522 43478 48536
rect 44354 48522 44436 48536
rect 44644 48522 44726 48536
rect 45602 48522 45684 48536
rect 45892 48522 45974 48536
rect 46850 48522 46932 48536
rect 47140 48522 47222 48536
rect 48098 48522 48180 48536
rect 48388 48522 48470 48536
rect 49346 48522 49428 48536
rect 49636 48522 49718 48536
rect 50594 48522 50676 48536
rect 50884 48522 50966 48536
rect 51842 48522 51924 48536
rect 52132 48522 52214 48536
rect 53090 48522 53172 48536
rect 53380 48522 53462 48536
rect 54338 48522 54420 48536
rect 54628 48522 54710 48536
rect 55586 48522 55668 48536
rect 55876 48522 55958 48536
rect 56834 48522 56916 48536
rect 57124 48522 57206 48536
rect 58082 48522 58164 48536
rect 58372 48522 58454 48536
rect 16418 48474 16864 48488
rect 17014 48474 17154 48488
rect 17304 48474 18112 48488
rect 18262 48474 18402 48488
rect 18552 48474 19360 48488
rect 19510 48474 19650 48488
rect 19800 48474 20608 48488
rect 20758 48474 20898 48488
rect 21048 48474 21856 48488
rect 22006 48474 22146 48488
rect 22296 48474 23104 48488
rect 23254 48474 23394 48488
rect 23544 48474 24352 48488
rect 24502 48474 24642 48488
rect 24792 48474 25600 48488
rect 25750 48474 25890 48488
rect 26040 48474 26848 48488
rect 26998 48474 27138 48488
rect 27288 48474 28096 48488
rect 28246 48474 28386 48488
rect 28536 48474 29344 48488
rect 29494 48474 29634 48488
rect 29784 48474 30592 48488
rect 30742 48474 30882 48488
rect 31032 48474 31840 48488
rect 31990 48474 32130 48488
rect 32280 48474 33088 48488
rect 33238 48474 33378 48488
rect 33528 48474 34336 48488
rect 34486 48474 34626 48488
rect 34776 48474 35584 48488
rect 35734 48474 35874 48488
rect 36024 48474 36832 48488
rect 36982 48474 37122 48488
rect 37272 48474 38080 48488
rect 38230 48474 38370 48488
rect 38520 48474 39328 48488
rect 39478 48474 39618 48488
rect 39768 48474 40576 48488
rect 40726 48474 40866 48488
rect 41016 48474 41824 48488
rect 41974 48474 42114 48488
rect 42264 48474 43072 48488
rect 43222 48474 43362 48488
rect 43512 48474 44320 48488
rect 44470 48474 44610 48488
rect 44760 48474 45568 48488
rect 45718 48474 45858 48488
rect 46008 48474 46816 48488
rect 46966 48474 47106 48488
rect 47256 48474 48064 48488
rect 48214 48474 48354 48488
rect 48504 48474 49312 48488
rect 49462 48474 49602 48488
rect 49752 48474 50560 48488
rect 50710 48474 50850 48488
rect 51000 48474 51808 48488
rect 51958 48474 52098 48488
rect 52248 48474 53056 48488
rect 53206 48474 53346 48488
rect 53496 48474 54304 48488
rect 54454 48474 54594 48488
rect 54744 48474 55552 48488
rect 55702 48474 55842 48488
rect 55992 48474 56800 48488
rect 56950 48474 57090 48488
rect 57240 48474 58048 48488
rect 58198 48474 58338 48488
rect 58488 48474 58934 48488
rect 16418 48426 58934 48474
rect 16418 48412 16864 48426
rect 17014 48412 17154 48426
rect 17304 48412 18112 48426
rect 18262 48412 18402 48426
rect 18552 48412 19360 48426
rect 19510 48412 19650 48426
rect 19800 48412 20608 48426
rect 20758 48412 20898 48426
rect 21048 48412 21856 48426
rect 22006 48412 22146 48426
rect 22296 48412 23104 48426
rect 23254 48412 23394 48426
rect 23544 48412 24352 48426
rect 24502 48412 24642 48426
rect 24792 48412 25600 48426
rect 25750 48412 25890 48426
rect 26040 48412 26848 48426
rect 26998 48412 27138 48426
rect 27288 48412 28096 48426
rect 28246 48412 28386 48426
rect 28536 48412 29344 48426
rect 29494 48412 29634 48426
rect 29784 48412 30592 48426
rect 30742 48412 30882 48426
rect 31032 48412 31840 48426
rect 31990 48412 32130 48426
rect 32280 48412 33088 48426
rect 33238 48412 33378 48426
rect 33528 48412 34336 48426
rect 34486 48412 34626 48426
rect 34776 48412 35584 48426
rect 35734 48412 35874 48426
rect 36024 48412 36832 48426
rect 36982 48412 37122 48426
rect 37272 48412 38080 48426
rect 38230 48412 38370 48426
rect 38520 48412 39328 48426
rect 39478 48412 39618 48426
rect 39768 48412 40576 48426
rect 40726 48412 40866 48426
rect 41016 48412 41824 48426
rect 41974 48412 42114 48426
rect 42264 48412 43072 48426
rect 43222 48412 43362 48426
rect 43512 48412 44320 48426
rect 44470 48412 44610 48426
rect 44760 48412 45568 48426
rect 45718 48412 45858 48426
rect 46008 48412 46816 48426
rect 46966 48412 47106 48426
rect 47256 48412 48064 48426
rect 48214 48412 48354 48426
rect 48504 48412 49312 48426
rect 49462 48412 49602 48426
rect 49752 48412 50560 48426
rect 50710 48412 50850 48426
rect 51000 48412 51808 48426
rect 51958 48412 52098 48426
rect 52248 48412 53056 48426
rect 53206 48412 53346 48426
rect 53496 48412 54304 48426
rect 54454 48412 54594 48426
rect 54744 48412 55552 48426
rect 55702 48412 55842 48426
rect 55992 48412 56800 48426
rect 56950 48412 57090 48426
rect 57240 48412 58048 48426
rect 58198 48412 58338 48426
rect 58488 48412 58934 48426
rect 16898 48364 16980 48378
rect 17188 48364 17270 48378
rect 18146 48364 18228 48378
rect 18436 48364 18518 48378
rect 19394 48364 19476 48378
rect 19684 48364 19766 48378
rect 20642 48364 20724 48378
rect 20932 48364 21014 48378
rect 21890 48364 21972 48378
rect 22180 48364 22262 48378
rect 23138 48364 23220 48378
rect 23428 48364 23510 48378
rect 24386 48364 24468 48378
rect 24676 48364 24758 48378
rect 25634 48364 25716 48378
rect 25924 48364 26006 48378
rect 26882 48364 26964 48378
rect 27172 48364 27254 48378
rect 28130 48364 28212 48378
rect 28420 48364 28502 48378
rect 29378 48364 29460 48378
rect 29668 48364 29750 48378
rect 30626 48364 30708 48378
rect 30916 48364 30998 48378
rect 31874 48364 31956 48378
rect 32164 48364 32246 48378
rect 33122 48364 33204 48378
rect 33412 48364 33494 48378
rect 34370 48364 34452 48378
rect 34660 48364 34742 48378
rect 35618 48364 35700 48378
rect 35908 48364 35990 48378
rect 36866 48364 36948 48378
rect 37156 48364 37238 48378
rect 38114 48364 38196 48378
rect 38404 48364 38486 48378
rect 39362 48364 39444 48378
rect 39652 48364 39734 48378
rect 40610 48364 40692 48378
rect 40900 48364 40982 48378
rect 41858 48364 41940 48378
rect 42148 48364 42230 48378
rect 43106 48364 43188 48378
rect 43396 48364 43478 48378
rect 44354 48364 44436 48378
rect 44644 48364 44726 48378
rect 45602 48364 45684 48378
rect 45892 48364 45974 48378
rect 46850 48364 46932 48378
rect 47140 48364 47222 48378
rect 48098 48364 48180 48378
rect 48388 48364 48470 48378
rect 49346 48364 49428 48378
rect 49636 48364 49718 48378
rect 50594 48364 50676 48378
rect 50884 48364 50966 48378
rect 51842 48364 51924 48378
rect 52132 48364 52214 48378
rect 53090 48364 53172 48378
rect 53380 48364 53462 48378
rect 54338 48364 54420 48378
rect 54628 48364 54710 48378
rect 55586 48364 55668 48378
rect 55876 48364 55958 48378
rect 56834 48364 56916 48378
rect 57124 48364 57206 48378
rect 58082 48364 58164 48378
rect 58372 48364 58454 48378
rect 16418 48316 58934 48364
rect 16418 48158 58934 48268
rect 16418 48062 58934 48110
rect 16898 48048 16980 48062
rect 17188 48048 17270 48062
rect 18146 48048 18228 48062
rect 18436 48048 18518 48062
rect 19394 48048 19476 48062
rect 19684 48048 19766 48062
rect 20642 48048 20724 48062
rect 20932 48048 21014 48062
rect 21890 48048 21972 48062
rect 22180 48048 22262 48062
rect 23138 48048 23220 48062
rect 23428 48048 23510 48062
rect 24386 48048 24468 48062
rect 24676 48048 24758 48062
rect 25634 48048 25716 48062
rect 25924 48048 26006 48062
rect 26882 48048 26964 48062
rect 27172 48048 27254 48062
rect 28130 48048 28212 48062
rect 28420 48048 28502 48062
rect 29378 48048 29460 48062
rect 29668 48048 29750 48062
rect 30626 48048 30708 48062
rect 30916 48048 30998 48062
rect 31874 48048 31956 48062
rect 32164 48048 32246 48062
rect 33122 48048 33204 48062
rect 33412 48048 33494 48062
rect 34370 48048 34452 48062
rect 34660 48048 34742 48062
rect 35618 48048 35700 48062
rect 35908 48048 35990 48062
rect 36866 48048 36948 48062
rect 37156 48048 37238 48062
rect 38114 48048 38196 48062
rect 38404 48048 38486 48062
rect 39362 48048 39444 48062
rect 39652 48048 39734 48062
rect 40610 48048 40692 48062
rect 40900 48048 40982 48062
rect 41858 48048 41940 48062
rect 42148 48048 42230 48062
rect 43106 48048 43188 48062
rect 43396 48048 43478 48062
rect 44354 48048 44436 48062
rect 44644 48048 44726 48062
rect 45602 48048 45684 48062
rect 45892 48048 45974 48062
rect 46850 48048 46932 48062
rect 47140 48048 47222 48062
rect 48098 48048 48180 48062
rect 48388 48048 48470 48062
rect 49346 48048 49428 48062
rect 49636 48048 49718 48062
rect 50594 48048 50676 48062
rect 50884 48048 50966 48062
rect 51842 48048 51924 48062
rect 52132 48048 52214 48062
rect 53090 48048 53172 48062
rect 53380 48048 53462 48062
rect 54338 48048 54420 48062
rect 54628 48048 54710 48062
rect 55586 48048 55668 48062
rect 55876 48048 55958 48062
rect 56834 48048 56916 48062
rect 57124 48048 57206 48062
rect 58082 48048 58164 48062
rect 58372 48048 58454 48062
rect 16418 48000 16864 48014
rect 17014 48000 17154 48014
rect 17304 48000 18112 48014
rect 18262 48000 18402 48014
rect 18552 48000 19360 48014
rect 19510 48000 19650 48014
rect 19800 48000 20608 48014
rect 20758 48000 20898 48014
rect 21048 48000 21856 48014
rect 22006 48000 22146 48014
rect 22296 48000 23104 48014
rect 23254 48000 23394 48014
rect 23544 48000 24352 48014
rect 24502 48000 24642 48014
rect 24792 48000 25600 48014
rect 25750 48000 25890 48014
rect 26040 48000 26848 48014
rect 26998 48000 27138 48014
rect 27288 48000 28096 48014
rect 28246 48000 28386 48014
rect 28536 48000 29344 48014
rect 29494 48000 29634 48014
rect 29784 48000 30592 48014
rect 30742 48000 30882 48014
rect 31032 48000 31840 48014
rect 31990 48000 32130 48014
rect 32280 48000 33088 48014
rect 33238 48000 33378 48014
rect 33528 48000 34336 48014
rect 34486 48000 34626 48014
rect 34776 48000 35584 48014
rect 35734 48000 35874 48014
rect 36024 48000 36832 48014
rect 36982 48000 37122 48014
rect 37272 48000 38080 48014
rect 38230 48000 38370 48014
rect 38520 48000 39328 48014
rect 39478 48000 39618 48014
rect 39768 48000 40576 48014
rect 40726 48000 40866 48014
rect 41016 48000 41824 48014
rect 41974 48000 42114 48014
rect 42264 48000 43072 48014
rect 43222 48000 43362 48014
rect 43512 48000 44320 48014
rect 44470 48000 44610 48014
rect 44760 48000 45568 48014
rect 45718 48000 45858 48014
rect 46008 48000 46816 48014
rect 46966 48000 47106 48014
rect 47256 48000 48064 48014
rect 48214 48000 48354 48014
rect 48504 48000 49312 48014
rect 49462 48000 49602 48014
rect 49752 48000 50560 48014
rect 50710 48000 50850 48014
rect 51000 48000 51808 48014
rect 51958 48000 52098 48014
rect 52248 48000 53056 48014
rect 53206 48000 53346 48014
rect 53496 48000 54304 48014
rect 54454 48000 54594 48014
rect 54744 48000 55552 48014
rect 55702 48000 55842 48014
rect 55992 48000 56800 48014
rect 56950 48000 57090 48014
rect 57240 48000 58048 48014
rect 58198 48000 58338 48014
rect 58488 48000 58934 48014
rect 16418 47952 58934 48000
rect 16418 47938 16864 47952
rect 17014 47938 17154 47952
rect 17304 47938 18112 47952
rect 18262 47938 18402 47952
rect 18552 47938 19360 47952
rect 19510 47938 19650 47952
rect 19800 47938 20608 47952
rect 20758 47938 20898 47952
rect 21048 47938 21856 47952
rect 22006 47938 22146 47952
rect 22296 47938 23104 47952
rect 23254 47938 23394 47952
rect 23544 47938 24352 47952
rect 24502 47938 24642 47952
rect 24792 47938 25600 47952
rect 25750 47938 25890 47952
rect 26040 47938 26848 47952
rect 26998 47938 27138 47952
rect 27288 47938 28096 47952
rect 28246 47938 28386 47952
rect 28536 47938 29344 47952
rect 29494 47938 29634 47952
rect 29784 47938 30592 47952
rect 30742 47938 30882 47952
rect 31032 47938 31840 47952
rect 31990 47938 32130 47952
rect 32280 47938 33088 47952
rect 33238 47938 33378 47952
rect 33528 47938 34336 47952
rect 34486 47938 34626 47952
rect 34776 47938 35584 47952
rect 35734 47938 35874 47952
rect 36024 47938 36832 47952
rect 36982 47938 37122 47952
rect 37272 47938 38080 47952
rect 38230 47938 38370 47952
rect 38520 47938 39328 47952
rect 39478 47938 39618 47952
rect 39768 47938 40576 47952
rect 40726 47938 40866 47952
rect 41016 47938 41824 47952
rect 41974 47938 42114 47952
rect 42264 47938 43072 47952
rect 43222 47938 43362 47952
rect 43512 47938 44320 47952
rect 44470 47938 44610 47952
rect 44760 47938 45568 47952
rect 45718 47938 45858 47952
rect 46008 47938 46816 47952
rect 46966 47938 47106 47952
rect 47256 47938 48064 47952
rect 48214 47938 48354 47952
rect 48504 47938 49312 47952
rect 49462 47938 49602 47952
rect 49752 47938 50560 47952
rect 50710 47938 50850 47952
rect 51000 47938 51808 47952
rect 51958 47938 52098 47952
rect 52248 47938 53056 47952
rect 53206 47938 53346 47952
rect 53496 47938 54304 47952
rect 54454 47938 54594 47952
rect 54744 47938 55552 47952
rect 55702 47938 55842 47952
rect 55992 47938 56800 47952
rect 56950 47938 57090 47952
rect 57240 47938 58048 47952
rect 58198 47938 58338 47952
rect 58488 47938 58934 47952
rect 16898 47890 16980 47904
rect 17188 47890 17270 47904
rect 18146 47890 18228 47904
rect 18436 47890 18518 47904
rect 19394 47890 19476 47904
rect 19684 47890 19766 47904
rect 20642 47890 20724 47904
rect 20932 47890 21014 47904
rect 21890 47890 21972 47904
rect 22180 47890 22262 47904
rect 23138 47890 23220 47904
rect 23428 47890 23510 47904
rect 24386 47890 24468 47904
rect 24676 47890 24758 47904
rect 25634 47890 25716 47904
rect 25924 47890 26006 47904
rect 26882 47890 26964 47904
rect 27172 47890 27254 47904
rect 28130 47890 28212 47904
rect 28420 47890 28502 47904
rect 29378 47890 29460 47904
rect 29668 47890 29750 47904
rect 30626 47890 30708 47904
rect 30916 47890 30998 47904
rect 31874 47890 31956 47904
rect 32164 47890 32246 47904
rect 33122 47890 33204 47904
rect 33412 47890 33494 47904
rect 34370 47890 34452 47904
rect 34660 47890 34742 47904
rect 35618 47890 35700 47904
rect 35908 47890 35990 47904
rect 36866 47890 36948 47904
rect 37156 47890 37238 47904
rect 38114 47890 38196 47904
rect 38404 47890 38486 47904
rect 39362 47890 39444 47904
rect 39652 47890 39734 47904
rect 40610 47890 40692 47904
rect 40900 47890 40982 47904
rect 41858 47890 41940 47904
rect 42148 47890 42230 47904
rect 43106 47890 43188 47904
rect 43396 47890 43478 47904
rect 44354 47890 44436 47904
rect 44644 47890 44726 47904
rect 45602 47890 45684 47904
rect 45892 47890 45974 47904
rect 46850 47890 46932 47904
rect 47140 47890 47222 47904
rect 48098 47890 48180 47904
rect 48388 47890 48470 47904
rect 49346 47890 49428 47904
rect 49636 47890 49718 47904
rect 50594 47890 50676 47904
rect 50884 47890 50966 47904
rect 51842 47890 51924 47904
rect 52132 47890 52214 47904
rect 53090 47890 53172 47904
rect 53380 47890 53462 47904
rect 54338 47890 54420 47904
rect 54628 47890 54710 47904
rect 55586 47890 55668 47904
rect 55876 47890 55958 47904
rect 56834 47890 56916 47904
rect 57124 47890 57206 47904
rect 58082 47890 58164 47904
rect 58372 47890 58454 47904
rect 16418 47842 58934 47890
rect 16418 47746 58934 47794
rect 16898 47732 16980 47746
rect 17188 47732 17270 47746
rect 18146 47732 18228 47746
rect 18436 47732 18518 47746
rect 19394 47732 19476 47746
rect 19684 47732 19766 47746
rect 20642 47732 20724 47746
rect 20932 47732 21014 47746
rect 21890 47732 21972 47746
rect 22180 47732 22262 47746
rect 23138 47732 23220 47746
rect 23428 47732 23510 47746
rect 24386 47732 24468 47746
rect 24676 47732 24758 47746
rect 25634 47732 25716 47746
rect 25924 47732 26006 47746
rect 26882 47732 26964 47746
rect 27172 47732 27254 47746
rect 28130 47732 28212 47746
rect 28420 47732 28502 47746
rect 29378 47732 29460 47746
rect 29668 47732 29750 47746
rect 30626 47732 30708 47746
rect 30916 47732 30998 47746
rect 31874 47732 31956 47746
rect 32164 47732 32246 47746
rect 33122 47732 33204 47746
rect 33412 47732 33494 47746
rect 34370 47732 34452 47746
rect 34660 47732 34742 47746
rect 35618 47732 35700 47746
rect 35908 47732 35990 47746
rect 36866 47732 36948 47746
rect 37156 47732 37238 47746
rect 38114 47732 38196 47746
rect 38404 47732 38486 47746
rect 39362 47732 39444 47746
rect 39652 47732 39734 47746
rect 40610 47732 40692 47746
rect 40900 47732 40982 47746
rect 41858 47732 41940 47746
rect 42148 47732 42230 47746
rect 43106 47732 43188 47746
rect 43396 47732 43478 47746
rect 44354 47732 44436 47746
rect 44644 47732 44726 47746
rect 45602 47732 45684 47746
rect 45892 47732 45974 47746
rect 46850 47732 46932 47746
rect 47140 47732 47222 47746
rect 48098 47732 48180 47746
rect 48388 47732 48470 47746
rect 49346 47732 49428 47746
rect 49636 47732 49718 47746
rect 50594 47732 50676 47746
rect 50884 47732 50966 47746
rect 51842 47732 51924 47746
rect 52132 47732 52214 47746
rect 53090 47732 53172 47746
rect 53380 47732 53462 47746
rect 54338 47732 54420 47746
rect 54628 47732 54710 47746
rect 55586 47732 55668 47746
rect 55876 47732 55958 47746
rect 56834 47732 56916 47746
rect 57124 47732 57206 47746
rect 58082 47732 58164 47746
rect 58372 47732 58454 47746
rect 16418 47684 16864 47698
rect 17014 47684 17154 47698
rect 17304 47684 18112 47698
rect 18262 47684 18402 47698
rect 18552 47684 19360 47698
rect 19510 47684 19650 47698
rect 19800 47684 20608 47698
rect 20758 47684 20898 47698
rect 21048 47684 21856 47698
rect 22006 47684 22146 47698
rect 22296 47684 23104 47698
rect 23254 47684 23394 47698
rect 23544 47684 24352 47698
rect 24502 47684 24642 47698
rect 24792 47684 25600 47698
rect 25750 47684 25890 47698
rect 26040 47684 26848 47698
rect 26998 47684 27138 47698
rect 27288 47684 28096 47698
rect 28246 47684 28386 47698
rect 28536 47684 29344 47698
rect 29494 47684 29634 47698
rect 29784 47684 30592 47698
rect 30742 47684 30882 47698
rect 31032 47684 31840 47698
rect 31990 47684 32130 47698
rect 32280 47684 33088 47698
rect 33238 47684 33378 47698
rect 33528 47684 34336 47698
rect 34486 47684 34626 47698
rect 34776 47684 35584 47698
rect 35734 47684 35874 47698
rect 36024 47684 36832 47698
rect 36982 47684 37122 47698
rect 37272 47684 38080 47698
rect 38230 47684 38370 47698
rect 38520 47684 39328 47698
rect 39478 47684 39618 47698
rect 39768 47684 40576 47698
rect 40726 47684 40866 47698
rect 41016 47684 41824 47698
rect 41974 47684 42114 47698
rect 42264 47684 43072 47698
rect 43222 47684 43362 47698
rect 43512 47684 44320 47698
rect 44470 47684 44610 47698
rect 44760 47684 45568 47698
rect 45718 47684 45858 47698
rect 46008 47684 46816 47698
rect 46966 47684 47106 47698
rect 47256 47684 48064 47698
rect 48214 47684 48354 47698
rect 48504 47684 49312 47698
rect 49462 47684 49602 47698
rect 49752 47684 50560 47698
rect 50710 47684 50850 47698
rect 51000 47684 51808 47698
rect 51958 47684 52098 47698
rect 52248 47684 53056 47698
rect 53206 47684 53346 47698
rect 53496 47684 54304 47698
rect 54454 47684 54594 47698
rect 54744 47684 55552 47698
rect 55702 47684 55842 47698
rect 55992 47684 56800 47698
rect 56950 47684 57090 47698
rect 57240 47684 58048 47698
rect 58198 47684 58338 47698
rect 58488 47684 58934 47698
rect 16418 47636 58934 47684
rect 16418 47622 16864 47636
rect 17014 47622 17154 47636
rect 17304 47622 18112 47636
rect 18262 47622 18402 47636
rect 18552 47622 19360 47636
rect 19510 47622 19650 47636
rect 19800 47622 20608 47636
rect 20758 47622 20898 47636
rect 21048 47622 21856 47636
rect 22006 47622 22146 47636
rect 22296 47622 23104 47636
rect 23254 47622 23394 47636
rect 23544 47622 24352 47636
rect 24502 47622 24642 47636
rect 24792 47622 25600 47636
rect 25750 47622 25890 47636
rect 26040 47622 26848 47636
rect 26998 47622 27138 47636
rect 27288 47622 28096 47636
rect 28246 47622 28386 47636
rect 28536 47622 29344 47636
rect 29494 47622 29634 47636
rect 29784 47622 30592 47636
rect 30742 47622 30882 47636
rect 31032 47622 31840 47636
rect 31990 47622 32130 47636
rect 32280 47622 33088 47636
rect 33238 47622 33378 47636
rect 33528 47622 34336 47636
rect 34486 47622 34626 47636
rect 34776 47622 35584 47636
rect 35734 47622 35874 47636
rect 36024 47622 36832 47636
rect 36982 47622 37122 47636
rect 37272 47622 38080 47636
rect 38230 47622 38370 47636
rect 38520 47622 39328 47636
rect 39478 47622 39618 47636
rect 39768 47622 40576 47636
rect 40726 47622 40866 47636
rect 41016 47622 41824 47636
rect 41974 47622 42114 47636
rect 42264 47622 43072 47636
rect 43222 47622 43362 47636
rect 43512 47622 44320 47636
rect 44470 47622 44610 47636
rect 44760 47622 45568 47636
rect 45718 47622 45858 47636
rect 46008 47622 46816 47636
rect 46966 47622 47106 47636
rect 47256 47622 48064 47636
rect 48214 47622 48354 47636
rect 48504 47622 49312 47636
rect 49462 47622 49602 47636
rect 49752 47622 50560 47636
rect 50710 47622 50850 47636
rect 51000 47622 51808 47636
rect 51958 47622 52098 47636
rect 52248 47622 53056 47636
rect 53206 47622 53346 47636
rect 53496 47622 54304 47636
rect 54454 47622 54594 47636
rect 54744 47622 55552 47636
rect 55702 47622 55842 47636
rect 55992 47622 56800 47636
rect 56950 47622 57090 47636
rect 57240 47622 58048 47636
rect 58198 47622 58338 47636
rect 58488 47622 58934 47636
rect 16898 47574 16980 47588
rect 17188 47574 17270 47588
rect 18146 47574 18228 47588
rect 18436 47574 18518 47588
rect 19394 47574 19476 47588
rect 19684 47574 19766 47588
rect 20642 47574 20724 47588
rect 20932 47574 21014 47588
rect 21890 47574 21972 47588
rect 22180 47574 22262 47588
rect 23138 47574 23220 47588
rect 23428 47574 23510 47588
rect 24386 47574 24468 47588
rect 24676 47574 24758 47588
rect 25634 47574 25716 47588
rect 25924 47574 26006 47588
rect 26882 47574 26964 47588
rect 27172 47574 27254 47588
rect 28130 47574 28212 47588
rect 28420 47574 28502 47588
rect 29378 47574 29460 47588
rect 29668 47574 29750 47588
rect 30626 47574 30708 47588
rect 30916 47574 30998 47588
rect 31874 47574 31956 47588
rect 32164 47574 32246 47588
rect 33122 47574 33204 47588
rect 33412 47574 33494 47588
rect 34370 47574 34452 47588
rect 34660 47574 34742 47588
rect 35618 47574 35700 47588
rect 35908 47574 35990 47588
rect 36866 47574 36948 47588
rect 37156 47574 37238 47588
rect 38114 47574 38196 47588
rect 38404 47574 38486 47588
rect 39362 47574 39444 47588
rect 39652 47574 39734 47588
rect 40610 47574 40692 47588
rect 40900 47574 40982 47588
rect 41858 47574 41940 47588
rect 42148 47574 42230 47588
rect 43106 47574 43188 47588
rect 43396 47574 43478 47588
rect 44354 47574 44436 47588
rect 44644 47574 44726 47588
rect 45602 47574 45684 47588
rect 45892 47574 45974 47588
rect 46850 47574 46932 47588
rect 47140 47574 47222 47588
rect 48098 47574 48180 47588
rect 48388 47574 48470 47588
rect 49346 47574 49428 47588
rect 49636 47574 49718 47588
rect 50594 47574 50676 47588
rect 50884 47574 50966 47588
rect 51842 47574 51924 47588
rect 52132 47574 52214 47588
rect 53090 47574 53172 47588
rect 53380 47574 53462 47588
rect 54338 47574 54420 47588
rect 54628 47574 54710 47588
rect 55586 47574 55668 47588
rect 55876 47574 55958 47588
rect 56834 47574 56916 47588
rect 57124 47574 57206 47588
rect 58082 47574 58164 47588
rect 58372 47574 58454 47588
rect 16418 47526 58934 47574
rect 16418 47368 58934 47478
rect 16418 47272 58934 47320
rect 16898 47258 16980 47272
rect 17188 47258 17270 47272
rect 18146 47258 18228 47272
rect 18436 47258 18518 47272
rect 19394 47258 19476 47272
rect 19684 47258 19766 47272
rect 20642 47258 20724 47272
rect 20932 47258 21014 47272
rect 21890 47258 21972 47272
rect 22180 47258 22262 47272
rect 23138 47258 23220 47272
rect 23428 47258 23510 47272
rect 24386 47258 24468 47272
rect 24676 47258 24758 47272
rect 25634 47258 25716 47272
rect 25924 47258 26006 47272
rect 26882 47258 26964 47272
rect 27172 47258 27254 47272
rect 28130 47258 28212 47272
rect 28420 47258 28502 47272
rect 29378 47258 29460 47272
rect 29668 47258 29750 47272
rect 30626 47258 30708 47272
rect 30916 47258 30998 47272
rect 31874 47258 31956 47272
rect 32164 47258 32246 47272
rect 33122 47258 33204 47272
rect 33412 47258 33494 47272
rect 34370 47258 34452 47272
rect 34660 47258 34742 47272
rect 35618 47258 35700 47272
rect 35908 47258 35990 47272
rect 36866 47258 36948 47272
rect 37156 47258 37238 47272
rect 38114 47258 38196 47272
rect 38404 47258 38486 47272
rect 39362 47258 39444 47272
rect 39652 47258 39734 47272
rect 40610 47258 40692 47272
rect 40900 47258 40982 47272
rect 41858 47258 41940 47272
rect 42148 47258 42230 47272
rect 43106 47258 43188 47272
rect 43396 47258 43478 47272
rect 44354 47258 44436 47272
rect 44644 47258 44726 47272
rect 45602 47258 45684 47272
rect 45892 47258 45974 47272
rect 46850 47258 46932 47272
rect 47140 47258 47222 47272
rect 48098 47258 48180 47272
rect 48388 47258 48470 47272
rect 49346 47258 49428 47272
rect 49636 47258 49718 47272
rect 50594 47258 50676 47272
rect 50884 47258 50966 47272
rect 51842 47258 51924 47272
rect 52132 47258 52214 47272
rect 53090 47258 53172 47272
rect 53380 47258 53462 47272
rect 54338 47258 54420 47272
rect 54628 47258 54710 47272
rect 55586 47258 55668 47272
rect 55876 47258 55958 47272
rect 56834 47258 56916 47272
rect 57124 47258 57206 47272
rect 58082 47258 58164 47272
rect 58372 47258 58454 47272
rect 16418 47210 16864 47224
rect 17014 47210 17154 47224
rect 17304 47210 18112 47224
rect 18262 47210 18402 47224
rect 18552 47210 19360 47224
rect 19510 47210 19650 47224
rect 19800 47210 20608 47224
rect 20758 47210 20898 47224
rect 21048 47210 21856 47224
rect 22006 47210 22146 47224
rect 22296 47210 23104 47224
rect 23254 47210 23394 47224
rect 23544 47210 24352 47224
rect 24502 47210 24642 47224
rect 24792 47210 25600 47224
rect 25750 47210 25890 47224
rect 26040 47210 26848 47224
rect 26998 47210 27138 47224
rect 27288 47210 28096 47224
rect 28246 47210 28386 47224
rect 28536 47210 29344 47224
rect 29494 47210 29634 47224
rect 29784 47210 30592 47224
rect 30742 47210 30882 47224
rect 31032 47210 31840 47224
rect 31990 47210 32130 47224
rect 32280 47210 33088 47224
rect 33238 47210 33378 47224
rect 33528 47210 34336 47224
rect 34486 47210 34626 47224
rect 34776 47210 35584 47224
rect 35734 47210 35874 47224
rect 36024 47210 36832 47224
rect 36982 47210 37122 47224
rect 37272 47210 38080 47224
rect 38230 47210 38370 47224
rect 38520 47210 39328 47224
rect 39478 47210 39618 47224
rect 39768 47210 40576 47224
rect 40726 47210 40866 47224
rect 41016 47210 41824 47224
rect 41974 47210 42114 47224
rect 42264 47210 43072 47224
rect 43222 47210 43362 47224
rect 43512 47210 44320 47224
rect 44470 47210 44610 47224
rect 44760 47210 45568 47224
rect 45718 47210 45858 47224
rect 46008 47210 46816 47224
rect 46966 47210 47106 47224
rect 47256 47210 48064 47224
rect 48214 47210 48354 47224
rect 48504 47210 49312 47224
rect 49462 47210 49602 47224
rect 49752 47210 50560 47224
rect 50710 47210 50850 47224
rect 51000 47210 51808 47224
rect 51958 47210 52098 47224
rect 52248 47210 53056 47224
rect 53206 47210 53346 47224
rect 53496 47210 54304 47224
rect 54454 47210 54594 47224
rect 54744 47210 55552 47224
rect 55702 47210 55842 47224
rect 55992 47210 56800 47224
rect 56950 47210 57090 47224
rect 57240 47210 58048 47224
rect 58198 47210 58338 47224
rect 58488 47210 58934 47224
rect 16418 47162 58934 47210
rect 16418 47148 16864 47162
rect 17014 47148 17154 47162
rect 17304 47148 18112 47162
rect 18262 47148 18402 47162
rect 18552 47148 19360 47162
rect 19510 47148 19650 47162
rect 19800 47148 20608 47162
rect 20758 47148 20898 47162
rect 21048 47148 21856 47162
rect 22006 47148 22146 47162
rect 22296 47148 23104 47162
rect 23254 47148 23394 47162
rect 23544 47148 24352 47162
rect 24502 47148 24642 47162
rect 24792 47148 25600 47162
rect 25750 47148 25890 47162
rect 26040 47148 26848 47162
rect 26998 47148 27138 47162
rect 27288 47148 28096 47162
rect 28246 47148 28386 47162
rect 28536 47148 29344 47162
rect 29494 47148 29634 47162
rect 29784 47148 30592 47162
rect 30742 47148 30882 47162
rect 31032 47148 31840 47162
rect 31990 47148 32130 47162
rect 32280 47148 33088 47162
rect 33238 47148 33378 47162
rect 33528 47148 34336 47162
rect 34486 47148 34626 47162
rect 34776 47148 35584 47162
rect 35734 47148 35874 47162
rect 36024 47148 36832 47162
rect 36982 47148 37122 47162
rect 37272 47148 38080 47162
rect 38230 47148 38370 47162
rect 38520 47148 39328 47162
rect 39478 47148 39618 47162
rect 39768 47148 40576 47162
rect 40726 47148 40866 47162
rect 41016 47148 41824 47162
rect 41974 47148 42114 47162
rect 42264 47148 43072 47162
rect 43222 47148 43362 47162
rect 43512 47148 44320 47162
rect 44470 47148 44610 47162
rect 44760 47148 45568 47162
rect 45718 47148 45858 47162
rect 46008 47148 46816 47162
rect 46966 47148 47106 47162
rect 47256 47148 48064 47162
rect 48214 47148 48354 47162
rect 48504 47148 49312 47162
rect 49462 47148 49602 47162
rect 49752 47148 50560 47162
rect 50710 47148 50850 47162
rect 51000 47148 51808 47162
rect 51958 47148 52098 47162
rect 52248 47148 53056 47162
rect 53206 47148 53346 47162
rect 53496 47148 54304 47162
rect 54454 47148 54594 47162
rect 54744 47148 55552 47162
rect 55702 47148 55842 47162
rect 55992 47148 56800 47162
rect 56950 47148 57090 47162
rect 57240 47148 58048 47162
rect 58198 47148 58338 47162
rect 58488 47148 58934 47162
rect 16898 47100 16980 47114
rect 17188 47100 17270 47114
rect 18146 47100 18228 47114
rect 18436 47100 18518 47114
rect 19394 47100 19476 47114
rect 19684 47100 19766 47114
rect 20642 47100 20724 47114
rect 20932 47100 21014 47114
rect 21890 47100 21972 47114
rect 22180 47100 22262 47114
rect 23138 47100 23220 47114
rect 23428 47100 23510 47114
rect 24386 47100 24468 47114
rect 24676 47100 24758 47114
rect 25634 47100 25716 47114
rect 25924 47100 26006 47114
rect 26882 47100 26964 47114
rect 27172 47100 27254 47114
rect 28130 47100 28212 47114
rect 28420 47100 28502 47114
rect 29378 47100 29460 47114
rect 29668 47100 29750 47114
rect 30626 47100 30708 47114
rect 30916 47100 30998 47114
rect 31874 47100 31956 47114
rect 32164 47100 32246 47114
rect 33122 47100 33204 47114
rect 33412 47100 33494 47114
rect 34370 47100 34452 47114
rect 34660 47100 34742 47114
rect 35618 47100 35700 47114
rect 35908 47100 35990 47114
rect 36866 47100 36948 47114
rect 37156 47100 37238 47114
rect 38114 47100 38196 47114
rect 38404 47100 38486 47114
rect 39362 47100 39444 47114
rect 39652 47100 39734 47114
rect 40610 47100 40692 47114
rect 40900 47100 40982 47114
rect 41858 47100 41940 47114
rect 42148 47100 42230 47114
rect 43106 47100 43188 47114
rect 43396 47100 43478 47114
rect 44354 47100 44436 47114
rect 44644 47100 44726 47114
rect 45602 47100 45684 47114
rect 45892 47100 45974 47114
rect 46850 47100 46932 47114
rect 47140 47100 47222 47114
rect 48098 47100 48180 47114
rect 48388 47100 48470 47114
rect 49346 47100 49428 47114
rect 49636 47100 49718 47114
rect 50594 47100 50676 47114
rect 50884 47100 50966 47114
rect 51842 47100 51924 47114
rect 52132 47100 52214 47114
rect 53090 47100 53172 47114
rect 53380 47100 53462 47114
rect 54338 47100 54420 47114
rect 54628 47100 54710 47114
rect 55586 47100 55668 47114
rect 55876 47100 55958 47114
rect 56834 47100 56916 47114
rect 57124 47100 57206 47114
rect 58082 47100 58164 47114
rect 58372 47100 58454 47114
rect 16418 47052 58934 47100
rect 16418 46956 58934 47004
rect 16898 46942 16980 46956
rect 17188 46942 17270 46956
rect 18146 46942 18228 46956
rect 18436 46942 18518 46956
rect 19394 46942 19476 46956
rect 19684 46942 19766 46956
rect 20642 46942 20724 46956
rect 20932 46942 21014 46956
rect 21890 46942 21972 46956
rect 22180 46942 22262 46956
rect 23138 46942 23220 46956
rect 23428 46942 23510 46956
rect 24386 46942 24468 46956
rect 24676 46942 24758 46956
rect 25634 46942 25716 46956
rect 25924 46942 26006 46956
rect 26882 46942 26964 46956
rect 27172 46942 27254 46956
rect 28130 46942 28212 46956
rect 28420 46942 28502 46956
rect 29378 46942 29460 46956
rect 29668 46942 29750 46956
rect 30626 46942 30708 46956
rect 30916 46942 30998 46956
rect 31874 46942 31956 46956
rect 32164 46942 32246 46956
rect 33122 46942 33204 46956
rect 33412 46942 33494 46956
rect 34370 46942 34452 46956
rect 34660 46942 34742 46956
rect 35618 46942 35700 46956
rect 35908 46942 35990 46956
rect 36866 46942 36948 46956
rect 37156 46942 37238 46956
rect 38114 46942 38196 46956
rect 38404 46942 38486 46956
rect 39362 46942 39444 46956
rect 39652 46942 39734 46956
rect 40610 46942 40692 46956
rect 40900 46942 40982 46956
rect 41858 46942 41940 46956
rect 42148 46942 42230 46956
rect 43106 46942 43188 46956
rect 43396 46942 43478 46956
rect 44354 46942 44436 46956
rect 44644 46942 44726 46956
rect 45602 46942 45684 46956
rect 45892 46942 45974 46956
rect 46850 46942 46932 46956
rect 47140 46942 47222 46956
rect 48098 46942 48180 46956
rect 48388 46942 48470 46956
rect 49346 46942 49428 46956
rect 49636 46942 49718 46956
rect 50594 46942 50676 46956
rect 50884 46942 50966 46956
rect 51842 46942 51924 46956
rect 52132 46942 52214 46956
rect 53090 46942 53172 46956
rect 53380 46942 53462 46956
rect 54338 46942 54420 46956
rect 54628 46942 54710 46956
rect 55586 46942 55668 46956
rect 55876 46942 55958 46956
rect 56834 46942 56916 46956
rect 57124 46942 57206 46956
rect 58082 46942 58164 46956
rect 58372 46942 58454 46956
rect 16418 46894 16864 46908
rect 17014 46894 17154 46908
rect 17304 46894 18112 46908
rect 18262 46894 18402 46908
rect 18552 46894 19360 46908
rect 19510 46894 19650 46908
rect 19800 46894 20608 46908
rect 20758 46894 20898 46908
rect 21048 46894 21856 46908
rect 22006 46894 22146 46908
rect 22296 46894 23104 46908
rect 23254 46894 23394 46908
rect 23544 46894 24352 46908
rect 24502 46894 24642 46908
rect 24792 46894 25600 46908
rect 25750 46894 25890 46908
rect 26040 46894 26848 46908
rect 26998 46894 27138 46908
rect 27288 46894 28096 46908
rect 28246 46894 28386 46908
rect 28536 46894 29344 46908
rect 29494 46894 29634 46908
rect 29784 46894 30592 46908
rect 30742 46894 30882 46908
rect 31032 46894 31840 46908
rect 31990 46894 32130 46908
rect 32280 46894 33088 46908
rect 33238 46894 33378 46908
rect 33528 46894 34336 46908
rect 34486 46894 34626 46908
rect 34776 46894 35584 46908
rect 35734 46894 35874 46908
rect 36024 46894 36832 46908
rect 36982 46894 37122 46908
rect 37272 46894 38080 46908
rect 38230 46894 38370 46908
rect 38520 46894 39328 46908
rect 39478 46894 39618 46908
rect 39768 46894 40576 46908
rect 40726 46894 40866 46908
rect 41016 46894 41824 46908
rect 41974 46894 42114 46908
rect 42264 46894 43072 46908
rect 43222 46894 43362 46908
rect 43512 46894 44320 46908
rect 44470 46894 44610 46908
rect 44760 46894 45568 46908
rect 45718 46894 45858 46908
rect 46008 46894 46816 46908
rect 46966 46894 47106 46908
rect 47256 46894 48064 46908
rect 48214 46894 48354 46908
rect 48504 46894 49312 46908
rect 49462 46894 49602 46908
rect 49752 46894 50560 46908
rect 50710 46894 50850 46908
rect 51000 46894 51808 46908
rect 51958 46894 52098 46908
rect 52248 46894 53056 46908
rect 53206 46894 53346 46908
rect 53496 46894 54304 46908
rect 54454 46894 54594 46908
rect 54744 46894 55552 46908
rect 55702 46894 55842 46908
rect 55992 46894 56800 46908
rect 56950 46894 57090 46908
rect 57240 46894 58048 46908
rect 58198 46894 58338 46908
rect 58488 46894 58934 46908
rect 16418 46846 58934 46894
rect 16418 46832 16864 46846
rect 17014 46832 17154 46846
rect 17304 46832 18112 46846
rect 18262 46832 18402 46846
rect 18552 46832 19360 46846
rect 19510 46832 19650 46846
rect 19800 46832 20608 46846
rect 20758 46832 20898 46846
rect 21048 46832 21856 46846
rect 22006 46832 22146 46846
rect 22296 46832 23104 46846
rect 23254 46832 23394 46846
rect 23544 46832 24352 46846
rect 24502 46832 24642 46846
rect 24792 46832 25600 46846
rect 25750 46832 25890 46846
rect 26040 46832 26848 46846
rect 26998 46832 27138 46846
rect 27288 46832 28096 46846
rect 28246 46832 28386 46846
rect 28536 46832 29344 46846
rect 29494 46832 29634 46846
rect 29784 46832 30592 46846
rect 30742 46832 30882 46846
rect 31032 46832 31840 46846
rect 31990 46832 32130 46846
rect 32280 46832 33088 46846
rect 33238 46832 33378 46846
rect 33528 46832 34336 46846
rect 34486 46832 34626 46846
rect 34776 46832 35584 46846
rect 35734 46832 35874 46846
rect 36024 46832 36832 46846
rect 36982 46832 37122 46846
rect 37272 46832 38080 46846
rect 38230 46832 38370 46846
rect 38520 46832 39328 46846
rect 39478 46832 39618 46846
rect 39768 46832 40576 46846
rect 40726 46832 40866 46846
rect 41016 46832 41824 46846
rect 41974 46832 42114 46846
rect 42264 46832 43072 46846
rect 43222 46832 43362 46846
rect 43512 46832 44320 46846
rect 44470 46832 44610 46846
rect 44760 46832 45568 46846
rect 45718 46832 45858 46846
rect 46008 46832 46816 46846
rect 46966 46832 47106 46846
rect 47256 46832 48064 46846
rect 48214 46832 48354 46846
rect 48504 46832 49312 46846
rect 49462 46832 49602 46846
rect 49752 46832 50560 46846
rect 50710 46832 50850 46846
rect 51000 46832 51808 46846
rect 51958 46832 52098 46846
rect 52248 46832 53056 46846
rect 53206 46832 53346 46846
rect 53496 46832 54304 46846
rect 54454 46832 54594 46846
rect 54744 46832 55552 46846
rect 55702 46832 55842 46846
rect 55992 46832 56800 46846
rect 56950 46832 57090 46846
rect 57240 46832 58048 46846
rect 58198 46832 58338 46846
rect 58488 46832 58934 46846
rect 16898 46784 16980 46798
rect 17188 46784 17270 46798
rect 18146 46784 18228 46798
rect 18436 46784 18518 46798
rect 19394 46784 19476 46798
rect 19684 46784 19766 46798
rect 20642 46784 20724 46798
rect 20932 46784 21014 46798
rect 21890 46784 21972 46798
rect 22180 46784 22262 46798
rect 23138 46784 23220 46798
rect 23428 46784 23510 46798
rect 24386 46784 24468 46798
rect 24676 46784 24758 46798
rect 25634 46784 25716 46798
rect 25924 46784 26006 46798
rect 26882 46784 26964 46798
rect 27172 46784 27254 46798
rect 28130 46784 28212 46798
rect 28420 46784 28502 46798
rect 29378 46784 29460 46798
rect 29668 46784 29750 46798
rect 30626 46784 30708 46798
rect 30916 46784 30998 46798
rect 31874 46784 31956 46798
rect 32164 46784 32246 46798
rect 33122 46784 33204 46798
rect 33412 46784 33494 46798
rect 34370 46784 34452 46798
rect 34660 46784 34742 46798
rect 35618 46784 35700 46798
rect 35908 46784 35990 46798
rect 36866 46784 36948 46798
rect 37156 46784 37238 46798
rect 38114 46784 38196 46798
rect 38404 46784 38486 46798
rect 39362 46784 39444 46798
rect 39652 46784 39734 46798
rect 40610 46784 40692 46798
rect 40900 46784 40982 46798
rect 41858 46784 41940 46798
rect 42148 46784 42230 46798
rect 43106 46784 43188 46798
rect 43396 46784 43478 46798
rect 44354 46784 44436 46798
rect 44644 46784 44726 46798
rect 45602 46784 45684 46798
rect 45892 46784 45974 46798
rect 46850 46784 46932 46798
rect 47140 46784 47222 46798
rect 48098 46784 48180 46798
rect 48388 46784 48470 46798
rect 49346 46784 49428 46798
rect 49636 46784 49718 46798
rect 50594 46784 50676 46798
rect 50884 46784 50966 46798
rect 51842 46784 51924 46798
rect 52132 46784 52214 46798
rect 53090 46784 53172 46798
rect 53380 46784 53462 46798
rect 54338 46784 54420 46798
rect 54628 46784 54710 46798
rect 55586 46784 55668 46798
rect 55876 46784 55958 46798
rect 56834 46784 56916 46798
rect 57124 46784 57206 46798
rect 58082 46784 58164 46798
rect 58372 46784 58454 46798
rect 16418 46736 58934 46784
rect 16418 46578 58934 46688
rect 16418 46482 58934 46530
rect 16898 46468 16980 46482
rect 17188 46468 17270 46482
rect 18146 46468 18228 46482
rect 18436 46468 18518 46482
rect 19394 46468 19476 46482
rect 19684 46468 19766 46482
rect 20642 46468 20724 46482
rect 20932 46468 21014 46482
rect 21890 46468 21972 46482
rect 22180 46468 22262 46482
rect 23138 46468 23220 46482
rect 23428 46468 23510 46482
rect 24386 46468 24468 46482
rect 24676 46468 24758 46482
rect 25634 46468 25716 46482
rect 25924 46468 26006 46482
rect 26882 46468 26964 46482
rect 27172 46468 27254 46482
rect 28130 46468 28212 46482
rect 28420 46468 28502 46482
rect 29378 46468 29460 46482
rect 29668 46468 29750 46482
rect 30626 46468 30708 46482
rect 30916 46468 30998 46482
rect 31874 46468 31956 46482
rect 32164 46468 32246 46482
rect 33122 46468 33204 46482
rect 33412 46468 33494 46482
rect 34370 46468 34452 46482
rect 34660 46468 34742 46482
rect 35618 46468 35700 46482
rect 35908 46468 35990 46482
rect 36866 46468 36948 46482
rect 37156 46468 37238 46482
rect 38114 46468 38196 46482
rect 38404 46468 38486 46482
rect 39362 46468 39444 46482
rect 39652 46468 39734 46482
rect 40610 46468 40692 46482
rect 40900 46468 40982 46482
rect 41858 46468 41940 46482
rect 42148 46468 42230 46482
rect 43106 46468 43188 46482
rect 43396 46468 43478 46482
rect 44354 46468 44436 46482
rect 44644 46468 44726 46482
rect 45602 46468 45684 46482
rect 45892 46468 45974 46482
rect 46850 46468 46932 46482
rect 47140 46468 47222 46482
rect 48098 46468 48180 46482
rect 48388 46468 48470 46482
rect 49346 46468 49428 46482
rect 49636 46468 49718 46482
rect 50594 46468 50676 46482
rect 50884 46468 50966 46482
rect 51842 46468 51924 46482
rect 52132 46468 52214 46482
rect 53090 46468 53172 46482
rect 53380 46468 53462 46482
rect 54338 46468 54420 46482
rect 54628 46468 54710 46482
rect 55586 46468 55668 46482
rect 55876 46468 55958 46482
rect 56834 46468 56916 46482
rect 57124 46468 57206 46482
rect 58082 46468 58164 46482
rect 58372 46468 58454 46482
rect 16418 46420 16864 46434
rect 17014 46420 17154 46434
rect 17304 46420 18112 46434
rect 18262 46420 18402 46434
rect 18552 46420 19360 46434
rect 19510 46420 19650 46434
rect 19800 46420 20608 46434
rect 20758 46420 20898 46434
rect 21048 46420 21856 46434
rect 22006 46420 22146 46434
rect 22296 46420 23104 46434
rect 23254 46420 23394 46434
rect 23544 46420 24352 46434
rect 24502 46420 24642 46434
rect 24792 46420 25600 46434
rect 25750 46420 25890 46434
rect 26040 46420 26848 46434
rect 26998 46420 27138 46434
rect 27288 46420 28096 46434
rect 28246 46420 28386 46434
rect 28536 46420 29344 46434
rect 29494 46420 29634 46434
rect 29784 46420 30592 46434
rect 30742 46420 30882 46434
rect 31032 46420 31840 46434
rect 31990 46420 32130 46434
rect 32280 46420 33088 46434
rect 33238 46420 33378 46434
rect 33528 46420 34336 46434
rect 34486 46420 34626 46434
rect 34776 46420 35584 46434
rect 35734 46420 35874 46434
rect 36024 46420 36832 46434
rect 36982 46420 37122 46434
rect 37272 46420 38080 46434
rect 38230 46420 38370 46434
rect 38520 46420 39328 46434
rect 39478 46420 39618 46434
rect 39768 46420 40576 46434
rect 40726 46420 40866 46434
rect 41016 46420 41824 46434
rect 41974 46420 42114 46434
rect 42264 46420 43072 46434
rect 43222 46420 43362 46434
rect 43512 46420 44320 46434
rect 44470 46420 44610 46434
rect 44760 46420 45568 46434
rect 45718 46420 45858 46434
rect 46008 46420 46816 46434
rect 46966 46420 47106 46434
rect 47256 46420 48064 46434
rect 48214 46420 48354 46434
rect 48504 46420 49312 46434
rect 49462 46420 49602 46434
rect 49752 46420 50560 46434
rect 50710 46420 50850 46434
rect 51000 46420 51808 46434
rect 51958 46420 52098 46434
rect 52248 46420 53056 46434
rect 53206 46420 53346 46434
rect 53496 46420 54304 46434
rect 54454 46420 54594 46434
rect 54744 46420 55552 46434
rect 55702 46420 55842 46434
rect 55992 46420 56800 46434
rect 56950 46420 57090 46434
rect 57240 46420 58048 46434
rect 58198 46420 58338 46434
rect 58488 46420 58934 46434
rect 16418 46372 58934 46420
rect 16418 46358 16864 46372
rect 17014 46358 17154 46372
rect 17304 46358 18112 46372
rect 18262 46358 18402 46372
rect 18552 46358 19360 46372
rect 19510 46358 19650 46372
rect 19800 46358 20608 46372
rect 20758 46358 20898 46372
rect 21048 46358 21856 46372
rect 22006 46358 22146 46372
rect 22296 46358 23104 46372
rect 23254 46358 23394 46372
rect 23544 46358 24352 46372
rect 24502 46358 24642 46372
rect 24792 46358 25600 46372
rect 25750 46358 25890 46372
rect 26040 46358 26848 46372
rect 26998 46358 27138 46372
rect 27288 46358 28096 46372
rect 28246 46358 28386 46372
rect 28536 46358 29344 46372
rect 29494 46358 29634 46372
rect 29784 46358 30592 46372
rect 30742 46358 30882 46372
rect 31032 46358 31840 46372
rect 31990 46358 32130 46372
rect 32280 46358 33088 46372
rect 33238 46358 33378 46372
rect 33528 46358 34336 46372
rect 34486 46358 34626 46372
rect 34776 46358 35584 46372
rect 35734 46358 35874 46372
rect 36024 46358 36832 46372
rect 36982 46358 37122 46372
rect 37272 46358 38080 46372
rect 38230 46358 38370 46372
rect 38520 46358 39328 46372
rect 39478 46358 39618 46372
rect 39768 46358 40576 46372
rect 40726 46358 40866 46372
rect 41016 46358 41824 46372
rect 41974 46358 42114 46372
rect 42264 46358 43072 46372
rect 43222 46358 43362 46372
rect 43512 46358 44320 46372
rect 44470 46358 44610 46372
rect 44760 46358 45568 46372
rect 45718 46358 45858 46372
rect 46008 46358 46816 46372
rect 46966 46358 47106 46372
rect 47256 46358 48064 46372
rect 48214 46358 48354 46372
rect 48504 46358 49312 46372
rect 49462 46358 49602 46372
rect 49752 46358 50560 46372
rect 50710 46358 50850 46372
rect 51000 46358 51808 46372
rect 51958 46358 52098 46372
rect 52248 46358 53056 46372
rect 53206 46358 53346 46372
rect 53496 46358 54304 46372
rect 54454 46358 54594 46372
rect 54744 46358 55552 46372
rect 55702 46358 55842 46372
rect 55992 46358 56800 46372
rect 56950 46358 57090 46372
rect 57240 46358 58048 46372
rect 58198 46358 58338 46372
rect 58488 46358 58934 46372
rect 16898 46310 16980 46324
rect 17188 46310 17270 46324
rect 18146 46310 18228 46324
rect 18436 46310 18518 46324
rect 19394 46310 19476 46324
rect 19684 46310 19766 46324
rect 20642 46310 20724 46324
rect 20932 46310 21014 46324
rect 21890 46310 21972 46324
rect 22180 46310 22262 46324
rect 23138 46310 23220 46324
rect 23428 46310 23510 46324
rect 24386 46310 24468 46324
rect 24676 46310 24758 46324
rect 25634 46310 25716 46324
rect 25924 46310 26006 46324
rect 26882 46310 26964 46324
rect 27172 46310 27254 46324
rect 28130 46310 28212 46324
rect 28420 46310 28502 46324
rect 29378 46310 29460 46324
rect 29668 46310 29750 46324
rect 30626 46310 30708 46324
rect 30916 46310 30998 46324
rect 31874 46310 31956 46324
rect 32164 46310 32246 46324
rect 33122 46310 33204 46324
rect 33412 46310 33494 46324
rect 34370 46310 34452 46324
rect 34660 46310 34742 46324
rect 35618 46310 35700 46324
rect 35908 46310 35990 46324
rect 36866 46310 36948 46324
rect 37156 46310 37238 46324
rect 38114 46310 38196 46324
rect 38404 46310 38486 46324
rect 39362 46310 39444 46324
rect 39652 46310 39734 46324
rect 40610 46310 40692 46324
rect 40900 46310 40982 46324
rect 41858 46310 41940 46324
rect 42148 46310 42230 46324
rect 43106 46310 43188 46324
rect 43396 46310 43478 46324
rect 44354 46310 44436 46324
rect 44644 46310 44726 46324
rect 45602 46310 45684 46324
rect 45892 46310 45974 46324
rect 46850 46310 46932 46324
rect 47140 46310 47222 46324
rect 48098 46310 48180 46324
rect 48388 46310 48470 46324
rect 49346 46310 49428 46324
rect 49636 46310 49718 46324
rect 50594 46310 50676 46324
rect 50884 46310 50966 46324
rect 51842 46310 51924 46324
rect 52132 46310 52214 46324
rect 53090 46310 53172 46324
rect 53380 46310 53462 46324
rect 54338 46310 54420 46324
rect 54628 46310 54710 46324
rect 55586 46310 55668 46324
rect 55876 46310 55958 46324
rect 56834 46310 56916 46324
rect 57124 46310 57206 46324
rect 58082 46310 58164 46324
rect 58372 46310 58454 46324
rect 16418 46262 58934 46310
rect 16418 46166 58934 46214
rect 16898 46152 16980 46166
rect 17188 46152 17270 46166
rect 18146 46152 18228 46166
rect 18436 46152 18518 46166
rect 19394 46152 19476 46166
rect 19684 46152 19766 46166
rect 20642 46152 20724 46166
rect 20932 46152 21014 46166
rect 21890 46152 21972 46166
rect 22180 46152 22262 46166
rect 23138 46152 23220 46166
rect 23428 46152 23510 46166
rect 24386 46152 24468 46166
rect 24676 46152 24758 46166
rect 25634 46152 25716 46166
rect 25924 46152 26006 46166
rect 26882 46152 26964 46166
rect 27172 46152 27254 46166
rect 28130 46152 28212 46166
rect 28420 46152 28502 46166
rect 29378 46152 29460 46166
rect 29668 46152 29750 46166
rect 30626 46152 30708 46166
rect 30916 46152 30998 46166
rect 31874 46152 31956 46166
rect 32164 46152 32246 46166
rect 33122 46152 33204 46166
rect 33412 46152 33494 46166
rect 34370 46152 34452 46166
rect 34660 46152 34742 46166
rect 35618 46152 35700 46166
rect 35908 46152 35990 46166
rect 36866 46152 36948 46166
rect 37156 46152 37238 46166
rect 38114 46152 38196 46166
rect 38404 46152 38486 46166
rect 39362 46152 39444 46166
rect 39652 46152 39734 46166
rect 40610 46152 40692 46166
rect 40900 46152 40982 46166
rect 41858 46152 41940 46166
rect 42148 46152 42230 46166
rect 43106 46152 43188 46166
rect 43396 46152 43478 46166
rect 44354 46152 44436 46166
rect 44644 46152 44726 46166
rect 45602 46152 45684 46166
rect 45892 46152 45974 46166
rect 46850 46152 46932 46166
rect 47140 46152 47222 46166
rect 48098 46152 48180 46166
rect 48388 46152 48470 46166
rect 49346 46152 49428 46166
rect 49636 46152 49718 46166
rect 50594 46152 50676 46166
rect 50884 46152 50966 46166
rect 51842 46152 51924 46166
rect 52132 46152 52214 46166
rect 53090 46152 53172 46166
rect 53380 46152 53462 46166
rect 54338 46152 54420 46166
rect 54628 46152 54710 46166
rect 55586 46152 55668 46166
rect 55876 46152 55958 46166
rect 56834 46152 56916 46166
rect 57124 46152 57206 46166
rect 58082 46152 58164 46166
rect 58372 46152 58454 46166
rect 16418 46104 16864 46118
rect 17014 46104 17154 46118
rect 17304 46104 18112 46118
rect 18262 46104 18402 46118
rect 18552 46104 19360 46118
rect 19510 46104 19650 46118
rect 19800 46104 20608 46118
rect 20758 46104 20898 46118
rect 21048 46104 21856 46118
rect 22006 46104 22146 46118
rect 22296 46104 23104 46118
rect 23254 46104 23394 46118
rect 23544 46104 24352 46118
rect 24502 46104 24642 46118
rect 24792 46104 25600 46118
rect 25750 46104 25890 46118
rect 26040 46104 26848 46118
rect 26998 46104 27138 46118
rect 27288 46104 28096 46118
rect 28246 46104 28386 46118
rect 28536 46104 29344 46118
rect 29494 46104 29634 46118
rect 29784 46104 30592 46118
rect 30742 46104 30882 46118
rect 31032 46104 31840 46118
rect 31990 46104 32130 46118
rect 32280 46104 33088 46118
rect 33238 46104 33378 46118
rect 33528 46104 34336 46118
rect 34486 46104 34626 46118
rect 34776 46104 35584 46118
rect 35734 46104 35874 46118
rect 36024 46104 36832 46118
rect 36982 46104 37122 46118
rect 37272 46104 38080 46118
rect 38230 46104 38370 46118
rect 38520 46104 39328 46118
rect 39478 46104 39618 46118
rect 39768 46104 40576 46118
rect 40726 46104 40866 46118
rect 41016 46104 41824 46118
rect 41974 46104 42114 46118
rect 42264 46104 43072 46118
rect 43222 46104 43362 46118
rect 43512 46104 44320 46118
rect 44470 46104 44610 46118
rect 44760 46104 45568 46118
rect 45718 46104 45858 46118
rect 46008 46104 46816 46118
rect 46966 46104 47106 46118
rect 47256 46104 48064 46118
rect 48214 46104 48354 46118
rect 48504 46104 49312 46118
rect 49462 46104 49602 46118
rect 49752 46104 50560 46118
rect 50710 46104 50850 46118
rect 51000 46104 51808 46118
rect 51958 46104 52098 46118
rect 52248 46104 53056 46118
rect 53206 46104 53346 46118
rect 53496 46104 54304 46118
rect 54454 46104 54594 46118
rect 54744 46104 55552 46118
rect 55702 46104 55842 46118
rect 55992 46104 56800 46118
rect 56950 46104 57090 46118
rect 57240 46104 58048 46118
rect 58198 46104 58338 46118
rect 58488 46104 58934 46118
rect 16418 46056 58934 46104
rect 16418 46042 16864 46056
rect 17014 46042 17154 46056
rect 17304 46042 18112 46056
rect 18262 46042 18402 46056
rect 18552 46042 19360 46056
rect 19510 46042 19650 46056
rect 19800 46042 20608 46056
rect 20758 46042 20898 46056
rect 21048 46042 21856 46056
rect 22006 46042 22146 46056
rect 22296 46042 23104 46056
rect 23254 46042 23394 46056
rect 23544 46042 24352 46056
rect 24502 46042 24642 46056
rect 24792 46042 25600 46056
rect 25750 46042 25890 46056
rect 26040 46042 26848 46056
rect 26998 46042 27138 46056
rect 27288 46042 28096 46056
rect 28246 46042 28386 46056
rect 28536 46042 29344 46056
rect 29494 46042 29634 46056
rect 29784 46042 30592 46056
rect 30742 46042 30882 46056
rect 31032 46042 31840 46056
rect 31990 46042 32130 46056
rect 32280 46042 33088 46056
rect 33238 46042 33378 46056
rect 33528 46042 34336 46056
rect 34486 46042 34626 46056
rect 34776 46042 35584 46056
rect 35734 46042 35874 46056
rect 36024 46042 36832 46056
rect 36982 46042 37122 46056
rect 37272 46042 38080 46056
rect 38230 46042 38370 46056
rect 38520 46042 39328 46056
rect 39478 46042 39618 46056
rect 39768 46042 40576 46056
rect 40726 46042 40866 46056
rect 41016 46042 41824 46056
rect 41974 46042 42114 46056
rect 42264 46042 43072 46056
rect 43222 46042 43362 46056
rect 43512 46042 44320 46056
rect 44470 46042 44610 46056
rect 44760 46042 45568 46056
rect 45718 46042 45858 46056
rect 46008 46042 46816 46056
rect 46966 46042 47106 46056
rect 47256 46042 48064 46056
rect 48214 46042 48354 46056
rect 48504 46042 49312 46056
rect 49462 46042 49602 46056
rect 49752 46042 50560 46056
rect 50710 46042 50850 46056
rect 51000 46042 51808 46056
rect 51958 46042 52098 46056
rect 52248 46042 53056 46056
rect 53206 46042 53346 46056
rect 53496 46042 54304 46056
rect 54454 46042 54594 46056
rect 54744 46042 55552 46056
rect 55702 46042 55842 46056
rect 55992 46042 56800 46056
rect 56950 46042 57090 46056
rect 57240 46042 58048 46056
rect 58198 46042 58338 46056
rect 58488 46042 58934 46056
rect 16898 45994 16980 46008
rect 17188 45994 17270 46008
rect 18146 45994 18228 46008
rect 18436 45994 18518 46008
rect 19394 45994 19476 46008
rect 19684 45994 19766 46008
rect 20642 45994 20724 46008
rect 20932 45994 21014 46008
rect 21890 45994 21972 46008
rect 22180 45994 22262 46008
rect 23138 45994 23220 46008
rect 23428 45994 23510 46008
rect 24386 45994 24468 46008
rect 24676 45994 24758 46008
rect 25634 45994 25716 46008
rect 25924 45994 26006 46008
rect 26882 45994 26964 46008
rect 27172 45994 27254 46008
rect 28130 45994 28212 46008
rect 28420 45994 28502 46008
rect 29378 45994 29460 46008
rect 29668 45994 29750 46008
rect 30626 45994 30708 46008
rect 30916 45994 30998 46008
rect 31874 45994 31956 46008
rect 32164 45994 32246 46008
rect 33122 45994 33204 46008
rect 33412 45994 33494 46008
rect 34370 45994 34452 46008
rect 34660 45994 34742 46008
rect 35618 45994 35700 46008
rect 35908 45994 35990 46008
rect 36866 45994 36948 46008
rect 37156 45994 37238 46008
rect 38114 45994 38196 46008
rect 38404 45994 38486 46008
rect 39362 45994 39444 46008
rect 39652 45994 39734 46008
rect 40610 45994 40692 46008
rect 40900 45994 40982 46008
rect 41858 45994 41940 46008
rect 42148 45994 42230 46008
rect 43106 45994 43188 46008
rect 43396 45994 43478 46008
rect 44354 45994 44436 46008
rect 44644 45994 44726 46008
rect 45602 45994 45684 46008
rect 45892 45994 45974 46008
rect 46850 45994 46932 46008
rect 47140 45994 47222 46008
rect 48098 45994 48180 46008
rect 48388 45994 48470 46008
rect 49346 45994 49428 46008
rect 49636 45994 49718 46008
rect 50594 45994 50676 46008
rect 50884 45994 50966 46008
rect 51842 45994 51924 46008
rect 52132 45994 52214 46008
rect 53090 45994 53172 46008
rect 53380 45994 53462 46008
rect 54338 45994 54420 46008
rect 54628 45994 54710 46008
rect 55586 45994 55668 46008
rect 55876 45994 55958 46008
rect 56834 45994 56916 46008
rect 57124 45994 57206 46008
rect 58082 45994 58164 46008
rect 58372 45994 58454 46008
rect 16418 45946 58934 45994
rect 16418 45788 58934 45898
rect 16418 45692 58934 45740
rect 16898 45678 16980 45692
rect 17188 45678 17270 45692
rect 18146 45678 18228 45692
rect 18436 45678 18518 45692
rect 19394 45678 19476 45692
rect 19684 45678 19766 45692
rect 20642 45678 20724 45692
rect 20932 45678 21014 45692
rect 21890 45678 21972 45692
rect 22180 45678 22262 45692
rect 23138 45678 23220 45692
rect 23428 45678 23510 45692
rect 24386 45678 24468 45692
rect 24676 45678 24758 45692
rect 25634 45678 25716 45692
rect 25924 45678 26006 45692
rect 26882 45678 26964 45692
rect 27172 45678 27254 45692
rect 28130 45678 28212 45692
rect 28420 45678 28502 45692
rect 29378 45678 29460 45692
rect 29668 45678 29750 45692
rect 30626 45678 30708 45692
rect 30916 45678 30998 45692
rect 31874 45678 31956 45692
rect 32164 45678 32246 45692
rect 33122 45678 33204 45692
rect 33412 45678 33494 45692
rect 34370 45678 34452 45692
rect 34660 45678 34742 45692
rect 35618 45678 35700 45692
rect 35908 45678 35990 45692
rect 36866 45678 36948 45692
rect 37156 45678 37238 45692
rect 38114 45678 38196 45692
rect 38404 45678 38486 45692
rect 39362 45678 39444 45692
rect 39652 45678 39734 45692
rect 40610 45678 40692 45692
rect 40900 45678 40982 45692
rect 41858 45678 41940 45692
rect 42148 45678 42230 45692
rect 43106 45678 43188 45692
rect 43396 45678 43478 45692
rect 44354 45678 44436 45692
rect 44644 45678 44726 45692
rect 45602 45678 45684 45692
rect 45892 45678 45974 45692
rect 46850 45678 46932 45692
rect 47140 45678 47222 45692
rect 48098 45678 48180 45692
rect 48388 45678 48470 45692
rect 49346 45678 49428 45692
rect 49636 45678 49718 45692
rect 50594 45678 50676 45692
rect 50884 45678 50966 45692
rect 51842 45678 51924 45692
rect 52132 45678 52214 45692
rect 53090 45678 53172 45692
rect 53380 45678 53462 45692
rect 54338 45678 54420 45692
rect 54628 45678 54710 45692
rect 55586 45678 55668 45692
rect 55876 45678 55958 45692
rect 56834 45678 56916 45692
rect 57124 45678 57206 45692
rect 58082 45678 58164 45692
rect 58372 45678 58454 45692
rect 16418 45630 16864 45644
rect 17014 45630 17154 45644
rect 17304 45630 18112 45644
rect 18262 45630 18402 45644
rect 18552 45630 19360 45644
rect 19510 45630 19650 45644
rect 19800 45630 20608 45644
rect 20758 45630 20898 45644
rect 21048 45630 21856 45644
rect 22006 45630 22146 45644
rect 22296 45630 23104 45644
rect 23254 45630 23394 45644
rect 23544 45630 24352 45644
rect 24502 45630 24642 45644
rect 24792 45630 25600 45644
rect 25750 45630 25890 45644
rect 26040 45630 26848 45644
rect 26998 45630 27138 45644
rect 27288 45630 28096 45644
rect 28246 45630 28386 45644
rect 28536 45630 29344 45644
rect 29494 45630 29634 45644
rect 29784 45630 30592 45644
rect 30742 45630 30882 45644
rect 31032 45630 31840 45644
rect 31990 45630 32130 45644
rect 32280 45630 33088 45644
rect 33238 45630 33378 45644
rect 33528 45630 34336 45644
rect 34486 45630 34626 45644
rect 34776 45630 35584 45644
rect 35734 45630 35874 45644
rect 36024 45630 36832 45644
rect 36982 45630 37122 45644
rect 37272 45630 38080 45644
rect 38230 45630 38370 45644
rect 38520 45630 39328 45644
rect 39478 45630 39618 45644
rect 39768 45630 40576 45644
rect 40726 45630 40866 45644
rect 41016 45630 41824 45644
rect 41974 45630 42114 45644
rect 42264 45630 43072 45644
rect 43222 45630 43362 45644
rect 43512 45630 44320 45644
rect 44470 45630 44610 45644
rect 44760 45630 45568 45644
rect 45718 45630 45858 45644
rect 46008 45630 46816 45644
rect 46966 45630 47106 45644
rect 47256 45630 48064 45644
rect 48214 45630 48354 45644
rect 48504 45630 49312 45644
rect 49462 45630 49602 45644
rect 49752 45630 50560 45644
rect 50710 45630 50850 45644
rect 51000 45630 51808 45644
rect 51958 45630 52098 45644
rect 52248 45630 53056 45644
rect 53206 45630 53346 45644
rect 53496 45630 54304 45644
rect 54454 45630 54594 45644
rect 54744 45630 55552 45644
rect 55702 45630 55842 45644
rect 55992 45630 56800 45644
rect 56950 45630 57090 45644
rect 57240 45630 58048 45644
rect 58198 45630 58338 45644
rect 58488 45630 58934 45644
rect 16418 45582 58934 45630
rect 16418 45568 16864 45582
rect 17014 45568 17154 45582
rect 17304 45568 18112 45582
rect 18262 45568 18402 45582
rect 18552 45568 19360 45582
rect 19510 45568 19650 45582
rect 19800 45568 20608 45582
rect 20758 45568 20898 45582
rect 21048 45568 21856 45582
rect 22006 45568 22146 45582
rect 22296 45568 23104 45582
rect 23254 45568 23394 45582
rect 23544 45568 24352 45582
rect 24502 45568 24642 45582
rect 24792 45568 25600 45582
rect 25750 45568 25890 45582
rect 26040 45568 26848 45582
rect 26998 45568 27138 45582
rect 27288 45568 28096 45582
rect 28246 45568 28386 45582
rect 28536 45568 29344 45582
rect 29494 45568 29634 45582
rect 29784 45568 30592 45582
rect 30742 45568 30882 45582
rect 31032 45568 31840 45582
rect 31990 45568 32130 45582
rect 32280 45568 33088 45582
rect 33238 45568 33378 45582
rect 33528 45568 34336 45582
rect 34486 45568 34626 45582
rect 34776 45568 35584 45582
rect 35734 45568 35874 45582
rect 36024 45568 36832 45582
rect 36982 45568 37122 45582
rect 37272 45568 38080 45582
rect 38230 45568 38370 45582
rect 38520 45568 39328 45582
rect 39478 45568 39618 45582
rect 39768 45568 40576 45582
rect 40726 45568 40866 45582
rect 41016 45568 41824 45582
rect 41974 45568 42114 45582
rect 42264 45568 43072 45582
rect 43222 45568 43362 45582
rect 43512 45568 44320 45582
rect 44470 45568 44610 45582
rect 44760 45568 45568 45582
rect 45718 45568 45858 45582
rect 46008 45568 46816 45582
rect 46966 45568 47106 45582
rect 47256 45568 48064 45582
rect 48214 45568 48354 45582
rect 48504 45568 49312 45582
rect 49462 45568 49602 45582
rect 49752 45568 50560 45582
rect 50710 45568 50850 45582
rect 51000 45568 51808 45582
rect 51958 45568 52098 45582
rect 52248 45568 53056 45582
rect 53206 45568 53346 45582
rect 53496 45568 54304 45582
rect 54454 45568 54594 45582
rect 54744 45568 55552 45582
rect 55702 45568 55842 45582
rect 55992 45568 56800 45582
rect 56950 45568 57090 45582
rect 57240 45568 58048 45582
rect 58198 45568 58338 45582
rect 58488 45568 58934 45582
rect 16898 45520 16980 45534
rect 17188 45520 17270 45534
rect 18146 45520 18228 45534
rect 18436 45520 18518 45534
rect 19394 45520 19476 45534
rect 19684 45520 19766 45534
rect 20642 45520 20724 45534
rect 20932 45520 21014 45534
rect 21890 45520 21972 45534
rect 22180 45520 22262 45534
rect 23138 45520 23220 45534
rect 23428 45520 23510 45534
rect 24386 45520 24468 45534
rect 24676 45520 24758 45534
rect 25634 45520 25716 45534
rect 25924 45520 26006 45534
rect 26882 45520 26964 45534
rect 27172 45520 27254 45534
rect 28130 45520 28212 45534
rect 28420 45520 28502 45534
rect 29378 45520 29460 45534
rect 29668 45520 29750 45534
rect 30626 45520 30708 45534
rect 30916 45520 30998 45534
rect 31874 45520 31956 45534
rect 32164 45520 32246 45534
rect 33122 45520 33204 45534
rect 33412 45520 33494 45534
rect 34370 45520 34452 45534
rect 34660 45520 34742 45534
rect 35618 45520 35700 45534
rect 35908 45520 35990 45534
rect 36866 45520 36948 45534
rect 37156 45520 37238 45534
rect 38114 45520 38196 45534
rect 38404 45520 38486 45534
rect 39362 45520 39444 45534
rect 39652 45520 39734 45534
rect 40610 45520 40692 45534
rect 40900 45520 40982 45534
rect 41858 45520 41940 45534
rect 42148 45520 42230 45534
rect 43106 45520 43188 45534
rect 43396 45520 43478 45534
rect 44354 45520 44436 45534
rect 44644 45520 44726 45534
rect 45602 45520 45684 45534
rect 45892 45520 45974 45534
rect 46850 45520 46932 45534
rect 47140 45520 47222 45534
rect 48098 45520 48180 45534
rect 48388 45520 48470 45534
rect 49346 45520 49428 45534
rect 49636 45520 49718 45534
rect 50594 45520 50676 45534
rect 50884 45520 50966 45534
rect 51842 45520 51924 45534
rect 52132 45520 52214 45534
rect 53090 45520 53172 45534
rect 53380 45520 53462 45534
rect 54338 45520 54420 45534
rect 54628 45520 54710 45534
rect 55586 45520 55668 45534
rect 55876 45520 55958 45534
rect 56834 45520 56916 45534
rect 57124 45520 57206 45534
rect 58082 45520 58164 45534
rect 58372 45520 58454 45534
rect 16418 45472 58934 45520
rect 16418 45376 58934 45424
rect 16898 45362 16980 45376
rect 17188 45362 17270 45376
rect 18146 45362 18228 45376
rect 18436 45362 18518 45376
rect 19394 45362 19476 45376
rect 19684 45362 19766 45376
rect 20642 45362 20724 45376
rect 20932 45362 21014 45376
rect 21890 45362 21972 45376
rect 22180 45362 22262 45376
rect 23138 45362 23220 45376
rect 23428 45362 23510 45376
rect 24386 45362 24468 45376
rect 24676 45362 24758 45376
rect 25634 45362 25716 45376
rect 25924 45362 26006 45376
rect 26882 45362 26964 45376
rect 27172 45362 27254 45376
rect 28130 45362 28212 45376
rect 28420 45362 28502 45376
rect 29378 45362 29460 45376
rect 29668 45362 29750 45376
rect 30626 45362 30708 45376
rect 30916 45362 30998 45376
rect 31874 45362 31956 45376
rect 32164 45362 32246 45376
rect 33122 45362 33204 45376
rect 33412 45362 33494 45376
rect 34370 45362 34452 45376
rect 34660 45362 34742 45376
rect 35618 45362 35700 45376
rect 35908 45362 35990 45376
rect 36866 45362 36948 45376
rect 37156 45362 37238 45376
rect 38114 45362 38196 45376
rect 38404 45362 38486 45376
rect 39362 45362 39444 45376
rect 39652 45362 39734 45376
rect 40610 45362 40692 45376
rect 40900 45362 40982 45376
rect 41858 45362 41940 45376
rect 42148 45362 42230 45376
rect 43106 45362 43188 45376
rect 43396 45362 43478 45376
rect 44354 45362 44436 45376
rect 44644 45362 44726 45376
rect 45602 45362 45684 45376
rect 45892 45362 45974 45376
rect 46850 45362 46932 45376
rect 47140 45362 47222 45376
rect 48098 45362 48180 45376
rect 48388 45362 48470 45376
rect 49346 45362 49428 45376
rect 49636 45362 49718 45376
rect 50594 45362 50676 45376
rect 50884 45362 50966 45376
rect 51842 45362 51924 45376
rect 52132 45362 52214 45376
rect 53090 45362 53172 45376
rect 53380 45362 53462 45376
rect 54338 45362 54420 45376
rect 54628 45362 54710 45376
rect 55586 45362 55668 45376
rect 55876 45362 55958 45376
rect 56834 45362 56916 45376
rect 57124 45362 57206 45376
rect 58082 45362 58164 45376
rect 58372 45362 58454 45376
rect 16418 45314 16864 45328
rect 17014 45314 17154 45328
rect 17304 45314 18112 45328
rect 18262 45314 18402 45328
rect 18552 45314 19360 45328
rect 19510 45314 19650 45328
rect 19800 45314 20608 45328
rect 20758 45314 20898 45328
rect 21048 45314 21856 45328
rect 22006 45314 22146 45328
rect 22296 45314 23104 45328
rect 23254 45314 23394 45328
rect 23544 45314 24352 45328
rect 24502 45314 24642 45328
rect 24792 45314 25600 45328
rect 25750 45314 25890 45328
rect 26040 45314 26848 45328
rect 26998 45314 27138 45328
rect 27288 45314 28096 45328
rect 28246 45314 28386 45328
rect 28536 45314 29344 45328
rect 29494 45314 29634 45328
rect 29784 45314 30592 45328
rect 30742 45314 30882 45328
rect 31032 45314 31840 45328
rect 31990 45314 32130 45328
rect 32280 45314 33088 45328
rect 33238 45314 33378 45328
rect 33528 45314 34336 45328
rect 34486 45314 34626 45328
rect 34776 45314 35584 45328
rect 35734 45314 35874 45328
rect 36024 45314 36832 45328
rect 36982 45314 37122 45328
rect 37272 45314 38080 45328
rect 38230 45314 38370 45328
rect 38520 45314 39328 45328
rect 39478 45314 39618 45328
rect 39768 45314 40576 45328
rect 40726 45314 40866 45328
rect 41016 45314 41824 45328
rect 41974 45314 42114 45328
rect 42264 45314 43072 45328
rect 43222 45314 43362 45328
rect 43512 45314 44320 45328
rect 44470 45314 44610 45328
rect 44760 45314 45568 45328
rect 45718 45314 45858 45328
rect 46008 45314 46816 45328
rect 46966 45314 47106 45328
rect 47256 45314 48064 45328
rect 48214 45314 48354 45328
rect 48504 45314 49312 45328
rect 49462 45314 49602 45328
rect 49752 45314 50560 45328
rect 50710 45314 50850 45328
rect 51000 45314 51808 45328
rect 51958 45314 52098 45328
rect 52248 45314 53056 45328
rect 53206 45314 53346 45328
rect 53496 45314 54304 45328
rect 54454 45314 54594 45328
rect 54744 45314 55552 45328
rect 55702 45314 55842 45328
rect 55992 45314 56800 45328
rect 56950 45314 57090 45328
rect 57240 45314 58048 45328
rect 58198 45314 58338 45328
rect 58488 45314 58934 45328
rect 16418 45266 58934 45314
rect 16418 45252 16864 45266
rect 17014 45252 17154 45266
rect 17304 45252 18112 45266
rect 18262 45252 18402 45266
rect 18552 45252 19360 45266
rect 19510 45252 19650 45266
rect 19800 45252 20608 45266
rect 20758 45252 20898 45266
rect 21048 45252 21856 45266
rect 22006 45252 22146 45266
rect 22296 45252 23104 45266
rect 23254 45252 23394 45266
rect 23544 45252 24352 45266
rect 24502 45252 24642 45266
rect 24792 45252 25600 45266
rect 25750 45252 25890 45266
rect 26040 45252 26848 45266
rect 26998 45252 27138 45266
rect 27288 45252 28096 45266
rect 28246 45252 28386 45266
rect 28536 45252 29344 45266
rect 29494 45252 29634 45266
rect 29784 45252 30592 45266
rect 30742 45252 30882 45266
rect 31032 45252 31840 45266
rect 31990 45252 32130 45266
rect 32280 45252 33088 45266
rect 33238 45252 33378 45266
rect 33528 45252 34336 45266
rect 34486 45252 34626 45266
rect 34776 45252 35584 45266
rect 35734 45252 35874 45266
rect 36024 45252 36832 45266
rect 36982 45252 37122 45266
rect 37272 45252 38080 45266
rect 38230 45252 38370 45266
rect 38520 45252 39328 45266
rect 39478 45252 39618 45266
rect 39768 45252 40576 45266
rect 40726 45252 40866 45266
rect 41016 45252 41824 45266
rect 41974 45252 42114 45266
rect 42264 45252 43072 45266
rect 43222 45252 43362 45266
rect 43512 45252 44320 45266
rect 44470 45252 44610 45266
rect 44760 45252 45568 45266
rect 45718 45252 45858 45266
rect 46008 45252 46816 45266
rect 46966 45252 47106 45266
rect 47256 45252 48064 45266
rect 48214 45252 48354 45266
rect 48504 45252 49312 45266
rect 49462 45252 49602 45266
rect 49752 45252 50560 45266
rect 50710 45252 50850 45266
rect 51000 45252 51808 45266
rect 51958 45252 52098 45266
rect 52248 45252 53056 45266
rect 53206 45252 53346 45266
rect 53496 45252 54304 45266
rect 54454 45252 54594 45266
rect 54744 45252 55552 45266
rect 55702 45252 55842 45266
rect 55992 45252 56800 45266
rect 56950 45252 57090 45266
rect 57240 45252 58048 45266
rect 58198 45252 58338 45266
rect 58488 45252 58934 45266
rect 16898 45204 16980 45218
rect 17188 45204 17270 45218
rect 18146 45204 18228 45218
rect 18436 45204 18518 45218
rect 19394 45204 19476 45218
rect 19684 45204 19766 45218
rect 20642 45204 20724 45218
rect 20932 45204 21014 45218
rect 21890 45204 21972 45218
rect 22180 45204 22262 45218
rect 23138 45204 23220 45218
rect 23428 45204 23510 45218
rect 24386 45204 24468 45218
rect 24676 45204 24758 45218
rect 25634 45204 25716 45218
rect 25924 45204 26006 45218
rect 26882 45204 26964 45218
rect 27172 45204 27254 45218
rect 28130 45204 28212 45218
rect 28420 45204 28502 45218
rect 29378 45204 29460 45218
rect 29668 45204 29750 45218
rect 30626 45204 30708 45218
rect 30916 45204 30998 45218
rect 31874 45204 31956 45218
rect 32164 45204 32246 45218
rect 33122 45204 33204 45218
rect 33412 45204 33494 45218
rect 34370 45204 34452 45218
rect 34660 45204 34742 45218
rect 35618 45204 35700 45218
rect 35908 45204 35990 45218
rect 36866 45204 36948 45218
rect 37156 45204 37238 45218
rect 38114 45204 38196 45218
rect 38404 45204 38486 45218
rect 39362 45204 39444 45218
rect 39652 45204 39734 45218
rect 40610 45204 40692 45218
rect 40900 45204 40982 45218
rect 41858 45204 41940 45218
rect 42148 45204 42230 45218
rect 43106 45204 43188 45218
rect 43396 45204 43478 45218
rect 44354 45204 44436 45218
rect 44644 45204 44726 45218
rect 45602 45204 45684 45218
rect 45892 45204 45974 45218
rect 46850 45204 46932 45218
rect 47140 45204 47222 45218
rect 48098 45204 48180 45218
rect 48388 45204 48470 45218
rect 49346 45204 49428 45218
rect 49636 45204 49718 45218
rect 50594 45204 50676 45218
rect 50884 45204 50966 45218
rect 51842 45204 51924 45218
rect 52132 45204 52214 45218
rect 53090 45204 53172 45218
rect 53380 45204 53462 45218
rect 54338 45204 54420 45218
rect 54628 45204 54710 45218
rect 55586 45204 55668 45218
rect 55876 45204 55958 45218
rect 56834 45204 56916 45218
rect 57124 45204 57206 45218
rect 58082 45204 58164 45218
rect 58372 45204 58454 45218
rect 16418 45156 58934 45204
rect 16418 44998 58934 45108
rect 16418 44902 58934 44950
rect 16898 44888 16980 44902
rect 17188 44888 17270 44902
rect 18146 44888 18228 44902
rect 18436 44888 18518 44902
rect 19394 44888 19476 44902
rect 19684 44888 19766 44902
rect 20642 44888 20724 44902
rect 20932 44888 21014 44902
rect 21890 44888 21972 44902
rect 22180 44888 22262 44902
rect 23138 44888 23220 44902
rect 23428 44888 23510 44902
rect 24386 44888 24468 44902
rect 24676 44888 24758 44902
rect 25634 44888 25716 44902
rect 25924 44888 26006 44902
rect 26882 44888 26964 44902
rect 27172 44888 27254 44902
rect 28130 44888 28212 44902
rect 28420 44888 28502 44902
rect 29378 44888 29460 44902
rect 29668 44888 29750 44902
rect 30626 44888 30708 44902
rect 30916 44888 30998 44902
rect 31874 44888 31956 44902
rect 32164 44888 32246 44902
rect 33122 44888 33204 44902
rect 33412 44888 33494 44902
rect 34370 44888 34452 44902
rect 34660 44888 34742 44902
rect 35618 44888 35700 44902
rect 35908 44888 35990 44902
rect 36866 44888 36948 44902
rect 37156 44888 37238 44902
rect 38114 44888 38196 44902
rect 38404 44888 38486 44902
rect 39362 44888 39444 44902
rect 39652 44888 39734 44902
rect 40610 44888 40692 44902
rect 40900 44888 40982 44902
rect 41858 44888 41940 44902
rect 42148 44888 42230 44902
rect 43106 44888 43188 44902
rect 43396 44888 43478 44902
rect 44354 44888 44436 44902
rect 44644 44888 44726 44902
rect 45602 44888 45684 44902
rect 45892 44888 45974 44902
rect 46850 44888 46932 44902
rect 47140 44888 47222 44902
rect 48098 44888 48180 44902
rect 48388 44888 48470 44902
rect 49346 44888 49428 44902
rect 49636 44888 49718 44902
rect 50594 44888 50676 44902
rect 50884 44888 50966 44902
rect 51842 44888 51924 44902
rect 52132 44888 52214 44902
rect 53090 44888 53172 44902
rect 53380 44888 53462 44902
rect 54338 44888 54420 44902
rect 54628 44888 54710 44902
rect 55586 44888 55668 44902
rect 55876 44888 55958 44902
rect 56834 44888 56916 44902
rect 57124 44888 57206 44902
rect 58082 44888 58164 44902
rect 58372 44888 58454 44902
rect 16418 44840 16864 44854
rect 17014 44840 17154 44854
rect 17304 44840 18112 44854
rect 18262 44840 18402 44854
rect 18552 44840 19360 44854
rect 19510 44840 19650 44854
rect 19800 44840 20608 44854
rect 20758 44840 20898 44854
rect 21048 44840 21856 44854
rect 22006 44840 22146 44854
rect 22296 44840 23104 44854
rect 23254 44840 23394 44854
rect 23544 44840 24352 44854
rect 24502 44840 24642 44854
rect 24792 44840 25600 44854
rect 25750 44840 25890 44854
rect 26040 44840 26848 44854
rect 26998 44840 27138 44854
rect 27288 44840 28096 44854
rect 28246 44840 28386 44854
rect 28536 44840 29344 44854
rect 29494 44840 29634 44854
rect 29784 44840 30592 44854
rect 30742 44840 30882 44854
rect 31032 44840 31840 44854
rect 31990 44840 32130 44854
rect 32280 44840 33088 44854
rect 33238 44840 33378 44854
rect 33528 44840 34336 44854
rect 34486 44840 34626 44854
rect 34776 44840 35584 44854
rect 35734 44840 35874 44854
rect 36024 44840 36832 44854
rect 36982 44840 37122 44854
rect 37272 44840 38080 44854
rect 38230 44840 38370 44854
rect 38520 44840 39328 44854
rect 39478 44840 39618 44854
rect 39768 44840 40576 44854
rect 40726 44840 40866 44854
rect 41016 44840 41824 44854
rect 41974 44840 42114 44854
rect 42264 44840 43072 44854
rect 43222 44840 43362 44854
rect 43512 44840 44320 44854
rect 44470 44840 44610 44854
rect 44760 44840 45568 44854
rect 45718 44840 45858 44854
rect 46008 44840 46816 44854
rect 46966 44840 47106 44854
rect 47256 44840 48064 44854
rect 48214 44840 48354 44854
rect 48504 44840 49312 44854
rect 49462 44840 49602 44854
rect 49752 44840 50560 44854
rect 50710 44840 50850 44854
rect 51000 44840 51808 44854
rect 51958 44840 52098 44854
rect 52248 44840 53056 44854
rect 53206 44840 53346 44854
rect 53496 44840 54304 44854
rect 54454 44840 54594 44854
rect 54744 44840 55552 44854
rect 55702 44840 55842 44854
rect 55992 44840 56800 44854
rect 56950 44840 57090 44854
rect 57240 44840 58048 44854
rect 58198 44840 58338 44854
rect 58488 44840 58934 44854
rect 16418 44792 58934 44840
rect 16418 44778 16864 44792
rect 17014 44778 17154 44792
rect 17304 44778 18112 44792
rect 18262 44778 18402 44792
rect 18552 44778 19360 44792
rect 19510 44778 19650 44792
rect 19800 44778 20608 44792
rect 20758 44778 20898 44792
rect 21048 44778 21856 44792
rect 22006 44778 22146 44792
rect 22296 44778 23104 44792
rect 23254 44778 23394 44792
rect 23544 44778 24352 44792
rect 24502 44778 24642 44792
rect 24792 44778 25600 44792
rect 25750 44778 25890 44792
rect 26040 44778 26848 44792
rect 26998 44778 27138 44792
rect 27288 44778 28096 44792
rect 28246 44778 28386 44792
rect 28536 44778 29344 44792
rect 29494 44778 29634 44792
rect 29784 44778 30592 44792
rect 30742 44778 30882 44792
rect 31032 44778 31840 44792
rect 31990 44778 32130 44792
rect 32280 44778 33088 44792
rect 33238 44778 33378 44792
rect 33528 44778 34336 44792
rect 34486 44778 34626 44792
rect 34776 44778 35584 44792
rect 35734 44778 35874 44792
rect 36024 44778 36832 44792
rect 36982 44778 37122 44792
rect 37272 44778 38080 44792
rect 38230 44778 38370 44792
rect 38520 44778 39328 44792
rect 39478 44778 39618 44792
rect 39768 44778 40576 44792
rect 40726 44778 40866 44792
rect 41016 44778 41824 44792
rect 41974 44778 42114 44792
rect 42264 44778 43072 44792
rect 43222 44778 43362 44792
rect 43512 44778 44320 44792
rect 44470 44778 44610 44792
rect 44760 44778 45568 44792
rect 45718 44778 45858 44792
rect 46008 44778 46816 44792
rect 46966 44778 47106 44792
rect 47256 44778 48064 44792
rect 48214 44778 48354 44792
rect 48504 44778 49312 44792
rect 49462 44778 49602 44792
rect 49752 44778 50560 44792
rect 50710 44778 50850 44792
rect 51000 44778 51808 44792
rect 51958 44778 52098 44792
rect 52248 44778 53056 44792
rect 53206 44778 53346 44792
rect 53496 44778 54304 44792
rect 54454 44778 54594 44792
rect 54744 44778 55552 44792
rect 55702 44778 55842 44792
rect 55992 44778 56800 44792
rect 56950 44778 57090 44792
rect 57240 44778 58048 44792
rect 58198 44778 58338 44792
rect 58488 44778 58934 44792
rect 16898 44730 16980 44744
rect 17188 44730 17270 44744
rect 18146 44730 18228 44744
rect 18436 44730 18518 44744
rect 19394 44730 19476 44744
rect 19684 44730 19766 44744
rect 20642 44730 20724 44744
rect 20932 44730 21014 44744
rect 21890 44730 21972 44744
rect 22180 44730 22262 44744
rect 23138 44730 23220 44744
rect 23428 44730 23510 44744
rect 24386 44730 24468 44744
rect 24676 44730 24758 44744
rect 25634 44730 25716 44744
rect 25924 44730 26006 44744
rect 26882 44730 26964 44744
rect 27172 44730 27254 44744
rect 28130 44730 28212 44744
rect 28420 44730 28502 44744
rect 29378 44730 29460 44744
rect 29668 44730 29750 44744
rect 30626 44730 30708 44744
rect 30916 44730 30998 44744
rect 31874 44730 31956 44744
rect 32164 44730 32246 44744
rect 33122 44730 33204 44744
rect 33412 44730 33494 44744
rect 34370 44730 34452 44744
rect 34660 44730 34742 44744
rect 35618 44730 35700 44744
rect 35908 44730 35990 44744
rect 36866 44730 36948 44744
rect 37156 44730 37238 44744
rect 38114 44730 38196 44744
rect 38404 44730 38486 44744
rect 39362 44730 39444 44744
rect 39652 44730 39734 44744
rect 40610 44730 40692 44744
rect 40900 44730 40982 44744
rect 41858 44730 41940 44744
rect 42148 44730 42230 44744
rect 43106 44730 43188 44744
rect 43396 44730 43478 44744
rect 44354 44730 44436 44744
rect 44644 44730 44726 44744
rect 45602 44730 45684 44744
rect 45892 44730 45974 44744
rect 46850 44730 46932 44744
rect 47140 44730 47222 44744
rect 48098 44730 48180 44744
rect 48388 44730 48470 44744
rect 49346 44730 49428 44744
rect 49636 44730 49718 44744
rect 50594 44730 50676 44744
rect 50884 44730 50966 44744
rect 51842 44730 51924 44744
rect 52132 44730 52214 44744
rect 53090 44730 53172 44744
rect 53380 44730 53462 44744
rect 54338 44730 54420 44744
rect 54628 44730 54710 44744
rect 55586 44730 55668 44744
rect 55876 44730 55958 44744
rect 56834 44730 56916 44744
rect 57124 44730 57206 44744
rect 58082 44730 58164 44744
rect 58372 44730 58454 44744
rect 16418 44682 58934 44730
rect 16418 44586 58934 44634
rect 16898 44572 16980 44586
rect 17188 44572 17270 44586
rect 18146 44572 18228 44586
rect 18436 44572 18518 44586
rect 19394 44572 19476 44586
rect 19684 44572 19766 44586
rect 20642 44572 20724 44586
rect 20932 44572 21014 44586
rect 21890 44572 21972 44586
rect 22180 44572 22262 44586
rect 23138 44572 23220 44586
rect 23428 44572 23510 44586
rect 24386 44572 24468 44586
rect 24676 44572 24758 44586
rect 25634 44572 25716 44586
rect 25924 44572 26006 44586
rect 26882 44572 26964 44586
rect 27172 44572 27254 44586
rect 28130 44572 28212 44586
rect 28420 44572 28502 44586
rect 29378 44572 29460 44586
rect 29668 44572 29750 44586
rect 30626 44572 30708 44586
rect 30916 44572 30998 44586
rect 31874 44572 31956 44586
rect 32164 44572 32246 44586
rect 33122 44572 33204 44586
rect 33412 44572 33494 44586
rect 34370 44572 34452 44586
rect 34660 44572 34742 44586
rect 35618 44572 35700 44586
rect 35908 44572 35990 44586
rect 36866 44572 36948 44586
rect 37156 44572 37238 44586
rect 38114 44572 38196 44586
rect 38404 44572 38486 44586
rect 39362 44572 39444 44586
rect 39652 44572 39734 44586
rect 40610 44572 40692 44586
rect 40900 44572 40982 44586
rect 41858 44572 41940 44586
rect 42148 44572 42230 44586
rect 43106 44572 43188 44586
rect 43396 44572 43478 44586
rect 44354 44572 44436 44586
rect 44644 44572 44726 44586
rect 45602 44572 45684 44586
rect 45892 44572 45974 44586
rect 46850 44572 46932 44586
rect 47140 44572 47222 44586
rect 48098 44572 48180 44586
rect 48388 44572 48470 44586
rect 49346 44572 49428 44586
rect 49636 44572 49718 44586
rect 50594 44572 50676 44586
rect 50884 44572 50966 44586
rect 51842 44572 51924 44586
rect 52132 44572 52214 44586
rect 53090 44572 53172 44586
rect 53380 44572 53462 44586
rect 54338 44572 54420 44586
rect 54628 44572 54710 44586
rect 55586 44572 55668 44586
rect 55876 44572 55958 44586
rect 56834 44572 56916 44586
rect 57124 44572 57206 44586
rect 58082 44572 58164 44586
rect 58372 44572 58454 44586
rect 16418 44524 16864 44538
rect 17014 44524 17154 44538
rect 17304 44524 18112 44538
rect 18262 44524 18402 44538
rect 18552 44524 19360 44538
rect 19510 44524 19650 44538
rect 19800 44524 20608 44538
rect 20758 44524 20898 44538
rect 21048 44524 21856 44538
rect 22006 44524 22146 44538
rect 22296 44524 23104 44538
rect 23254 44524 23394 44538
rect 23544 44524 24352 44538
rect 24502 44524 24642 44538
rect 24792 44524 25600 44538
rect 25750 44524 25890 44538
rect 26040 44524 26848 44538
rect 26998 44524 27138 44538
rect 27288 44524 28096 44538
rect 28246 44524 28386 44538
rect 28536 44524 29344 44538
rect 29494 44524 29634 44538
rect 29784 44524 30592 44538
rect 30742 44524 30882 44538
rect 31032 44524 31840 44538
rect 31990 44524 32130 44538
rect 32280 44524 33088 44538
rect 33238 44524 33378 44538
rect 33528 44524 34336 44538
rect 34486 44524 34626 44538
rect 34776 44524 35584 44538
rect 35734 44524 35874 44538
rect 36024 44524 36832 44538
rect 36982 44524 37122 44538
rect 37272 44524 38080 44538
rect 38230 44524 38370 44538
rect 38520 44524 39328 44538
rect 39478 44524 39618 44538
rect 39768 44524 40576 44538
rect 40726 44524 40866 44538
rect 41016 44524 41824 44538
rect 41974 44524 42114 44538
rect 42264 44524 43072 44538
rect 43222 44524 43362 44538
rect 43512 44524 44320 44538
rect 44470 44524 44610 44538
rect 44760 44524 45568 44538
rect 45718 44524 45858 44538
rect 46008 44524 46816 44538
rect 46966 44524 47106 44538
rect 47256 44524 48064 44538
rect 48214 44524 48354 44538
rect 48504 44524 49312 44538
rect 49462 44524 49602 44538
rect 49752 44524 50560 44538
rect 50710 44524 50850 44538
rect 51000 44524 51808 44538
rect 51958 44524 52098 44538
rect 52248 44524 53056 44538
rect 53206 44524 53346 44538
rect 53496 44524 54304 44538
rect 54454 44524 54594 44538
rect 54744 44524 55552 44538
rect 55702 44524 55842 44538
rect 55992 44524 56800 44538
rect 56950 44524 57090 44538
rect 57240 44524 58048 44538
rect 58198 44524 58338 44538
rect 58488 44524 58934 44538
rect 16418 44476 58934 44524
rect 16418 44462 16864 44476
rect 17014 44462 17154 44476
rect 17304 44462 18112 44476
rect 18262 44462 18402 44476
rect 18552 44462 19360 44476
rect 19510 44462 19650 44476
rect 19800 44462 20608 44476
rect 20758 44462 20898 44476
rect 21048 44462 21856 44476
rect 22006 44462 22146 44476
rect 22296 44462 23104 44476
rect 23254 44462 23394 44476
rect 23544 44462 24352 44476
rect 24502 44462 24642 44476
rect 24792 44462 25600 44476
rect 25750 44462 25890 44476
rect 26040 44462 26848 44476
rect 26998 44462 27138 44476
rect 27288 44462 28096 44476
rect 28246 44462 28386 44476
rect 28536 44462 29344 44476
rect 29494 44462 29634 44476
rect 29784 44462 30592 44476
rect 30742 44462 30882 44476
rect 31032 44462 31840 44476
rect 31990 44462 32130 44476
rect 32280 44462 33088 44476
rect 33238 44462 33378 44476
rect 33528 44462 34336 44476
rect 34486 44462 34626 44476
rect 34776 44462 35584 44476
rect 35734 44462 35874 44476
rect 36024 44462 36832 44476
rect 36982 44462 37122 44476
rect 37272 44462 38080 44476
rect 38230 44462 38370 44476
rect 38520 44462 39328 44476
rect 39478 44462 39618 44476
rect 39768 44462 40576 44476
rect 40726 44462 40866 44476
rect 41016 44462 41824 44476
rect 41974 44462 42114 44476
rect 42264 44462 43072 44476
rect 43222 44462 43362 44476
rect 43512 44462 44320 44476
rect 44470 44462 44610 44476
rect 44760 44462 45568 44476
rect 45718 44462 45858 44476
rect 46008 44462 46816 44476
rect 46966 44462 47106 44476
rect 47256 44462 48064 44476
rect 48214 44462 48354 44476
rect 48504 44462 49312 44476
rect 49462 44462 49602 44476
rect 49752 44462 50560 44476
rect 50710 44462 50850 44476
rect 51000 44462 51808 44476
rect 51958 44462 52098 44476
rect 52248 44462 53056 44476
rect 53206 44462 53346 44476
rect 53496 44462 54304 44476
rect 54454 44462 54594 44476
rect 54744 44462 55552 44476
rect 55702 44462 55842 44476
rect 55992 44462 56800 44476
rect 56950 44462 57090 44476
rect 57240 44462 58048 44476
rect 58198 44462 58338 44476
rect 58488 44462 58934 44476
rect 16898 44414 16980 44428
rect 17188 44414 17270 44428
rect 18146 44414 18228 44428
rect 18436 44414 18518 44428
rect 19394 44414 19476 44428
rect 19684 44414 19766 44428
rect 20642 44414 20724 44428
rect 20932 44414 21014 44428
rect 21890 44414 21972 44428
rect 22180 44414 22262 44428
rect 23138 44414 23220 44428
rect 23428 44414 23510 44428
rect 24386 44414 24468 44428
rect 24676 44414 24758 44428
rect 25634 44414 25716 44428
rect 25924 44414 26006 44428
rect 26882 44414 26964 44428
rect 27172 44414 27254 44428
rect 28130 44414 28212 44428
rect 28420 44414 28502 44428
rect 29378 44414 29460 44428
rect 29668 44414 29750 44428
rect 30626 44414 30708 44428
rect 30916 44414 30998 44428
rect 31874 44414 31956 44428
rect 32164 44414 32246 44428
rect 33122 44414 33204 44428
rect 33412 44414 33494 44428
rect 34370 44414 34452 44428
rect 34660 44414 34742 44428
rect 35618 44414 35700 44428
rect 35908 44414 35990 44428
rect 36866 44414 36948 44428
rect 37156 44414 37238 44428
rect 38114 44414 38196 44428
rect 38404 44414 38486 44428
rect 39362 44414 39444 44428
rect 39652 44414 39734 44428
rect 40610 44414 40692 44428
rect 40900 44414 40982 44428
rect 41858 44414 41940 44428
rect 42148 44414 42230 44428
rect 43106 44414 43188 44428
rect 43396 44414 43478 44428
rect 44354 44414 44436 44428
rect 44644 44414 44726 44428
rect 45602 44414 45684 44428
rect 45892 44414 45974 44428
rect 46850 44414 46932 44428
rect 47140 44414 47222 44428
rect 48098 44414 48180 44428
rect 48388 44414 48470 44428
rect 49346 44414 49428 44428
rect 49636 44414 49718 44428
rect 50594 44414 50676 44428
rect 50884 44414 50966 44428
rect 51842 44414 51924 44428
rect 52132 44414 52214 44428
rect 53090 44414 53172 44428
rect 53380 44414 53462 44428
rect 54338 44414 54420 44428
rect 54628 44414 54710 44428
rect 55586 44414 55668 44428
rect 55876 44414 55958 44428
rect 56834 44414 56916 44428
rect 57124 44414 57206 44428
rect 58082 44414 58164 44428
rect 58372 44414 58454 44428
rect 16418 44366 58934 44414
rect 16418 44208 58934 44318
rect 16418 44112 58934 44160
rect 16898 44098 16980 44112
rect 17188 44098 17270 44112
rect 18146 44098 18228 44112
rect 18436 44098 18518 44112
rect 19394 44098 19476 44112
rect 19684 44098 19766 44112
rect 20642 44098 20724 44112
rect 20932 44098 21014 44112
rect 21890 44098 21972 44112
rect 22180 44098 22262 44112
rect 23138 44098 23220 44112
rect 23428 44098 23510 44112
rect 24386 44098 24468 44112
rect 24676 44098 24758 44112
rect 25634 44098 25716 44112
rect 25924 44098 26006 44112
rect 26882 44098 26964 44112
rect 27172 44098 27254 44112
rect 28130 44098 28212 44112
rect 28420 44098 28502 44112
rect 29378 44098 29460 44112
rect 29668 44098 29750 44112
rect 30626 44098 30708 44112
rect 30916 44098 30998 44112
rect 31874 44098 31956 44112
rect 32164 44098 32246 44112
rect 33122 44098 33204 44112
rect 33412 44098 33494 44112
rect 34370 44098 34452 44112
rect 34660 44098 34742 44112
rect 35618 44098 35700 44112
rect 35908 44098 35990 44112
rect 36866 44098 36948 44112
rect 37156 44098 37238 44112
rect 38114 44098 38196 44112
rect 38404 44098 38486 44112
rect 39362 44098 39444 44112
rect 39652 44098 39734 44112
rect 40610 44098 40692 44112
rect 40900 44098 40982 44112
rect 41858 44098 41940 44112
rect 42148 44098 42230 44112
rect 43106 44098 43188 44112
rect 43396 44098 43478 44112
rect 44354 44098 44436 44112
rect 44644 44098 44726 44112
rect 45602 44098 45684 44112
rect 45892 44098 45974 44112
rect 46850 44098 46932 44112
rect 47140 44098 47222 44112
rect 48098 44098 48180 44112
rect 48388 44098 48470 44112
rect 49346 44098 49428 44112
rect 49636 44098 49718 44112
rect 50594 44098 50676 44112
rect 50884 44098 50966 44112
rect 51842 44098 51924 44112
rect 52132 44098 52214 44112
rect 53090 44098 53172 44112
rect 53380 44098 53462 44112
rect 54338 44098 54420 44112
rect 54628 44098 54710 44112
rect 55586 44098 55668 44112
rect 55876 44098 55958 44112
rect 56834 44098 56916 44112
rect 57124 44098 57206 44112
rect 58082 44098 58164 44112
rect 58372 44098 58454 44112
rect 16418 44050 16864 44064
rect 17014 44050 17154 44064
rect 17304 44050 18112 44064
rect 18262 44050 18402 44064
rect 18552 44050 19360 44064
rect 19510 44050 19650 44064
rect 19800 44050 20608 44064
rect 20758 44050 20898 44064
rect 21048 44050 21856 44064
rect 22006 44050 22146 44064
rect 22296 44050 23104 44064
rect 23254 44050 23394 44064
rect 23544 44050 24352 44064
rect 24502 44050 24642 44064
rect 24792 44050 25600 44064
rect 25750 44050 25890 44064
rect 26040 44050 26848 44064
rect 26998 44050 27138 44064
rect 27288 44050 28096 44064
rect 28246 44050 28386 44064
rect 28536 44050 29344 44064
rect 29494 44050 29634 44064
rect 29784 44050 30592 44064
rect 30742 44050 30882 44064
rect 31032 44050 31840 44064
rect 31990 44050 32130 44064
rect 32280 44050 33088 44064
rect 33238 44050 33378 44064
rect 33528 44050 34336 44064
rect 34486 44050 34626 44064
rect 34776 44050 35584 44064
rect 35734 44050 35874 44064
rect 36024 44050 36832 44064
rect 36982 44050 37122 44064
rect 37272 44050 38080 44064
rect 38230 44050 38370 44064
rect 38520 44050 39328 44064
rect 39478 44050 39618 44064
rect 39768 44050 40576 44064
rect 40726 44050 40866 44064
rect 41016 44050 41824 44064
rect 41974 44050 42114 44064
rect 42264 44050 43072 44064
rect 43222 44050 43362 44064
rect 43512 44050 44320 44064
rect 44470 44050 44610 44064
rect 44760 44050 45568 44064
rect 45718 44050 45858 44064
rect 46008 44050 46816 44064
rect 46966 44050 47106 44064
rect 47256 44050 48064 44064
rect 48214 44050 48354 44064
rect 48504 44050 49312 44064
rect 49462 44050 49602 44064
rect 49752 44050 50560 44064
rect 50710 44050 50850 44064
rect 51000 44050 51808 44064
rect 51958 44050 52098 44064
rect 52248 44050 53056 44064
rect 53206 44050 53346 44064
rect 53496 44050 54304 44064
rect 54454 44050 54594 44064
rect 54744 44050 55552 44064
rect 55702 44050 55842 44064
rect 55992 44050 56800 44064
rect 56950 44050 57090 44064
rect 57240 44050 58048 44064
rect 58198 44050 58338 44064
rect 58488 44050 58934 44064
rect 16418 44002 58934 44050
rect 16418 43988 16864 44002
rect 17014 43988 17154 44002
rect 17304 43988 18112 44002
rect 18262 43988 18402 44002
rect 18552 43988 19360 44002
rect 19510 43988 19650 44002
rect 19800 43988 20608 44002
rect 20758 43988 20898 44002
rect 21048 43988 21856 44002
rect 22006 43988 22146 44002
rect 22296 43988 23104 44002
rect 23254 43988 23394 44002
rect 23544 43988 24352 44002
rect 24502 43988 24642 44002
rect 24792 43988 25600 44002
rect 25750 43988 25890 44002
rect 26040 43988 26848 44002
rect 26998 43988 27138 44002
rect 27288 43988 28096 44002
rect 28246 43988 28386 44002
rect 28536 43988 29344 44002
rect 29494 43988 29634 44002
rect 29784 43988 30592 44002
rect 30742 43988 30882 44002
rect 31032 43988 31840 44002
rect 31990 43988 32130 44002
rect 32280 43988 33088 44002
rect 33238 43988 33378 44002
rect 33528 43988 34336 44002
rect 34486 43988 34626 44002
rect 34776 43988 35584 44002
rect 35734 43988 35874 44002
rect 36024 43988 36832 44002
rect 36982 43988 37122 44002
rect 37272 43988 38080 44002
rect 38230 43988 38370 44002
rect 38520 43988 39328 44002
rect 39478 43988 39618 44002
rect 39768 43988 40576 44002
rect 40726 43988 40866 44002
rect 41016 43988 41824 44002
rect 41974 43988 42114 44002
rect 42264 43988 43072 44002
rect 43222 43988 43362 44002
rect 43512 43988 44320 44002
rect 44470 43988 44610 44002
rect 44760 43988 45568 44002
rect 45718 43988 45858 44002
rect 46008 43988 46816 44002
rect 46966 43988 47106 44002
rect 47256 43988 48064 44002
rect 48214 43988 48354 44002
rect 48504 43988 49312 44002
rect 49462 43988 49602 44002
rect 49752 43988 50560 44002
rect 50710 43988 50850 44002
rect 51000 43988 51808 44002
rect 51958 43988 52098 44002
rect 52248 43988 53056 44002
rect 53206 43988 53346 44002
rect 53496 43988 54304 44002
rect 54454 43988 54594 44002
rect 54744 43988 55552 44002
rect 55702 43988 55842 44002
rect 55992 43988 56800 44002
rect 56950 43988 57090 44002
rect 57240 43988 58048 44002
rect 58198 43988 58338 44002
rect 58488 43988 58934 44002
rect 16898 43940 16980 43954
rect 17188 43940 17270 43954
rect 18146 43940 18228 43954
rect 18436 43940 18518 43954
rect 19394 43940 19476 43954
rect 19684 43940 19766 43954
rect 20642 43940 20724 43954
rect 20932 43940 21014 43954
rect 21890 43940 21972 43954
rect 22180 43940 22262 43954
rect 23138 43940 23220 43954
rect 23428 43940 23510 43954
rect 24386 43940 24468 43954
rect 24676 43940 24758 43954
rect 25634 43940 25716 43954
rect 25924 43940 26006 43954
rect 26882 43940 26964 43954
rect 27172 43940 27254 43954
rect 28130 43940 28212 43954
rect 28420 43940 28502 43954
rect 29378 43940 29460 43954
rect 29668 43940 29750 43954
rect 30626 43940 30708 43954
rect 30916 43940 30998 43954
rect 31874 43940 31956 43954
rect 32164 43940 32246 43954
rect 33122 43940 33204 43954
rect 33412 43940 33494 43954
rect 34370 43940 34452 43954
rect 34660 43940 34742 43954
rect 35618 43940 35700 43954
rect 35908 43940 35990 43954
rect 36866 43940 36948 43954
rect 37156 43940 37238 43954
rect 38114 43940 38196 43954
rect 38404 43940 38486 43954
rect 39362 43940 39444 43954
rect 39652 43940 39734 43954
rect 40610 43940 40692 43954
rect 40900 43940 40982 43954
rect 41858 43940 41940 43954
rect 42148 43940 42230 43954
rect 43106 43940 43188 43954
rect 43396 43940 43478 43954
rect 44354 43940 44436 43954
rect 44644 43940 44726 43954
rect 45602 43940 45684 43954
rect 45892 43940 45974 43954
rect 46850 43940 46932 43954
rect 47140 43940 47222 43954
rect 48098 43940 48180 43954
rect 48388 43940 48470 43954
rect 49346 43940 49428 43954
rect 49636 43940 49718 43954
rect 50594 43940 50676 43954
rect 50884 43940 50966 43954
rect 51842 43940 51924 43954
rect 52132 43940 52214 43954
rect 53090 43940 53172 43954
rect 53380 43940 53462 43954
rect 54338 43940 54420 43954
rect 54628 43940 54710 43954
rect 55586 43940 55668 43954
rect 55876 43940 55958 43954
rect 56834 43940 56916 43954
rect 57124 43940 57206 43954
rect 58082 43940 58164 43954
rect 58372 43940 58454 43954
rect 16418 43892 58934 43940
rect 16418 43796 58934 43844
rect 16898 43782 16980 43796
rect 17188 43782 17270 43796
rect 18146 43782 18228 43796
rect 18436 43782 18518 43796
rect 19394 43782 19476 43796
rect 19684 43782 19766 43796
rect 20642 43782 20724 43796
rect 20932 43782 21014 43796
rect 21890 43782 21972 43796
rect 22180 43782 22262 43796
rect 23138 43782 23220 43796
rect 23428 43782 23510 43796
rect 24386 43782 24468 43796
rect 24676 43782 24758 43796
rect 25634 43782 25716 43796
rect 25924 43782 26006 43796
rect 26882 43782 26964 43796
rect 27172 43782 27254 43796
rect 28130 43782 28212 43796
rect 28420 43782 28502 43796
rect 29378 43782 29460 43796
rect 29668 43782 29750 43796
rect 30626 43782 30708 43796
rect 30916 43782 30998 43796
rect 31874 43782 31956 43796
rect 32164 43782 32246 43796
rect 33122 43782 33204 43796
rect 33412 43782 33494 43796
rect 34370 43782 34452 43796
rect 34660 43782 34742 43796
rect 35618 43782 35700 43796
rect 35908 43782 35990 43796
rect 36866 43782 36948 43796
rect 37156 43782 37238 43796
rect 38114 43782 38196 43796
rect 38404 43782 38486 43796
rect 39362 43782 39444 43796
rect 39652 43782 39734 43796
rect 40610 43782 40692 43796
rect 40900 43782 40982 43796
rect 41858 43782 41940 43796
rect 42148 43782 42230 43796
rect 43106 43782 43188 43796
rect 43396 43782 43478 43796
rect 44354 43782 44436 43796
rect 44644 43782 44726 43796
rect 45602 43782 45684 43796
rect 45892 43782 45974 43796
rect 46850 43782 46932 43796
rect 47140 43782 47222 43796
rect 48098 43782 48180 43796
rect 48388 43782 48470 43796
rect 49346 43782 49428 43796
rect 49636 43782 49718 43796
rect 50594 43782 50676 43796
rect 50884 43782 50966 43796
rect 51842 43782 51924 43796
rect 52132 43782 52214 43796
rect 53090 43782 53172 43796
rect 53380 43782 53462 43796
rect 54338 43782 54420 43796
rect 54628 43782 54710 43796
rect 55586 43782 55668 43796
rect 55876 43782 55958 43796
rect 56834 43782 56916 43796
rect 57124 43782 57206 43796
rect 58082 43782 58164 43796
rect 58372 43782 58454 43796
rect 16418 43734 16864 43748
rect 17014 43734 17154 43748
rect 17304 43734 18112 43748
rect 18262 43734 18402 43748
rect 18552 43734 19360 43748
rect 19510 43734 19650 43748
rect 19800 43734 20608 43748
rect 20758 43734 20898 43748
rect 21048 43734 21856 43748
rect 22006 43734 22146 43748
rect 22296 43734 23104 43748
rect 23254 43734 23394 43748
rect 23544 43734 24352 43748
rect 24502 43734 24642 43748
rect 24792 43734 25600 43748
rect 25750 43734 25890 43748
rect 26040 43734 26848 43748
rect 26998 43734 27138 43748
rect 27288 43734 28096 43748
rect 28246 43734 28386 43748
rect 28536 43734 29344 43748
rect 29494 43734 29634 43748
rect 29784 43734 30592 43748
rect 30742 43734 30882 43748
rect 31032 43734 31840 43748
rect 31990 43734 32130 43748
rect 32280 43734 33088 43748
rect 33238 43734 33378 43748
rect 33528 43734 34336 43748
rect 34486 43734 34626 43748
rect 34776 43734 35584 43748
rect 35734 43734 35874 43748
rect 36024 43734 36832 43748
rect 36982 43734 37122 43748
rect 37272 43734 38080 43748
rect 38230 43734 38370 43748
rect 38520 43734 39328 43748
rect 39478 43734 39618 43748
rect 39768 43734 40576 43748
rect 40726 43734 40866 43748
rect 41016 43734 41824 43748
rect 41974 43734 42114 43748
rect 42264 43734 43072 43748
rect 43222 43734 43362 43748
rect 43512 43734 44320 43748
rect 44470 43734 44610 43748
rect 44760 43734 45568 43748
rect 45718 43734 45858 43748
rect 46008 43734 46816 43748
rect 46966 43734 47106 43748
rect 47256 43734 48064 43748
rect 48214 43734 48354 43748
rect 48504 43734 49312 43748
rect 49462 43734 49602 43748
rect 49752 43734 50560 43748
rect 50710 43734 50850 43748
rect 51000 43734 51808 43748
rect 51958 43734 52098 43748
rect 52248 43734 53056 43748
rect 53206 43734 53346 43748
rect 53496 43734 54304 43748
rect 54454 43734 54594 43748
rect 54744 43734 55552 43748
rect 55702 43734 55842 43748
rect 55992 43734 56800 43748
rect 56950 43734 57090 43748
rect 57240 43734 58048 43748
rect 58198 43734 58338 43748
rect 58488 43734 58934 43748
rect 16418 43686 58934 43734
rect 16418 43672 16864 43686
rect 17014 43672 17154 43686
rect 17304 43672 18112 43686
rect 18262 43672 18402 43686
rect 18552 43672 19360 43686
rect 19510 43672 19650 43686
rect 19800 43672 20608 43686
rect 20758 43672 20898 43686
rect 21048 43672 21856 43686
rect 22006 43672 22146 43686
rect 22296 43672 23104 43686
rect 23254 43672 23394 43686
rect 23544 43672 24352 43686
rect 24502 43672 24642 43686
rect 24792 43672 25600 43686
rect 25750 43672 25890 43686
rect 26040 43672 26848 43686
rect 26998 43672 27138 43686
rect 27288 43672 28096 43686
rect 28246 43672 28386 43686
rect 28536 43672 29344 43686
rect 29494 43672 29634 43686
rect 29784 43672 30592 43686
rect 30742 43672 30882 43686
rect 31032 43672 31840 43686
rect 31990 43672 32130 43686
rect 32280 43672 33088 43686
rect 33238 43672 33378 43686
rect 33528 43672 34336 43686
rect 34486 43672 34626 43686
rect 34776 43672 35584 43686
rect 35734 43672 35874 43686
rect 36024 43672 36832 43686
rect 36982 43672 37122 43686
rect 37272 43672 38080 43686
rect 38230 43672 38370 43686
rect 38520 43672 39328 43686
rect 39478 43672 39618 43686
rect 39768 43672 40576 43686
rect 40726 43672 40866 43686
rect 41016 43672 41824 43686
rect 41974 43672 42114 43686
rect 42264 43672 43072 43686
rect 43222 43672 43362 43686
rect 43512 43672 44320 43686
rect 44470 43672 44610 43686
rect 44760 43672 45568 43686
rect 45718 43672 45858 43686
rect 46008 43672 46816 43686
rect 46966 43672 47106 43686
rect 47256 43672 48064 43686
rect 48214 43672 48354 43686
rect 48504 43672 49312 43686
rect 49462 43672 49602 43686
rect 49752 43672 50560 43686
rect 50710 43672 50850 43686
rect 51000 43672 51808 43686
rect 51958 43672 52098 43686
rect 52248 43672 53056 43686
rect 53206 43672 53346 43686
rect 53496 43672 54304 43686
rect 54454 43672 54594 43686
rect 54744 43672 55552 43686
rect 55702 43672 55842 43686
rect 55992 43672 56800 43686
rect 56950 43672 57090 43686
rect 57240 43672 58048 43686
rect 58198 43672 58338 43686
rect 58488 43672 58934 43686
rect 16898 43624 16980 43638
rect 17188 43624 17270 43638
rect 18146 43624 18228 43638
rect 18436 43624 18518 43638
rect 19394 43624 19476 43638
rect 19684 43624 19766 43638
rect 20642 43624 20724 43638
rect 20932 43624 21014 43638
rect 21890 43624 21972 43638
rect 22180 43624 22262 43638
rect 23138 43624 23220 43638
rect 23428 43624 23510 43638
rect 24386 43624 24468 43638
rect 24676 43624 24758 43638
rect 25634 43624 25716 43638
rect 25924 43624 26006 43638
rect 26882 43624 26964 43638
rect 27172 43624 27254 43638
rect 28130 43624 28212 43638
rect 28420 43624 28502 43638
rect 29378 43624 29460 43638
rect 29668 43624 29750 43638
rect 30626 43624 30708 43638
rect 30916 43624 30998 43638
rect 31874 43624 31956 43638
rect 32164 43624 32246 43638
rect 33122 43624 33204 43638
rect 33412 43624 33494 43638
rect 34370 43624 34452 43638
rect 34660 43624 34742 43638
rect 35618 43624 35700 43638
rect 35908 43624 35990 43638
rect 36866 43624 36948 43638
rect 37156 43624 37238 43638
rect 38114 43624 38196 43638
rect 38404 43624 38486 43638
rect 39362 43624 39444 43638
rect 39652 43624 39734 43638
rect 40610 43624 40692 43638
rect 40900 43624 40982 43638
rect 41858 43624 41940 43638
rect 42148 43624 42230 43638
rect 43106 43624 43188 43638
rect 43396 43624 43478 43638
rect 44354 43624 44436 43638
rect 44644 43624 44726 43638
rect 45602 43624 45684 43638
rect 45892 43624 45974 43638
rect 46850 43624 46932 43638
rect 47140 43624 47222 43638
rect 48098 43624 48180 43638
rect 48388 43624 48470 43638
rect 49346 43624 49428 43638
rect 49636 43624 49718 43638
rect 50594 43624 50676 43638
rect 50884 43624 50966 43638
rect 51842 43624 51924 43638
rect 52132 43624 52214 43638
rect 53090 43624 53172 43638
rect 53380 43624 53462 43638
rect 54338 43624 54420 43638
rect 54628 43624 54710 43638
rect 55586 43624 55668 43638
rect 55876 43624 55958 43638
rect 56834 43624 56916 43638
rect 57124 43624 57206 43638
rect 58082 43624 58164 43638
rect 58372 43624 58454 43638
rect 16418 43576 58934 43624
rect 16418 43418 58934 43528
rect 16418 43322 58934 43370
rect 16898 43308 16980 43322
rect 17188 43308 17270 43322
rect 18146 43308 18228 43322
rect 18436 43308 18518 43322
rect 19394 43308 19476 43322
rect 19684 43308 19766 43322
rect 20642 43308 20724 43322
rect 20932 43308 21014 43322
rect 21890 43308 21972 43322
rect 22180 43308 22262 43322
rect 23138 43308 23220 43322
rect 23428 43308 23510 43322
rect 24386 43308 24468 43322
rect 24676 43308 24758 43322
rect 25634 43308 25716 43322
rect 25924 43308 26006 43322
rect 26882 43308 26964 43322
rect 27172 43308 27254 43322
rect 28130 43308 28212 43322
rect 28420 43308 28502 43322
rect 29378 43308 29460 43322
rect 29668 43308 29750 43322
rect 30626 43308 30708 43322
rect 30916 43308 30998 43322
rect 31874 43308 31956 43322
rect 32164 43308 32246 43322
rect 33122 43308 33204 43322
rect 33412 43308 33494 43322
rect 34370 43308 34452 43322
rect 34660 43308 34742 43322
rect 35618 43308 35700 43322
rect 35908 43308 35990 43322
rect 36866 43308 36948 43322
rect 37156 43308 37238 43322
rect 38114 43308 38196 43322
rect 38404 43308 38486 43322
rect 39362 43308 39444 43322
rect 39652 43308 39734 43322
rect 40610 43308 40692 43322
rect 40900 43308 40982 43322
rect 41858 43308 41940 43322
rect 42148 43308 42230 43322
rect 43106 43308 43188 43322
rect 43396 43308 43478 43322
rect 44354 43308 44436 43322
rect 44644 43308 44726 43322
rect 45602 43308 45684 43322
rect 45892 43308 45974 43322
rect 46850 43308 46932 43322
rect 47140 43308 47222 43322
rect 48098 43308 48180 43322
rect 48388 43308 48470 43322
rect 49346 43308 49428 43322
rect 49636 43308 49718 43322
rect 50594 43308 50676 43322
rect 50884 43308 50966 43322
rect 51842 43308 51924 43322
rect 52132 43308 52214 43322
rect 53090 43308 53172 43322
rect 53380 43308 53462 43322
rect 54338 43308 54420 43322
rect 54628 43308 54710 43322
rect 55586 43308 55668 43322
rect 55876 43308 55958 43322
rect 56834 43308 56916 43322
rect 57124 43308 57206 43322
rect 58082 43308 58164 43322
rect 58372 43308 58454 43322
rect 16418 43260 16864 43274
rect 17014 43260 17154 43274
rect 17304 43260 18112 43274
rect 18262 43260 18402 43274
rect 18552 43260 19360 43274
rect 19510 43260 19650 43274
rect 19800 43260 20608 43274
rect 20758 43260 20898 43274
rect 21048 43260 21856 43274
rect 22006 43260 22146 43274
rect 22296 43260 23104 43274
rect 23254 43260 23394 43274
rect 23544 43260 24352 43274
rect 24502 43260 24642 43274
rect 24792 43260 25600 43274
rect 25750 43260 25890 43274
rect 26040 43260 26848 43274
rect 26998 43260 27138 43274
rect 27288 43260 28096 43274
rect 28246 43260 28386 43274
rect 28536 43260 29344 43274
rect 29494 43260 29634 43274
rect 29784 43260 30592 43274
rect 30742 43260 30882 43274
rect 31032 43260 31840 43274
rect 31990 43260 32130 43274
rect 32280 43260 33088 43274
rect 33238 43260 33378 43274
rect 33528 43260 34336 43274
rect 34486 43260 34626 43274
rect 34776 43260 35584 43274
rect 35734 43260 35874 43274
rect 36024 43260 36832 43274
rect 36982 43260 37122 43274
rect 37272 43260 38080 43274
rect 38230 43260 38370 43274
rect 38520 43260 39328 43274
rect 39478 43260 39618 43274
rect 39768 43260 40576 43274
rect 40726 43260 40866 43274
rect 41016 43260 41824 43274
rect 41974 43260 42114 43274
rect 42264 43260 43072 43274
rect 43222 43260 43362 43274
rect 43512 43260 44320 43274
rect 44470 43260 44610 43274
rect 44760 43260 45568 43274
rect 45718 43260 45858 43274
rect 46008 43260 46816 43274
rect 46966 43260 47106 43274
rect 47256 43260 48064 43274
rect 48214 43260 48354 43274
rect 48504 43260 49312 43274
rect 49462 43260 49602 43274
rect 49752 43260 50560 43274
rect 50710 43260 50850 43274
rect 51000 43260 51808 43274
rect 51958 43260 52098 43274
rect 52248 43260 53056 43274
rect 53206 43260 53346 43274
rect 53496 43260 54304 43274
rect 54454 43260 54594 43274
rect 54744 43260 55552 43274
rect 55702 43260 55842 43274
rect 55992 43260 56800 43274
rect 56950 43260 57090 43274
rect 57240 43260 58048 43274
rect 58198 43260 58338 43274
rect 58488 43260 58934 43274
rect 16418 43212 58934 43260
rect 16418 43198 16864 43212
rect 17014 43198 17154 43212
rect 17304 43198 18112 43212
rect 18262 43198 18402 43212
rect 18552 43198 19360 43212
rect 19510 43198 19650 43212
rect 19800 43198 20608 43212
rect 20758 43198 20898 43212
rect 21048 43198 21856 43212
rect 22006 43198 22146 43212
rect 22296 43198 23104 43212
rect 23254 43198 23394 43212
rect 23544 43198 24352 43212
rect 24502 43198 24642 43212
rect 24792 43198 25600 43212
rect 25750 43198 25890 43212
rect 26040 43198 26848 43212
rect 26998 43198 27138 43212
rect 27288 43198 28096 43212
rect 28246 43198 28386 43212
rect 28536 43198 29344 43212
rect 29494 43198 29634 43212
rect 29784 43198 30592 43212
rect 30742 43198 30882 43212
rect 31032 43198 31840 43212
rect 31990 43198 32130 43212
rect 32280 43198 33088 43212
rect 33238 43198 33378 43212
rect 33528 43198 34336 43212
rect 34486 43198 34626 43212
rect 34776 43198 35584 43212
rect 35734 43198 35874 43212
rect 36024 43198 36832 43212
rect 36982 43198 37122 43212
rect 37272 43198 38080 43212
rect 38230 43198 38370 43212
rect 38520 43198 39328 43212
rect 39478 43198 39618 43212
rect 39768 43198 40576 43212
rect 40726 43198 40866 43212
rect 41016 43198 41824 43212
rect 41974 43198 42114 43212
rect 42264 43198 43072 43212
rect 43222 43198 43362 43212
rect 43512 43198 44320 43212
rect 44470 43198 44610 43212
rect 44760 43198 45568 43212
rect 45718 43198 45858 43212
rect 46008 43198 46816 43212
rect 46966 43198 47106 43212
rect 47256 43198 48064 43212
rect 48214 43198 48354 43212
rect 48504 43198 49312 43212
rect 49462 43198 49602 43212
rect 49752 43198 50560 43212
rect 50710 43198 50850 43212
rect 51000 43198 51808 43212
rect 51958 43198 52098 43212
rect 52248 43198 53056 43212
rect 53206 43198 53346 43212
rect 53496 43198 54304 43212
rect 54454 43198 54594 43212
rect 54744 43198 55552 43212
rect 55702 43198 55842 43212
rect 55992 43198 56800 43212
rect 56950 43198 57090 43212
rect 57240 43198 58048 43212
rect 58198 43198 58338 43212
rect 58488 43198 58934 43212
rect 16898 43150 16980 43164
rect 17188 43150 17270 43164
rect 18146 43150 18228 43164
rect 18436 43150 18518 43164
rect 19394 43150 19476 43164
rect 19684 43150 19766 43164
rect 20642 43150 20724 43164
rect 20932 43150 21014 43164
rect 21890 43150 21972 43164
rect 22180 43150 22262 43164
rect 23138 43150 23220 43164
rect 23428 43150 23510 43164
rect 24386 43150 24468 43164
rect 24676 43150 24758 43164
rect 25634 43150 25716 43164
rect 25924 43150 26006 43164
rect 26882 43150 26964 43164
rect 27172 43150 27254 43164
rect 28130 43150 28212 43164
rect 28420 43150 28502 43164
rect 29378 43150 29460 43164
rect 29668 43150 29750 43164
rect 30626 43150 30708 43164
rect 30916 43150 30998 43164
rect 31874 43150 31956 43164
rect 32164 43150 32246 43164
rect 33122 43150 33204 43164
rect 33412 43150 33494 43164
rect 34370 43150 34452 43164
rect 34660 43150 34742 43164
rect 35618 43150 35700 43164
rect 35908 43150 35990 43164
rect 36866 43150 36948 43164
rect 37156 43150 37238 43164
rect 38114 43150 38196 43164
rect 38404 43150 38486 43164
rect 39362 43150 39444 43164
rect 39652 43150 39734 43164
rect 40610 43150 40692 43164
rect 40900 43150 40982 43164
rect 41858 43150 41940 43164
rect 42148 43150 42230 43164
rect 43106 43150 43188 43164
rect 43396 43150 43478 43164
rect 44354 43150 44436 43164
rect 44644 43150 44726 43164
rect 45602 43150 45684 43164
rect 45892 43150 45974 43164
rect 46850 43150 46932 43164
rect 47140 43150 47222 43164
rect 48098 43150 48180 43164
rect 48388 43150 48470 43164
rect 49346 43150 49428 43164
rect 49636 43150 49718 43164
rect 50594 43150 50676 43164
rect 50884 43150 50966 43164
rect 51842 43150 51924 43164
rect 52132 43150 52214 43164
rect 53090 43150 53172 43164
rect 53380 43150 53462 43164
rect 54338 43150 54420 43164
rect 54628 43150 54710 43164
rect 55586 43150 55668 43164
rect 55876 43150 55958 43164
rect 56834 43150 56916 43164
rect 57124 43150 57206 43164
rect 58082 43150 58164 43164
rect 58372 43150 58454 43164
rect 16418 43102 58934 43150
rect 16418 43006 58934 43054
rect 16898 42992 16980 43006
rect 17188 42992 17270 43006
rect 18146 42992 18228 43006
rect 18436 42992 18518 43006
rect 19394 42992 19476 43006
rect 19684 42992 19766 43006
rect 20642 42992 20724 43006
rect 20932 42992 21014 43006
rect 21890 42992 21972 43006
rect 22180 42992 22262 43006
rect 23138 42992 23220 43006
rect 23428 42992 23510 43006
rect 24386 42992 24468 43006
rect 24676 42992 24758 43006
rect 25634 42992 25716 43006
rect 25924 42992 26006 43006
rect 26882 42992 26964 43006
rect 27172 42992 27254 43006
rect 28130 42992 28212 43006
rect 28420 42992 28502 43006
rect 29378 42992 29460 43006
rect 29668 42992 29750 43006
rect 30626 42992 30708 43006
rect 30916 42992 30998 43006
rect 31874 42992 31956 43006
rect 32164 42992 32246 43006
rect 33122 42992 33204 43006
rect 33412 42992 33494 43006
rect 34370 42992 34452 43006
rect 34660 42992 34742 43006
rect 35618 42992 35700 43006
rect 35908 42992 35990 43006
rect 36866 42992 36948 43006
rect 37156 42992 37238 43006
rect 38114 42992 38196 43006
rect 38404 42992 38486 43006
rect 39362 42992 39444 43006
rect 39652 42992 39734 43006
rect 40610 42992 40692 43006
rect 40900 42992 40982 43006
rect 41858 42992 41940 43006
rect 42148 42992 42230 43006
rect 43106 42992 43188 43006
rect 43396 42992 43478 43006
rect 44354 42992 44436 43006
rect 44644 42992 44726 43006
rect 45602 42992 45684 43006
rect 45892 42992 45974 43006
rect 46850 42992 46932 43006
rect 47140 42992 47222 43006
rect 48098 42992 48180 43006
rect 48388 42992 48470 43006
rect 49346 42992 49428 43006
rect 49636 42992 49718 43006
rect 50594 42992 50676 43006
rect 50884 42992 50966 43006
rect 51842 42992 51924 43006
rect 52132 42992 52214 43006
rect 53090 42992 53172 43006
rect 53380 42992 53462 43006
rect 54338 42992 54420 43006
rect 54628 42992 54710 43006
rect 55586 42992 55668 43006
rect 55876 42992 55958 43006
rect 56834 42992 56916 43006
rect 57124 42992 57206 43006
rect 58082 42992 58164 43006
rect 58372 42992 58454 43006
rect 16418 42944 16864 42958
rect 17014 42944 17154 42958
rect 17304 42944 18112 42958
rect 18262 42944 18402 42958
rect 18552 42944 19360 42958
rect 19510 42944 19650 42958
rect 19800 42944 20608 42958
rect 20758 42944 20898 42958
rect 21048 42944 21856 42958
rect 22006 42944 22146 42958
rect 22296 42944 23104 42958
rect 23254 42944 23394 42958
rect 23544 42944 24352 42958
rect 24502 42944 24642 42958
rect 24792 42944 25600 42958
rect 25750 42944 25890 42958
rect 26040 42944 26848 42958
rect 26998 42944 27138 42958
rect 27288 42944 28096 42958
rect 28246 42944 28386 42958
rect 28536 42944 29344 42958
rect 29494 42944 29634 42958
rect 29784 42944 30592 42958
rect 30742 42944 30882 42958
rect 31032 42944 31840 42958
rect 31990 42944 32130 42958
rect 32280 42944 33088 42958
rect 33238 42944 33378 42958
rect 33528 42944 34336 42958
rect 34486 42944 34626 42958
rect 34776 42944 35584 42958
rect 35734 42944 35874 42958
rect 36024 42944 36832 42958
rect 36982 42944 37122 42958
rect 37272 42944 38080 42958
rect 38230 42944 38370 42958
rect 38520 42944 39328 42958
rect 39478 42944 39618 42958
rect 39768 42944 40576 42958
rect 40726 42944 40866 42958
rect 41016 42944 41824 42958
rect 41974 42944 42114 42958
rect 42264 42944 43072 42958
rect 43222 42944 43362 42958
rect 43512 42944 44320 42958
rect 44470 42944 44610 42958
rect 44760 42944 45568 42958
rect 45718 42944 45858 42958
rect 46008 42944 46816 42958
rect 46966 42944 47106 42958
rect 47256 42944 48064 42958
rect 48214 42944 48354 42958
rect 48504 42944 49312 42958
rect 49462 42944 49602 42958
rect 49752 42944 50560 42958
rect 50710 42944 50850 42958
rect 51000 42944 51808 42958
rect 51958 42944 52098 42958
rect 52248 42944 53056 42958
rect 53206 42944 53346 42958
rect 53496 42944 54304 42958
rect 54454 42944 54594 42958
rect 54744 42944 55552 42958
rect 55702 42944 55842 42958
rect 55992 42944 56800 42958
rect 56950 42944 57090 42958
rect 57240 42944 58048 42958
rect 58198 42944 58338 42958
rect 58488 42944 58934 42958
rect 16418 42896 58934 42944
rect 16418 42882 16864 42896
rect 17014 42882 17154 42896
rect 17304 42882 18112 42896
rect 18262 42882 18402 42896
rect 18552 42882 19360 42896
rect 19510 42882 19650 42896
rect 19800 42882 20608 42896
rect 20758 42882 20898 42896
rect 21048 42882 21856 42896
rect 22006 42882 22146 42896
rect 22296 42882 23104 42896
rect 23254 42882 23394 42896
rect 23544 42882 24352 42896
rect 24502 42882 24642 42896
rect 24792 42882 25600 42896
rect 25750 42882 25890 42896
rect 26040 42882 26848 42896
rect 26998 42882 27138 42896
rect 27288 42882 28096 42896
rect 28246 42882 28386 42896
rect 28536 42882 29344 42896
rect 29494 42882 29634 42896
rect 29784 42882 30592 42896
rect 30742 42882 30882 42896
rect 31032 42882 31840 42896
rect 31990 42882 32130 42896
rect 32280 42882 33088 42896
rect 33238 42882 33378 42896
rect 33528 42882 34336 42896
rect 34486 42882 34626 42896
rect 34776 42882 35584 42896
rect 35734 42882 35874 42896
rect 36024 42882 36832 42896
rect 36982 42882 37122 42896
rect 37272 42882 38080 42896
rect 38230 42882 38370 42896
rect 38520 42882 39328 42896
rect 39478 42882 39618 42896
rect 39768 42882 40576 42896
rect 40726 42882 40866 42896
rect 41016 42882 41824 42896
rect 41974 42882 42114 42896
rect 42264 42882 43072 42896
rect 43222 42882 43362 42896
rect 43512 42882 44320 42896
rect 44470 42882 44610 42896
rect 44760 42882 45568 42896
rect 45718 42882 45858 42896
rect 46008 42882 46816 42896
rect 46966 42882 47106 42896
rect 47256 42882 48064 42896
rect 48214 42882 48354 42896
rect 48504 42882 49312 42896
rect 49462 42882 49602 42896
rect 49752 42882 50560 42896
rect 50710 42882 50850 42896
rect 51000 42882 51808 42896
rect 51958 42882 52098 42896
rect 52248 42882 53056 42896
rect 53206 42882 53346 42896
rect 53496 42882 54304 42896
rect 54454 42882 54594 42896
rect 54744 42882 55552 42896
rect 55702 42882 55842 42896
rect 55992 42882 56800 42896
rect 56950 42882 57090 42896
rect 57240 42882 58048 42896
rect 58198 42882 58338 42896
rect 58488 42882 58934 42896
rect 16898 42834 16980 42848
rect 17188 42834 17270 42848
rect 18146 42834 18228 42848
rect 18436 42834 18518 42848
rect 19394 42834 19476 42848
rect 19684 42834 19766 42848
rect 20642 42834 20724 42848
rect 20932 42834 21014 42848
rect 21890 42834 21972 42848
rect 22180 42834 22262 42848
rect 23138 42834 23220 42848
rect 23428 42834 23510 42848
rect 24386 42834 24468 42848
rect 24676 42834 24758 42848
rect 25634 42834 25716 42848
rect 25924 42834 26006 42848
rect 26882 42834 26964 42848
rect 27172 42834 27254 42848
rect 28130 42834 28212 42848
rect 28420 42834 28502 42848
rect 29378 42834 29460 42848
rect 29668 42834 29750 42848
rect 30626 42834 30708 42848
rect 30916 42834 30998 42848
rect 31874 42834 31956 42848
rect 32164 42834 32246 42848
rect 33122 42834 33204 42848
rect 33412 42834 33494 42848
rect 34370 42834 34452 42848
rect 34660 42834 34742 42848
rect 35618 42834 35700 42848
rect 35908 42834 35990 42848
rect 36866 42834 36948 42848
rect 37156 42834 37238 42848
rect 38114 42834 38196 42848
rect 38404 42834 38486 42848
rect 39362 42834 39444 42848
rect 39652 42834 39734 42848
rect 40610 42834 40692 42848
rect 40900 42834 40982 42848
rect 41858 42834 41940 42848
rect 42148 42834 42230 42848
rect 43106 42834 43188 42848
rect 43396 42834 43478 42848
rect 44354 42834 44436 42848
rect 44644 42834 44726 42848
rect 45602 42834 45684 42848
rect 45892 42834 45974 42848
rect 46850 42834 46932 42848
rect 47140 42834 47222 42848
rect 48098 42834 48180 42848
rect 48388 42834 48470 42848
rect 49346 42834 49428 42848
rect 49636 42834 49718 42848
rect 50594 42834 50676 42848
rect 50884 42834 50966 42848
rect 51842 42834 51924 42848
rect 52132 42834 52214 42848
rect 53090 42834 53172 42848
rect 53380 42834 53462 42848
rect 54338 42834 54420 42848
rect 54628 42834 54710 42848
rect 55586 42834 55668 42848
rect 55876 42834 55958 42848
rect 56834 42834 56916 42848
rect 57124 42834 57206 42848
rect 58082 42834 58164 42848
rect 58372 42834 58454 42848
rect 16418 42786 58934 42834
rect 16418 42628 58934 42738
rect 16418 42532 58934 42580
rect 16898 42518 16980 42532
rect 17188 42518 17270 42532
rect 18146 42518 18228 42532
rect 18436 42518 18518 42532
rect 19394 42518 19476 42532
rect 19684 42518 19766 42532
rect 20642 42518 20724 42532
rect 20932 42518 21014 42532
rect 21890 42518 21972 42532
rect 22180 42518 22262 42532
rect 23138 42518 23220 42532
rect 23428 42518 23510 42532
rect 24386 42518 24468 42532
rect 24676 42518 24758 42532
rect 25634 42518 25716 42532
rect 25924 42518 26006 42532
rect 26882 42518 26964 42532
rect 27172 42518 27254 42532
rect 28130 42518 28212 42532
rect 28420 42518 28502 42532
rect 29378 42518 29460 42532
rect 29668 42518 29750 42532
rect 30626 42518 30708 42532
rect 30916 42518 30998 42532
rect 31874 42518 31956 42532
rect 32164 42518 32246 42532
rect 33122 42518 33204 42532
rect 33412 42518 33494 42532
rect 34370 42518 34452 42532
rect 34660 42518 34742 42532
rect 35618 42518 35700 42532
rect 35908 42518 35990 42532
rect 36866 42518 36948 42532
rect 37156 42518 37238 42532
rect 38114 42518 38196 42532
rect 38404 42518 38486 42532
rect 39362 42518 39444 42532
rect 39652 42518 39734 42532
rect 40610 42518 40692 42532
rect 40900 42518 40982 42532
rect 41858 42518 41940 42532
rect 42148 42518 42230 42532
rect 43106 42518 43188 42532
rect 43396 42518 43478 42532
rect 44354 42518 44436 42532
rect 44644 42518 44726 42532
rect 45602 42518 45684 42532
rect 45892 42518 45974 42532
rect 46850 42518 46932 42532
rect 47140 42518 47222 42532
rect 48098 42518 48180 42532
rect 48388 42518 48470 42532
rect 49346 42518 49428 42532
rect 49636 42518 49718 42532
rect 50594 42518 50676 42532
rect 50884 42518 50966 42532
rect 51842 42518 51924 42532
rect 52132 42518 52214 42532
rect 53090 42518 53172 42532
rect 53380 42518 53462 42532
rect 54338 42518 54420 42532
rect 54628 42518 54710 42532
rect 55586 42518 55668 42532
rect 55876 42518 55958 42532
rect 56834 42518 56916 42532
rect 57124 42518 57206 42532
rect 58082 42518 58164 42532
rect 58372 42518 58454 42532
rect 16418 42470 16864 42484
rect 17014 42470 17154 42484
rect 17304 42470 18112 42484
rect 18262 42470 18402 42484
rect 18552 42470 19360 42484
rect 19510 42470 19650 42484
rect 19800 42470 20608 42484
rect 20758 42470 20898 42484
rect 21048 42470 21856 42484
rect 22006 42470 22146 42484
rect 22296 42470 23104 42484
rect 23254 42470 23394 42484
rect 23544 42470 24352 42484
rect 24502 42470 24642 42484
rect 24792 42470 25600 42484
rect 25750 42470 25890 42484
rect 26040 42470 26848 42484
rect 26998 42470 27138 42484
rect 27288 42470 28096 42484
rect 28246 42470 28386 42484
rect 28536 42470 29344 42484
rect 29494 42470 29634 42484
rect 29784 42470 30592 42484
rect 30742 42470 30882 42484
rect 31032 42470 31840 42484
rect 31990 42470 32130 42484
rect 32280 42470 33088 42484
rect 33238 42470 33378 42484
rect 33528 42470 34336 42484
rect 34486 42470 34626 42484
rect 34776 42470 35584 42484
rect 35734 42470 35874 42484
rect 36024 42470 36832 42484
rect 36982 42470 37122 42484
rect 37272 42470 38080 42484
rect 38230 42470 38370 42484
rect 38520 42470 39328 42484
rect 39478 42470 39618 42484
rect 39768 42470 40576 42484
rect 40726 42470 40866 42484
rect 41016 42470 41824 42484
rect 41974 42470 42114 42484
rect 42264 42470 43072 42484
rect 43222 42470 43362 42484
rect 43512 42470 44320 42484
rect 44470 42470 44610 42484
rect 44760 42470 45568 42484
rect 45718 42470 45858 42484
rect 46008 42470 46816 42484
rect 46966 42470 47106 42484
rect 47256 42470 48064 42484
rect 48214 42470 48354 42484
rect 48504 42470 49312 42484
rect 49462 42470 49602 42484
rect 49752 42470 50560 42484
rect 50710 42470 50850 42484
rect 51000 42470 51808 42484
rect 51958 42470 52098 42484
rect 52248 42470 53056 42484
rect 53206 42470 53346 42484
rect 53496 42470 54304 42484
rect 54454 42470 54594 42484
rect 54744 42470 55552 42484
rect 55702 42470 55842 42484
rect 55992 42470 56800 42484
rect 56950 42470 57090 42484
rect 57240 42470 58048 42484
rect 58198 42470 58338 42484
rect 58488 42470 58934 42484
rect 16418 42422 58934 42470
rect 16418 42408 16864 42422
rect 17014 42408 17154 42422
rect 17304 42408 18112 42422
rect 18262 42408 18402 42422
rect 18552 42408 19360 42422
rect 19510 42408 19650 42422
rect 19800 42408 20608 42422
rect 20758 42408 20898 42422
rect 21048 42408 21856 42422
rect 22006 42408 22146 42422
rect 22296 42408 23104 42422
rect 23254 42408 23394 42422
rect 23544 42408 24352 42422
rect 24502 42408 24642 42422
rect 24792 42408 25600 42422
rect 25750 42408 25890 42422
rect 26040 42408 26848 42422
rect 26998 42408 27138 42422
rect 27288 42408 28096 42422
rect 28246 42408 28386 42422
rect 28536 42408 29344 42422
rect 29494 42408 29634 42422
rect 29784 42408 30592 42422
rect 30742 42408 30882 42422
rect 31032 42408 31840 42422
rect 31990 42408 32130 42422
rect 32280 42408 33088 42422
rect 33238 42408 33378 42422
rect 33528 42408 34336 42422
rect 34486 42408 34626 42422
rect 34776 42408 35584 42422
rect 35734 42408 35874 42422
rect 36024 42408 36832 42422
rect 36982 42408 37122 42422
rect 37272 42408 38080 42422
rect 38230 42408 38370 42422
rect 38520 42408 39328 42422
rect 39478 42408 39618 42422
rect 39768 42408 40576 42422
rect 40726 42408 40866 42422
rect 41016 42408 41824 42422
rect 41974 42408 42114 42422
rect 42264 42408 43072 42422
rect 43222 42408 43362 42422
rect 43512 42408 44320 42422
rect 44470 42408 44610 42422
rect 44760 42408 45568 42422
rect 45718 42408 45858 42422
rect 46008 42408 46816 42422
rect 46966 42408 47106 42422
rect 47256 42408 48064 42422
rect 48214 42408 48354 42422
rect 48504 42408 49312 42422
rect 49462 42408 49602 42422
rect 49752 42408 50560 42422
rect 50710 42408 50850 42422
rect 51000 42408 51808 42422
rect 51958 42408 52098 42422
rect 52248 42408 53056 42422
rect 53206 42408 53346 42422
rect 53496 42408 54304 42422
rect 54454 42408 54594 42422
rect 54744 42408 55552 42422
rect 55702 42408 55842 42422
rect 55992 42408 56800 42422
rect 56950 42408 57090 42422
rect 57240 42408 58048 42422
rect 58198 42408 58338 42422
rect 58488 42408 58934 42422
rect 16898 42360 16980 42374
rect 17188 42360 17270 42374
rect 18146 42360 18228 42374
rect 18436 42360 18518 42374
rect 19394 42360 19476 42374
rect 19684 42360 19766 42374
rect 20642 42360 20724 42374
rect 20932 42360 21014 42374
rect 21890 42360 21972 42374
rect 22180 42360 22262 42374
rect 23138 42360 23220 42374
rect 23428 42360 23510 42374
rect 24386 42360 24468 42374
rect 24676 42360 24758 42374
rect 25634 42360 25716 42374
rect 25924 42360 26006 42374
rect 26882 42360 26964 42374
rect 27172 42360 27254 42374
rect 28130 42360 28212 42374
rect 28420 42360 28502 42374
rect 29378 42360 29460 42374
rect 29668 42360 29750 42374
rect 30626 42360 30708 42374
rect 30916 42360 30998 42374
rect 31874 42360 31956 42374
rect 32164 42360 32246 42374
rect 33122 42360 33204 42374
rect 33412 42360 33494 42374
rect 34370 42360 34452 42374
rect 34660 42360 34742 42374
rect 35618 42360 35700 42374
rect 35908 42360 35990 42374
rect 36866 42360 36948 42374
rect 37156 42360 37238 42374
rect 38114 42360 38196 42374
rect 38404 42360 38486 42374
rect 39362 42360 39444 42374
rect 39652 42360 39734 42374
rect 40610 42360 40692 42374
rect 40900 42360 40982 42374
rect 41858 42360 41940 42374
rect 42148 42360 42230 42374
rect 43106 42360 43188 42374
rect 43396 42360 43478 42374
rect 44354 42360 44436 42374
rect 44644 42360 44726 42374
rect 45602 42360 45684 42374
rect 45892 42360 45974 42374
rect 46850 42360 46932 42374
rect 47140 42360 47222 42374
rect 48098 42360 48180 42374
rect 48388 42360 48470 42374
rect 49346 42360 49428 42374
rect 49636 42360 49718 42374
rect 50594 42360 50676 42374
rect 50884 42360 50966 42374
rect 51842 42360 51924 42374
rect 52132 42360 52214 42374
rect 53090 42360 53172 42374
rect 53380 42360 53462 42374
rect 54338 42360 54420 42374
rect 54628 42360 54710 42374
rect 55586 42360 55668 42374
rect 55876 42360 55958 42374
rect 56834 42360 56916 42374
rect 57124 42360 57206 42374
rect 58082 42360 58164 42374
rect 58372 42360 58454 42374
rect 16418 42312 58934 42360
rect 16418 42216 58934 42264
rect 16898 42202 16980 42216
rect 17188 42202 17270 42216
rect 18146 42202 18228 42216
rect 18436 42202 18518 42216
rect 19394 42202 19476 42216
rect 19684 42202 19766 42216
rect 20642 42202 20724 42216
rect 20932 42202 21014 42216
rect 21890 42202 21972 42216
rect 22180 42202 22262 42216
rect 23138 42202 23220 42216
rect 23428 42202 23510 42216
rect 24386 42202 24468 42216
rect 24676 42202 24758 42216
rect 25634 42202 25716 42216
rect 25924 42202 26006 42216
rect 26882 42202 26964 42216
rect 27172 42202 27254 42216
rect 28130 42202 28212 42216
rect 28420 42202 28502 42216
rect 29378 42202 29460 42216
rect 29668 42202 29750 42216
rect 30626 42202 30708 42216
rect 30916 42202 30998 42216
rect 31874 42202 31956 42216
rect 32164 42202 32246 42216
rect 33122 42202 33204 42216
rect 33412 42202 33494 42216
rect 34370 42202 34452 42216
rect 34660 42202 34742 42216
rect 35618 42202 35700 42216
rect 35908 42202 35990 42216
rect 36866 42202 36948 42216
rect 37156 42202 37238 42216
rect 38114 42202 38196 42216
rect 38404 42202 38486 42216
rect 39362 42202 39444 42216
rect 39652 42202 39734 42216
rect 40610 42202 40692 42216
rect 40900 42202 40982 42216
rect 41858 42202 41940 42216
rect 42148 42202 42230 42216
rect 43106 42202 43188 42216
rect 43396 42202 43478 42216
rect 44354 42202 44436 42216
rect 44644 42202 44726 42216
rect 45602 42202 45684 42216
rect 45892 42202 45974 42216
rect 46850 42202 46932 42216
rect 47140 42202 47222 42216
rect 48098 42202 48180 42216
rect 48388 42202 48470 42216
rect 49346 42202 49428 42216
rect 49636 42202 49718 42216
rect 50594 42202 50676 42216
rect 50884 42202 50966 42216
rect 51842 42202 51924 42216
rect 52132 42202 52214 42216
rect 53090 42202 53172 42216
rect 53380 42202 53462 42216
rect 54338 42202 54420 42216
rect 54628 42202 54710 42216
rect 55586 42202 55668 42216
rect 55876 42202 55958 42216
rect 56834 42202 56916 42216
rect 57124 42202 57206 42216
rect 58082 42202 58164 42216
rect 58372 42202 58454 42216
rect 16418 42154 16864 42168
rect 17014 42154 17154 42168
rect 17304 42154 18112 42168
rect 18262 42154 18402 42168
rect 18552 42154 19360 42168
rect 19510 42154 19650 42168
rect 19800 42154 20608 42168
rect 20758 42154 20898 42168
rect 21048 42154 21856 42168
rect 22006 42154 22146 42168
rect 22296 42154 23104 42168
rect 23254 42154 23394 42168
rect 23544 42154 24352 42168
rect 24502 42154 24642 42168
rect 24792 42154 25600 42168
rect 25750 42154 25890 42168
rect 26040 42154 26848 42168
rect 26998 42154 27138 42168
rect 27288 42154 28096 42168
rect 28246 42154 28386 42168
rect 28536 42154 29344 42168
rect 29494 42154 29634 42168
rect 29784 42154 30592 42168
rect 30742 42154 30882 42168
rect 31032 42154 31840 42168
rect 31990 42154 32130 42168
rect 32280 42154 33088 42168
rect 33238 42154 33378 42168
rect 33528 42154 34336 42168
rect 34486 42154 34626 42168
rect 34776 42154 35584 42168
rect 35734 42154 35874 42168
rect 36024 42154 36832 42168
rect 36982 42154 37122 42168
rect 37272 42154 38080 42168
rect 38230 42154 38370 42168
rect 38520 42154 39328 42168
rect 39478 42154 39618 42168
rect 39768 42154 40576 42168
rect 40726 42154 40866 42168
rect 41016 42154 41824 42168
rect 41974 42154 42114 42168
rect 42264 42154 43072 42168
rect 43222 42154 43362 42168
rect 43512 42154 44320 42168
rect 44470 42154 44610 42168
rect 44760 42154 45568 42168
rect 45718 42154 45858 42168
rect 46008 42154 46816 42168
rect 46966 42154 47106 42168
rect 47256 42154 48064 42168
rect 48214 42154 48354 42168
rect 48504 42154 49312 42168
rect 49462 42154 49602 42168
rect 49752 42154 50560 42168
rect 50710 42154 50850 42168
rect 51000 42154 51808 42168
rect 51958 42154 52098 42168
rect 52248 42154 53056 42168
rect 53206 42154 53346 42168
rect 53496 42154 54304 42168
rect 54454 42154 54594 42168
rect 54744 42154 55552 42168
rect 55702 42154 55842 42168
rect 55992 42154 56800 42168
rect 56950 42154 57090 42168
rect 57240 42154 58048 42168
rect 58198 42154 58338 42168
rect 58488 42154 58934 42168
rect 16418 42106 58934 42154
rect 16418 42092 16864 42106
rect 17014 42092 17154 42106
rect 17304 42092 18112 42106
rect 18262 42092 18402 42106
rect 18552 42092 19360 42106
rect 19510 42092 19650 42106
rect 19800 42092 20608 42106
rect 20758 42092 20898 42106
rect 21048 42092 21856 42106
rect 22006 42092 22146 42106
rect 22296 42092 23104 42106
rect 23254 42092 23394 42106
rect 23544 42092 24352 42106
rect 24502 42092 24642 42106
rect 24792 42092 25600 42106
rect 25750 42092 25890 42106
rect 26040 42092 26848 42106
rect 26998 42092 27138 42106
rect 27288 42092 28096 42106
rect 28246 42092 28386 42106
rect 28536 42092 29344 42106
rect 29494 42092 29634 42106
rect 29784 42092 30592 42106
rect 30742 42092 30882 42106
rect 31032 42092 31840 42106
rect 31990 42092 32130 42106
rect 32280 42092 33088 42106
rect 33238 42092 33378 42106
rect 33528 42092 34336 42106
rect 34486 42092 34626 42106
rect 34776 42092 35584 42106
rect 35734 42092 35874 42106
rect 36024 42092 36832 42106
rect 36982 42092 37122 42106
rect 37272 42092 38080 42106
rect 38230 42092 38370 42106
rect 38520 42092 39328 42106
rect 39478 42092 39618 42106
rect 39768 42092 40576 42106
rect 40726 42092 40866 42106
rect 41016 42092 41824 42106
rect 41974 42092 42114 42106
rect 42264 42092 43072 42106
rect 43222 42092 43362 42106
rect 43512 42092 44320 42106
rect 44470 42092 44610 42106
rect 44760 42092 45568 42106
rect 45718 42092 45858 42106
rect 46008 42092 46816 42106
rect 46966 42092 47106 42106
rect 47256 42092 48064 42106
rect 48214 42092 48354 42106
rect 48504 42092 49312 42106
rect 49462 42092 49602 42106
rect 49752 42092 50560 42106
rect 50710 42092 50850 42106
rect 51000 42092 51808 42106
rect 51958 42092 52098 42106
rect 52248 42092 53056 42106
rect 53206 42092 53346 42106
rect 53496 42092 54304 42106
rect 54454 42092 54594 42106
rect 54744 42092 55552 42106
rect 55702 42092 55842 42106
rect 55992 42092 56800 42106
rect 56950 42092 57090 42106
rect 57240 42092 58048 42106
rect 58198 42092 58338 42106
rect 58488 42092 58934 42106
rect 16898 42044 16980 42058
rect 17188 42044 17270 42058
rect 18146 42044 18228 42058
rect 18436 42044 18518 42058
rect 19394 42044 19476 42058
rect 19684 42044 19766 42058
rect 20642 42044 20724 42058
rect 20932 42044 21014 42058
rect 21890 42044 21972 42058
rect 22180 42044 22262 42058
rect 23138 42044 23220 42058
rect 23428 42044 23510 42058
rect 24386 42044 24468 42058
rect 24676 42044 24758 42058
rect 25634 42044 25716 42058
rect 25924 42044 26006 42058
rect 26882 42044 26964 42058
rect 27172 42044 27254 42058
rect 28130 42044 28212 42058
rect 28420 42044 28502 42058
rect 29378 42044 29460 42058
rect 29668 42044 29750 42058
rect 30626 42044 30708 42058
rect 30916 42044 30998 42058
rect 31874 42044 31956 42058
rect 32164 42044 32246 42058
rect 33122 42044 33204 42058
rect 33412 42044 33494 42058
rect 34370 42044 34452 42058
rect 34660 42044 34742 42058
rect 35618 42044 35700 42058
rect 35908 42044 35990 42058
rect 36866 42044 36948 42058
rect 37156 42044 37238 42058
rect 38114 42044 38196 42058
rect 38404 42044 38486 42058
rect 39362 42044 39444 42058
rect 39652 42044 39734 42058
rect 40610 42044 40692 42058
rect 40900 42044 40982 42058
rect 41858 42044 41940 42058
rect 42148 42044 42230 42058
rect 43106 42044 43188 42058
rect 43396 42044 43478 42058
rect 44354 42044 44436 42058
rect 44644 42044 44726 42058
rect 45602 42044 45684 42058
rect 45892 42044 45974 42058
rect 46850 42044 46932 42058
rect 47140 42044 47222 42058
rect 48098 42044 48180 42058
rect 48388 42044 48470 42058
rect 49346 42044 49428 42058
rect 49636 42044 49718 42058
rect 50594 42044 50676 42058
rect 50884 42044 50966 42058
rect 51842 42044 51924 42058
rect 52132 42044 52214 42058
rect 53090 42044 53172 42058
rect 53380 42044 53462 42058
rect 54338 42044 54420 42058
rect 54628 42044 54710 42058
rect 55586 42044 55668 42058
rect 55876 42044 55958 42058
rect 56834 42044 56916 42058
rect 57124 42044 57206 42058
rect 58082 42044 58164 42058
rect 58372 42044 58454 42058
rect 16418 41996 58934 42044
rect 16418 41838 58934 41948
rect 16418 41742 58934 41790
rect 16898 41728 16980 41742
rect 17188 41728 17270 41742
rect 18146 41728 18228 41742
rect 18436 41728 18518 41742
rect 19394 41728 19476 41742
rect 19684 41728 19766 41742
rect 20642 41728 20724 41742
rect 20932 41728 21014 41742
rect 21890 41728 21972 41742
rect 22180 41728 22262 41742
rect 23138 41728 23220 41742
rect 23428 41728 23510 41742
rect 24386 41728 24468 41742
rect 24676 41728 24758 41742
rect 25634 41728 25716 41742
rect 25924 41728 26006 41742
rect 26882 41728 26964 41742
rect 27172 41728 27254 41742
rect 28130 41728 28212 41742
rect 28420 41728 28502 41742
rect 29378 41728 29460 41742
rect 29668 41728 29750 41742
rect 30626 41728 30708 41742
rect 30916 41728 30998 41742
rect 31874 41728 31956 41742
rect 32164 41728 32246 41742
rect 33122 41728 33204 41742
rect 33412 41728 33494 41742
rect 34370 41728 34452 41742
rect 34660 41728 34742 41742
rect 35618 41728 35700 41742
rect 35908 41728 35990 41742
rect 36866 41728 36948 41742
rect 37156 41728 37238 41742
rect 38114 41728 38196 41742
rect 38404 41728 38486 41742
rect 39362 41728 39444 41742
rect 39652 41728 39734 41742
rect 40610 41728 40692 41742
rect 40900 41728 40982 41742
rect 41858 41728 41940 41742
rect 42148 41728 42230 41742
rect 43106 41728 43188 41742
rect 43396 41728 43478 41742
rect 44354 41728 44436 41742
rect 44644 41728 44726 41742
rect 45602 41728 45684 41742
rect 45892 41728 45974 41742
rect 46850 41728 46932 41742
rect 47140 41728 47222 41742
rect 48098 41728 48180 41742
rect 48388 41728 48470 41742
rect 49346 41728 49428 41742
rect 49636 41728 49718 41742
rect 50594 41728 50676 41742
rect 50884 41728 50966 41742
rect 51842 41728 51924 41742
rect 52132 41728 52214 41742
rect 53090 41728 53172 41742
rect 53380 41728 53462 41742
rect 54338 41728 54420 41742
rect 54628 41728 54710 41742
rect 55586 41728 55668 41742
rect 55876 41728 55958 41742
rect 56834 41728 56916 41742
rect 57124 41728 57206 41742
rect 58082 41728 58164 41742
rect 58372 41728 58454 41742
rect 16418 41680 16864 41694
rect 17014 41680 17154 41694
rect 17304 41680 18112 41694
rect 18262 41680 18402 41694
rect 18552 41680 19360 41694
rect 19510 41680 19650 41694
rect 19800 41680 20608 41694
rect 20758 41680 20898 41694
rect 21048 41680 21856 41694
rect 22006 41680 22146 41694
rect 22296 41680 23104 41694
rect 23254 41680 23394 41694
rect 23544 41680 24352 41694
rect 24502 41680 24642 41694
rect 24792 41680 25600 41694
rect 25750 41680 25890 41694
rect 26040 41680 26848 41694
rect 26998 41680 27138 41694
rect 27288 41680 28096 41694
rect 28246 41680 28386 41694
rect 28536 41680 29344 41694
rect 29494 41680 29634 41694
rect 29784 41680 30592 41694
rect 30742 41680 30882 41694
rect 31032 41680 31840 41694
rect 31990 41680 32130 41694
rect 32280 41680 33088 41694
rect 33238 41680 33378 41694
rect 33528 41680 34336 41694
rect 34486 41680 34626 41694
rect 34776 41680 35584 41694
rect 35734 41680 35874 41694
rect 36024 41680 36832 41694
rect 36982 41680 37122 41694
rect 37272 41680 38080 41694
rect 38230 41680 38370 41694
rect 38520 41680 39328 41694
rect 39478 41680 39618 41694
rect 39768 41680 40576 41694
rect 40726 41680 40866 41694
rect 41016 41680 41824 41694
rect 41974 41680 42114 41694
rect 42264 41680 43072 41694
rect 43222 41680 43362 41694
rect 43512 41680 44320 41694
rect 44470 41680 44610 41694
rect 44760 41680 45568 41694
rect 45718 41680 45858 41694
rect 46008 41680 46816 41694
rect 46966 41680 47106 41694
rect 47256 41680 48064 41694
rect 48214 41680 48354 41694
rect 48504 41680 49312 41694
rect 49462 41680 49602 41694
rect 49752 41680 50560 41694
rect 50710 41680 50850 41694
rect 51000 41680 51808 41694
rect 51958 41680 52098 41694
rect 52248 41680 53056 41694
rect 53206 41680 53346 41694
rect 53496 41680 54304 41694
rect 54454 41680 54594 41694
rect 54744 41680 55552 41694
rect 55702 41680 55842 41694
rect 55992 41680 56800 41694
rect 56950 41680 57090 41694
rect 57240 41680 58048 41694
rect 58198 41680 58338 41694
rect 58488 41680 58934 41694
rect 16418 41632 58934 41680
rect 16418 41618 16864 41632
rect 17014 41618 17154 41632
rect 17304 41618 18112 41632
rect 18262 41618 18402 41632
rect 18552 41618 19360 41632
rect 19510 41618 19650 41632
rect 19800 41618 20608 41632
rect 20758 41618 20898 41632
rect 21048 41618 21856 41632
rect 22006 41618 22146 41632
rect 22296 41618 23104 41632
rect 23254 41618 23394 41632
rect 23544 41618 24352 41632
rect 24502 41618 24642 41632
rect 24792 41618 25600 41632
rect 25750 41618 25890 41632
rect 26040 41618 26848 41632
rect 26998 41618 27138 41632
rect 27288 41618 28096 41632
rect 28246 41618 28386 41632
rect 28536 41618 29344 41632
rect 29494 41618 29634 41632
rect 29784 41618 30592 41632
rect 30742 41618 30882 41632
rect 31032 41618 31840 41632
rect 31990 41618 32130 41632
rect 32280 41618 33088 41632
rect 33238 41618 33378 41632
rect 33528 41618 34336 41632
rect 34486 41618 34626 41632
rect 34776 41618 35584 41632
rect 35734 41618 35874 41632
rect 36024 41618 36832 41632
rect 36982 41618 37122 41632
rect 37272 41618 38080 41632
rect 38230 41618 38370 41632
rect 38520 41618 39328 41632
rect 39478 41618 39618 41632
rect 39768 41618 40576 41632
rect 40726 41618 40866 41632
rect 41016 41618 41824 41632
rect 41974 41618 42114 41632
rect 42264 41618 43072 41632
rect 43222 41618 43362 41632
rect 43512 41618 44320 41632
rect 44470 41618 44610 41632
rect 44760 41618 45568 41632
rect 45718 41618 45858 41632
rect 46008 41618 46816 41632
rect 46966 41618 47106 41632
rect 47256 41618 48064 41632
rect 48214 41618 48354 41632
rect 48504 41618 49312 41632
rect 49462 41618 49602 41632
rect 49752 41618 50560 41632
rect 50710 41618 50850 41632
rect 51000 41618 51808 41632
rect 51958 41618 52098 41632
rect 52248 41618 53056 41632
rect 53206 41618 53346 41632
rect 53496 41618 54304 41632
rect 54454 41618 54594 41632
rect 54744 41618 55552 41632
rect 55702 41618 55842 41632
rect 55992 41618 56800 41632
rect 56950 41618 57090 41632
rect 57240 41618 58048 41632
rect 58198 41618 58338 41632
rect 58488 41618 58934 41632
rect 16898 41570 16980 41584
rect 17188 41570 17270 41584
rect 18146 41570 18228 41584
rect 18436 41570 18518 41584
rect 19394 41570 19476 41584
rect 19684 41570 19766 41584
rect 20642 41570 20724 41584
rect 20932 41570 21014 41584
rect 21890 41570 21972 41584
rect 22180 41570 22262 41584
rect 23138 41570 23220 41584
rect 23428 41570 23510 41584
rect 24386 41570 24468 41584
rect 24676 41570 24758 41584
rect 25634 41570 25716 41584
rect 25924 41570 26006 41584
rect 26882 41570 26964 41584
rect 27172 41570 27254 41584
rect 28130 41570 28212 41584
rect 28420 41570 28502 41584
rect 29378 41570 29460 41584
rect 29668 41570 29750 41584
rect 30626 41570 30708 41584
rect 30916 41570 30998 41584
rect 31874 41570 31956 41584
rect 32164 41570 32246 41584
rect 33122 41570 33204 41584
rect 33412 41570 33494 41584
rect 34370 41570 34452 41584
rect 34660 41570 34742 41584
rect 35618 41570 35700 41584
rect 35908 41570 35990 41584
rect 36866 41570 36948 41584
rect 37156 41570 37238 41584
rect 38114 41570 38196 41584
rect 38404 41570 38486 41584
rect 39362 41570 39444 41584
rect 39652 41570 39734 41584
rect 40610 41570 40692 41584
rect 40900 41570 40982 41584
rect 41858 41570 41940 41584
rect 42148 41570 42230 41584
rect 43106 41570 43188 41584
rect 43396 41570 43478 41584
rect 44354 41570 44436 41584
rect 44644 41570 44726 41584
rect 45602 41570 45684 41584
rect 45892 41570 45974 41584
rect 46850 41570 46932 41584
rect 47140 41570 47222 41584
rect 48098 41570 48180 41584
rect 48388 41570 48470 41584
rect 49346 41570 49428 41584
rect 49636 41570 49718 41584
rect 50594 41570 50676 41584
rect 50884 41570 50966 41584
rect 51842 41570 51924 41584
rect 52132 41570 52214 41584
rect 53090 41570 53172 41584
rect 53380 41570 53462 41584
rect 54338 41570 54420 41584
rect 54628 41570 54710 41584
rect 55586 41570 55668 41584
rect 55876 41570 55958 41584
rect 56834 41570 56916 41584
rect 57124 41570 57206 41584
rect 58082 41570 58164 41584
rect 58372 41570 58454 41584
rect 16418 41522 58934 41570
rect 16418 41426 58934 41474
rect 16898 41412 16980 41426
rect 17188 41412 17270 41426
rect 18146 41412 18228 41426
rect 18436 41412 18518 41426
rect 19394 41412 19476 41426
rect 19684 41412 19766 41426
rect 20642 41412 20724 41426
rect 20932 41412 21014 41426
rect 21890 41412 21972 41426
rect 22180 41412 22262 41426
rect 23138 41412 23220 41426
rect 23428 41412 23510 41426
rect 24386 41412 24468 41426
rect 24676 41412 24758 41426
rect 25634 41412 25716 41426
rect 25924 41412 26006 41426
rect 26882 41412 26964 41426
rect 27172 41412 27254 41426
rect 28130 41412 28212 41426
rect 28420 41412 28502 41426
rect 29378 41412 29460 41426
rect 29668 41412 29750 41426
rect 30626 41412 30708 41426
rect 30916 41412 30998 41426
rect 31874 41412 31956 41426
rect 32164 41412 32246 41426
rect 33122 41412 33204 41426
rect 33412 41412 33494 41426
rect 34370 41412 34452 41426
rect 34660 41412 34742 41426
rect 35618 41412 35700 41426
rect 35908 41412 35990 41426
rect 36866 41412 36948 41426
rect 37156 41412 37238 41426
rect 38114 41412 38196 41426
rect 38404 41412 38486 41426
rect 39362 41412 39444 41426
rect 39652 41412 39734 41426
rect 40610 41412 40692 41426
rect 40900 41412 40982 41426
rect 41858 41412 41940 41426
rect 42148 41412 42230 41426
rect 43106 41412 43188 41426
rect 43396 41412 43478 41426
rect 44354 41412 44436 41426
rect 44644 41412 44726 41426
rect 45602 41412 45684 41426
rect 45892 41412 45974 41426
rect 46850 41412 46932 41426
rect 47140 41412 47222 41426
rect 48098 41412 48180 41426
rect 48388 41412 48470 41426
rect 49346 41412 49428 41426
rect 49636 41412 49718 41426
rect 50594 41412 50676 41426
rect 50884 41412 50966 41426
rect 51842 41412 51924 41426
rect 52132 41412 52214 41426
rect 53090 41412 53172 41426
rect 53380 41412 53462 41426
rect 54338 41412 54420 41426
rect 54628 41412 54710 41426
rect 55586 41412 55668 41426
rect 55876 41412 55958 41426
rect 56834 41412 56916 41426
rect 57124 41412 57206 41426
rect 58082 41412 58164 41426
rect 58372 41412 58454 41426
rect 16418 41364 16864 41378
rect 17014 41364 17154 41378
rect 17304 41364 18112 41378
rect 18262 41364 18402 41378
rect 18552 41364 19360 41378
rect 19510 41364 19650 41378
rect 19800 41364 20608 41378
rect 20758 41364 20898 41378
rect 21048 41364 21856 41378
rect 22006 41364 22146 41378
rect 22296 41364 23104 41378
rect 23254 41364 23394 41378
rect 23544 41364 24352 41378
rect 24502 41364 24642 41378
rect 24792 41364 25600 41378
rect 25750 41364 25890 41378
rect 26040 41364 26848 41378
rect 26998 41364 27138 41378
rect 27288 41364 28096 41378
rect 28246 41364 28386 41378
rect 28536 41364 29344 41378
rect 29494 41364 29634 41378
rect 29784 41364 30592 41378
rect 30742 41364 30882 41378
rect 31032 41364 31840 41378
rect 31990 41364 32130 41378
rect 32280 41364 33088 41378
rect 33238 41364 33378 41378
rect 33528 41364 34336 41378
rect 34486 41364 34626 41378
rect 34776 41364 35584 41378
rect 35734 41364 35874 41378
rect 36024 41364 36832 41378
rect 36982 41364 37122 41378
rect 37272 41364 38080 41378
rect 38230 41364 38370 41378
rect 38520 41364 39328 41378
rect 39478 41364 39618 41378
rect 39768 41364 40576 41378
rect 40726 41364 40866 41378
rect 41016 41364 41824 41378
rect 41974 41364 42114 41378
rect 42264 41364 43072 41378
rect 43222 41364 43362 41378
rect 43512 41364 44320 41378
rect 44470 41364 44610 41378
rect 44760 41364 45568 41378
rect 45718 41364 45858 41378
rect 46008 41364 46816 41378
rect 46966 41364 47106 41378
rect 47256 41364 48064 41378
rect 48214 41364 48354 41378
rect 48504 41364 49312 41378
rect 49462 41364 49602 41378
rect 49752 41364 50560 41378
rect 50710 41364 50850 41378
rect 51000 41364 51808 41378
rect 51958 41364 52098 41378
rect 52248 41364 53056 41378
rect 53206 41364 53346 41378
rect 53496 41364 54304 41378
rect 54454 41364 54594 41378
rect 54744 41364 55552 41378
rect 55702 41364 55842 41378
rect 55992 41364 56800 41378
rect 56950 41364 57090 41378
rect 57240 41364 58048 41378
rect 58198 41364 58338 41378
rect 58488 41364 58934 41378
rect 16418 41316 58934 41364
rect 16418 41302 16864 41316
rect 17014 41302 17154 41316
rect 17304 41302 18112 41316
rect 18262 41302 18402 41316
rect 18552 41302 19360 41316
rect 19510 41302 19650 41316
rect 19800 41302 20608 41316
rect 20758 41302 20898 41316
rect 21048 41302 21856 41316
rect 22006 41302 22146 41316
rect 22296 41302 23104 41316
rect 23254 41302 23394 41316
rect 23544 41302 24352 41316
rect 24502 41302 24642 41316
rect 24792 41302 25600 41316
rect 25750 41302 25890 41316
rect 26040 41302 26848 41316
rect 26998 41302 27138 41316
rect 27288 41302 28096 41316
rect 28246 41302 28386 41316
rect 28536 41302 29344 41316
rect 29494 41302 29634 41316
rect 29784 41302 30592 41316
rect 30742 41302 30882 41316
rect 31032 41302 31840 41316
rect 31990 41302 32130 41316
rect 32280 41302 33088 41316
rect 33238 41302 33378 41316
rect 33528 41302 34336 41316
rect 34486 41302 34626 41316
rect 34776 41302 35584 41316
rect 35734 41302 35874 41316
rect 36024 41302 36832 41316
rect 36982 41302 37122 41316
rect 37272 41302 38080 41316
rect 38230 41302 38370 41316
rect 38520 41302 39328 41316
rect 39478 41302 39618 41316
rect 39768 41302 40576 41316
rect 40726 41302 40866 41316
rect 41016 41302 41824 41316
rect 41974 41302 42114 41316
rect 42264 41302 43072 41316
rect 43222 41302 43362 41316
rect 43512 41302 44320 41316
rect 44470 41302 44610 41316
rect 44760 41302 45568 41316
rect 45718 41302 45858 41316
rect 46008 41302 46816 41316
rect 46966 41302 47106 41316
rect 47256 41302 48064 41316
rect 48214 41302 48354 41316
rect 48504 41302 49312 41316
rect 49462 41302 49602 41316
rect 49752 41302 50560 41316
rect 50710 41302 50850 41316
rect 51000 41302 51808 41316
rect 51958 41302 52098 41316
rect 52248 41302 53056 41316
rect 53206 41302 53346 41316
rect 53496 41302 54304 41316
rect 54454 41302 54594 41316
rect 54744 41302 55552 41316
rect 55702 41302 55842 41316
rect 55992 41302 56800 41316
rect 56950 41302 57090 41316
rect 57240 41302 58048 41316
rect 58198 41302 58338 41316
rect 58488 41302 58934 41316
rect 16898 41254 16980 41268
rect 17188 41254 17270 41268
rect 18146 41254 18228 41268
rect 18436 41254 18518 41268
rect 19394 41254 19476 41268
rect 19684 41254 19766 41268
rect 20642 41254 20724 41268
rect 20932 41254 21014 41268
rect 21890 41254 21972 41268
rect 22180 41254 22262 41268
rect 23138 41254 23220 41268
rect 23428 41254 23510 41268
rect 24386 41254 24468 41268
rect 24676 41254 24758 41268
rect 25634 41254 25716 41268
rect 25924 41254 26006 41268
rect 26882 41254 26964 41268
rect 27172 41254 27254 41268
rect 28130 41254 28212 41268
rect 28420 41254 28502 41268
rect 29378 41254 29460 41268
rect 29668 41254 29750 41268
rect 30626 41254 30708 41268
rect 30916 41254 30998 41268
rect 31874 41254 31956 41268
rect 32164 41254 32246 41268
rect 33122 41254 33204 41268
rect 33412 41254 33494 41268
rect 34370 41254 34452 41268
rect 34660 41254 34742 41268
rect 35618 41254 35700 41268
rect 35908 41254 35990 41268
rect 36866 41254 36948 41268
rect 37156 41254 37238 41268
rect 38114 41254 38196 41268
rect 38404 41254 38486 41268
rect 39362 41254 39444 41268
rect 39652 41254 39734 41268
rect 40610 41254 40692 41268
rect 40900 41254 40982 41268
rect 41858 41254 41940 41268
rect 42148 41254 42230 41268
rect 43106 41254 43188 41268
rect 43396 41254 43478 41268
rect 44354 41254 44436 41268
rect 44644 41254 44726 41268
rect 45602 41254 45684 41268
rect 45892 41254 45974 41268
rect 46850 41254 46932 41268
rect 47140 41254 47222 41268
rect 48098 41254 48180 41268
rect 48388 41254 48470 41268
rect 49346 41254 49428 41268
rect 49636 41254 49718 41268
rect 50594 41254 50676 41268
rect 50884 41254 50966 41268
rect 51842 41254 51924 41268
rect 52132 41254 52214 41268
rect 53090 41254 53172 41268
rect 53380 41254 53462 41268
rect 54338 41254 54420 41268
rect 54628 41254 54710 41268
rect 55586 41254 55668 41268
rect 55876 41254 55958 41268
rect 56834 41254 56916 41268
rect 57124 41254 57206 41268
rect 58082 41254 58164 41268
rect 58372 41254 58454 41268
rect 16418 41206 58934 41254
rect 16418 41048 58934 41158
rect 16418 40952 58934 41000
rect 16898 40938 16980 40952
rect 17188 40938 17270 40952
rect 18146 40938 18228 40952
rect 18436 40938 18518 40952
rect 19394 40938 19476 40952
rect 19684 40938 19766 40952
rect 20642 40938 20724 40952
rect 20932 40938 21014 40952
rect 21890 40938 21972 40952
rect 22180 40938 22262 40952
rect 23138 40938 23220 40952
rect 23428 40938 23510 40952
rect 24386 40938 24468 40952
rect 24676 40938 24758 40952
rect 25634 40938 25716 40952
rect 25924 40938 26006 40952
rect 26882 40938 26964 40952
rect 27172 40938 27254 40952
rect 28130 40938 28212 40952
rect 28420 40938 28502 40952
rect 29378 40938 29460 40952
rect 29668 40938 29750 40952
rect 30626 40938 30708 40952
rect 30916 40938 30998 40952
rect 31874 40938 31956 40952
rect 32164 40938 32246 40952
rect 33122 40938 33204 40952
rect 33412 40938 33494 40952
rect 34370 40938 34452 40952
rect 34660 40938 34742 40952
rect 35618 40938 35700 40952
rect 35908 40938 35990 40952
rect 36866 40938 36948 40952
rect 37156 40938 37238 40952
rect 38114 40938 38196 40952
rect 38404 40938 38486 40952
rect 39362 40938 39444 40952
rect 39652 40938 39734 40952
rect 40610 40938 40692 40952
rect 40900 40938 40982 40952
rect 41858 40938 41940 40952
rect 42148 40938 42230 40952
rect 43106 40938 43188 40952
rect 43396 40938 43478 40952
rect 44354 40938 44436 40952
rect 44644 40938 44726 40952
rect 45602 40938 45684 40952
rect 45892 40938 45974 40952
rect 46850 40938 46932 40952
rect 47140 40938 47222 40952
rect 48098 40938 48180 40952
rect 48388 40938 48470 40952
rect 49346 40938 49428 40952
rect 49636 40938 49718 40952
rect 50594 40938 50676 40952
rect 50884 40938 50966 40952
rect 51842 40938 51924 40952
rect 52132 40938 52214 40952
rect 53090 40938 53172 40952
rect 53380 40938 53462 40952
rect 54338 40938 54420 40952
rect 54628 40938 54710 40952
rect 55586 40938 55668 40952
rect 55876 40938 55958 40952
rect 56834 40938 56916 40952
rect 57124 40938 57206 40952
rect 58082 40938 58164 40952
rect 58372 40938 58454 40952
rect 16418 40890 16864 40904
rect 17014 40890 17154 40904
rect 17304 40890 18112 40904
rect 18262 40890 18402 40904
rect 18552 40890 19360 40904
rect 19510 40890 19650 40904
rect 19800 40890 20608 40904
rect 20758 40890 20898 40904
rect 21048 40890 21856 40904
rect 22006 40890 22146 40904
rect 22296 40890 23104 40904
rect 23254 40890 23394 40904
rect 23544 40890 24352 40904
rect 24502 40890 24642 40904
rect 24792 40890 25600 40904
rect 25750 40890 25890 40904
rect 26040 40890 26848 40904
rect 26998 40890 27138 40904
rect 27288 40890 28096 40904
rect 28246 40890 28386 40904
rect 28536 40890 29344 40904
rect 29494 40890 29634 40904
rect 29784 40890 30592 40904
rect 30742 40890 30882 40904
rect 31032 40890 31840 40904
rect 31990 40890 32130 40904
rect 32280 40890 33088 40904
rect 33238 40890 33378 40904
rect 33528 40890 34336 40904
rect 34486 40890 34626 40904
rect 34776 40890 35584 40904
rect 35734 40890 35874 40904
rect 36024 40890 36832 40904
rect 36982 40890 37122 40904
rect 37272 40890 38080 40904
rect 38230 40890 38370 40904
rect 38520 40890 39328 40904
rect 39478 40890 39618 40904
rect 39768 40890 40576 40904
rect 40726 40890 40866 40904
rect 41016 40890 41824 40904
rect 41974 40890 42114 40904
rect 42264 40890 43072 40904
rect 43222 40890 43362 40904
rect 43512 40890 44320 40904
rect 44470 40890 44610 40904
rect 44760 40890 45568 40904
rect 45718 40890 45858 40904
rect 46008 40890 46816 40904
rect 46966 40890 47106 40904
rect 47256 40890 48064 40904
rect 48214 40890 48354 40904
rect 48504 40890 49312 40904
rect 49462 40890 49602 40904
rect 49752 40890 50560 40904
rect 50710 40890 50850 40904
rect 51000 40890 51808 40904
rect 51958 40890 52098 40904
rect 52248 40890 53056 40904
rect 53206 40890 53346 40904
rect 53496 40890 54304 40904
rect 54454 40890 54594 40904
rect 54744 40890 55552 40904
rect 55702 40890 55842 40904
rect 55992 40890 56800 40904
rect 56950 40890 57090 40904
rect 57240 40890 58048 40904
rect 58198 40890 58338 40904
rect 58488 40890 58934 40904
rect 16418 40842 58934 40890
rect 16418 40828 16864 40842
rect 17014 40828 17154 40842
rect 17304 40828 18112 40842
rect 18262 40828 18402 40842
rect 18552 40828 19360 40842
rect 19510 40828 19650 40842
rect 19800 40828 20608 40842
rect 20758 40828 20898 40842
rect 21048 40828 21856 40842
rect 22006 40828 22146 40842
rect 22296 40828 23104 40842
rect 23254 40828 23394 40842
rect 23544 40828 24352 40842
rect 24502 40828 24642 40842
rect 24792 40828 25600 40842
rect 25750 40828 25890 40842
rect 26040 40828 26848 40842
rect 26998 40828 27138 40842
rect 27288 40828 28096 40842
rect 28246 40828 28386 40842
rect 28536 40828 29344 40842
rect 29494 40828 29634 40842
rect 29784 40828 30592 40842
rect 30742 40828 30882 40842
rect 31032 40828 31840 40842
rect 31990 40828 32130 40842
rect 32280 40828 33088 40842
rect 33238 40828 33378 40842
rect 33528 40828 34336 40842
rect 34486 40828 34626 40842
rect 34776 40828 35584 40842
rect 35734 40828 35874 40842
rect 36024 40828 36832 40842
rect 36982 40828 37122 40842
rect 37272 40828 38080 40842
rect 38230 40828 38370 40842
rect 38520 40828 39328 40842
rect 39478 40828 39618 40842
rect 39768 40828 40576 40842
rect 40726 40828 40866 40842
rect 41016 40828 41824 40842
rect 41974 40828 42114 40842
rect 42264 40828 43072 40842
rect 43222 40828 43362 40842
rect 43512 40828 44320 40842
rect 44470 40828 44610 40842
rect 44760 40828 45568 40842
rect 45718 40828 45858 40842
rect 46008 40828 46816 40842
rect 46966 40828 47106 40842
rect 47256 40828 48064 40842
rect 48214 40828 48354 40842
rect 48504 40828 49312 40842
rect 49462 40828 49602 40842
rect 49752 40828 50560 40842
rect 50710 40828 50850 40842
rect 51000 40828 51808 40842
rect 51958 40828 52098 40842
rect 52248 40828 53056 40842
rect 53206 40828 53346 40842
rect 53496 40828 54304 40842
rect 54454 40828 54594 40842
rect 54744 40828 55552 40842
rect 55702 40828 55842 40842
rect 55992 40828 56800 40842
rect 56950 40828 57090 40842
rect 57240 40828 58048 40842
rect 58198 40828 58338 40842
rect 58488 40828 58934 40842
rect 16898 40780 16980 40794
rect 17188 40780 17270 40794
rect 18146 40780 18228 40794
rect 18436 40780 18518 40794
rect 19394 40780 19476 40794
rect 19684 40780 19766 40794
rect 20642 40780 20724 40794
rect 20932 40780 21014 40794
rect 21890 40780 21972 40794
rect 22180 40780 22262 40794
rect 23138 40780 23220 40794
rect 23428 40780 23510 40794
rect 24386 40780 24468 40794
rect 24676 40780 24758 40794
rect 25634 40780 25716 40794
rect 25924 40780 26006 40794
rect 26882 40780 26964 40794
rect 27172 40780 27254 40794
rect 28130 40780 28212 40794
rect 28420 40780 28502 40794
rect 29378 40780 29460 40794
rect 29668 40780 29750 40794
rect 30626 40780 30708 40794
rect 30916 40780 30998 40794
rect 31874 40780 31956 40794
rect 32164 40780 32246 40794
rect 33122 40780 33204 40794
rect 33412 40780 33494 40794
rect 34370 40780 34452 40794
rect 34660 40780 34742 40794
rect 35618 40780 35700 40794
rect 35908 40780 35990 40794
rect 36866 40780 36948 40794
rect 37156 40780 37238 40794
rect 38114 40780 38196 40794
rect 38404 40780 38486 40794
rect 39362 40780 39444 40794
rect 39652 40780 39734 40794
rect 40610 40780 40692 40794
rect 40900 40780 40982 40794
rect 41858 40780 41940 40794
rect 42148 40780 42230 40794
rect 43106 40780 43188 40794
rect 43396 40780 43478 40794
rect 44354 40780 44436 40794
rect 44644 40780 44726 40794
rect 45602 40780 45684 40794
rect 45892 40780 45974 40794
rect 46850 40780 46932 40794
rect 47140 40780 47222 40794
rect 48098 40780 48180 40794
rect 48388 40780 48470 40794
rect 49346 40780 49428 40794
rect 49636 40780 49718 40794
rect 50594 40780 50676 40794
rect 50884 40780 50966 40794
rect 51842 40780 51924 40794
rect 52132 40780 52214 40794
rect 53090 40780 53172 40794
rect 53380 40780 53462 40794
rect 54338 40780 54420 40794
rect 54628 40780 54710 40794
rect 55586 40780 55668 40794
rect 55876 40780 55958 40794
rect 56834 40780 56916 40794
rect 57124 40780 57206 40794
rect 58082 40780 58164 40794
rect 58372 40780 58454 40794
rect 16418 40732 58934 40780
rect 16418 40636 58934 40684
rect 16898 40622 16980 40636
rect 17188 40622 17270 40636
rect 18146 40622 18228 40636
rect 18436 40622 18518 40636
rect 19394 40622 19476 40636
rect 19684 40622 19766 40636
rect 20642 40622 20724 40636
rect 20932 40622 21014 40636
rect 21890 40622 21972 40636
rect 22180 40622 22262 40636
rect 23138 40622 23220 40636
rect 23428 40622 23510 40636
rect 24386 40622 24468 40636
rect 24676 40622 24758 40636
rect 25634 40622 25716 40636
rect 25924 40622 26006 40636
rect 26882 40622 26964 40636
rect 27172 40622 27254 40636
rect 28130 40622 28212 40636
rect 28420 40622 28502 40636
rect 29378 40622 29460 40636
rect 29668 40622 29750 40636
rect 30626 40622 30708 40636
rect 30916 40622 30998 40636
rect 31874 40622 31956 40636
rect 32164 40622 32246 40636
rect 33122 40622 33204 40636
rect 33412 40622 33494 40636
rect 34370 40622 34452 40636
rect 34660 40622 34742 40636
rect 35618 40622 35700 40636
rect 35908 40622 35990 40636
rect 36866 40622 36948 40636
rect 37156 40622 37238 40636
rect 38114 40622 38196 40636
rect 38404 40622 38486 40636
rect 39362 40622 39444 40636
rect 39652 40622 39734 40636
rect 40610 40622 40692 40636
rect 40900 40622 40982 40636
rect 41858 40622 41940 40636
rect 42148 40622 42230 40636
rect 43106 40622 43188 40636
rect 43396 40622 43478 40636
rect 44354 40622 44436 40636
rect 44644 40622 44726 40636
rect 45602 40622 45684 40636
rect 45892 40622 45974 40636
rect 46850 40622 46932 40636
rect 47140 40622 47222 40636
rect 48098 40622 48180 40636
rect 48388 40622 48470 40636
rect 49346 40622 49428 40636
rect 49636 40622 49718 40636
rect 50594 40622 50676 40636
rect 50884 40622 50966 40636
rect 51842 40622 51924 40636
rect 52132 40622 52214 40636
rect 53090 40622 53172 40636
rect 53380 40622 53462 40636
rect 54338 40622 54420 40636
rect 54628 40622 54710 40636
rect 55586 40622 55668 40636
rect 55876 40622 55958 40636
rect 56834 40622 56916 40636
rect 57124 40622 57206 40636
rect 58082 40622 58164 40636
rect 58372 40622 58454 40636
rect 16418 40574 16864 40588
rect 17014 40574 17154 40588
rect 17304 40574 18112 40588
rect 18262 40574 18402 40588
rect 18552 40574 19360 40588
rect 19510 40574 19650 40588
rect 19800 40574 20608 40588
rect 20758 40574 20898 40588
rect 21048 40574 21856 40588
rect 22006 40574 22146 40588
rect 22296 40574 23104 40588
rect 23254 40574 23394 40588
rect 23544 40574 24352 40588
rect 24502 40574 24642 40588
rect 24792 40574 25600 40588
rect 25750 40574 25890 40588
rect 26040 40574 26848 40588
rect 26998 40574 27138 40588
rect 27288 40574 28096 40588
rect 28246 40574 28386 40588
rect 28536 40574 29344 40588
rect 29494 40574 29634 40588
rect 29784 40574 30592 40588
rect 30742 40574 30882 40588
rect 31032 40574 31840 40588
rect 31990 40574 32130 40588
rect 32280 40574 33088 40588
rect 33238 40574 33378 40588
rect 33528 40574 34336 40588
rect 34486 40574 34626 40588
rect 34776 40574 35584 40588
rect 35734 40574 35874 40588
rect 36024 40574 36832 40588
rect 36982 40574 37122 40588
rect 37272 40574 38080 40588
rect 38230 40574 38370 40588
rect 38520 40574 39328 40588
rect 39478 40574 39618 40588
rect 39768 40574 40576 40588
rect 40726 40574 40866 40588
rect 41016 40574 41824 40588
rect 41974 40574 42114 40588
rect 42264 40574 43072 40588
rect 43222 40574 43362 40588
rect 43512 40574 44320 40588
rect 44470 40574 44610 40588
rect 44760 40574 45568 40588
rect 45718 40574 45858 40588
rect 46008 40574 46816 40588
rect 46966 40574 47106 40588
rect 47256 40574 48064 40588
rect 48214 40574 48354 40588
rect 48504 40574 49312 40588
rect 49462 40574 49602 40588
rect 49752 40574 50560 40588
rect 50710 40574 50850 40588
rect 51000 40574 51808 40588
rect 51958 40574 52098 40588
rect 52248 40574 53056 40588
rect 53206 40574 53346 40588
rect 53496 40574 54304 40588
rect 54454 40574 54594 40588
rect 54744 40574 55552 40588
rect 55702 40574 55842 40588
rect 55992 40574 56800 40588
rect 56950 40574 57090 40588
rect 57240 40574 58048 40588
rect 58198 40574 58338 40588
rect 58488 40574 58934 40588
rect 16418 40526 58934 40574
rect 16418 40512 16864 40526
rect 17014 40512 17154 40526
rect 17304 40512 18112 40526
rect 18262 40512 18402 40526
rect 18552 40512 19360 40526
rect 19510 40512 19650 40526
rect 19800 40512 20608 40526
rect 20758 40512 20898 40526
rect 21048 40512 21856 40526
rect 22006 40512 22146 40526
rect 22296 40512 23104 40526
rect 23254 40512 23394 40526
rect 23544 40512 24352 40526
rect 24502 40512 24642 40526
rect 24792 40512 25600 40526
rect 25750 40512 25890 40526
rect 26040 40512 26848 40526
rect 26998 40512 27138 40526
rect 27288 40512 28096 40526
rect 28246 40512 28386 40526
rect 28536 40512 29344 40526
rect 29494 40512 29634 40526
rect 29784 40512 30592 40526
rect 30742 40512 30882 40526
rect 31032 40512 31840 40526
rect 31990 40512 32130 40526
rect 32280 40512 33088 40526
rect 33238 40512 33378 40526
rect 33528 40512 34336 40526
rect 34486 40512 34626 40526
rect 34776 40512 35584 40526
rect 35734 40512 35874 40526
rect 36024 40512 36832 40526
rect 36982 40512 37122 40526
rect 37272 40512 38080 40526
rect 38230 40512 38370 40526
rect 38520 40512 39328 40526
rect 39478 40512 39618 40526
rect 39768 40512 40576 40526
rect 40726 40512 40866 40526
rect 41016 40512 41824 40526
rect 41974 40512 42114 40526
rect 42264 40512 43072 40526
rect 43222 40512 43362 40526
rect 43512 40512 44320 40526
rect 44470 40512 44610 40526
rect 44760 40512 45568 40526
rect 45718 40512 45858 40526
rect 46008 40512 46816 40526
rect 46966 40512 47106 40526
rect 47256 40512 48064 40526
rect 48214 40512 48354 40526
rect 48504 40512 49312 40526
rect 49462 40512 49602 40526
rect 49752 40512 50560 40526
rect 50710 40512 50850 40526
rect 51000 40512 51808 40526
rect 51958 40512 52098 40526
rect 52248 40512 53056 40526
rect 53206 40512 53346 40526
rect 53496 40512 54304 40526
rect 54454 40512 54594 40526
rect 54744 40512 55552 40526
rect 55702 40512 55842 40526
rect 55992 40512 56800 40526
rect 56950 40512 57090 40526
rect 57240 40512 58048 40526
rect 58198 40512 58338 40526
rect 58488 40512 58934 40526
rect 16898 40464 16980 40478
rect 17188 40464 17270 40478
rect 18146 40464 18228 40478
rect 18436 40464 18518 40478
rect 19394 40464 19476 40478
rect 19684 40464 19766 40478
rect 20642 40464 20724 40478
rect 20932 40464 21014 40478
rect 21890 40464 21972 40478
rect 22180 40464 22262 40478
rect 23138 40464 23220 40478
rect 23428 40464 23510 40478
rect 24386 40464 24468 40478
rect 24676 40464 24758 40478
rect 25634 40464 25716 40478
rect 25924 40464 26006 40478
rect 26882 40464 26964 40478
rect 27172 40464 27254 40478
rect 28130 40464 28212 40478
rect 28420 40464 28502 40478
rect 29378 40464 29460 40478
rect 29668 40464 29750 40478
rect 30626 40464 30708 40478
rect 30916 40464 30998 40478
rect 31874 40464 31956 40478
rect 32164 40464 32246 40478
rect 33122 40464 33204 40478
rect 33412 40464 33494 40478
rect 34370 40464 34452 40478
rect 34660 40464 34742 40478
rect 35618 40464 35700 40478
rect 35908 40464 35990 40478
rect 36866 40464 36948 40478
rect 37156 40464 37238 40478
rect 38114 40464 38196 40478
rect 38404 40464 38486 40478
rect 39362 40464 39444 40478
rect 39652 40464 39734 40478
rect 40610 40464 40692 40478
rect 40900 40464 40982 40478
rect 41858 40464 41940 40478
rect 42148 40464 42230 40478
rect 43106 40464 43188 40478
rect 43396 40464 43478 40478
rect 44354 40464 44436 40478
rect 44644 40464 44726 40478
rect 45602 40464 45684 40478
rect 45892 40464 45974 40478
rect 46850 40464 46932 40478
rect 47140 40464 47222 40478
rect 48098 40464 48180 40478
rect 48388 40464 48470 40478
rect 49346 40464 49428 40478
rect 49636 40464 49718 40478
rect 50594 40464 50676 40478
rect 50884 40464 50966 40478
rect 51842 40464 51924 40478
rect 52132 40464 52214 40478
rect 53090 40464 53172 40478
rect 53380 40464 53462 40478
rect 54338 40464 54420 40478
rect 54628 40464 54710 40478
rect 55586 40464 55668 40478
rect 55876 40464 55958 40478
rect 56834 40464 56916 40478
rect 57124 40464 57206 40478
rect 58082 40464 58164 40478
rect 58372 40464 58454 40478
rect 16418 40416 58934 40464
rect 16418 40258 58934 40368
rect 16418 40162 58934 40210
rect 16898 40148 16980 40162
rect 17188 40148 17270 40162
rect 18146 40148 18228 40162
rect 18436 40148 18518 40162
rect 19394 40148 19476 40162
rect 19684 40148 19766 40162
rect 20642 40148 20724 40162
rect 20932 40148 21014 40162
rect 21890 40148 21972 40162
rect 22180 40148 22262 40162
rect 23138 40148 23220 40162
rect 23428 40148 23510 40162
rect 24386 40148 24468 40162
rect 24676 40148 24758 40162
rect 25634 40148 25716 40162
rect 25924 40148 26006 40162
rect 26882 40148 26964 40162
rect 27172 40148 27254 40162
rect 28130 40148 28212 40162
rect 28420 40148 28502 40162
rect 29378 40148 29460 40162
rect 29668 40148 29750 40162
rect 30626 40148 30708 40162
rect 30916 40148 30998 40162
rect 31874 40148 31956 40162
rect 32164 40148 32246 40162
rect 33122 40148 33204 40162
rect 33412 40148 33494 40162
rect 34370 40148 34452 40162
rect 34660 40148 34742 40162
rect 35618 40148 35700 40162
rect 35908 40148 35990 40162
rect 36866 40148 36948 40162
rect 37156 40148 37238 40162
rect 38114 40148 38196 40162
rect 38404 40148 38486 40162
rect 39362 40148 39444 40162
rect 39652 40148 39734 40162
rect 40610 40148 40692 40162
rect 40900 40148 40982 40162
rect 41858 40148 41940 40162
rect 42148 40148 42230 40162
rect 43106 40148 43188 40162
rect 43396 40148 43478 40162
rect 44354 40148 44436 40162
rect 44644 40148 44726 40162
rect 45602 40148 45684 40162
rect 45892 40148 45974 40162
rect 46850 40148 46932 40162
rect 47140 40148 47222 40162
rect 48098 40148 48180 40162
rect 48388 40148 48470 40162
rect 49346 40148 49428 40162
rect 49636 40148 49718 40162
rect 50594 40148 50676 40162
rect 50884 40148 50966 40162
rect 51842 40148 51924 40162
rect 52132 40148 52214 40162
rect 53090 40148 53172 40162
rect 53380 40148 53462 40162
rect 54338 40148 54420 40162
rect 54628 40148 54710 40162
rect 55586 40148 55668 40162
rect 55876 40148 55958 40162
rect 56834 40148 56916 40162
rect 57124 40148 57206 40162
rect 58082 40148 58164 40162
rect 58372 40148 58454 40162
rect 16418 40100 16864 40114
rect 17014 40100 17154 40114
rect 17304 40100 18112 40114
rect 18262 40100 18402 40114
rect 18552 40100 19360 40114
rect 19510 40100 19650 40114
rect 19800 40100 20608 40114
rect 20758 40100 20898 40114
rect 21048 40100 21856 40114
rect 22006 40100 22146 40114
rect 22296 40100 23104 40114
rect 23254 40100 23394 40114
rect 23544 40100 24352 40114
rect 24502 40100 24642 40114
rect 24792 40100 25600 40114
rect 25750 40100 25890 40114
rect 26040 40100 26848 40114
rect 26998 40100 27138 40114
rect 27288 40100 28096 40114
rect 28246 40100 28386 40114
rect 28536 40100 29344 40114
rect 29494 40100 29634 40114
rect 29784 40100 30592 40114
rect 30742 40100 30882 40114
rect 31032 40100 31840 40114
rect 31990 40100 32130 40114
rect 32280 40100 33088 40114
rect 33238 40100 33378 40114
rect 33528 40100 34336 40114
rect 34486 40100 34626 40114
rect 34776 40100 35584 40114
rect 35734 40100 35874 40114
rect 36024 40100 36832 40114
rect 36982 40100 37122 40114
rect 37272 40100 38080 40114
rect 38230 40100 38370 40114
rect 38520 40100 39328 40114
rect 39478 40100 39618 40114
rect 39768 40100 40576 40114
rect 40726 40100 40866 40114
rect 41016 40100 41824 40114
rect 41974 40100 42114 40114
rect 42264 40100 43072 40114
rect 43222 40100 43362 40114
rect 43512 40100 44320 40114
rect 44470 40100 44610 40114
rect 44760 40100 45568 40114
rect 45718 40100 45858 40114
rect 46008 40100 46816 40114
rect 46966 40100 47106 40114
rect 47256 40100 48064 40114
rect 48214 40100 48354 40114
rect 48504 40100 49312 40114
rect 49462 40100 49602 40114
rect 49752 40100 50560 40114
rect 50710 40100 50850 40114
rect 51000 40100 51808 40114
rect 51958 40100 52098 40114
rect 52248 40100 53056 40114
rect 53206 40100 53346 40114
rect 53496 40100 54304 40114
rect 54454 40100 54594 40114
rect 54744 40100 55552 40114
rect 55702 40100 55842 40114
rect 55992 40100 56800 40114
rect 56950 40100 57090 40114
rect 57240 40100 58048 40114
rect 58198 40100 58338 40114
rect 58488 40100 58934 40114
rect 16418 40052 58934 40100
rect 16418 40038 16864 40052
rect 17014 40038 17154 40052
rect 17304 40038 18112 40052
rect 18262 40038 18402 40052
rect 18552 40038 19360 40052
rect 19510 40038 19650 40052
rect 19800 40038 20608 40052
rect 20758 40038 20898 40052
rect 21048 40038 21856 40052
rect 22006 40038 22146 40052
rect 22296 40038 23104 40052
rect 23254 40038 23394 40052
rect 23544 40038 24352 40052
rect 24502 40038 24642 40052
rect 24792 40038 25600 40052
rect 25750 40038 25890 40052
rect 26040 40038 26848 40052
rect 26998 40038 27138 40052
rect 27288 40038 28096 40052
rect 28246 40038 28386 40052
rect 28536 40038 29344 40052
rect 29494 40038 29634 40052
rect 29784 40038 30592 40052
rect 30742 40038 30882 40052
rect 31032 40038 31840 40052
rect 31990 40038 32130 40052
rect 32280 40038 33088 40052
rect 33238 40038 33378 40052
rect 33528 40038 34336 40052
rect 34486 40038 34626 40052
rect 34776 40038 35584 40052
rect 35734 40038 35874 40052
rect 36024 40038 36832 40052
rect 36982 40038 37122 40052
rect 37272 40038 38080 40052
rect 38230 40038 38370 40052
rect 38520 40038 39328 40052
rect 39478 40038 39618 40052
rect 39768 40038 40576 40052
rect 40726 40038 40866 40052
rect 41016 40038 41824 40052
rect 41974 40038 42114 40052
rect 42264 40038 43072 40052
rect 43222 40038 43362 40052
rect 43512 40038 44320 40052
rect 44470 40038 44610 40052
rect 44760 40038 45568 40052
rect 45718 40038 45858 40052
rect 46008 40038 46816 40052
rect 46966 40038 47106 40052
rect 47256 40038 48064 40052
rect 48214 40038 48354 40052
rect 48504 40038 49312 40052
rect 49462 40038 49602 40052
rect 49752 40038 50560 40052
rect 50710 40038 50850 40052
rect 51000 40038 51808 40052
rect 51958 40038 52098 40052
rect 52248 40038 53056 40052
rect 53206 40038 53346 40052
rect 53496 40038 54304 40052
rect 54454 40038 54594 40052
rect 54744 40038 55552 40052
rect 55702 40038 55842 40052
rect 55992 40038 56800 40052
rect 56950 40038 57090 40052
rect 57240 40038 58048 40052
rect 58198 40038 58338 40052
rect 58488 40038 58934 40052
rect 16898 39990 16980 40004
rect 17188 39990 17270 40004
rect 18146 39990 18228 40004
rect 18436 39990 18518 40004
rect 19394 39990 19476 40004
rect 19684 39990 19766 40004
rect 20642 39990 20724 40004
rect 20932 39990 21014 40004
rect 21890 39990 21972 40004
rect 22180 39990 22262 40004
rect 23138 39990 23220 40004
rect 23428 39990 23510 40004
rect 24386 39990 24468 40004
rect 24676 39990 24758 40004
rect 25634 39990 25716 40004
rect 25924 39990 26006 40004
rect 26882 39990 26964 40004
rect 27172 39990 27254 40004
rect 28130 39990 28212 40004
rect 28420 39990 28502 40004
rect 29378 39990 29460 40004
rect 29668 39990 29750 40004
rect 30626 39990 30708 40004
rect 30916 39990 30998 40004
rect 31874 39990 31956 40004
rect 32164 39990 32246 40004
rect 33122 39990 33204 40004
rect 33412 39990 33494 40004
rect 34370 39990 34452 40004
rect 34660 39990 34742 40004
rect 35618 39990 35700 40004
rect 35908 39990 35990 40004
rect 36866 39990 36948 40004
rect 37156 39990 37238 40004
rect 38114 39990 38196 40004
rect 38404 39990 38486 40004
rect 39362 39990 39444 40004
rect 39652 39990 39734 40004
rect 40610 39990 40692 40004
rect 40900 39990 40982 40004
rect 41858 39990 41940 40004
rect 42148 39990 42230 40004
rect 43106 39990 43188 40004
rect 43396 39990 43478 40004
rect 44354 39990 44436 40004
rect 44644 39990 44726 40004
rect 45602 39990 45684 40004
rect 45892 39990 45974 40004
rect 46850 39990 46932 40004
rect 47140 39990 47222 40004
rect 48098 39990 48180 40004
rect 48388 39990 48470 40004
rect 49346 39990 49428 40004
rect 49636 39990 49718 40004
rect 50594 39990 50676 40004
rect 50884 39990 50966 40004
rect 51842 39990 51924 40004
rect 52132 39990 52214 40004
rect 53090 39990 53172 40004
rect 53380 39990 53462 40004
rect 54338 39990 54420 40004
rect 54628 39990 54710 40004
rect 55586 39990 55668 40004
rect 55876 39990 55958 40004
rect 56834 39990 56916 40004
rect 57124 39990 57206 40004
rect 58082 39990 58164 40004
rect 58372 39990 58454 40004
rect 16418 39942 58934 39990
rect 16418 39846 58934 39894
rect 16898 39832 16980 39846
rect 17188 39832 17270 39846
rect 18146 39832 18228 39846
rect 18436 39832 18518 39846
rect 19394 39832 19476 39846
rect 19684 39832 19766 39846
rect 20642 39832 20724 39846
rect 20932 39832 21014 39846
rect 21890 39832 21972 39846
rect 22180 39832 22262 39846
rect 23138 39832 23220 39846
rect 23428 39832 23510 39846
rect 24386 39832 24468 39846
rect 24676 39832 24758 39846
rect 25634 39832 25716 39846
rect 25924 39832 26006 39846
rect 26882 39832 26964 39846
rect 27172 39832 27254 39846
rect 28130 39832 28212 39846
rect 28420 39832 28502 39846
rect 29378 39832 29460 39846
rect 29668 39832 29750 39846
rect 30626 39832 30708 39846
rect 30916 39832 30998 39846
rect 31874 39832 31956 39846
rect 32164 39832 32246 39846
rect 33122 39832 33204 39846
rect 33412 39832 33494 39846
rect 34370 39832 34452 39846
rect 34660 39832 34742 39846
rect 35618 39832 35700 39846
rect 35908 39832 35990 39846
rect 36866 39832 36948 39846
rect 37156 39832 37238 39846
rect 38114 39832 38196 39846
rect 38404 39832 38486 39846
rect 39362 39832 39444 39846
rect 39652 39832 39734 39846
rect 40610 39832 40692 39846
rect 40900 39832 40982 39846
rect 41858 39832 41940 39846
rect 42148 39832 42230 39846
rect 43106 39832 43188 39846
rect 43396 39832 43478 39846
rect 44354 39832 44436 39846
rect 44644 39832 44726 39846
rect 45602 39832 45684 39846
rect 45892 39832 45974 39846
rect 46850 39832 46932 39846
rect 47140 39832 47222 39846
rect 48098 39832 48180 39846
rect 48388 39832 48470 39846
rect 49346 39832 49428 39846
rect 49636 39832 49718 39846
rect 50594 39832 50676 39846
rect 50884 39832 50966 39846
rect 51842 39832 51924 39846
rect 52132 39832 52214 39846
rect 53090 39832 53172 39846
rect 53380 39832 53462 39846
rect 54338 39832 54420 39846
rect 54628 39832 54710 39846
rect 55586 39832 55668 39846
rect 55876 39832 55958 39846
rect 56834 39832 56916 39846
rect 57124 39832 57206 39846
rect 58082 39832 58164 39846
rect 58372 39832 58454 39846
rect 16418 39784 16864 39798
rect 17014 39784 17154 39798
rect 17304 39784 18112 39798
rect 18262 39784 18402 39798
rect 18552 39784 19360 39798
rect 19510 39784 19650 39798
rect 19800 39784 20608 39798
rect 20758 39784 20898 39798
rect 21048 39784 21856 39798
rect 22006 39784 22146 39798
rect 22296 39784 23104 39798
rect 23254 39784 23394 39798
rect 23544 39784 24352 39798
rect 24502 39784 24642 39798
rect 24792 39784 25600 39798
rect 25750 39784 25890 39798
rect 26040 39784 26848 39798
rect 26998 39784 27138 39798
rect 27288 39784 28096 39798
rect 28246 39784 28386 39798
rect 28536 39784 29344 39798
rect 29494 39784 29634 39798
rect 29784 39784 30592 39798
rect 30742 39784 30882 39798
rect 31032 39784 31840 39798
rect 31990 39784 32130 39798
rect 32280 39784 33088 39798
rect 33238 39784 33378 39798
rect 33528 39784 34336 39798
rect 34486 39784 34626 39798
rect 34776 39784 35584 39798
rect 35734 39784 35874 39798
rect 36024 39784 36832 39798
rect 36982 39784 37122 39798
rect 37272 39784 38080 39798
rect 38230 39784 38370 39798
rect 38520 39784 39328 39798
rect 39478 39784 39618 39798
rect 39768 39784 40576 39798
rect 40726 39784 40866 39798
rect 41016 39784 41824 39798
rect 41974 39784 42114 39798
rect 42264 39784 43072 39798
rect 43222 39784 43362 39798
rect 43512 39784 44320 39798
rect 44470 39784 44610 39798
rect 44760 39784 45568 39798
rect 45718 39784 45858 39798
rect 46008 39784 46816 39798
rect 46966 39784 47106 39798
rect 47256 39784 48064 39798
rect 48214 39784 48354 39798
rect 48504 39784 49312 39798
rect 49462 39784 49602 39798
rect 49752 39784 50560 39798
rect 50710 39784 50850 39798
rect 51000 39784 51808 39798
rect 51958 39784 52098 39798
rect 52248 39784 53056 39798
rect 53206 39784 53346 39798
rect 53496 39784 54304 39798
rect 54454 39784 54594 39798
rect 54744 39784 55552 39798
rect 55702 39784 55842 39798
rect 55992 39784 56800 39798
rect 56950 39784 57090 39798
rect 57240 39784 58048 39798
rect 58198 39784 58338 39798
rect 58488 39784 58934 39798
rect 16418 39736 58934 39784
rect 16418 39722 16864 39736
rect 17014 39722 17154 39736
rect 17304 39722 18112 39736
rect 18262 39722 18402 39736
rect 18552 39722 19360 39736
rect 19510 39722 19650 39736
rect 19800 39722 20608 39736
rect 20758 39722 20898 39736
rect 21048 39722 21856 39736
rect 22006 39722 22146 39736
rect 22296 39722 23104 39736
rect 23254 39722 23394 39736
rect 23544 39722 24352 39736
rect 24502 39722 24642 39736
rect 24792 39722 25600 39736
rect 25750 39722 25890 39736
rect 26040 39722 26848 39736
rect 26998 39722 27138 39736
rect 27288 39722 28096 39736
rect 28246 39722 28386 39736
rect 28536 39722 29344 39736
rect 29494 39722 29634 39736
rect 29784 39722 30592 39736
rect 30742 39722 30882 39736
rect 31032 39722 31840 39736
rect 31990 39722 32130 39736
rect 32280 39722 33088 39736
rect 33238 39722 33378 39736
rect 33528 39722 34336 39736
rect 34486 39722 34626 39736
rect 34776 39722 35584 39736
rect 35734 39722 35874 39736
rect 36024 39722 36832 39736
rect 36982 39722 37122 39736
rect 37272 39722 38080 39736
rect 38230 39722 38370 39736
rect 38520 39722 39328 39736
rect 39478 39722 39618 39736
rect 39768 39722 40576 39736
rect 40726 39722 40866 39736
rect 41016 39722 41824 39736
rect 41974 39722 42114 39736
rect 42264 39722 43072 39736
rect 43222 39722 43362 39736
rect 43512 39722 44320 39736
rect 44470 39722 44610 39736
rect 44760 39722 45568 39736
rect 45718 39722 45858 39736
rect 46008 39722 46816 39736
rect 46966 39722 47106 39736
rect 47256 39722 48064 39736
rect 48214 39722 48354 39736
rect 48504 39722 49312 39736
rect 49462 39722 49602 39736
rect 49752 39722 50560 39736
rect 50710 39722 50850 39736
rect 51000 39722 51808 39736
rect 51958 39722 52098 39736
rect 52248 39722 53056 39736
rect 53206 39722 53346 39736
rect 53496 39722 54304 39736
rect 54454 39722 54594 39736
rect 54744 39722 55552 39736
rect 55702 39722 55842 39736
rect 55992 39722 56800 39736
rect 56950 39722 57090 39736
rect 57240 39722 58048 39736
rect 58198 39722 58338 39736
rect 58488 39722 58934 39736
rect 16898 39674 16980 39688
rect 17188 39674 17270 39688
rect 18146 39674 18228 39688
rect 18436 39674 18518 39688
rect 19394 39674 19476 39688
rect 19684 39674 19766 39688
rect 20642 39674 20724 39688
rect 20932 39674 21014 39688
rect 21890 39674 21972 39688
rect 22180 39674 22262 39688
rect 23138 39674 23220 39688
rect 23428 39674 23510 39688
rect 24386 39674 24468 39688
rect 24676 39674 24758 39688
rect 25634 39674 25716 39688
rect 25924 39674 26006 39688
rect 26882 39674 26964 39688
rect 27172 39674 27254 39688
rect 28130 39674 28212 39688
rect 28420 39674 28502 39688
rect 29378 39674 29460 39688
rect 29668 39674 29750 39688
rect 30626 39674 30708 39688
rect 30916 39674 30998 39688
rect 31874 39674 31956 39688
rect 32164 39674 32246 39688
rect 33122 39674 33204 39688
rect 33412 39674 33494 39688
rect 34370 39674 34452 39688
rect 34660 39674 34742 39688
rect 35618 39674 35700 39688
rect 35908 39674 35990 39688
rect 36866 39674 36948 39688
rect 37156 39674 37238 39688
rect 38114 39674 38196 39688
rect 38404 39674 38486 39688
rect 39362 39674 39444 39688
rect 39652 39674 39734 39688
rect 40610 39674 40692 39688
rect 40900 39674 40982 39688
rect 41858 39674 41940 39688
rect 42148 39674 42230 39688
rect 43106 39674 43188 39688
rect 43396 39674 43478 39688
rect 44354 39674 44436 39688
rect 44644 39674 44726 39688
rect 45602 39674 45684 39688
rect 45892 39674 45974 39688
rect 46850 39674 46932 39688
rect 47140 39674 47222 39688
rect 48098 39674 48180 39688
rect 48388 39674 48470 39688
rect 49346 39674 49428 39688
rect 49636 39674 49718 39688
rect 50594 39674 50676 39688
rect 50884 39674 50966 39688
rect 51842 39674 51924 39688
rect 52132 39674 52214 39688
rect 53090 39674 53172 39688
rect 53380 39674 53462 39688
rect 54338 39674 54420 39688
rect 54628 39674 54710 39688
rect 55586 39674 55668 39688
rect 55876 39674 55958 39688
rect 56834 39674 56916 39688
rect 57124 39674 57206 39688
rect 58082 39674 58164 39688
rect 58372 39674 58454 39688
rect 16418 39626 58934 39674
rect 16418 39468 58934 39578
rect 16418 39372 58934 39420
rect 16898 39358 16980 39372
rect 17188 39358 17270 39372
rect 18146 39358 18228 39372
rect 18436 39358 18518 39372
rect 19394 39358 19476 39372
rect 19684 39358 19766 39372
rect 20642 39358 20724 39372
rect 20932 39358 21014 39372
rect 21890 39358 21972 39372
rect 22180 39358 22262 39372
rect 23138 39358 23220 39372
rect 23428 39358 23510 39372
rect 24386 39358 24468 39372
rect 24676 39358 24758 39372
rect 25634 39358 25716 39372
rect 25924 39358 26006 39372
rect 26882 39358 26964 39372
rect 27172 39358 27254 39372
rect 28130 39358 28212 39372
rect 28420 39358 28502 39372
rect 29378 39358 29460 39372
rect 29668 39358 29750 39372
rect 30626 39358 30708 39372
rect 30916 39358 30998 39372
rect 31874 39358 31956 39372
rect 32164 39358 32246 39372
rect 33122 39358 33204 39372
rect 33412 39358 33494 39372
rect 34370 39358 34452 39372
rect 34660 39358 34742 39372
rect 35618 39358 35700 39372
rect 35908 39358 35990 39372
rect 36866 39358 36948 39372
rect 37156 39358 37238 39372
rect 38114 39358 38196 39372
rect 38404 39358 38486 39372
rect 39362 39358 39444 39372
rect 39652 39358 39734 39372
rect 40610 39358 40692 39372
rect 40900 39358 40982 39372
rect 41858 39358 41940 39372
rect 42148 39358 42230 39372
rect 43106 39358 43188 39372
rect 43396 39358 43478 39372
rect 44354 39358 44436 39372
rect 44644 39358 44726 39372
rect 45602 39358 45684 39372
rect 45892 39358 45974 39372
rect 46850 39358 46932 39372
rect 47140 39358 47222 39372
rect 48098 39358 48180 39372
rect 48388 39358 48470 39372
rect 49346 39358 49428 39372
rect 49636 39358 49718 39372
rect 50594 39358 50676 39372
rect 50884 39358 50966 39372
rect 51842 39358 51924 39372
rect 52132 39358 52214 39372
rect 53090 39358 53172 39372
rect 53380 39358 53462 39372
rect 54338 39358 54420 39372
rect 54628 39358 54710 39372
rect 55586 39358 55668 39372
rect 55876 39358 55958 39372
rect 56834 39358 56916 39372
rect 57124 39358 57206 39372
rect 58082 39358 58164 39372
rect 58372 39358 58454 39372
rect 16418 39310 16864 39324
rect 17014 39310 17154 39324
rect 17304 39310 18112 39324
rect 18262 39310 18402 39324
rect 18552 39310 19360 39324
rect 19510 39310 19650 39324
rect 19800 39310 20608 39324
rect 20758 39310 20898 39324
rect 21048 39310 21856 39324
rect 22006 39310 22146 39324
rect 22296 39310 23104 39324
rect 23254 39310 23394 39324
rect 23544 39310 24352 39324
rect 24502 39310 24642 39324
rect 24792 39310 25600 39324
rect 25750 39310 25890 39324
rect 26040 39310 26848 39324
rect 26998 39310 27138 39324
rect 27288 39310 28096 39324
rect 28246 39310 28386 39324
rect 28536 39310 29344 39324
rect 29494 39310 29634 39324
rect 29784 39310 30592 39324
rect 30742 39310 30882 39324
rect 31032 39310 31840 39324
rect 31990 39310 32130 39324
rect 32280 39310 33088 39324
rect 33238 39310 33378 39324
rect 33528 39310 34336 39324
rect 34486 39310 34626 39324
rect 34776 39310 35584 39324
rect 35734 39310 35874 39324
rect 36024 39310 36832 39324
rect 36982 39310 37122 39324
rect 37272 39310 38080 39324
rect 38230 39310 38370 39324
rect 38520 39310 39328 39324
rect 39478 39310 39618 39324
rect 39768 39310 40576 39324
rect 40726 39310 40866 39324
rect 41016 39310 41824 39324
rect 41974 39310 42114 39324
rect 42264 39310 43072 39324
rect 43222 39310 43362 39324
rect 43512 39310 44320 39324
rect 44470 39310 44610 39324
rect 44760 39310 45568 39324
rect 45718 39310 45858 39324
rect 46008 39310 46816 39324
rect 46966 39310 47106 39324
rect 47256 39310 48064 39324
rect 48214 39310 48354 39324
rect 48504 39310 49312 39324
rect 49462 39310 49602 39324
rect 49752 39310 50560 39324
rect 50710 39310 50850 39324
rect 51000 39310 51808 39324
rect 51958 39310 52098 39324
rect 52248 39310 53056 39324
rect 53206 39310 53346 39324
rect 53496 39310 54304 39324
rect 54454 39310 54594 39324
rect 54744 39310 55552 39324
rect 55702 39310 55842 39324
rect 55992 39310 56800 39324
rect 56950 39310 57090 39324
rect 57240 39310 58048 39324
rect 58198 39310 58338 39324
rect 58488 39310 58934 39324
rect 16418 39262 58934 39310
rect 16418 39248 16864 39262
rect 17014 39248 17154 39262
rect 17304 39248 18112 39262
rect 18262 39248 18402 39262
rect 18552 39248 19360 39262
rect 19510 39248 19650 39262
rect 19800 39248 20608 39262
rect 20758 39248 20898 39262
rect 21048 39248 21856 39262
rect 22006 39248 22146 39262
rect 22296 39248 23104 39262
rect 23254 39248 23394 39262
rect 23544 39248 24352 39262
rect 24502 39248 24642 39262
rect 24792 39248 25600 39262
rect 25750 39248 25890 39262
rect 26040 39248 26848 39262
rect 26998 39248 27138 39262
rect 27288 39248 28096 39262
rect 28246 39248 28386 39262
rect 28536 39248 29344 39262
rect 29494 39248 29634 39262
rect 29784 39248 30592 39262
rect 30742 39248 30882 39262
rect 31032 39248 31840 39262
rect 31990 39248 32130 39262
rect 32280 39248 33088 39262
rect 33238 39248 33378 39262
rect 33528 39248 34336 39262
rect 34486 39248 34626 39262
rect 34776 39248 35584 39262
rect 35734 39248 35874 39262
rect 36024 39248 36832 39262
rect 36982 39248 37122 39262
rect 37272 39248 38080 39262
rect 38230 39248 38370 39262
rect 38520 39248 39328 39262
rect 39478 39248 39618 39262
rect 39768 39248 40576 39262
rect 40726 39248 40866 39262
rect 41016 39248 41824 39262
rect 41974 39248 42114 39262
rect 42264 39248 43072 39262
rect 43222 39248 43362 39262
rect 43512 39248 44320 39262
rect 44470 39248 44610 39262
rect 44760 39248 45568 39262
rect 45718 39248 45858 39262
rect 46008 39248 46816 39262
rect 46966 39248 47106 39262
rect 47256 39248 48064 39262
rect 48214 39248 48354 39262
rect 48504 39248 49312 39262
rect 49462 39248 49602 39262
rect 49752 39248 50560 39262
rect 50710 39248 50850 39262
rect 51000 39248 51808 39262
rect 51958 39248 52098 39262
rect 52248 39248 53056 39262
rect 53206 39248 53346 39262
rect 53496 39248 54304 39262
rect 54454 39248 54594 39262
rect 54744 39248 55552 39262
rect 55702 39248 55842 39262
rect 55992 39248 56800 39262
rect 56950 39248 57090 39262
rect 57240 39248 58048 39262
rect 58198 39248 58338 39262
rect 58488 39248 58934 39262
rect 16898 39200 16980 39214
rect 17188 39200 17270 39214
rect 18146 39200 18228 39214
rect 18436 39200 18518 39214
rect 19394 39200 19476 39214
rect 19684 39200 19766 39214
rect 20642 39200 20724 39214
rect 20932 39200 21014 39214
rect 21890 39200 21972 39214
rect 22180 39200 22262 39214
rect 23138 39200 23220 39214
rect 23428 39200 23510 39214
rect 24386 39200 24468 39214
rect 24676 39200 24758 39214
rect 25634 39200 25716 39214
rect 25924 39200 26006 39214
rect 26882 39200 26964 39214
rect 27172 39200 27254 39214
rect 28130 39200 28212 39214
rect 28420 39200 28502 39214
rect 29378 39200 29460 39214
rect 29668 39200 29750 39214
rect 30626 39200 30708 39214
rect 30916 39200 30998 39214
rect 31874 39200 31956 39214
rect 32164 39200 32246 39214
rect 33122 39200 33204 39214
rect 33412 39200 33494 39214
rect 34370 39200 34452 39214
rect 34660 39200 34742 39214
rect 35618 39200 35700 39214
rect 35908 39200 35990 39214
rect 36866 39200 36948 39214
rect 37156 39200 37238 39214
rect 38114 39200 38196 39214
rect 38404 39200 38486 39214
rect 39362 39200 39444 39214
rect 39652 39200 39734 39214
rect 40610 39200 40692 39214
rect 40900 39200 40982 39214
rect 41858 39200 41940 39214
rect 42148 39200 42230 39214
rect 43106 39200 43188 39214
rect 43396 39200 43478 39214
rect 44354 39200 44436 39214
rect 44644 39200 44726 39214
rect 45602 39200 45684 39214
rect 45892 39200 45974 39214
rect 46850 39200 46932 39214
rect 47140 39200 47222 39214
rect 48098 39200 48180 39214
rect 48388 39200 48470 39214
rect 49346 39200 49428 39214
rect 49636 39200 49718 39214
rect 50594 39200 50676 39214
rect 50884 39200 50966 39214
rect 51842 39200 51924 39214
rect 52132 39200 52214 39214
rect 53090 39200 53172 39214
rect 53380 39200 53462 39214
rect 54338 39200 54420 39214
rect 54628 39200 54710 39214
rect 55586 39200 55668 39214
rect 55876 39200 55958 39214
rect 56834 39200 56916 39214
rect 57124 39200 57206 39214
rect 58082 39200 58164 39214
rect 58372 39200 58454 39214
rect 16418 39152 58934 39200
rect 16418 39056 58934 39104
rect 16898 39042 16980 39056
rect 17188 39042 17270 39056
rect 18146 39042 18228 39056
rect 18436 39042 18518 39056
rect 19394 39042 19476 39056
rect 19684 39042 19766 39056
rect 20642 39042 20724 39056
rect 20932 39042 21014 39056
rect 21890 39042 21972 39056
rect 22180 39042 22262 39056
rect 23138 39042 23220 39056
rect 23428 39042 23510 39056
rect 24386 39042 24468 39056
rect 24676 39042 24758 39056
rect 25634 39042 25716 39056
rect 25924 39042 26006 39056
rect 26882 39042 26964 39056
rect 27172 39042 27254 39056
rect 28130 39042 28212 39056
rect 28420 39042 28502 39056
rect 29378 39042 29460 39056
rect 29668 39042 29750 39056
rect 30626 39042 30708 39056
rect 30916 39042 30998 39056
rect 31874 39042 31956 39056
rect 32164 39042 32246 39056
rect 33122 39042 33204 39056
rect 33412 39042 33494 39056
rect 34370 39042 34452 39056
rect 34660 39042 34742 39056
rect 35618 39042 35700 39056
rect 35908 39042 35990 39056
rect 36866 39042 36948 39056
rect 37156 39042 37238 39056
rect 38114 39042 38196 39056
rect 38404 39042 38486 39056
rect 39362 39042 39444 39056
rect 39652 39042 39734 39056
rect 40610 39042 40692 39056
rect 40900 39042 40982 39056
rect 41858 39042 41940 39056
rect 42148 39042 42230 39056
rect 43106 39042 43188 39056
rect 43396 39042 43478 39056
rect 44354 39042 44436 39056
rect 44644 39042 44726 39056
rect 45602 39042 45684 39056
rect 45892 39042 45974 39056
rect 46850 39042 46932 39056
rect 47140 39042 47222 39056
rect 48098 39042 48180 39056
rect 48388 39042 48470 39056
rect 49346 39042 49428 39056
rect 49636 39042 49718 39056
rect 50594 39042 50676 39056
rect 50884 39042 50966 39056
rect 51842 39042 51924 39056
rect 52132 39042 52214 39056
rect 53090 39042 53172 39056
rect 53380 39042 53462 39056
rect 54338 39042 54420 39056
rect 54628 39042 54710 39056
rect 55586 39042 55668 39056
rect 55876 39042 55958 39056
rect 56834 39042 56916 39056
rect 57124 39042 57206 39056
rect 58082 39042 58164 39056
rect 58372 39042 58454 39056
rect 16418 38994 16864 39008
rect 17014 38994 17154 39008
rect 17304 38994 18112 39008
rect 18262 38994 18402 39008
rect 18552 38994 19360 39008
rect 19510 38994 19650 39008
rect 19800 38994 20608 39008
rect 20758 38994 20898 39008
rect 21048 38994 21856 39008
rect 22006 38994 22146 39008
rect 22296 38994 23104 39008
rect 23254 38994 23394 39008
rect 23544 38994 24352 39008
rect 24502 38994 24642 39008
rect 24792 38994 25600 39008
rect 25750 38994 25890 39008
rect 26040 38994 26848 39008
rect 26998 38994 27138 39008
rect 27288 38994 28096 39008
rect 28246 38994 28386 39008
rect 28536 38994 29344 39008
rect 29494 38994 29634 39008
rect 29784 38994 30592 39008
rect 30742 38994 30882 39008
rect 31032 38994 31840 39008
rect 31990 38994 32130 39008
rect 32280 38994 33088 39008
rect 33238 38994 33378 39008
rect 33528 38994 34336 39008
rect 34486 38994 34626 39008
rect 34776 38994 35584 39008
rect 35734 38994 35874 39008
rect 36024 38994 36832 39008
rect 36982 38994 37122 39008
rect 37272 38994 38080 39008
rect 38230 38994 38370 39008
rect 38520 38994 39328 39008
rect 39478 38994 39618 39008
rect 39768 38994 40576 39008
rect 40726 38994 40866 39008
rect 41016 38994 41824 39008
rect 41974 38994 42114 39008
rect 42264 38994 43072 39008
rect 43222 38994 43362 39008
rect 43512 38994 44320 39008
rect 44470 38994 44610 39008
rect 44760 38994 45568 39008
rect 45718 38994 45858 39008
rect 46008 38994 46816 39008
rect 46966 38994 47106 39008
rect 47256 38994 48064 39008
rect 48214 38994 48354 39008
rect 48504 38994 49312 39008
rect 49462 38994 49602 39008
rect 49752 38994 50560 39008
rect 50710 38994 50850 39008
rect 51000 38994 51808 39008
rect 51958 38994 52098 39008
rect 52248 38994 53056 39008
rect 53206 38994 53346 39008
rect 53496 38994 54304 39008
rect 54454 38994 54594 39008
rect 54744 38994 55552 39008
rect 55702 38994 55842 39008
rect 55992 38994 56800 39008
rect 56950 38994 57090 39008
rect 57240 38994 58048 39008
rect 58198 38994 58338 39008
rect 58488 38994 58934 39008
rect 16418 38946 58934 38994
rect 16418 38932 16864 38946
rect 17014 38932 17154 38946
rect 17304 38932 18112 38946
rect 18262 38932 18402 38946
rect 18552 38932 19360 38946
rect 19510 38932 19650 38946
rect 19800 38932 20608 38946
rect 20758 38932 20898 38946
rect 21048 38932 21856 38946
rect 22006 38932 22146 38946
rect 22296 38932 23104 38946
rect 23254 38932 23394 38946
rect 23544 38932 24352 38946
rect 24502 38932 24642 38946
rect 24792 38932 25600 38946
rect 25750 38932 25890 38946
rect 26040 38932 26848 38946
rect 26998 38932 27138 38946
rect 27288 38932 28096 38946
rect 28246 38932 28386 38946
rect 28536 38932 29344 38946
rect 29494 38932 29634 38946
rect 29784 38932 30592 38946
rect 30742 38932 30882 38946
rect 31032 38932 31840 38946
rect 31990 38932 32130 38946
rect 32280 38932 33088 38946
rect 33238 38932 33378 38946
rect 33528 38932 34336 38946
rect 34486 38932 34626 38946
rect 34776 38932 35584 38946
rect 35734 38932 35874 38946
rect 36024 38932 36832 38946
rect 36982 38932 37122 38946
rect 37272 38932 38080 38946
rect 38230 38932 38370 38946
rect 38520 38932 39328 38946
rect 39478 38932 39618 38946
rect 39768 38932 40576 38946
rect 40726 38932 40866 38946
rect 41016 38932 41824 38946
rect 41974 38932 42114 38946
rect 42264 38932 43072 38946
rect 43222 38932 43362 38946
rect 43512 38932 44320 38946
rect 44470 38932 44610 38946
rect 44760 38932 45568 38946
rect 45718 38932 45858 38946
rect 46008 38932 46816 38946
rect 46966 38932 47106 38946
rect 47256 38932 48064 38946
rect 48214 38932 48354 38946
rect 48504 38932 49312 38946
rect 49462 38932 49602 38946
rect 49752 38932 50560 38946
rect 50710 38932 50850 38946
rect 51000 38932 51808 38946
rect 51958 38932 52098 38946
rect 52248 38932 53056 38946
rect 53206 38932 53346 38946
rect 53496 38932 54304 38946
rect 54454 38932 54594 38946
rect 54744 38932 55552 38946
rect 55702 38932 55842 38946
rect 55992 38932 56800 38946
rect 56950 38932 57090 38946
rect 57240 38932 58048 38946
rect 58198 38932 58338 38946
rect 58488 38932 58934 38946
rect 16898 38884 16980 38898
rect 17188 38884 17270 38898
rect 18146 38884 18228 38898
rect 18436 38884 18518 38898
rect 19394 38884 19476 38898
rect 19684 38884 19766 38898
rect 20642 38884 20724 38898
rect 20932 38884 21014 38898
rect 21890 38884 21972 38898
rect 22180 38884 22262 38898
rect 23138 38884 23220 38898
rect 23428 38884 23510 38898
rect 24386 38884 24468 38898
rect 24676 38884 24758 38898
rect 25634 38884 25716 38898
rect 25924 38884 26006 38898
rect 26882 38884 26964 38898
rect 27172 38884 27254 38898
rect 28130 38884 28212 38898
rect 28420 38884 28502 38898
rect 29378 38884 29460 38898
rect 29668 38884 29750 38898
rect 30626 38884 30708 38898
rect 30916 38884 30998 38898
rect 31874 38884 31956 38898
rect 32164 38884 32246 38898
rect 33122 38884 33204 38898
rect 33412 38884 33494 38898
rect 34370 38884 34452 38898
rect 34660 38884 34742 38898
rect 35618 38884 35700 38898
rect 35908 38884 35990 38898
rect 36866 38884 36948 38898
rect 37156 38884 37238 38898
rect 38114 38884 38196 38898
rect 38404 38884 38486 38898
rect 39362 38884 39444 38898
rect 39652 38884 39734 38898
rect 40610 38884 40692 38898
rect 40900 38884 40982 38898
rect 41858 38884 41940 38898
rect 42148 38884 42230 38898
rect 43106 38884 43188 38898
rect 43396 38884 43478 38898
rect 44354 38884 44436 38898
rect 44644 38884 44726 38898
rect 45602 38884 45684 38898
rect 45892 38884 45974 38898
rect 46850 38884 46932 38898
rect 47140 38884 47222 38898
rect 48098 38884 48180 38898
rect 48388 38884 48470 38898
rect 49346 38884 49428 38898
rect 49636 38884 49718 38898
rect 50594 38884 50676 38898
rect 50884 38884 50966 38898
rect 51842 38884 51924 38898
rect 52132 38884 52214 38898
rect 53090 38884 53172 38898
rect 53380 38884 53462 38898
rect 54338 38884 54420 38898
rect 54628 38884 54710 38898
rect 55586 38884 55668 38898
rect 55876 38884 55958 38898
rect 56834 38884 56916 38898
rect 57124 38884 57206 38898
rect 58082 38884 58164 38898
rect 58372 38884 58454 38898
rect 16418 38836 58934 38884
rect 16418 38678 58934 38788
rect 16418 38582 58934 38630
rect 16898 38568 16980 38582
rect 17188 38568 17270 38582
rect 18146 38568 18228 38582
rect 18436 38568 18518 38582
rect 19394 38568 19476 38582
rect 19684 38568 19766 38582
rect 20642 38568 20724 38582
rect 20932 38568 21014 38582
rect 21890 38568 21972 38582
rect 22180 38568 22262 38582
rect 23138 38568 23220 38582
rect 23428 38568 23510 38582
rect 24386 38568 24468 38582
rect 24676 38568 24758 38582
rect 25634 38568 25716 38582
rect 25924 38568 26006 38582
rect 26882 38568 26964 38582
rect 27172 38568 27254 38582
rect 28130 38568 28212 38582
rect 28420 38568 28502 38582
rect 29378 38568 29460 38582
rect 29668 38568 29750 38582
rect 30626 38568 30708 38582
rect 30916 38568 30998 38582
rect 31874 38568 31956 38582
rect 32164 38568 32246 38582
rect 33122 38568 33204 38582
rect 33412 38568 33494 38582
rect 34370 38568 34452 38582
rect 34660 38568 34742 38582
rect 35618 38568 35700 38582
rect 35908 38568 35990 38582
rect 36866 38568 36948 38582
rect 37156 38568 37238 38582
rect 38114 38568 38196 38582
rect 38404 38568 38486 38582
rect 39362 38568 39444 38582
rect 39652 38568 39734 38582
rect 40610 38568 40692 38582
rect 40900 38568 40982 38582
rect 41858 38568 41940 38582
rect 42148 38568 42230 38582
rect 43106 38568 43188 38582
rect 43396 38568 43478 38582
rect 44354 38568 44436 38582
rect 44644 38568 44726 38582
rect 45602 38568 45684 38582
rect 45892 38568 45974 38582
rect 46850 38568 46932 38582
rect 47140 38568 47222 38582
rect 48098 38568 48180 38582
rect 48388 38568 48470 38582
rect 49346 38568 49428 38582
rect 49636 38568 49718 38582
rect 50594 38568 50676 38582
rect 50884 38568 50966 38582
rect 51842 38568 51924 38582
rect 52132 38568 52214 38582
rect 53090 38568 53172 38582
rect 53380 38568 53462 38582
rect 54338 38568 54420 38582
rect 54628 38568 54710 38582
rect 55586 38568 55668 38582
rect 55876 38568 55958 38582
rect 56834 38568 56916 38582
rect 57124 38568 57206 38582
rect 58082 38568 58164 38582
rect 58372 38568 58454 38582
rect 16418 38520 16864 38534
rect 17014 38520 17154 38534
rect 17304 38520 18112 38534
rect 18262 38520 18402 38534
rect 18552 38520 19360 38534
rect 19510 38520 19650 38534
rect 19800 38520 20608 38534
rect 20758 38520 20898 38534
rect 21048 38520 21856 38534
rect 22006 38520 22146 38534
rect 22296 38520 23104 38534
rect 23254 38520 23394 38534
rect 23544 38520 24352 38534
rect 24502 38520 24642 38534
rect 24792 38520 25600 38534
rect 25750 38520 25890 38534
rect 26040 38520 26848 38534
rect 26998 38520 27138 38534
rect 27288 38520 28096 38534
rect 28246 38520 28386 38534
rect 28536 38520 29344 38534
rect 29494 38520 29634 38534
rect 29784 38520 30592 38534
rect 30742 38520 30882 38534
rect 31032 38520 31840 38534
rect 31990 38520 32130 38534
rect 32280 38520 33088 38534
rect 33238 38520 33378 38534
rect 33528 38520 34336 38534
rect 34486 38520 34626 38534
rect 34776 38520 35584 38534
rect 35734 38520 35874 38534
rect 36024 38520 36832 38534
rect 36982 38520 37122 38534
rect 37272 38520 38080 38534
rect 38230 38520 38370 38534
rect 38520 38520 39328 38534
rect 39478 38520 39618 38534
rect 39768 38520 40576 38534
rect 40726 38520 40866 38534
rect 41016 38520 41824 38534
rect 41974 38520 42114 38534
rect 42264 38520 43072 38534
rect 43222 38520 43362 38534
rect 43512 38520 44320 38534
rect 44470 38520 44610 38534
rect 44760 38520 45568 38534
rect 45718 38520 45858 38534
rect 46008 38520 46816 38534
rect 46966 38520 47106 38534
rect 47256 38520 48064 38534
rect 48214 38520 48354 38534
rect 48504 38520 49312 38534
rect 49462 38520 49602 38534
rect 49752 38520 50560 38534
rect 50710 38520 50850 38534
rect 51000 38520 51808 38534
rect 51958 38520 52098 38534
rect 52248 38520 53056 38534
rect 53206 38520 53346 38534
rect 53496 38520 54304 38534
rect 54454 38520 54594 38534
rect 54744 38520 55552 38534
rect 55702 38520 55842 38534
rect 55992 38520 56800 38534
rect 56950 38520 57090 38534
rect 57240 38520 58048 38534
rect 58198 38520 58338 38534
rect 58488 38520 58934 38534
rect 16418 38472 58934 38520
rect 16418 38458 16864 38472
rect 17014 38458 17154 38472
rect 17304 38458 18112 38472
rect 18262 38458 18402 38472
rect 18552 38458 19360 38472
rect 19510 38458 19650 38472
rect 19800 38458 20608 38472
rect 20758 38458 20898 38472
rect 21048 38458 21856 38472
rect 22006 38458 22146 38472
rect 22296 38458 23104 38472
rect 23254 38458 23394 38472
rect 23544 38458 24352 38472
rect 24502 38458 24642 38472
rect 24792 38458 25600 38472
rect 25750 38458 25890 38472
rect 26040 38458 26848 38472
rect 26998 38458 27138 38472
rect 27288 38458 28096 38472
rect 28246 38458 28386 38472
rect 28536 38458 29344 38472
rect 29494 38458 29634 38472
rect 29784 38458 30592 38472
rect 30742 38458 30882 38472
rect 31032 38458 31840 38472
rect 31990 38458 32130 38472
rect 32280 38458 33088 38472
rect 33238 38458 33378 38472
rect 33528 38458 34336 38472
rect 34486 38458 34626 38472
rect 34776 38458 35584 38472
rect 35734 38458 35874 38472
rect 36024 38458 36832 38472
rect 36982 38458 37122 38472
rect 37272 38458 38080 38472
rect 38230 38458 38370 38472
rect 38520 38458 39328 38472
rect 39478 38458 39618 38472
rect 39768 38458 40576 38472
rect 40726 38458 40866 38472
rect 41016 38458 41824 38472
rect 41974 38458 42114 38472
rect 42264 38458 43072 38472
rect 43222 38458 43362 38472
rect 43512 38458 44320 38472
rect 44470 38458 44610 38472
rect 44760 38458 45568 38472
rect 45718 38458 45858 38472
rect 46008 38458 46816 38472
rect 46966 38458 47106 38472
rect 47256 38458 48064 38472
rect 48214 38458 48354 38472
rect 48504 38458 49312 38472
rect 49462 38458 49602 38472
rect 49752 38458 50560 38472
rect 50710 38458 50850 38472
rect 51000 38458 51808 38472
rect 51958 38458 52098 38472
rect 52248 38458 53056 38472
rect 53206 38458 53346 38472
rect 53496 38458 54304 38472
rect 54454 38458 54594 38472
rect 54744 38458 55552 38472
rect 55702 38458 55842 38472
rect 55992 38458 56800 38472
rect 56950 38458 57090 38472
rect 57240 38458 58048 38472
rect 58198 38458 58338 38472
rect 58488 38458 58934 38472
rect 16898 38410 16980 38424
rect 17188 38410 17270 38424
rect 18146 38410 18228 38424
rect 18436 38410 18518 38424
rect 19394 38410 19476 38424
rect 19684 38410 19766 38424
rect 20642 38410 20724 38424
rect 20932 38410 21014 38424
rect 21890 38410 21972 38424
rect 22180 38410 22262 38424
rect 23138 38410 23220 38424
rect 23428 38410 23510 38424
rect 24386 38410 24468 38424
rect 24676 38410 24758 38424
rect 25634 38410 25716 38424
rect 25924 38410 26006 38424
rect 26882 38410 26964 38424
rect 27172 38410 27254 38424
rect 28130 38410 28212 38424
rect 28420 38410 28502 38424
rect 29378 38410 29460 38424
rect 29668 38410 29750 38424
rect 30626 38410 30708 38424
rect 30916 38410 30998 38424
rect 31874 38410 31956 38424
rect 32164 38410 32246 38424
rect 33122 38410 33204 38424
rect 33412 38410 33494 38424
rect 34370 38410 34452 38424
rect 34660 38410 34742 38424
rect 35618 38410 35700 38424
rect 35908 38410 35990 38424
rect 36866 38410 36948 38424
rect 37156 38410 37238 38424
rect 38114 38410 38196 38424
rect 38404 38410 38486 38424
rect 39362 38410 39444 38424
rect 39652 38410 39734 38424
rect 40610 38410 40692 38424
rect 40900 38410 40982 38424
rect 41858 38410 41940 38424
rect 42148 38410 42230 38424
rect 43106 38410 43188 38424
rect 43396 38410 43478 38424
rect 44354 38410 44436 38424
rect 44644 38410 44726 38424
rect 45602 38410 45684 38424
rect 45892 38410 45974 38424
rect 46850 38410 46932 38424
rect 47140 38410 47222 38424
rect 48098 38410 48180 38424
rect 48388 38410 48470 38424
rect 49346 38410 49428 38424
rect 49636 38410 49718 38424
rect 50594 38410 50676 38424
rect 50884 38410 50966 38424
rect 51842 38410 51924 38424
rect 52132 38410 52214 38424
rect 53090 38410 53172 38424
rect 53380 38410 53462 38424
rect 54338 38410 54420 38424
rect 54628 38410 54710 38424
rect 55586 38410 55668 38424
rect 55876 38410 55958 38424
rect 56834 38410 56916 38424
rect 57124 38410 57206 38424
rect 58082 38410 58164 38424
rect 58372 38410 58454 38424
rect 16418 38362 58934 38410
rect 16418 38266 58934 38314
rect 16898 38252 16980 38266
rect 17188 38252 17270 38266
rect 18146 38252 18228 38266
rect 18436 38252 18518 38266
rect 19394 38252 19476 38266
rect 19684 38252 19766 38266
rect 20642 38252 20724 38266
rect 20932 38252 21014 38266
rect 21890 38252 21972 38266
rect 22180 38252 22262 38266
rect 23138 38252 23220 38266
rect 23428 38252 23510 38266
rect 24386 38252 24468 38266
rect 24676 38252 24758 38266
rect 25634 38252 25716 38266
rect 25924 38252 26006 38266
rect 26882 38252 26964 38266
rect 27172 38252 27254 38266
rect 28130 38252 28212 38266
rect 28420 38252 28502 38266
rect 29378 38252 29460 38266
rect 29668 38252 29750 38266
rect 30626 38252 30708 38266
rect 30916 38252 30998 38266
rect 31874 38252 31956 38266
rect 32164 38252 32246 38266
rect 33122 38252 33204 38266
rect 33412 38252 33494 38266
rect 34370 38252 34452 38266
rect 34660 38252 34742 38266
rect 35618 38252 35700 38266
rect 35908 38252 35990 38266
rect 36866 38252 36948 38266
rect 37156 38252 37238 38266
rect 38114 38252 38196 38266
rect 38404 38252 38486 38266
rect 39362 38252 39444 38266
rect 39652 38252 39734 38266
rect 40610 38252 40692 38266
rect 40900 38252 40982 38266
rect 41858 38252 41940 38266
rect 42148 38252 42230 38266
rect 43106 38252 43188 38266
rect 43396 38252 43478 38266
rect 44354 38252 44436 38266
rect 44644 38252 44726 38266
rect 45602 38252 45684 38266
rect 45892 38252 45974 38266
rect 46850 38252 46932 38266
rect 47140 38252 47222 38266
rect 48098 38252 48180 38266
rect 48388 38252 48470 38266
rect 49346 38252 49428 38266
rect 49636 38252 49718 38266
rect 50594 38252 50676 38266
rect 50884 38252 50966 38266
rect 51842 38252 51924 38266
rect 52132 38252 52214 38266
rect 53090 38252 53172 38266
rect 53380 38252 53462 38266
rect 54338 38252 54420 38266
rect 54628 38252 54710 38266
rect 55586 38252 55668 38266
rect 55876 38252 55958 38266
rect 56834 38252 56916 38266
rect 57124 38252 57206 38266
rect 58082 38252 58164 38266
rect 58372 38252 58454 38266
rect 16418 38204 16864 38218
rect 17014 38204 17154 38218
rect 17304 38204 18112 38218
rect 18262 38204 18402 38218
rect 18552 38204 19360 38218
rect 19510 38204 19650 38218
rect 19800 38204 20608 38218
rect 20758 38204 20898 38218
rect 21048 38204 21856 38218
rect 22006 38204 22146 38218
rect 22296 38204 23104 38218
rect 23254 38204 23394 38218
rect 23544 38204 24352 38218
rect 24502 38204 24642 38218
rect 24792 38204 25600 38218
rect 25750 38204 25890 38218
rect 26040 38204 26848 38218
rect 26998 38204 27138 38218
rect 27288 38204 28096 38218
rect 28246 38204 28386 38218
rect 28536 38204 29344 38218
rect 29494 38204 29634 38218
rect 29784 38204 30592 38218
rect 30742 38204 30882 38218
rect 31032 38204 31840 38218
rect 31990 38204 32130 38218
rect 32280 38204 33088 38218
rect 33238 38204 33378 38218
rect 33528 38204 34336 38218
rect 34486 38204 34626 38218
rect 34776 38204 35584 38218
rect 35734 38204 35874 38218
rect 36024 38204 36832 38218
rect 36982 38204 37122 38218
rect 37272 38204 38080 38218
rect 38230 38204 38370 38218
rect 38520 38204 39328 38218
rect 39478 38204 39618 38218
rect 39768 38204 40576 38218
rect 40726 38204 40866 38218
rect 41016 38204 41824 38218
rect 41974 38204 42114 38218
rect 42264 38204 43072 38218
rect 43222 38204 43362 38218
rect 43512 38204 44320 38218
rect 44470 38204 44610 38218
rect 44760 38204 45568 38218
rect 45718 38204 45858 38218
rect 46008 38204 46816 38218
rect 46966 38204 47106 38218
rect 47256 38204 48064 38218
rect 48214 38204 48354 38218
rect 48504 38204 49312 38218
rect 49462 38204 49602 38218
rect 49752 38204 50560 38218
rect 50710 38204 50850 38218
rect 51000 38204 51808 38218
rect 51958 38204 52098 38218
rect 52248 38204 53056 38218
rect 53206 38204 53346 38218
rect 53496 38204 54304 38218
rect 54454 38204 54594 38218
rect 54744 38204 55552 38218
rect 55702 38204 55842 38218
rect 55992 38204 56800 38218
rect 56950 38204 57090 38218
rect 57240 38204 58048 38218
rect 58198 38204 58338 38218
rect 58488 38204 58934 38218
rect 16418 38156 58934 38204
rect 16418 38142 16864 38156
rect 17014 38142 17154 38156
rect 17304 38142 18112 38156
rect 18262 38142 18402 38156
rect 18552 38142 19360 38156
rect 19510 38142 19650 38156
rect 19800 38142 20608 38156
rect 20758 38142 20898 38156
rect 21048 38142 21856 38156
rect 22006 38142 22146 38156
rect 22296 38142 23104 38156
rect 23254 38142 23394 38156
rect 23544 38142 24352 38156
rect 24502 38142 24642 38156
rect 24792 38142 25600 38156
rect 25750 38142 25890 38156
rect 26040 38142 26848 38156
rect 26998 38142 27138 38156
rect 27288 38142 28096 38156
rect 28246 38142 28386 38156
rect 28536 38142 29344 38156
rect 29494 38142 29634 38156
rect 29784 38142 30592 38156
rect 30742 38142 30882 38156
rect 31032 38142 31840 38156
rect 31990 38142 32130 38156
rect 32280 38142 33088 38156
rect 33238 38142 33378 38156
rect 33528 38142 34336 38156
rect 34486 38142 34626 38156
rect 34776 38142 35584 38156
rect 35734 38142 35874 38156
rect 36024 38142 36832 38156
rect 36982 38142 37122 38156
rect 37272 38142 38080 38156
rect 38230 38142 38370 38156
rect 38520 38142 39328 38156
rect 39478 38142 39618 38156
rect 39768 38142 40576 38156
rect 40726 38142 40866 38156
rect 41016 38142 41824 38156
rect 41974 38142 42114 38156
rect 42264 38142 43072 38156
rect 43222 38142 43362 38156
rect 43512 38142 44320 38156
rect 44470 38142 44610 38156
rect 44760 38142 45568 38156
rect 45718 38142 45858 38156
rect 46008 38142 46816 38156
rect 46966 38142 47106 38156
rect 47256 38142 48064 38156
rect 48214 38142 48354 38156
rect 48504 38142 49312 38156
rect 49462 38142 49602 38156
rect 49752 38142 50560 38156
rect 50710 38142 50850 38156
rect 51000 38142 51808 38156
rect 51958 38142 52098 38156
rect 52248 38142 53056 38156
rect 53206 38142 53346 38156
rect 53496 38142 54304 38156
rect 54454 38142 54594 38156
rect 54744 38142 55552 38156
rect 55702 38142 55842 38156
rect 55992 38142 56800 38156
rect 56950 38142 57090 38156
rect 57240 38142 58048 38156
rect 58198 38142 58338 38156
rect 58488 38142 58934 38156
rect 16898 38094 16980 38108
rect 17188 38094 17270 38108
rect 18146 38094 18228 38108
rect 18436 38094 18518 38108
rect 19394 38094 19476 38108
rect 19684 38094 19766 38108
rect 20642 38094 20724 38108
rect 20932 38094 21014 38108
rect 21890 38094 21972 38108
rect 22180 38094 22262 38108
rect 23138 38094 23220 38108
rect 23428 38094 23510 38108
rect 24386 38094 24468 38108
rect 24676 38094 24758 38108
rect 25634 38094 25716 38108
rect 25924 38094 26006 38108
rect 26882 38094 26964 38108
rect 27172 38094 27254 38108
rect 28130 38094 28212 38108
rect 28420 38094 28502 38108
rect 29378 38094 29460 38108
rect 29668 38094 29750 38108
rect 30626 38094 30708 38108
rect 30916 38094 30998 38108
rect 31874 38094 31956 38108
rect 32164 38094 32246 38108
rect 33122 38094 33204 38108
rect 33412 38094 33494 38108
rect 34370 38094 34452 38108
rect 34660 38094 34742 38108
rect 35618 38094 35700 38108
rect 35908 38094 35990 38108
rect 36866 38094 36948 38108
rect 37156 38094 37238 38108
rect 38114 38094 38196 38108
rect 38404 38094 38486 38108
rect 39362 38094 39444 38108
rect 39652 38094 39734 38108
rect 40610 38094 40692 38108
rect 40900 38094 40982 38108
rect 41858 38094 41940 38108
rect 42148 38094 42230 38108
rect 43106 38094 43188 38108
rect 43396 38094 43478 38108
rect 44354 38094 44436 38108
rect 44644 38094 44726 38108
rect 45602 38094 45684 38108
rect 45892 38094 45974 38108
rect 46850 38094 46932 38108
rect 47140 38094 47222 38108
rect 48098 38094 48180 38108
rect 48388 38094 48470 38108
rect 49346 38094 49428 38108
rect 49636 38094 49718 38108
rect 50594 38094 50676 38108
rect 50884 38094 50966 38108
rect 51842 38094 51924 38108
rect 52132 38094 52214 38108
rect 53090 38094 53172 38108
rect 53380 38094 53462 38108
rect 54338 38094 54420 38108
rect 54628 38094 54710 38108
rect 55586 38094 55668 38108
rect 55876 38094 55958 38108
rect 56834 38094 56916 38108
rect 57124 38094 57206 38108
rect 58082 38094 58164 38108
rect 58372 38094 58454 38108
rect 16418 38046 58934 38094
rect 16418 37888 58934 37998
rect 16418 37792 58934 37840
rect 16898 37778 16980 37792
rect 17188 37778 17270 37792
rect 18146 37778 18228 37792
rect 18436 37778 18518 37792
rect 19394 37778 19476 37792
rect 19684 37778 19766 37792
rect 20642 37778 20724 37792
rect 20932 37778 21014 37792
rect 21890 37778 21972 37792
rect 22180 37778 22262 37792
rect 23138 37778 23220 37792
rect 23428 37778 23510 37792
rect 24386 37778 24468 37792
rect 24676 37778 24758 37792
rect 25634 37778 25716 37792
rect 25924 37778 26006 37792
rect 26882 37778 26964 37792
rect 27172 37778 27254 37792
rect 28130 37778 28212 37792
rect 28420 37778 28502 37792
rect 29378 37778 29460 37792
rect 29668 37778 29750 37792
rect 30626 37778 30708 37792
rect 30916 37778 30998 37792
rect 31874 37778 31956 37792
rect 32164 37778 32246 37792
rect 33122 37778 33204 37792
rect 33412 37778 33494 37792
rect 34370 37778 34452 37792
rect 34660 37778 34742 37792
rect 35618 37778 35700 37792
rect 35908 37778 35990 37792
rect 36866 37778 36948 37792
rect 37156 37778 37238 37792
rect 38114 37778 38196 37792
rect 38404 37778 38486 37792
rect 39362 37778 39444 37792
rect 39652 37778 39734 37792
rect 40610 37778 40692 37792
rect 40900 37778 40982 37792
rect 41858 37778 41940 37792
rect 42148 37778 42230 37792
rect 43106 37778 43188 37792
rect 43396 37778 43478 37792
rect 44354 37778 44436 37792
rect 44644 37778 44726 37792
rect 45602 37778 45684 37792
rect 45892 37778 45974 37792
rect 46850 37778 46932 37792
rect 47140 37778 47222 37792
rect 48098 37778 48180 37792
rect 48388 37778 48470 37792
rect 49346 37778 49428 37792
rect 49636 37778 49718 37792
rect 50594 37778 50676 37792
rect 50884 37778 50966 37792
rect 51842 37778 51924 37792
rect 52132 37778 52214 37792
rect 53090 37778 53172 37792
rect 53380 37778 53462 37792
rect 54338 37778 54420 37792
rect 54628 37778 54710 37792
rect 55586 37778 55668 37792
rect 55876 37778 55958 37792
rect 56834 37778 56916 37792
rect 57124 37778 57206 37792
rect 58082 37778 58164 37792
rect 58372 37778 58454 37792
rect 16418 37730 16864 37744
rect 17014 37730 17154 37744
rect 17304 37730 18112 37744
rect 18262 37730 18402 37744
rect 18552 37730 19360 37744
rect 19510 37730 19650 37744
rect 19800 37730 20608 37744
rect 20758 37730 20898 37744
rect 21048 37730 21856 37744
rect 22006 37730 22146 37744
rect 22296 37730 23104 37744
rect 23254 37730 23394 37744
rect 23544 37730 24352 37744
rect 24502 37730 24642 37744
rect 24792 37730 25600 37744
rect 25750 37730 25890 37744
rect 26040 37730 26848 37744
rect 26998 37730 27138 37744
rect 27288 37730 28096 37744
rect 28246 37730 28386 37744
rect 28536 37730 29344 37744
rect 29494 37730 29634 37744
rect 29784 37730 30592 37744
rect 30742 37730 30882 37744
rect 31032 37730 31840 37744
rect 31990 37730 32130 37744
rect 32280 37730 33088 37744
rect 33238 37730 33378 37744
rect 33528 37730 34336 37744
rect 34486 37730 34626 37744
rect 34776 37730 35584 37744
rect 35734 37730 35874 37744
rect 36024 37730 36832 37744
rect 36982 37730 37122 37744
rect 37272 37730 38080 37744
rect 38230 37730 38370 37744
rect 38520 37730 39328 37744
rect 39478 37730 39618 37744
rect 39768 37730 40576 37744
rect 40726 37730 40866 37744
rect 41016 37730 41824 37744
rect 41974 37730 42114 37744
rect 42264 37730 43072 37744
rect 43222 37730 43362 37744
rect 43512 37730 44320 37744
rect 44470 37730 44610 37744
rect 44760 37730 45568 37744
rect 45718 37730 45858 37744
rect 46008 37730 46816 37744
rect 46966 37730 47106 37744
rect 47256 37730 48064 37744
rect 48214 37730 48354 37744
rect 48504 37730 49312 37744
rect 49462 37730 49602 37744
rect 49752 37730 50560 37744
rect 50710 37730 50850 37744
rect 51000 37730 51808 37744
rect 51958 37730 52098 37744
rect 52248 37730 53056 37744
rect 53206 37730 53346 37744
rect 53496 37730 54304 37744
rect 54454 37730 54594 37744
rect 54744 37730 55552 37744
rect 55702 37730 55842 37744
rect 55992 37730 56800 37744
rect 56950 37730 57090 37744
rect 57240 37730 58048 37744
rect 58198 37730 58338 37744
rect 58488 37730 58934 37744
rect 16418 37682 58934 37730
rect 16418 37668 16864 37682
rect 17014 37668 17154 37682
rect 17304 37668 18112 37682
rect 18262 37668 18402 37682
rect 18552 37668 19360 37682
rect 19510 37668 19650 37682
rect 19800 37668 20608 37682
rect 20758 37668 20898 37682
rect 21048 37668 21856 37682
rect 22006 37668 22146 37682
rect 22296 37668 23104 37682
rect 23254 37668 23394 37682
rect 23544 37668 24352 37682
rect 24502 37668 24642 37682
rect 24792 37668 25600 37682
rect 25750 37668 25890 37682
rect 26040 37668 26848 37682
rect 26998 37668 27138 37682
rect 27288 37668 28096 37682
rect 28246 37668 28386 37682
rect 28536 37668 29344 37682
rect 29494 37668 29634 37682
rect 29784 37668 30592 37682
rect 30742 37668 30882 37682
rect 31032 37668 31840 37682
rect 31990 37668 32130 37682
rect 32280 37668 33088 37682
rect 33238 37668 33378 37682
rect 33528 37668 34336 37682
rect 34486 37668 34626 37682
rect 34776 37668 35584 37682
rect 35734 37668 35874 37682
rect 36024 37668 36832 37682
rect 36982 37668 37122 37682
rect 37272 37668 38080 37682
rect 38230 37668 38370 37682
rect 38520 37668 39328 37682
rect 39478 37668 39618 37682
rect 39768 37668 40576 37682
rect 40726 37668 40866 37682
rect 41016 37668 41824 37682
rect 41974 37668 42114 37682
rect 42264 37668 43072 37682
rect 43222 37668 43362 37682
rect 43512 37668 44320 37682
rect 44470 37668 44610 37682
rect 44760 37668 45568 37682
rect 45718 37668 45858 37682
rect 46008 37668 46816 37682
rect 46966 37668 47106 37682
rect 47256 37668 48064 37682
rect 48214 37668 48354 37682
rect 48504 37668 49312 37682
rect 49462 37668 49602 37682
rect 49752 37668 50560 37682
rect 50710 37668 50850 37682
rect 51000 37668 51808 37682
rect 51958 37668 52098 37682
rect 52248 37668 53056 37682
rect 53206 37668 53346 37682
rect 53496 37668 54304 37682
rect 54454 37668 54594 37682
rect 54744 37668 55552 37682
rect 55702 37668 55842 37682
rect 55992 37668 56800 37682
rect 56950 37668 57090 37682
rect 57240 37668 58048 37682
rect 58198 37668 58338 37682
rect 58488 37668 58934 37682
rect 16898 37620 16980 37634
rect 17188 37620 17270 37634
rect 18146 37620 18228 37634
rect 18436 37620 18518 37634
rect 19394 37620 19476 37634
rect 19684 37620 19766 37634
rect 20642 37620 20724 37634
rect 20932 37620 21014 37634
rect 21890 37620 21972 37634
rect 22180 37620 22262 37634
rect 23138 37620 23220 37634
rect 23428 37620 23510 37634
rect 24386 37620 24468 37634
rect 24676 37620 24758 37634
rect 25634 37620 25716 37634
rect 25924 37620 26006 37634
rect 26882 37620 26964 37634
rect 27172 37620 27254 37634
rect 28130 37620 28212 37634
rect 28420 37620 28502 37634
rect 29378 37620 29460 37634
rect 29668 37620 29750 37634
rect 30626 37620 30708 37634
rect 30916 37620 30998 37634
rect 31874 37620 31956 37634
rect 32164 37620 32246 37634
rect 33122 37620 33204 37634
rect 33412 37620 33494 37634
rect 34370 37620 34452 37634
rect 34660 37620 34742 37634
rect 35618 37620 35700 37634
rect 35908 37620 35990 37634
rect 36866 37620 36948 37634
rect 37156 37620 37238 37634
rect 38114 37620 38196 37634
rect 38404 37620 38486 37634
rect 39362 37620 39444 37634
rect 39652 37620 39734 37634
rect 40610 37620 40692 37634
rect 40900 37620 40982 37634
rect 41858 37620 41940 37634
rect 42148 37620 42230 37634
rect 43106 37620 43188 37634
rect 43396 37620 43478 37634
rect 44354 37620 44436 37634
rect 44644 37620 44726 37634
rect 45602 37620 45684 37634
rect 45892 37620 45974 37634
rect 46850 37620 46932 37634
rect 47140 37620 47222 37634
rect 48098 37620 48180 37634
rect 48388 37620 48470 37634
rect 49346 37620 49428 37634
rect 49636 37620 49718 37634
rect 50594 37620 50676 37634
rect 50884 37620 50966 37634
rect 51842 37620 51924 37634
rect 52132 37620 52214 37634
rect 53090 37620 53172 37634
rect 53380 37620 53462 37634
rect 54338 37620 54420 37634
rect 54628 37620 54710 37634
rect 55586 37620 55668 37634
rect 55876 37620 55958 37634
rect 56834 37620 56916 37634
rect 57124 37620 57206 37634
rect 58082 37620 58164 37634
rect 58372 37620 58454 37634
rect 16418 37572 58934 37620
rect 16418 37476 58934 37524
rect 16898 37462 16980 37476
rect 17188 37462 17270 37476
rect 18146 37462 18228 37476
rect 18436 37462 18518 37476
rect 19394 37462 19476 37476
rect 19684 37462 19766 37476
rect 20642 37462 20724 37476
rect 20932 37462 21014 37476
rect 21890 37462 21972 37476
rect 22180 37462 22262 37476
rect 23138 37462 23220 37476
rect 23428 37462 23510 37476
rect 24386 37462 24468 37476
rect 24676 37462 24758 37476
rect 25634 37462 25716 37476
rect 25924 37462 26006 37476
rect 26882 37462 26964 37476
rect 27172 37462 27254 37476
rect 28130 37462 28212 37476
rect 28420 37462 28502 37476
rect 29378 37462 29460 37476
rect 29668 37462 29750 37476
rect 30626 37462 30708 37476
rect 30916 37462 30998 37476
rect 31874 37462 31956 37476
rect 32164 37462 32246 37476
rect 33122 37462 33204 37476
rect 33412 37462 33494 37476
rect 34370 37462 34452 37476
rect 34660 37462 34742 37476
rect 35618 37462 35700 37476
rect 35908 37462 35990 37476
rect 36866 37462 36948 37476
rect 37156 37462 37238 37476
rect 38114 37462 38196 37476
rect 38404 37462 38486 37476
rect 39362 37462 39444 37476
rect 39652 37462 39734 37476
rect 40610 37462 40692 37476
rect 40900 37462 40982 37476
rect 41858 37462 41940 37476
rect 42148 37462 42230 37476
rect 43106 37462 43188 37476
rect 43396 37462 43478 37476
rect 44354 37462 44436 37476
rect 44644 37462 44726 37476
rect 45602 37462 45684 37476
rect 45892 37462 45974 37476
rect 46850 37462 46932 37476
rect 47140 37462 47222 37476
rect 48098 37462 48180 37476
rect 48388 37462 48470 37476
rect 49346 37462 49428 37476
rect 49636 37462 49718 37476
rect 50594 37462 50676 37476
rect 50884 37462 50966 37476
rect 51842 37462 51924 37476
rect 52132 37462 52214 37476
rect 53090 37462 53172 37476
rect 53380 37462 53462 37476
rect 54338 37462 54420 37476
rect 54628 37462 54710 37476
rect 55586 37462 55668 37476
rect 55876 37462 55958 37476
rect 56834 37462 56916 37476
rect 57124 37462 57206 37476
rect 58082 37462 58164 37476
rect 58372 37462 58454 37476
rect 16418 37414 16864 37428
rect 17014 37414 17154 37428
rect 17304 37414 18112 37428
rect 18262 37414 18402 37428
rect 18552 37414 19360 37428
rect 19510 37414 19650 37428
rect 19800 37414 20608 37428
rect 20758 37414 20898 37428
rect 21048 37414 21856 37428
rect 22006 37414 22146 37428
rect 22296 37414 23104 37428
rect 23254 37414 23394 37428
rect 23544 37414 24352 37428
rect 24502 37414 24642 37428
rect 24792 37414 25600 37428
rect 25750 37414 25890 37428
rect 26040 37414 26848 37428
rect 26998 37414 27138 37428
rect 27288 37414 28096 37428
rect 28246 37414 28386 37428
rect 28536 37414 29344 37428
rect 29494 37414 29634 37428
rect 29784 37414 30592 37428
rect 30742 37414 30882 37428
rect 31032 37414 31840 37428
rect 31990 37414 32130 37428
rect 32280 37414 33088 37428
rect 33238 37414 33378 37428
rect 33528 37414 34336 37428
rect 34486 37414 34626 37428
rect 34776 37414 35584 37428
rect 35734 37414 35874 37428
rect 36024 37414 36832 37428
rect 36982 37414 37122 37428
rect 37272 37414 38080 37428
rect 38230 37414 38370 37428
rect 38520 37414 39328 37428
rect 39478 37414 39618 37428
rect 39768 37414 40576 37428
rect 40726 37414 40866 37428
rect 41016 37414 41824 37428
rect 41974 37414 42114 37428
rect 42264 37414 43072 37428
rect 43222 37414 43362 37428
rect 43512 37414 44320 37428
rect 44470 37414 44610 37428
rect 44760 37414 45568 37428
rect 45718 37414 45858 37428
rect 46008 37414 46816 37428
rect 46966 37414 47106 37428
rect 47256 37414 48064 37428
rect 48214 37414 48354 37428
rect 48504 37414 49312 37428
rect 49462 37414 49602 37428
rect 49752 37414 50560 37428
rect 50710 37414 50850 37428
rect 51000 37414 51808 37428
rect 51958 37414 52098 37428
rect 52248 37414 53056 37428
rect 53206 37414 53346 37428
rect 53496 37414 54304 37428
rect 54454 37414 54594 37428
rect 54744 37414 55552 37428
rect 55702 37414 55842 37428
rect 55992 37414 56800 37428
rect 56950 37414 57090 37428
rect 57240 37414 58048 37428
rect 58198 37414 58338 37428
rect 58488 37414 58934 37428
rect 16418 37366 58934 37414
rect 16418 37352 16864 37366
rect 17014 37352 17154 37366
rect 17304 37352 18112 37366
rect 18262 37352 18402 37366
rect 18552 37352 19360 37366
rect 19510 37352 19650 37366
rect 19800 37352 20608 37366
rect 20758 37352 20898 37366
rect 21048 37352 21856 37366
rect 22006 37352 22146 37366
rect 22296 37352 23104 37366
rect 23254 37352 23394 37366
rect 23544 37352 24352 37366
rect 24502 37352 24642 37366
rect 24792 37352 25600 37366
rect 25750 37352 25890 37366
rect 26040 37352 26848 37366
rect 26998 37352 27138 37366
rect 27288 37352 28096 37366
rect 28246 37352 28386 37366
rect 28536 37352 29344 37366
rect 29494 37352 29634 37366
rect 29784 37352 30592 37366
rect 30742 37352 30882 37366
rect 31032 37352 31840 37366
rect 31990 37352 32130 37366
rect 32280 37352 33088 37366
rect 33238 37352 33378 37366
rect 33528 37352 34336 37366
rect 34486 37352 34626 37366
rect 34776 37352 35584 37366
rect 35734 37352 35874 37366
rect 36024 37352 36832 37366
rect 36982 37352 37122 37366
rect 37272 37352 38080 37366
rect 38230 37352 38370 37366
rect 38520 37352 39328 37366
rect 39478 37352 39618 37366
rect 39768 37352 40576 37366
rect 40726 37352 40866 37366
rect 41016 37352 41824 37366
rect 41974 37352 42114 37366
rect 42264 37352 43072 37366
rect 43222 37352 43362 37366
rect 43512 37352 44320 37366
rect 44470 37352 44610 37366
rect 44760 37352 45568 37366
rect 45718 37352 45858 37366
rect 46008 37352 46816 37366
rect 46966 37352 47106 37366
rect 47256 37352 48064 37366
rect 48214 37352 48354 37366
rect 48504 37352 49312 37366
rect 49462 37352 49602 37366
rect 49752 37352 50560 37366
rect 50710 37352 50850 37366
rect 51000 37352 51808 37366
rect 51958 37352 52098 37366
rect 52248 37352 53056 37366
rect 53206 37352 53346 37366
rect 53496 37352 54304 37366
rect 54454 37352 54594 37366
rect 54744 37352 55552 37366
rect 55702 37352 55842 37366
rect 55992 37352 56800 37366
rect 56950 37352 57090 37366
rect 57240 37352 58048 37366
rect 58198 37352 58338 37366
rect 58488 37352 58934 37366
rect 16898 37304 16980 37318
rect 17188 37304 17270 37318
rect 18146 37304 18228 37318
rect 18436 37304 18518 37318
rect 19394 37304 19476 37318
rect 19684 37304 19766 37318
rect 20642 37304 20724 37318
rect 20932 37304 21014 37318
rect 21890 37304 21972 37318
rect 22180 37304 22262 37318
rect 23138 37304 23220 37318
rect 23428 37304 23510 37318
rect 24386 37304 24468 37318
rect 24676 37304 24758 37318
rect 25634 37304 25716 37318
rect 25924 37304 26006 37318
rect 26882 37304 26964 37318
rect 27172 37304 27254 37318
rect 28130 37304 28212 37318
rect 28420 37304 28502 37318
rect 29378 37304 29460 37318
rect 29668 37304 29750 37318
rect 30626 37304 30708 37318
rect 30916 37304 30998 37318
rect 31874 37304 31956 37318
rect 32164 37304 32246 37318
rect 33122 37304 33204 37318
rect 33412 37304 33494 37318
rect 34370 37304 34452 37318
rect 34660 37304 34742 37318
rect 35618 37304 35700 37318
rect 35908 37304 35990 37318
rect 36866 37304 36948 37318
rect 37156 37304 37238 37318
rect 38114 37304 38196 37318
rect 38404 37304 38486 37318
rect 39362 37304 39444 37318
rect 39652 37304 39734 37318
rect 40610 37304 40692 37318
rect 40900 37304 40982 37318
rect 41858 37304 41940 37318
rect 42148 37304 42230 37318
rect 43106 37304 43188 37318
rect 43396 37304 43478 37318
rect 44354 37304 44436 37318
rect 44644 37304 44726 37318
rect 45602 37304 45684 37318
rect 45892 37304 45974 37318
rect 46850 37304 46932 37318
rect 47140 37304 47222 37318
rect 48098 37304 48180 37318
rect 48388 37304 48470 37318
rect 49346 37304 49428 37318
rect 49636 37304 49718 37318
rect 50594 37304 50676 37318
rect 50884 37304 50966 37318
rect 51842 37304 51924 37318
rect 52132 37304 52214 37318
rect 53090 37304 53172 37318
rect 53380 37304 53462 37318
rect 54338 37304 54420 37318
rect 54628 37304 54710 37318
rect 55586 37304 55668 37318
rect 55876 37304 55958 37318
rect 56834 37304 56916 37318
rect 57124 37304 57206 37318
rect 58082 37304 58164 37318
rect 58372 37304 58454 37318
rect 16418 37256 58934 37304
rect 16418 37098 58934 37208
rect 16418 37002 58934 37050
rect 16898 36988 16980 37002
rect 17188 36988 17270 37002
rect 18146 36988 18228 37002
rect 18436 36988 18518 37002
rect 19394 36988 19476 37002
rect 19684 36988 19766 37002
rect 20642 36988 20724 37002
rect 20932 36988 21014 37002
rect 21890 36988 21972 37002
rect 22180 36988 22262 37002
rect 23138 36988 23220 37002
rect 23428 36988 23510 37002
rect 24386 36988 24468 37002
rect 24676 36988 24758 37002
rect 25634 36988 25716 37002
rect 25924 36988 26006 37002
rect 26882 36988 26964 37002
rect 27172 36988 27254 37002
rect 28130 36988 28212 37002
rect 28420 36988 28502 37002
rect 29378 36988 29460 37002
rect 29668 36988 29750 37002
rect 30626 36988 30708 37002
rect 30916 36988 30998 37002
rect 31874 36988 31956 37002
rect 32164 36988 32246 37002
rect 33122 36988 33204 37002
rect 33412 36988 33494 37002
rect 34370 36988 34452 37002
rect 34660 36988 34742 37002
rect 35618 36988 35700 37002
rect 35908 36988 35990 37002
rect 36866 36988 36948 37002
rect 37156 36988 37238 37002
rect 38114 36988 38196 37002
rect 38404 36988 38486 37002
rect 39362 36988 39444 37002
rect 39652 36988 39734 37002
rect 40610 36988 40692 37002
rect 40900 36988 40982 37002
rect 41858 36988 41940 37002
rect 42148 36988 42230 37002
rect 43106 36988 43188 37002
rect 43396 36988 43478 37002
rect 44354 36988 44436 37002
rect 44644 36988 44726 37002
rect 45602 36988 45684 37002
rect 45892 36988 45974 37002
rect 46850 36988 46932 37002
rect 47140 36988 47222 37002
rect 48098 36988 48180 37002
rect 48388 36988 48470 37002
rect 49346 36988 49428 37002
rect 49636 36988 49718 37002
rect 50594 36988 50676 37002
rect 50884 36988 50966 37002
rect 51842 36988 51924 37002
rect 52132 36988 52214 37002
rect 53090 36988 53172 37002
rect 53380 36988 53462 37002
rect 54338 36988 54420 37002
rect 54628 36988 54710 37002
rect 55586 36988 55668 37002
rect 55876 36988 55958 37002
rect 56834 36988 56916 37002
rect 57124 36988 57206 37002
rect 58082 36988 58164 37002
rect 58372 36988 58454 37002
rect 16418 36940 16864 36954
rect 17014 36940 17154 36954
rect 17304 36940 18112 36954
rect 18262 36940 18402 36954
rect 18552 36940 19360 36954
rect 19510 36940 19650 36954
rect 19800 36940 20608 36954
rect 20758 36940 20898 36954
rect 21048 36940 21856 36954
rect 22006 36940 22146 36954
rect 22296 36940 23104 36954
rect 23254 36940 23394 36954
rect 23544 36940 24352 36954
rect 24502 36940 24642 36954
rect 24792 36940 25600 36954
rect 25750 36940 25890 36954
rect 26040 36940 26848 36954
rect 26998 36940 27138 36954
rect 27288 36940 28096 36954
rect 28246 36940 28386 36954
rect 28536 36940 29344 36954
rect 29494 36940 29634 36954
rect 29784 36940 30592 36954
rect 30742 36940 30882 36954
rect 31032 36940 31840 36954
rect 31990 36940 32130 36954
rect 32280 36940 33088 36954
rect 33238 36940 33378 36954
rect 33528 36940 34336 36954
rect 34486 36940 34626 36954
rect 34776 36940 35584 36954
rect 35734 36940 35874 36954
rect 36024 36940 36832 36954
rect 36982 36940 37122 36954
rect 37272 36940 38080 36954
rect 38230 36940 38370 36954
rect 38520 36940 39328 36954
rect 39478 36940 39618 36954
rect 39768 36940 40576 36954
rect 40726 36940 40866 36954
rect 41016 36940 41824 36954
rect 41974 36940 42114 36954
rect 42264 36940 43072 36954
rect 43222 36940 43362 36954
rect 43512 36940 44320 36954
rect 44470 36940 44610 36954
rect 44760 36940 45568 36954
rect 45718 36940 45858 36954
rect 46008 36940 46816 36954
rect 46966 36940 47106 36954
rect 47256 36940 48064 36954
rect 48214 36940 48354 36954
rect 48504 36940 49312 36954
rect 49462 36940 49602 36954
rect 49752 36940 50560 36954
rect 50710 36940 50850 36954
rect 51000 36940 51808 36954
rect 51958 36940 52098 36954
rect 52248 36940 53056 36954
rect 53206 36940 53346 36954
rect 53496 36940 54304 36954
rect 54454 36940 54594 36954
rect 54744 36940 55552 36954
rect 55702 36940 55842 36954
rect 55992 36940 56800 36954
rect 56950 36940 57090 36954
rect 57240 36940 58048 36954
rect 58198 36940 58338 36954
rect 58488 36940 58934 36954
rect 16418 36892 58934 36940
rect 16418 36878 16864 36892
rect 17014 36878 17154 36892
rect 17304 36878 18112 36892
rect 18262 36878 18402 36892
rect 18552 36878 19360 36892
rect 19510 36878 19650 36892
rect 19800 36878 20608 36892
rect 20758 36878 20898 36892
rect 21048 36878 21856 36892
rect 22006 36878 22146 36892
rect 22296 36878 23104 36892
rect 23254 36878 23394 36892
rect 23544 36878 24352 36892
rect 24502 36878 24642 36892
rect 24792 36878 25600 36892
rect 25750 36878 25890 36892
rect 26040 36878 26848 36892
rect 26998 36878 27138 36892
rect 27288 36878 28096 36892
rect 28246 36878 28386 36892
rect 28536 36878 29344 36892
rect 29494 36878 29634 36892
rect 29784 36878 30592 36892
rect 30742 36878 30882 36892
rect 31032 36878 31840 36892
rect 31990 36878 32130 36892
rect 32280 36878 33088 36892
rect 33238 36878 33378 36892
rect 33528 36878 34336 36892
rect 34486 36878 34626 36892
rect 34776 36878 35584 36892
rect 35734 36878 35874 36892
rect 36024 36878 36832 36892
rect 36982 36878 37122 36892
rect 37272 36878 38080 36892
rect 38230 36878 38370 36892
rect 38520 36878 39328 36892
rect 39478 36878 39618 36892
rect 39768 36878 40576 36892
rect 40726 36878 40866 36892
rect 41016 36878 41824 36892
rect 41974 36878 42114 36892
rect 42264 36878 43072 36892
rect 43222 36878 43362 36892
rect 43512 36878 44320 36892
rect 44470 36878 44610 36892
rect 44760 36878 45568 36892
rect 45718 36878 45858 36892
rect 46008 36878 46816 36892
rect 46966 36878 47106 36892
rect 47256 36878 48064 36892
rect 48214 36878 48354 36892
rect 48504 36878 49312 36892
rect 49462 36878 49602 36892
rect 49752 36878 50560 36892
rect 50710 36878 50850 36892
rect 51000 36878 51808 36892
rect 51958 36878 52098 36892
rect 52248 36878 53056 36892
rect 53206 36878 53346 36892
rect 53496 36878 54304 36892
rect 54454 36878 54594 36892
rect 54744 36878 55552 36892
rect 55702 36878 55842 36892
rect 55992 36878 56800 36892
rect 56950 36878 57090 36892
rect 57240 36878 58048 36892
rect 58198 36878 58338 36892
rect 58488 36878 58934 36892
rect 16898 36830 16980 36844
rect 17188 36830 17270 36844
rect 18146 36830 18228 36844
rect 18436 36830 18518 36844
rect 19394 36830 19476 36844
rect 19684 36830 19766 36844
rect 20642 36830 20724 36844
rect 20932 36830 21014 36844
rect 21890 36830 21972 36844
rect 22180 36830 22262 36844
rect 23138 36830 23220 36844
rect 23428 36830 23510 36844
rect 24386 36830 24468 36844
rect 24676 36830 24758 36844
rect 25634 36830 25716 36844
rect 25924 36830 26006 36844
rect 26882 36830 26964 36844
rect 27172 36830 27254 36844
rect 28130 36830 28212 36844
rect 28420 36830 28502 36844
rect 29378 36830 29460 36844
rect 29668 36830 29750 36844
rect 30626 36830 30708 36844
rect 30916 36830 30998 36844
rect 31874 36830 31956 36844
rect 32164 36830 32246 36844
rect 33122 36830 33204 36844
rect 33412 36830 33494 36844
rect 34370 36830 34452 36844
rect 34660 36830 34742 36844
rect 35618 36830 35700 36844
rect 35908 36830 35990 36844
rect 36866 36830 36948 36844
rect 37156 36830 37238 36844
rect 38114 36830 38196 36844
rect 38404 36830 38486 36844
rect 39362 36830 39444 36844
rect 39652 36830 39734 36844
rect 40610 36830 40692 36844
rect 40900 36830 40982 36844
rect 41858 36830 41940 36844
rect 42148 36830 42230 36844
rect 43106 36830 43188 36844
rect 43396 36830 43478 36844
rect 44354 36830 44436 36844
rect 44644 36830 44726 36844
rect 45602 36830 45684 36844
rect 45892 36830 45974 36844
rect 46850 36830 46932 36844
rect 47140 36830 47222 36844
rect 48098 36830 48180 36844
rect 48388 36830 48470 36844
rect 49346 36830 49428 36844
rect 49636 36830 49718 36844
rect 50594 36830 50676 36844
rect 50884 36830 50966 36844
rect 51842 36830 51924 36844
rect 52132 36830 52214 36844
rect 53090 36830 53172 36844
rect 53380 36830 53462 36844
rect 54338 36830 54420 36844
rect 54628 36830 54710 36844
rect 55586 36830 55668 36844
rect 55876 36830 55958 36844
rect 56834 36830 56916 36844
rect 57124 36830 57206 36844
rect 58082 36830 58164 36844
rect 58372 36830 58454 36844
rect 16418 36782 58934 36830
rect 16418 36686 58934 36734
rect 16898 36672 16980 36686
rect 17188 36672 17270 36686
rect 18146 36672 18228 36686
rect 18436 36672 18518 36686
rect 19394 36672 19476 36686
rect 19684 36672 19766 36686
rect 20642 36672 20724 36686
rect 20932 36672 21014 36686
rect 21890 36672 21972 36686
rect 22180 36672 22262 36686
rect 23138 36672 23220 36686
rect 23428 36672 23510 36686
rect 24386 36672 24468 36686
rect 24676 36672 24758 36686
rect 25634 36672 25716 36686
rect 25924 36672 26006 36686
rect 26882 36672 26964 36686
rect 27172 36672 27254 36686
rect 28130 36672 28212 36686
rect 28420 36672 28502 36686
rect 29378 36672 29460 36686
rect 29668 36672 29750 36686
rect 30626 36672 30708 36686
rect 30916 36672 30998 36686
rect 31874 36672 31956 36686
rect 32164 36672 32246 36686
rect 33122 36672 33204 36686
rect 33412 36672 33494 36686
rect 34370 36672 34452 36686
rect 34660 36672 34742 36686
rect 35618 36672 35700 36686
rect 35908 36672 35990 36686
rect 36866 36672 36948 36686
rect 37156 36672 37238 36686
rect 38114 36672 38196 36686
rect 38404 36672 38486 36686
rect 39362 36672 39444 36686
rect 39652 36672 39734 36686
rect 40610 36672 40692 36686
rect 40900 36672 40982 36686
rect 41858 36672 41940 36686
rect 42148 36672 42230 36686
rect 43106 36672 43188 36686
rect 43396 36672 43478 36686
rect 44354 36672 44436 36686
rect 44644 36672 44726 36686
rect 45602 36672 45684 36686
rect 45892 36672 45974 36686
rect 46850 36672 46932 36686
rect 47140 36672 47222 36686
rect 48098 36672 48180 36686
rect 48388 36672 48470 36686
rect 49346 36672 49428 36686
rect 49636 36672 49718 36686
rect 50594 36672 50676 36686
rect 50884 36672 50966 36686
rect 51842 36672 51924 36686
rect 52132 36672 52214 36686
rect 53090 36672 53172 36686
rect 53380 36672 53462 36686
rect 54338 36672 54420 36686
rect 54628 36672 54710 36686
rect 55586 36672 55668 36686
rect 55876 36672 55958 36686
rect 56834 36672 56916 36686
rect 57124 36672 57206 36686
rect 58082 36672 58164 36686
rect 58372 36672 58454 36686
rect 16418 36624 16864 36638
rect 17014 36624 17154 36638
rect 17304 36624 18112 36638
rect 18262 36624 18402 36638
rect 18552 36624 19360 36638
rect 19510 36624 19650 36638
rect 19800 36624 20608 36638
rect 20758 36624 20898 36638
rect 21048 36624 21856 36638
rect 22006 36624 22146 36638
rect 22296 36624 23104 36638
rect 23254 36624 23394 36638
rect 23544 36624 24352 36638
rect 24502 36624 24642 36638
rect 24792 36624 25600 36638
rect 25750 36624 25890 36638
rect 26040 36624 26848 36638
rect 26998 36624 27138 36638
rect 27288 36624 28096 36638
rect 28246 36624 28386 36638
rect 28536 36624 29344 36638
rect 29494 36624 29634 36638
rect 29784 36624 30592 36638
rect 30742 36624 30882 36638
rect 31032 36624 31840 36638
rect 31990 36624 32130 36638
rect 32280 36624 33088 36638
rect 33238 36624 33378 36638
rect 33528 36624 34336 36638
rect 34486 36624 34626 36638
rect 34776 36624 35584 36638
rect 35734 36624 35874 36638
rect 36024 36624 36832 36638
rect 36982 36624 37122 36638
rect 37272 36624 38080 36638
rect 38230 36624 38370 36638
rect 38520 36624 39328 36638
rect 39478 36624 39618 36638
rect 39768 36624 40576 36638
rect 40726 36624 40866 36638
rect 41016 36624 41824 36638
rect 41974 36624 42114 36638
rect 42264 36624 43072 36638
rect 43222 36624 43362 36638
rect 43512 36624 44320 36638
rect 44470 36624 44610 36638
rect 44760 36624 45568 36638
rect 45718 36624 45858 36638
rect 46008 36624 46816 36638
rect 46966 36624 47106 36638
rect 47256 36624 48064 36638
rect 48214 36624 48354 36638
rect 48504 36624 49312 36638
rect 49462 36624 49602 36638
rect 49752 36624 50560 36638
rect 50710 36624 50850 36638
rect 51000 36624 51808 36638
rect 51958 36624 52098 36638
rect 52248 36624 53056 36638
rect 53206 36624 53346 36638
rect 53496 36624 54304 36638
rect 54454 36624 54594 36638
rect 54744 36624 55552 36638
rect 55702 36624 55842 36638
rect 55992 36624 56800 36638
rect 56950 36624 57090 36638
rect 57240 36624 58048 36638
rect 58198 36624 58338 36638
rect 58488 36624 58934 36638
rect 16418 36576 58934 36624
rect 16418 36562 16864 36576
rect 17014 36562 17154 36576
rect 17304 36562 18112 36576
rect 18262 36562 18402 36576
rect 18552 36562 19360 36576
rect 19510 36562 19650 36576
rect 19800 36562 20608 36576
rect 20758 36562 20898 36576
rect 21048 36562 21856 36576
rect 22006 36562 22146 36576
rect 22296 36562 23104 36576
rect 23254 36562 23394 36576
rect 23544 36562 24352 36576
rect 24502 36562 24642 36576
rect 24792 36562 25600 36576
rect 25750 36562 25890 36576
rect 26040 36562 26848 36576
rect 26998 36562 27138 36576
rect 27288 36562 28096 36576
rect 28246 36562 28386 36576
rect 28536 36562 29344 36576
rect 29494 36562 29634 36576
rect 29784 36562 30592 36576
rect 30742 36562 30882 36576
rect 31032 36562 31840 36576
rect 31990 36562 32130 36576
rect 32280 36562 33088 36576
rect 33238 36562 33378 36576
rect 33528 36562 34336 36576
rect 34486 36562 34626 36576
rect 34776 36562 35584 36576
rect 35734 36562 35874 36576
rect 36024 36562 36832 36576
rect 36982 36562 37122 36576
rect 37272 36562 38080 36576
rect 38230 36562 38370 36576
rect 38520 36562 39328 36576
rect 39478 36562 39618 36576
rect 39768 36562 40576 36576
rect 40726 36562 40866 36576
rect 41016 36562 41824 36576
rect 41974 36562 42114 36576
rect 42264 36562 43072 36576
rect 43222 36562 43362 36576
rect 43512 36562 44320 36576
rect 44470 36562 44610 36576
rect 44760 36562 45568 36576
rect 45718 36562 45858 36576
rect 46008 36562 46816 36576
rect 46966 36562 47106 36576
rect 47256 36562 48064 36576
rect 48214 36562 48354 36576
rect 48504 36562 49312 36576
rect 49462 36562 49602 36576
rect 49752 36562 50560 36576
rect 50710 36562 50850 36576
rect 51000 36562 51808 36576
rect 51958 36562 52098 36576
rect 52248 36562 53056 36576
rect 53206 36562 53346 36576
rect 53496 36562 54304 36576
rect 54454 36562 54594 36576
rect 54744 36562 55552 36576
rect 55702 36562 55842 36576
rect 55992 36562 56800 36576
rect 56950 36562 57090 36576
rect 57240 36562 58048 36576
rect 58198 36562 58338 36576
rect 58488 36562 58934 36576
rect 16898 36514 16980 36528
rect 17188 36514 17270 36528
rect 18146 36514 18228 36528
rect 18436 36514 18518 36528
rect 19394 36514 19476 36528
rect 19684 36514 19766 36528
rect 20642 36514 20724 36528
rect 20932 36514 21014 36528
rect 21890 36514 21972 36528
rect 22180 36514 22262 36528
rect 23138 36514 23220 36528
rect 23428 36514 23510 36528
rect 24386 36514 24468 36528
rect 24676 36514 24758 36528
rect 25634 36514 25716 36528
rect 25924 36514 26006 36528
rect 26882 36514 26964 36528
rect 27172 36514 27254 36528
rect 28130 36514 28212 36528
rect 28420 36514 28502 36528
rect 29378 36514 29460 36528
rect 29668 36514 29750 36528
rect 30626 36514 30708 36528
rect 30916 36514 30998 36528
rect 31874 36514 31956 36528
rect 32164 36514 32246 36528
rect 33122 36514 33204 36528
rect 33412 36514 33494 36528
rect 34370 36514 34452 36528
rect 34660 36514 34742 36528
rect 35618 36514 35700 36528
rect 35908 36514 35990 36528
rect 36866 36514 36948 36528
rect 37156 36514 37238 36528
rect 38114 36514 38196 36528
rect 38404 36514 38486 36528
rect 39362 36514 39444 36528
rect 39652 36514 39734 36528
rect 40610 36514 40692 36528
rect 40900 36514 40982 36528
rect 41858 36514 41940 36528
rect 42148 36514 42230 36528
rect 43106 36514 43188 36528
rect 43396 36514 43478 36528
rect 44354 36514 44436 36528
rect 44644 36514 44726 36528
rect 45602 36514 45684 36528
rect 45892 36514 45974 36528
rect 46850 36514 46932 36528
rect 47140 36514 47222 36528
rect 48098 36514 48180 36528
rect 48388 36514 48470 36528
rect 49346 36514 49428 36528
rect 49636 36514 49718 36528
rect 50594 36514 50676 36528
rect 50884 36514 50966 36528
rect 51842 36514 51924 36528
rect 52132 36514 52214 36528
rect 53090 36514 53172 36528
rect 53380 36514 53462 36528
rect 54338 36514 54420 36528
rect 54628 36514 54710 36528
rect 55586 36514 55668 36528
rect 55876 36514 55958 36528
rect 56834 36514 56916 36528
rect 57124 36514 57206 36528
rect 58082 36514 58164 36528
rect 58372 36514 58454 36528
rect 16418 36466 58934 36514
rect 16418 36308 58934 36418
rect 16418 36212 58934 36260
rect 16898 36198 16980 36212
rect 17188 36198 17270 36212
rect 18146 36198 18228 36212
rect 18436 36198 18518 36212
rect 19394 36198 19476 36212
rect 19684 36198 19766 36212
rect 20642 36198 20724 36212
rect 20932 36198 21014 36212
rect 21890 36198 21972 36212
rect 22180 36198 22262 36212
rect 23138 36198 23220 36212
rect 23428 36198 23510 36212
rect 24386 36198 24468 36212
rect 24676 36198 24758 36212
rect 25634 36198 25716 36212
rect 25924 36198 26006 36212
rect 26882 36198 26964 36212
rect 27172 36198 27254 36212
rect 28130 36198 28212 36212
rect 28420 36198 28502 36212
rect 29378 36198 29460 36212
rect 29668 36198 29750 36212
rect 30626 36198 30708 36212
rect 30916 36198 30998 36212
rect 31874 36198 31956 36212
rect 32164 36198 32246 36212
rect 33122 36198 33204 36212
rect 33412 36198 33494 36212
rect 34370 36198 34452 36212
rect 34660 36198 34742 36212
rect 35618 36198 35700 36212
rect 35908 36198 35990 36212
rect 36866 36198 36948 36212
rect 37156 36198 37238 36212
rect 38114 36198 38196 36212
rect 38404 36198 38486 36212
rect 39362 36198 39444 36212
rect 39652 36198 39734 36212
rect 40610 36198 40692 36212
rect 40900 36198 40982 36212
rect 41858 36198 41940 36212
rect 42148 36198 42230 36212
rect 43106 36198 43188 36212
rect 43396 36198 43478 36212
rect 44354 36198 44436 36212
rect 44644 36198 44726 36212
rect 45602 36198 45684 36212
rect 45892 36198 45974 36212
rect 46850 36198 46932 36212
rect 47140 36198 47222 36212
rect 48098 36198 48180 36212
rect 48388 36198 48470 36212
rect 49346 36198 49428 36212
rect 49636 36198 49718 36212
rect 50594 36198 50676 36212
rect 50884 36198 50966 36212
rect 51842 36198 51924 36212
rect 52132 36198 52214 36212
rect 53090 36198 53172 36212
rect 53380 36198 53462 36212
rect 54338 36198 54420 36212
rect 54628 36198 54710 36212
rect 55586 36198 55668 36212
rect 55876 36198 55958 36212
rect 56834 36198 56916 36212
rect 57124 36198 57206 36212
rect 58082 36198 58164 36212
rect 58372 36198 58454 36212
rect 16418 36150 16864 36164
rect 17014 36150 17154 36164
rect 17304 36150 18112 36164
rect 18262 36150 18402 36164
rect 18552 36150 19360 36164
rect 19510 36150 19650 36164
rect 19800 36150 20608 36164
rect 20758 36150 20898 36164
rect 21048 36150 21856 36164
rect 22006 36150 22146 36164
rect 22296 36150 23104 36164
rect 23254 36150 23394 36164
rect 23544 36150 24352 36164
rect 24502 36150 24642 36164
rect 24792 36150 25600 36164
rect 25750 36150 25890 36164
rect 26040 36150 26848 36164
rect 26998 36150 27138 36164
rect 27288 36150 28096 36164
rect 28246 36150 28386 36164
rect 28536 36150 29344 36164
rect 29494 36150 29634 36164
rect 29784 36150 30592 36164
rect 30742 36150 30882 36164
rect 31032 36150 31840 36164
rect 31990 36150 32130 36164
rect 32280 36150 33088 36164
rect 33238 36150 33378 36164
rect 33528 36150 34336 36164
rect 34486 36150 34626 36164
rect 34776 36150 35584 36164
rect 35734 36150 35874 36164
rect 36024 36150 36832 36164
rect 36982 36150 37122 36164
rect 37272 36150 38080 36164
rect 38230 36150 38370 36164
rect 38520 36150 39328 36164
rect 39478 36150 39618 36164
rect 39768 36150 40576 36164
rect 40726 36150 40866 36164
rect 41016 36150 41824 36164
rect 41974 36150 42114 36164
rect 42264 36150 43072 36164
rect 43222 36150 43362 36164
rect 43512 36150 44320 36164
rect 44470 36150 44610 36164
rect 44760 36150 45568 36164
rect 45718 36150 45858 36164
rect 46008 36150 46816 36164
rect 46966 36150 47106 36164
rect 47256 36150 48064 36164
rect 48214 36150 48354 36164
rect 48504 36150 49312 36164
rect 49462 36150 49602 36164
rect 49752 36150 50560 36164
rect 50710 36150 50850 36164
rect 51000 36150 51808 36164
rect 51958 36150 52098 36164
rect 52248 36150 53056 36164
rect 53206 36150 53346 36164
rect 53496 36150 54304 36164
rect 54454 36150 54594 36164
rect 54744 36150 55552 36164
rect 55702 36150 55842 36164
rect 55992 36150 56800 36164
rect 56950 36150 57090 36164
rect 57240 36150 58048 36164
rect 58198 36150 58338 36164
rect 58488 36150 58934 36164
rect 16418 36102 58934 36150
rect 16418 36088 16864 36102
rect 17014 36088 17154 36102
rect 17304 36088 18112 36102
rect 18262 36088 18402 36102
rect 18552 36088 19360 36102
rect 19510 36088 19650 36102
rect 19800 36088 20608 36102
rect 20758 36088 20898 36102
rect 21048 36088 21856 36102
rect 22006 36088 22146 36102
rect 22296 36088 23104 36102
rect 23254 36088 23394 36102
rect 23544 36088 24352 36102
rect 24502 36088 24642 36102
rect 24792 36088 25600 36102
rect 25750 36088 25890 36102
rect 26040 36088 26848 36102
rect 26998 36088 27138 36102
rect 27288 36088 28096 36102
rect 28246 36088 28386 36102
rect 28536 36088 29344 36102
rect 29494 36088 29634 36102
rect 29784 36088 30592 36102
rect 30742 36088 30882 36102
rect 31032 36088 31840 36102
rect 31990 36088 32130 36102
rect 32280 36088 33088 36102
rect 33238 36088 33378 36102
rect 33528 36088 34336 36102
rect 34486 36088 34626 36102
rect 34776 36088 35584 36102
rect 35734 36088 35874 36102
rect 36024 36088 36832 36102
rect 36982 36088 37122 36102
rect 37272 36088 38080 36102
rect 38230 36088 38370 36102
rect 38520 36088 39328 36102
rect 39478 36088 39618 36102
rect 39768 36088 40576 36102
rect 40726 36088 40866 36102
rect 41016 36088 41824 36102
rect 41974 36088 42114 36102
rect 42264 36088 43072 36102
rect 43222 36088 43362 36102
rect 43512 36088 44320 36102
rect 44470 36088 44610 36102
rect 44760 36088 45568 36102
rect 45718 36088 45858 36102
rect 46008 36088 46816 36102
rect 46966 36088 47106 36102
rect 47256 36088 48064 36102
rect 48214 36088 48354 36102
rect 48504 36088 49312 36102
rect 49462 36088 49602 36102
rect 49752 36088 50560 36102
rect 50710 36088 50850 36102
rect 51000 36088 51808 36102
rect 51958 36088 52098 36102
rect 52248 36088 53056 36102
rect 53206 36088 53346 36102
rect 53496 36088 54304 36102
rect 54454 36088 54594 36102
rect 54744 36088 55552 36102
rect 55702 36088 55842 36102
rect 55992 36088 56800 36102
rect 56950 36088 57090 36102
rect 57240 36088 58048 36102
rect 58198 36088 58338 36102
rect 58488 36088 58934 36102
rect 16898 36040 16980 36054
rect 17188 36040 17270 36054
rect 18146 36040 18228 36054
rect 18436 36040 18518 36054
rect 19394 36040 19476 36054
rect 19684 36040 19766 36054
rect 20642 36040 20724 36054
rect 20932 36040 21014 36054
rect 21890 36040 21972 36054
rect 22180 36040 22262 36054
rect 23138 36040 23220 36054
rect 23428 36040 23510 36054
rect 24386 36040 24468 36054
rect 24676 36040 24758 36054
rect 25634 36040 25716 36054
rect 25924 36040 26006 36054
rect 26882 36040 26964 36054
rect 27172 36040 27254 36054
rect 28130 36040 28212 36054
rect 28420 36040 28502 36054
rect 29378 36040 29460 36054
rect 29668 36040 29750 36054
rect 30626 36040 30708 36054
rect 30916 36040 30998 36054
rect 31874 36040 31956 36054
rect 32164 36040 32246 36054
rect 33122 36040 33204 36054
rect 33412 36040 33494 36054
rect 34370 36040 34452 36054
rect 34660 36040 34742 36054
rect 35618 36040 35700 36054
rect 35908 36040 35990 36054
rect 36866 36040 36948 36054
rect 37156 36040 37238 36054
rect 38114 36040 38196 36054
rect 38404 36040 38486 36054
rect 39362 36040 39444 36054
rect 39652 36040 39734 36054
rect 40610 36040 40692 36054
rect 40900 36040 40982 36054
rect 41858 36040 41940 36054
rect 42148 36040 42230 36054
rect 43106 36040 43188 36054
rect 43396 36040 43478 36054
rect 44354 36040 44436 36054
rect 44644 36040 44726 36054
rect 45602 36040 45684 36054
rect 45892 36040 45974 36054
rect 46850 36040 46932 36054
rect 47140 36040 47222 36054
rect 48098 36040 48180 36054
rect 48388 36040 48470 36054
rect 49346 36040 49428 36054
rect 49636 36040 49718 36054
rect 50594 36040 50676 36054
rect 50884 36040 50966 36054
rect 51842 36040 51924 36054
rect 52132 36040 52214 36054
rect 53090 36040 53172 36054
rect 53380 36040 53462 36054
rect 54338 36040 54420 36054
rect 54628 36040 54710 36054
rect 55586 36040 55668 36054
rect 55876 36040 55958 36054
rect 56834 36040 56916 36054
rect 57124 36040 57206 36054
rect 58082 36040 58164 36054
rect 58372 36040 58454 36054
rect 16418 35992 58934 36040
rect 16418 35896 58934 35944
rect 16898 35882 16980 35896
rect 17188 35882 17270 35896
rect 18146 35882 18228 35896
rect 18436 35882 18518 35896
rect 19394 35882 19476 35896
rect 19684 35882 19766 35896
rect 20642 35882 20724 35896
rect 20932 35882 21014 35896
rect 21890 35882 21972 35896
rect 22180 35882 22262 35896
rect 23138 35882 23220 35896
rect 23428 35882 23510 35896
rect 24386 35882 24468 35896
rect 24676 35882 24758 35896
rect 25634 35882 25716 35896
rect 25924 35882 26006 35896
rect 26882 35882 26964 35896
rect 27172 35882 27254 35896
rect 28130 35882 28212 35896
rect 28420 35882 28502 35896
rect 29378 35882 29460 35896
rect 29668 35882 29750 35896
rect 30626 35882 30708 35896
rect 30916 35882 30998 35896
rect 31874 35882 31956 35896
rect 32164 35882 32246 35896
rect 33122 35882 33204 35896
rect 33412 35882 33494 35896
rect 34370 35882 34452 35896
rect 34660 35882 34742 35896
rect 35618 35882 35700 35896
rect 35908 35882 35990 35896
rect 36866 35882 36948 35896
rect 37156 35882 37238 35896
rect 38114 35882 38196 35896
rect 38404 35882 38486 35896
rect 39362 35882 39444 35896
rect 39652 35882 39734 35896
rect 40610 35882 40692 35896
rect 40900 35882 40982 35896
rect 41858 35882 41940 35896
rect 42148 35882 42230 35896
rect 43106 35882 43188 35896
rect 43396 35882 43478 35896
rect 44354 35882 44436 35896
rect 44644 35882 44726 35896
rect 45602 35882 45684 35896
rect 45892 35882 45974 35896
rect 46850 35882 46932 35896
rect 47140 35882 47222 35896
rect 48098 35882 48180 35896
rect 48388 35882 48470 35896
rect 49346 35882 49428 35896
rect 49636 35882 49718 35896
rect 50594 35882 50676 35896
rect 50884 35882 50966 35896
rect 51842 35882 51924 35896
rect 52132 35882 52214 35896
rect 53090 35882 53172 35896
rect 53380 35882 53462 35896
rect 54338 35882 54420 35896
rect 54628 35882 54710 35896
rect 55586 35882 55668 35896
rect 55876 35882 55958 35896
rect 56834 35882 56916 35896
rect 57124 35882 57206 35896
rect 58082 35882 58164 35896
rect 58372 35882 58454 35896
rect 16418 35834 16864 35848
rect 17014 35834 17154 35848
rect 17304 35834 18112 35848
rect 18262 35834 18402 35848
rect 18552 35834 19360 35848
rect 19510 35834 19650 35848
rect 19800 35834 20608 35848
rect 20758 35834 20898 35848
rect 21048 35834 21856 35848
rect 22006 35834 22146 35848
rect 22296 35834 23104 35848
rect 23254 35834 23394 35848
rect 23544 35834 24352 35848
rect 24502 35834 24642 35848
rect 24792 35834 25600 35848
rect 25750 35834 25890 35848
rect 26040 35834 26848 35848
rect 26998 35834 27138 35848
rect 27288 35834 28096 35848
rect 28246 35834 28386 35848
rect 28536 35834 29344 35848
rect 29494 35834 29634 35848
rect 29784 35834 30592 35848
rect 30742 35834 30882 35848
rect 31032 35834 31840 35848
rect 31990 35834 32130 35848
rect 32280 35834 33088 35848
rect 33238 35834 33378 35848
rect 33528 35834 34336 35848
rect 34486 35834 34626 35848
rect 34776 35834 35584 35848
rect 35734 35834 35874 35848
rect 36024 35834 36832 35848
rect 36982 35834 37122 35848
rect 37272 35834 38080 35848
rect 38230 35834 38370 35848
rect 38520 35834 39328 35848
rect 39478 35834 39618 35848
rect 39768 35834 40576 35848
rect 40726 35834 40866 35848
rect 41016 35834 41824 35848
rect 41974 35834 42114 35848
rect 42264 35834 43072 35848
rect 43222 35834 43362 35848
rect 43512 35834 44320 35848
rect 44470 35834 44610 35848
rect 44760 35834 45568 35848
rect 45718 35834 45858 35848
rect 46008 35834 46816 35848
rect 46966 35834 47106 35848
rect 47256 35834 48064 35848
rect 48214 35834 48354 35848
rect 48504 35834 49312 35848
rect 49462 35834 49602 35848
rect 49752 35834 50560 35848
rect 50710 35834 50850 35848
rect 51000 35834 51808 35848
rect 51958 35834 52098 35848
rect 52248 35834 53056 35848
rect 53206 35834 53346 35848
rect 53496 35834 54304 35848
rect 54454 35834 54594 35848
rect 54744 35834 55552 35848
rect 55702 35834 55842 35848
rect 55992 35834 56800 35848
rect 56950 35834 57090 35848
rect 57240 35834 58048 35848
rect 58198 35834 58338 35848
rect 58488 35834 58934 35848
rect 16418 35786 58934 35834
rect 16418 35772 16864 35786
rect 17014 35772 17154 35786
rect 17304 35772 18112 35786
rect 18262 35772 18402 35786
rect 18552 35772 19360 35786
rect 19510 35772 19650 35786
rect 19800 35772 20608 35786
rect 20758 35772 20898 35786
rect 21048 35772 21856 35786
rect 22006 35772 22146 35786
rect 22296 35772 23104 35786
rect 23254 35772 23394 35786
rect 23544 35772 24352 35786
rect 24502 35772 24642 35786
rect 24792 35772 25600 35786
rect 25750 35772 25890 35786
rect 26040 35772 26848 35786
rect 26998 35772 27138 35786
rect 27288 35772 28096 35786
rect 28246 35772 28386 35786
rect 28536 35772 29344 35786
rect 29494 35772 29634 35786
rect 29784 35772 30592 35786
rect 30742 35772 30882 35786
rect 31032 35772 31840 35786
rect 31990 35772 32130 35786
rect 32280 35772 33088 35786
rect 33238 35772 33378 35786
rect 33528 35772 34336 35786
rect 34486 35772 34626 35786
rect 34776 35772 35584 35786
rect 35734 35772 35874 35786
rect 36024 35772 36832 35786
rect 36982 35772 37122 35786
rect 37272 35772 38080 35786
rect 38230 35772 38370 35786
rect 38520 35772 39328 35786
rect 39478 35772 39618 35786
rect 39768 35772 40576 35786
rect 40726 35772 40866 35786
rect 41016 35772 41824 35786
rect 41974 35772 42114 35786
rect 42264 35772 43072 35786
rect 43222 35772 43362 35786
rect 43512 35772 44320 35786
rect 44470 35772 44610 35786
rect 44760 35772 45568 35786
rect 45718 35772 45858 35786
rect 46008 35772 46816 35786
rect 46966 35772 47106 35786
rect 47256 35772 48064 35786
rect 48214 35772 48354 35786
rect 48504 35772 49312 35786
rect 49462 35772 49602 35786
rect 49752 35772 50560 35786
rect 50710 35772 50850 35786
rect 51000 35772 51808 35786
rect 51958 35772 52098 35786
rect 52248 35772 53056 35786
rect 53206 35772 53346 35786
rect 53496 35772 54304 35786
rect 54454 35772 54594 35786
rect 54744 35772 55552 35786
rect 55702 35772 55842 35786
rect 55992 35772 56800 35786
rect 56950 35772 57090 35786
rect 57240 35772 58048 35786
rect 58198 35772 58338 35786
rect 58488 35772 58934 35786
rect 16898 35724 16980 35738
rect 17188 35724 17270 35738
rect 18146 35724 18228 35738
rect 18436 35724 18518 35738
rect 19394 35724 19476 35738
rect 19684 35724 19766 35738
rect 20642 35724 20724 35738
rect 20932 35724 21014 35738
rect 21890 35724 21972 35738
rect 22180 35724 22262 35738
rect 23138 35724 23220 35738
rect 23428 35724 23510 35738
rect 24386 35724 24468 35738
rect 24676 35724 24758 35738
rect 25634 35724 25716 35738
rect 25924 35724 26006 35738
rect 26882 35724 26964 35738
rect 27172 35724 27254 35738
rect 28130 35724 28212 35738
rect 28420 35724 28502 35738
rect 29378 35724 29460 35738
rect 29668 35724 29750 35738
rect 30626 35724 30708 35738
rect 30916 35724 30998 35738
rect 31874 35724 31956 35738
rect 32164 35724 32246 35738
rect 33122 35724 33204 35738
rect 33412 35724 33494 35738
rect 34370 35724 34452 35738
rect 34660 35724 34742 35738
rect 35618 35724 35700 35738
rect 35908 35724 35990 35738
rect 36866 35724 36948 35738
rect 37156 35724 37238 35738
rect 38114 35724 38196 35738
rect 38404 35724 38486 35738
rect 39362 35724 39444 35738
rect 39652 35724 39734 35738
rect 40610 35724 40692 35738
rect 40900 35724 40982 35738
rect 41858 35724 41940 35738
rect 42148 35724 42230 35738
rect 43106 35724 43188 35738
rect 43396 35724 43478 35738
rect 44354 35724 44436 35738
rect 44644 35724 44726 35738
rect 45602 35724 45684 35738
rect 45892 35724 45974 35738
rect 46850 35724 46932 35738
rect 47140 35724 47222 35738
rect 48098 35724 48180 35738
rect 48388 35724 48470 35738
rect 49346 35724 49428 35738
rect 49636 35724 49718 35738
rect 50594 35724 50676 35738
rect 50884 35724 50966 35738
rect 51842 35724 51924 35738
rect 52132 35724 52214 35738
rect 53090 35724 53172 35738
rect 53380 35724 53462 35738
rect 54338 35724 54420 35738
rect 54628 35724 54710 35738
rect 55586 35724 55668 35738
rect 55876 35724 55958 35738
rect 56834 35724 56916 35738
rect 57124 35724 57206 35738
rect 58082 35724 58164 35738
rect 58372 35724 58454 35738
rect 16418 35676 58934 35724
rect 16418 35518 58934 35628
rect 16418 35422 58934 35470
rect 16898 35408 16980 35422
rect 17188 35408 17270 35422
rect 18146 35408 18228 35422
rect 18436 35408 18518 35422
rect 19394 35408 19476 35422
rect 19684 35408 19766 35422
rect 20642 35408 20724 35422
rect 20932 35408 21014 35422
rect 21890 35408 21972 35422
rect 22180 35408 22262 35422
rect 23138 35408 23220 35422
rect 23428 35408 23510 35422
rect 24386 35408 24468 35422
rect 24676 35408 24758 35422
rect 25634 35408 25716 35422
rect 25924 35408 26006 35422
rect 26882 35408 26964 35422
rect 27172 35408 27254 35422
rect 28130 35408 28212 35422
rect 28420 35408 28502 35422
rect 29378 35408 29460 35422
rect 29668 35408 29750 35422
rect 30626 35408 30708 35422
rect 30916 35408 30998 35422
rect 31874 35408 31956 35422
rect 32164 35408 32246 35422
rect 33122 35408 33204 35422
rect 33412 35408 33494 35422
rect 34370 35408 34452 35422
rect 34660 35408 34742 35422
rect 35618 35408 35700 35422
rect 35908 35408 35990 35422
rect 36866 35408 36948 35422
rect 37156 35408 37238 35422
rect 38114 35408 38196 35422
rect 38404 35408 38486 35422
rect 39362 35408 39444 35422
rect 39652 35408 39734 35422
rect 40610 35408 40692 35422
rect 40900 35408 40982 35422
rect 41858 35408 41940 35422
rect 42148 35408 42230 35422
rect 43106 35408 43188 35422
rect 43396 35408 43478 35422
rect 44354 35408 44436 35422
rect 44644 35408 44726 35422
rect 45602 35408 45684 35422
rect 45892 35408 45974 35422
rect 46850 35408 46932 35422
rect 47140 35408 47222 35422
rect 48098 35408 48180 35422
rect 48388 35408 48470 35422
rect 49346 35408 49428 35422
rect 49636 35408 49718 35422
rect 50594 35408 50676 35422
rect 50884 35408 50966 35422
rect 51842 35408 51924 35422
rect 52132 35408 52214 35422
rect 53090 35408 53172 35422
rect 53380 35408 53462 35422
rect 54338 35408 54420 35422
rect 54628 35408 54710 35422
rect 55586 35408 55668 35422
rect 55876 35408 55958 35422
rect 56834 35408 56916 35422
rect 57124 35408 57206 35422
rect 58082 35408 58164 35422
rect 58372 35408 58454 35422
rect 16418 35360 16864 35374
rect 17014 35360 17154 35374
rect 17304 35360 18112 35374
rect 18262 35360 18402 35374
rect 18552 35360 19360 35374
rect 19510 35360 19650 35374
rect 19800 35360 20608 35374
rect 20758 35360 20898 35374
rect 21048 35360 21856 35374
rect 22006 35360 22146 35374
rect 22296 35360 23104 35374
rect 23254 35360 23394 35374
rect 23544 35360 24352 35374
rect 24502 35360 24642 35374
rect 24792 35360 25600 35374
rect 25750 35360 25890 35374
rect 26040 35360 26848 35374
rect 26998 35360 27138 35374
rect 27288 35360 28096 35374
rect 28246 35360 28386 35374
rect 28536 35360 29344 35374
rect 29494 35360 29634 35374
rect 29784 35360 30592 35374
rect 30742 35360 30882 35374
rect 31032 35360 31840 35374
rect 31990 35360 32130 35374
rect 32280 35360 33088 35374
rect 33238 35360 33378 35374
rect 33528 35360 34336 35374
rect 34486 35360 34626 35374
rect 34776 35360 35584 35374
rect 35734 35360 35874 35374
rect 36024 35360 36832 35374
rect 36982 35360 37122 35374
rect 37272 35360 38080 35374
rect 38230 35360 38370 35374
rect 38520 35360 39328 35374
rect 39478 35360 39618 35374
rect 39768 35360 40576 35374
rect 40726 35360 40866 35374
rect 41016 35360 41824 35374
rect 41974 35360 42114 35374
rect 42264 35360 43072 35374
rect 43222 35360 43362 35374
rect 43512 35360 44320 35374
rect 44470 35360 44610 35374
rect 44760 35360 45568 35374
rect 45718 35360 45858 35374
rect 46008 35360 46816 35374
rect 46966 35360 47106 35374
rect 47256 35360 48064 35374
rect 48214 35360 48354 35374
rect 48504 35360 49312 35374
rect 49462 35360 49602 35374
rect 49752 35360 50560 35374
rect 50710 35360 50850 35374
rect 51000 35360 51808 35374
rect 51958 35360 52098 35374
rect 52248 35360 53056 35374
rect 53206 35360 53346 35374
rect 53496 35360 54304 35374
rect 54454 35360 54594 35374
rect 54744 35360 55552 35374
rect 55702 35360 55842 35374
rect 55992 35360 56800 35374
rect 56950 35360 57090 35374
rect 57240 35360 58048 35374
rect 58198 35360 58338 35374
rect 58488 35360 58934 35374
rect 16418 35312 58934 35360
rect 16418 35298 16864 35312
rect 17014 35298 17154 35312
rect 17304 35298 18112 35312
rect 18262 35298 18402 35312
rect 18552 35298 19360 35312
rect 19510 35298 19650 35312
rect 19800 35298 20608 35312
rect 20758 35298 20898 35312
rect 21048 35298 21856 35312
rect 22006 35298 22146 35312
rect 22296 35298 23104 35312
rect 23254 35298 23394 35312
rect 23544 35298 24352 35312
rect 24502 35298 24642 35312
rect 24792 35298 25600 35312
rect 25750 35298 25890 35312
rect 26040 35298 26848 35312
rect 26998 35298 27138 35312
rect 27288 35298 28096 35312
rect 28246 35298 28386 35312
rect 28536 35298 29344 35312
rect 29494 35298 29634 35312
rect 29784 35298 30592 35312
rect 30742 35298 30882 35312
rect 31032 35298 31840 35312
rect 31990 35298 32130 35312
rect 32280 35298 33088 35312
rect 33238 35298 33378 35312
rect 33528 35298 34336 35312
rect 34486 35298 34626 35312
rect 34776 35298 35584 35312
rect 35734 35298 35874 35312
rect 36024 35298 36832 35312
rect 36982 35298 37122 35312
rect 37272 35298 38080 35312
rect 38230 35298 38370 35312
rect 38520 35298 39328 35312
rect 39478 35298 39618 35312
rect 39768 35298 40576 35312
rect 40726 35298 40866 35312
rect 41016 35298 41824 35312
rect 41974 35298 42114 35312
rect 42264 35298 43072 35312
rect 43222 35298 43362 35312
rect 43512 35298 44320 35312
rect 44470 35298 44610 35312
rect 44760 35298 45568 35312
rect 45718 35298 45858 35312
rect 46008 35298 46816 35312
rect 46966 35298 47106 35312
rect 47256 35298 48064 35312
rect 48214 35298 48354 35312
rect 48504 35298 49312 35312
rect 49462 35298 49602 35312
rect 49752 35298 50560 35312
rect 50710 35298 50850 35312
rect 51000 35298 51808 35312
rect 51958 35298 52098 35312
rect 52248 35298 53056 35312
rect 53206 35298 53346 35312
rect 53496 35298 54304 35312
rect 54454 35298 54594 35312
rect 54744 35298 55552 35312
rect 55702 35298 55842 35312
rect 55992 35298 56800 35312
rect 56950 35298 57090 35312
rect 57240 35298 58048 35312
rect 58198 35298 58338 35312
rect 58488 35298 58934 35312
rect 16898 35250 16980 35264
rect 17188 35250 17270 35264
rect 18146 35250 18228 35264
rect 18436 35250 18518 35264
rect 19394 35250 19476 35264
rect 19684 35250 19766 35264
rect 20642 35250 20724 35264
rect 20932 35250 21014 35264
rect 21890 35250 21972 35264
rect 22180 35250 22262 35264
rect 23138 35250 23220 35264
rect 23428 35250 23510 35264
rect 24386 35250 24468 35264
rect 24676 35250 24758 35264
rect 25634 35250 25716 35264
rect 25924 35250 26006 35264
rect 26882 35250 26964 35264
rect 27172 35250 27254 35264
rect 28130 35250 28212 35264
rect 28420 35250 28502 35264
rect 29378 35250 29460 35264
rect 29668 35250 29750 35264
rect 30626 35250 30708 35264
rect 30916 35250 30998 35264
rect 31874 35250 31956 35264
rect 32164 35250 32246 35264
rect 33122 35250 33204 35264
rect 33412 35250 33494 35264
rect 34370 35250 34452 35264
rect 34660 35250 34742 35264
rect 35618 35250 35700 35264
rect 35908 35250 35990 35264
rect 36866 35250 36948 35264
rect 37156 35250 37238 35264
rect 38114 35250 38196 35264
rect 38404 35250 38486 35264
rect 39362 35250 39444 35264
rect 39652 35250 39734 35264
rect 40610 35250 40692 35264
rect 40900 35250 40982 35264
rect 41858 35250 41940 35264
rect 42148 35250 42230 35264
rect 43106 35250 43188 35264
rect 43396 35250 43478 35264
rect 44354 35250 44436 35264
rect 44644 35250 44726 35264
rect 45602 35250 45684 35264
rect 45892 35250 45974 35264
rect 46850 35250 46932 35264
rect 47140 35250 47222 35264
rect 48098 35250 48180 35264
rect 48388 35250 48470 35264
rect 49346 35250 49428 35264
rect 49636 35250 49718 35264
rect 50594 35250 50676 35264
rect 50884 35250 50966 35264
rect 51842 35250 51924 35264
rect 52132 35250 52214 35264
rect 53090 35250 53172 35264
rect 53380 35250 53462 35264
rect 54338 35250 54420 35264
rect 54628 35250 54710 35264
rect 55586 35250 55668 35264
rect 55876 35250 55958 35264
rect 56834 35250 56916 35264
rect 57124 35250 57206 35264
rect 58082 35250 58164 35264
rect 58372 35250 58454 35264
rect 16418 35202 58934 35250
rect 16418 35106 58934 35154
rect 16898 35092 16980 35106
rect 17188 35092 17270 35106
rect 18146 35092 18228 35106
rect 18436 35092 18518 35106
rect 19394 35092 19476 35106
rect 19684 35092 19766 35106
rect 20642 35092 20724 35106
rect 20932 35092 21014 35106
rect 21890 35092 21972 35106
rect 22180 35092 22262 35106
rect 23138 35092 23220 35106
rect 23428 35092 23510 35106
rect 24386 35092 24468 35106
rect 24676 35092 24758 35106
rect 25634 35092 25716 35106
rect 25924 35092 26006 35106
rect 26882 35092 26964 35106
rect 27172 35092 27254 35106
rect 28130 35092 28212 35106
rect 28420 35092 28502 35106
rect 29378 35092 29460 35106
rect 29668 35092 29750 35106
rect 30626 35092 30708 35106
rect 30916 35092 30998 35106
rect 31874 35092 31956 35106
rect 32164 35092 32246 35106
rect 33122 35092 33204 35106
rect 33412 35092 33494 35106
rect 34370 35092 34452 35106
rect 34660 35092 34742 35106
rect 35618 35092 35700 35106
rect 35908 35092 35990 35106
rect 36866 35092 36948 35106
rect 37156 35092 37238 35106
rect 38114 35092 38196 35106
rect 38404 35092 38486 35106
rect 39362 35092 39444 35106
rect 39652 35092 39734 35106
rect 40610 35092 40692 35106
rect 40900 35092 40982 35106
rect 41858 35092 41940 35106
rect 42148 35092 42230 35106
rect 43106 35092 43188 35106
rect 43396 35092 43478 35106
rect 44354 35092 44436 35106
rect 44644 35092 44726 35106
rect 45602 35092 45684 35106
rect 45892 35092 45974 35106
rect 46850 35092 46932 35106
rect 47140 35092 47222 35106
rect 48098 35092 48180 35106
rect 48388 35092 48470 35106
rect 49346 35092 49428 35106
rect 49636 35092 49718 35106
rect 50594 35092 50676 35106
rect 50884 35092 50966 35106
rect 51842 35092 51924 35106
rect 52132 35092 52214 35106
rect 53090 35092 53172 35106
rect 53380 35092 53462 35106
rect 54338 35092 54420 35106
rect 54628 35092 54710 35106
rect 55586 35092 55668 35106
rect 55876 35092 55958 35106
rect 56834 35092 56916 35106
rect 57124 35092 57206 35106
rect 58082 35092 58164 35106
rect 58372 35092 58454 35106
rect 16418 35044 16864 35058
rect 17014 35044 17154 35058
rect 17304 35044 18112 35058
rect 18262 35044 18402 35058
rect 18552 35044 19360 35058
rect 19510 35044 19650 35058
rect 19800 35044 20608 35058
rect 20758 35044 20898 35058
rect 21048 35044 21856 35058
rect 22006 35044 22146 35058
rect 22296 35044 23104 35058
rect 23254 35044 23394 35058
rect 23544 35044 24352 35058
rect 24502 35044 24642 35058
rect 24792 35044 25600 35058
rect 25750 35044 25890 35058
rect 26040 35044 26848 35058
rect 26998 35044 27138 35058
rect 27288 35044 28096 35058
rect 28246 35044 28386 35058
rect 28536 35044 29344 35058
rect 29494 35044 29634 35058
rect 29784 35044 30592 35058
rect 30742 35044 30882 35058
rect 31032 35044 31840 35058
rect 31990 35044 32130 35058
rect 32280 35044 33088 35058
rect 33238 35044 33378 35058
rect 33528 35044 34336 35058
rect 34486 35044 34626 35058
rect 34776 35044 35584 35058
rect 35734 35044 35874 35058
rect 36024 35044 36832 35058
rect 36982 35044 37122 35058
rect 37272 35044 38080 35058
rect 38230 35044 38370 35058
rect 38520 35044 39328 35058
rect 39478 35044 39618 35058
rect 39768 35044 40576 35058
rect 40726 35044 40866 35058
rect 41016 35044 41824 35058
rect 41974 35044 42114 35058
rect 42264 35044 43072 35058
rect 43222 35044 43362 35058
rect 43512 35044 44320 35058
rect 44470 35044 44610 35058
rect 44760 35044 45568 35058
rect 45718 35044 45858 35058
rect 46008 35044 46816 35058
rect 46966 35044 47106 35058
rect 47256 35044 48064 35058
rect 48214 35044 48354 35058
rect 48504 35044 49312 35058
rect 49462 35044 49602 35058
rect 49752 35044 50560 35058
rect 50710 35044 50850 35058
rect 51000 35044 51808 35058
rect 51958 35044 52098 35058
rect 52248 35044 53056 35058
rect 53206 35044 53346 35058
rect 53496 35044 54304 35058
rect 54454 35044 54594 35058
rect 54744 35044 55552 35058
rect 55702 35044 55842 35058
rect 55992 35044 56800 35058
rect 56950 35044 57090 35058
rect 57240 35044 58048 35058
rect 58198 35044 58338 35058
rect 58488 35044 58934 35058
rect 16418 34996 58934 35044
rect 16418 34982 16864 34996
rect 17014 34982 17154 34996
rect 17304 34982 18112 34996
rect 18262 34982 18402 34996
rect 18552 34982 19360 34996
rect 19510 34982 19650 34996
rect 19800 34982 20608 34996
rect 20758 34982 20898 34996
rect 21048 34982 21856 34996
rect 22006 34982 22146 34996
rect 22296 34982 23104 34996
rect 23254 34982 23394 34996
rect 23544 34982 24352 34996
rect 24502 34982 24642 34996
rect 24792 34982 25600 34996
rect 25750 34982 25890 34996
rect 26040 34982 26848 34996
rect 26998 34982 27138 34996
rect 27288 34982 28096 34996
rect 28246 34982 28386 34996
rect 28536 34982 29344 34996
rect 29494 34982 29634 34996
rect 29784 34982 30592 34996
rect 30742 34982 30882 34996
rect 31032 34982 31840 34996
rect 31990 34982 32130 34996
rect 32280 34982 33088 34996
rect 33238 34982 33378 34996
rect 33528 34982 34336 34996
rect 34486 34982 34626 34996
rect 34776 34982 35584 34996
rect 35734 34982 35874 34996
rect 36024 34982 36832 34996
rect 36982 34982 37122 34996
rect 37272 34982 38080 34996
rect 38230 34982 38370 34996
rect 38520 34982 39328 34996
rect 39478 34982 39618 34996
rect 39768 34982 40576 34996
rect 40726 34982 40866 34996
rect 41016 34982 41824 34996
rect 41974 34982 42114 34996
rect 42264 34982 43072 34996
rect 43222 34982 43362 34996
rect 43512 34982 44320 34996
rect 44470 34982 44610 34996
rect 44760 34982 45568 34996
rect 45718 34982 45858 34996
rect 46008 34982 46816 34996
rect 46966 34982 47106 34996
rect 47256 34982 48064 34996
rect 48214 34982 48354 34996
rect 48504 34982 49312 34996
rect 49462 34982 49602 34996
rect 49752 34982 50560 34996
rect 50710 34982 50850 34996
rect 51000 34982 51808 34996
rect 51958 34982 52098 34996
rect 52248 34982 53056 34996
rect 53206 34982 53346 34996
rect 53496 34982 54304 34996
rect 54454 34982 54594 34996
rect 54744 34982 55552 34996
rect 55702 34982 55842 34996
rect 55992 34982 56800 34996
rect 56950 34982 57090 34996
rect 57240 34982 58048 34996
rect 58198 34982 58338 34996
rect 58488 34982 58934 34996
rect 16898 34934 16980 34948
rect 17188 34934 17270 34948
rect 18146 34934 18228 34948
rect 18436 34934 18518 34948
rect 19394 34934 19476 34948
rect 19684 34934 19766 34948
rect 20642 34934 20724 34948
rect 20932 34934 21014 34948
rect 21890 34934 21972 34948
rect 22180 34934 22262 34948
rect 23138 34934 23220 34948
rect 23428 34934 23510 34948
rect 24386 34934 24468 34948
rect 24676 34934 24758 34948
rect 25634 34934 25716 34948
rect 25924 34934 26006 34948
rect 26882 34934 26964 34948
rect 27172 34934 27254 34948
rect 28130 34934 28212 34948
rect 28420 34934 28502 34948
rect 29378 34934 29460 34948
rect 29668 34934 29750 34948
rect 30626 34934 30708 34948
rect 30916 34934 30998 34948
rect 31874 34934 31956 34948
rect 32164 34934 32246 34948
rect 33122 34934 33204 34948
rect 33412 34934 33494 34948
rect 34370 34934 34452 34948
rect 34660 34934 34742 34948
rect 35618 34934 35700 34948
rect 35908 34934 35990 34948
rect 36866 34934 36948 34948
rect 37156 34934 37238 34948
rect 38114 34934 38196 34948
rect 38404 34934 38486 34948
rect 39362 34934 39444 34948
rect 39652 34934 39734 34948
rect 40610 34934 40692 34948
rect 40900 34934 40982 34948
rect 41858 34934 41940 34948
rect 42148 34934 42230 34948
rect 43106 34934 43188 34948
rect 43396 34934 43478 34948
rect 44354 34934 44436 34948
rect 44644 34934 44726 34948
rect 45602 34934 45684 34948
rect 45892 34934 45974 34948
rect 46850 34934 46932 34948
rect 47140 34934 47222 34948
rect 48098 34934 48180 34948
rect 48388 34934 48470 34948
rect 49346 34934 49428 34948
rect 49636 34934 49718 34948
rect 50594 34934 50676 34948
rect 50884 34934 50966 34948
rect 51842 34934 51924 34948
rect 52132 34934 52214 34948
rect 53090 34934 53172 34948
rect 53380 34934 53462 34948
rect 54338 34934 54420 34948
rect 54628 34934 54710 34948
rect 55586 34934 55668 34948
rect 55876 34934 55958 34948
rect 56834 34934 56916 34948
rect 57124 34934 57206 34948
rect 58082 34934 58164 34948
rect 58372 34934 58454 34948
rect 16418 34886 58934 34934
rect 16418 34728 58934 34838
rect 16418 34632 58934 34680
rect 16898 34618 16980 34632
rect 17188 34618 17270 34632
rect 18146 34618 18228 34632
rect 18436 34618 18518 34632
rect 19394 34618 19476 34632
rect 19684 34618 19766 34632
rect 20642 34618 20724 34632
rect 20932 34618 21014 34632
rect 21890 34618 21972 34632
rect 22180 34618 22262 34632
rect 23138 34618 23220 34632
rect 23428 34618 23510 34632
rect 24386 34618 24468 34632
rect 24676 34618 24758 34632
rect 25634 34618 25716 34632
rect 25924 34618 26006 34632
rect 26882 34618 26964 34632
rect 27172 34618 27254 34632
rect 28130 34618 28212 34632
rect 28420 34618 28502 34632
rect 29378 34618 29460 34632
rect 29668 34618 29750 34632
rect 30626 34618 30708 34632
rect 30916 34618 30998 34632
rect 31874 34618 31956 34632
rect 32164 34618 32246 34632
rect 33122 34618 33204 34632
rect 33412 34618 33494 34632
rect 34370 34618 34452 34632
rect 34660 34618 34742 34632
rect 35618 34618 35700 34632
rect 35908 34618 35990 34632
rect 36866 34618 36948 34632
rect 37156 34618 37238 34632
rect 38114 34618 38196 34632
rect 38404 34618 38486 34632
rect 39362 34618 39444 34632
rect 39652 34618 39734 34632
rect 40610 34618 40692 34632
rect 40900 34618 40982 34632
rect 41858 34618 41940 34632
rect 42148 34618 42230 34632
rect 43106 34618 43188 34632
rect 43396 34618 43478 34632
rect 44354 34618 44436 34632
rect 44644 34618 44726 34632
rect 45602 34618 45684 34632
rect 45892 34618 45974 34632
rect 46850 34618 46932 34632
rect 47140 34618 47222 34632
rect 48098 34618 48180 34632
rect 48388 34618 48470 34632
rect 49346 34618 49428 34632
rect 49636 34618 49718 34632
rect 50594 34618 50676 34632
rect 50884 34618 50966 34632
rect 51842 34618 51924 34632
rect 52132 34618 52214 34632
rect 53090 34618 53172 34632
rect 53380 34618 53462 34632
rect 54338 34618 54420 34632
rect 54628 34618 54710 34632
rect 55586 34618 55668 34632
rect 55876 34618 55958 34632
rect 56834 34618 56916 34632
rect 57124 34618 57206 34632
rect 58082 34618 58164 34632
rect 58372 34618 58454 34632
rect 16418 34570 16864 34584
rect 17014 34570 17154 34584
rect 17304 34570 18112 34584
rect 18262 34570 18402 34584
rect 18552 34570 19360 34584
rect 19510 34570 19650 34584
rect 19800 34570 20608 34584
rect 20758 34570 20898 34584
rect 21048 34570 21856 34584
rect 22006 34570 22146 34584
rect 22296 34570 23104 34584
rect 23254 34570 23394 34584
rect 23544 34570 24352 34584
rect 24502 34570 24642 34584
rect 24792 34570 25600 34584
rect 25750 34570 25890 34584
rect 26040 34570 26848 34584
rect 26998 34570 27138 34584
rect 27288 34570 28096 34584
rect 28246 34570 28386 34584
rect 28536 34570 29344 34584
rect 29494 34570 29634 34584
rect 29784 34570 30592 34584
rect 30742 34570 30882 34584
rect 31032 34570 31840 34584
rect 31990 34570 32130 34584
rect 32280 34570 33088 34584
rect 33238 34570 33378 34584
rect 33528 34570 34336 34584
rect 34486 34570 34626 34584
rect 34776 34570 35584 34584
rect 35734 34570 35874 34584
rect 36024 34570 36832 34584
rect 36982 34570 37122 34584
rect 37272 34570 38080 34584
rect 38230 34570 38370 34584
rect 38520 34570 39328 34584
rect 39478 34570 39618 34584
rect 39768 34570 40576 34584
rect 40726 34570 40866 34584
rect 41016 34570 41824 34584
rect 41974 34570 42114 34584
rect 42264 34570 43072 34584
rect 43222 34570 43362 34584
rect 43512 34570 44320 34584
rect 44470 34570 44610 34584
rect 44760 34570 45568 34584
rect 45718 34570 45858 34584
rect 46008 34570 46816 34584
rect 46966 34570 47106 34584
rect 47256 34570 48064 34584
rect 48214 34570 48354 34584
rect 48504 34570 49312 34584
rect 49462 34570 49602 34584
rect 49752 34570 50560 34584
rect 50710 34570 50850 34584
rect 51000 34570 51808 34584
rect 51958 34570 52098 34584
rect 52248 34570 53056 34584
rect 53206 34570 53346 34584
rect 53496 34570 54304 34584
rect 54454 34570 54594 34584
rect 54744 34570 55552 34584
rect 55702 34570 55842 34584
rect 55992 34570 56800 34584
rect 56950 34570 57090 34584
rect 57240 34570 58048 34584
rect 58198 34570 58338 34584
rect 58488 34570 58934 34584
rect 16418 34522 58934 34570
rect 16418 34508 16864 34522
rect 17014 34508 17154 34522
rect 17304 34508 18112 34522
rect 18262 34508 18402 34522
rect 18552 34508 19360 34522
rect 19510 34508 19650 34522
rect 19800 34508 20608 34522
rect 20758 34508 20898 34522
rect 21048 34508 21856 34522
rect 22006 34508 22146 34522
rect 22296 34508 23104 34522
rect 23254 34508 23394 34522
rect 23544 34508 24352 34522
rect 24502 34508 24642 34522
rect 24792 34508 25600 34522
rect 25750 34508 25890 34522
rect 26040 34508 26848 34522
rect 26998 34508 27138 34522
rect 27288 34508 28096 34522
rect 28246 34508 28386 34522
rect 28536 34508 29344 34522
rect 29494 34508 29634 34522
rect 29784 34508 30592 34522
rect 30742 34508 30882 34522
rect 31032 34508 31840 34522
rect 31990 34508 32130 34522
rect 32280 34508 33088 34522
rect 33238 34508 33378 34522
rect 33528 34508 34336 34522
rect 34486 34508 34626 34522
rect 34776 34508 35584 34522
rect 35734 34508 35874 34522
rect 36024 34508 36832 34522
rect 36982 34508 37122 34522
rect 37272 34508 38080 34522
rect 38230 34508 38370 34522
rect 38520 34508 39328 34522
rect 39478 34508 39618 34522
rect 39768 34508 40576 34522
rect 40726 34508 40866 34522
rect 41016 34508 41824 34522
rect 41974 34508 42114 34522
rect 42264 34508 43072 34522
rect 43222 34508 43362 34522
rect 43512 34508 44320 34522
rect 44470 34508 44610 34522
rect 44760 34508 45568 34522
rect 45718 34508 45858 34522
rect 46008 34508 46816 34522
rect 46966 34508 47106 34522
rect 47256 34508 48064 34522
rect 48214 34508 48354 34522
rect 48504 34508 49312 34522
rect 49462 34508 49602 34522
rect 49752 34508 50560 34522
rect 50710 34508 50850 34522
rect 51000 34508 51808 34522
rect 51958 34508 52098 34522
rect 52248 34508 53056 34522
rect 53206 34508 53346 34522
rect 53496 34508 54304 34522
rect 54454 34508 54594 34522
rect 54744 34508 55552 34522
rect 55702 34508 55842 34522
rect 55992 34508 56800 34522
rect 56950 34508 57090 34522
rect 57240 34508 58048 34522
rect 58198 34508 58338 34522
rect 58488 34508 58934 34522
rect 16898 34460 16980 34474
rect 17188 34460 17270 34474
rect 18146 34460 18228 34474
rect 18436 34460 18518 34474
rect 19394 34460 19476 34474
rect 19684 34460 19766 34474
rect 20642 34460 20724 34474
rect 20932 34460 21014 34474
rect 21890 34460 21972 34474
rect 22180 34460 22262 34474
rect 23138 34460 23220 34474
rect 23428 34460 23510 34474
rect 24386 34460 24468 34474
rect 24676 34460 24758 34474
rect 25634 34460 25716 34474
rect 25924 34460 26006 34474
rect 26882 34460 26964 34474
rect 27172 34460 27254 34474
rect 28130 34460 28212 34474
rect 28420 34460 28502 34474
rect 29378 34460 29460 34474
rect 29668 34460 29750 34474
rect 30626 34460 30708 34474
rect 30916 34460 30998 34474
rect 31874 34460 31956 34474
rect 32164 34460 32246 34474
rect 33122 34460 33204 34474
rect 33412 34460 33494 34474
rect 34370 34460 34452 34474
rect 34660 34460 34742 34474
rect 35618 34460 35700 34474
rect 35908 34460 35990 34474
rect 36866 34460 36948 34474
rect 37156 34460 37238 34474
rect 38114 34460 38196 34474
rect 38404 34460 38486 34474
rect 39362 34460 39444 34474
rect 39652 34460 39734 34474
rect 40610 34460 40692 34474
rect 40900 34460 40982 34474
rect 41858 34460 41940 34474
rect 42148 34460 42230 34474
rect 43106 34460 43188 34474
rect 43396 34460 43478 34474
rect 44354 34460 44436 34474
rect 44644 34460 44726 34474
rect 45602 34460 45684 34474
rect 45892 34460 45974 34474
rect 46850 34460 46932 34474
rect 47140 34460 47222 34474
rect 48098 34460 48180 34474
rect 48388 34460 48470 34474
rect 49346 34460 49428 34474
rect 49636 34460 49718 34474
rect 50594 34460 50676 34474
rect 50884 34460 50966 34474
rect 51842 34460 51924 34474
rect 52132 34460 52214 34474
rect 53090 34460 53172 34474
rect 53380 34460 53462 34474
rect 54338 34460 54420 34474
rect 54628 34460 54710 34474
rect 55586 34460 55668 34474
rect 55876 34460 55958 34474
rect 56834 34460 56916 34474
rect 57124 34460 57206 34474
rect 58082 34460 58164 34474
rect 58372 34460 58454 34474
rect 16418 34412 58934 34460
rect 16418 34316 58934 34364
rect 16898 34302 16980 34316
rect 17188 34302 17270 34316
rect 18146 34302 18228 34316
rect 18436 34302 18518 34316
rect 19394 34302 19476 34316
rect 19684 34302 19766 34316
rect 20642 34302 20724 34316
rect 20932 34302 21014 34316
rect 21890 34302 21972 34316
rect 22180 34302 22262 34316
rect 23138 34302 23220 34316
rect 23428 34302 23510 34316
rect 24386 34302 24468 34316
rect 24676 34302 24758 34316
rect 25634 34302 25716 34316
rect 25924 34302 26006 34316
rect 26882 34302 26964 34316
rect 27172 34302 27254 34316
rect 28130 34302 28212 34316
rect 28420 34302 28502 34316
rect 29378 34302 29460 34316
rect 29668 34302 29750 34316
rect 30626 34302 30708 34316
rect 30916 34302 30998 34316
rect 31874 34302 31956 34316
rect 32164 34302 32246 34316
rect 33122 34302 33204 34316
rect 33412 34302 33494 34316
rect 34370 34302 34452 34316
rect 34660 34302 34742 34316
rect 35618 34302 35700 34316
rect 35908 34302 35990 34316
rect 36866 34302 36948 34316
rect 37156 34302 37238 34316
rect 38114 34302 38196 34316
rect 38404 34302 38486 34316
rect 39362 34302 39444 34316
rect 39652 34302 39734 34316
rect 40610 34302 40692 34316
rect 40900 34302 40982 34316
rect 41858 34302 41940 34316
rect 42148 34302 42230 34316
rect 43106 34302 43188 34316
rect 43396 34302 43478 34316
rect 44354 34302 44436 34316
rect 44644 34302 44726 34316
rect 45602 34302 45684 34316
rect 45892 34302 45974 34316
rect 46850 34302 46932 34316
rect 47140 34302 47222 34316
rect 48098 34302 48180 34316
rect 48388 34302 48470 34316
rect 49346 34302 49428 34316
rect 49636 34302 49718 34316
rect 50594 34302 50676 34316
rect 50884 34302 50966 34316
rect 51842 34302 51924 34316
rect 52132 34302 52214 34316
rect 53090 34302 53172 34316
rect 53380 34302 53462 34316
rect 54338 34302 54420 34316
rect 54628 34302 54710 34316
rect 55586 34302 55668 34316
rect 55876 34302 55958 34316
rect 56834 34302 56916 34316
rect 57124 34302 57206 34316
rect 58082 34302 58164 34316
rect 58372 34302 58454 34316
rect 16418 34254 16864 34268
rect 17014 34254 17154 34268
rect 17304 34254 18112 34268
rect 18262 34254 18402 34268
rect 18552 34254 19360 34268
rect 19510 34254 19650 34268
rect 19800 34254 20608 34268
rect 20758 34254 20898 34268
rect 21048 34254 21856 34268
rect 22006 34254 22146 34268
rect 22296 34254 23104 34268
rect 23254 34254 23394 34268
rect 23544 34254 24352 34268
rect 24502 34254 24642 34268
rect 24792 34254 25600 34268
rect 25750 34254 25890 34268
rect 26040 34254 26848 34268
rect 26998 34254 27138 34268
rect 27288 34254 28096 34268
rect 28246 34254 28386 34268
rect 28536 34254 29344 34268
rect 29494 34254 29634 34268
rect 29784 34254 30592 34268
rect 30742 34254 30882 34268
rect 31032 34254 31840 34268
rect 31990 34254 32130 34268
rect 32280 34254 33088 34268
rect 33238 34254 33378 34268
rect 33528 34254 34336 34268
rect 34486 34254 34626 34268
rect 34776 34254 35584 34268
rect 35734 34254 35874 34268
rect 36024 34254 36832 34268
rect 36982 34254 37122 34268
rect 37272 34254 38080 34268
rect 38230 34254 38370 34268
rect 38520 34254 39328 34268
rect 39478 34254 39618 34268
rect 39768 34254 40576 34268
rect 40726 34254 40866 34268
rect 41016 34254 41824 34268
rect 41974 34254 42114 34268
rect 42264 34254 43072 34268
rect 43222 34254 43362 34268
rect 43512 34254 44320 34268
rect 44470 34254 44610 34268
rect 44760 34254 45568 34268
rect 45718 34254 45858 34268
rect 46008 34254 46816 34268
rect 46966 34254 47106 34268
rect 47256 34254 48064 34268
rect 48214 34254 48354 34268
rect 48504 34254 49312 34268
rect 49462 34254 49602 34268
rect 49752 34254 50560 34268
rect 50710 34254 50850 34268
rect 51000 34254 51808 34268
rect 51958 34254 52098 34268
rect 52248 34254 53056 34268
rect 53206 34254 53346 34268
rect 53496 34254 54304 34268
rect 54454 34254 54594 34268
rect 54744 34254 55552 34268
rect 55702 34254 55842 34268
rect 55992 34254 56800 34268
rect 56950 34254 57090 34268
rect 57240 34254 58048 34268
rect 58198 34254 58338 34268
rect 58488 34254 58934 34268
rect 16418 34206 58934 34254
rect 16418 34192 16864 34206
rect 17014 34192 17154 34206
rect 17304 34192 18112 34206
rect 18262 34192 18402 34206
rect 18552 34192 19360 34206
rect 19510 34192 19650 34206
rect 19800 34192 20608 34206
rect 20758 34192 20898 34206
rect 21048 34192 21856 34206
rect 22006 34192 22146 34206
rect 22296 34192 23104 34206
rect 23254 34192 23394 34206
rect 23544 34192 24352 34206
rect 24502 34192 24642 34206
rect 24792 34192 25600 34206
rect 25750 34192 25890 34206
rect 26040 34192 26848 34206
rect 26998 34192 27138 34206
rect 27288 34192 28096 34206
rect 28246 34192 28386 34206
rect 28536 34192 29344 34206
rect 29494 34192 29634 34206
rect 29784 34192 30592 34206
rect 30742 34192 30882 34206
rect 31032 34192 31840 34206
rect 31990 34192 32130 34206
rect 32280 34192 33088 34206
rect 33238 34192 33378 34206
rect 33528 34192 34336 34206
rect 34486 34192 34626 34206
rect 34776 34192 35584 34206
rect 35734 34192 35874 34206
rect 36024 34192 36832 34206
rect 36982 34192 37122 34206
rect 37272 34192 38080 34206
rect 38230 34192 38370 34206
rect 38520 34192 39328 34206
rect 39478 34192 39618 34206
rect 39768 34192 40576 34206
rect 40726 34192 40866 34206
rect 41016 34192 41824 34206
rect 41974 34192 42114 34206
rect 42264 34192 43072 34206
rect 43222 34192 43362 34206
rect 43512 34192 44320 34206
rect 44470 34192 44610 34206
rect 44760 34192 45568 34206
rect 45718 34192 45858 34206
rect 46008 34192 46816 34206
rect 46966 34192 47106 34206
rect 47256 34192 48064 34206
rect 48214 34192 48354 34206
rect 48504 34192 49312 34206
rect 49462 34192 49602 34206
rect 49752 34192 50560 34206
rect 50710 34192 50850 34206
rect 51000 34192 51808 34206
rect 51958 34192 52098 34206
rect 52248 34192 53056 34206
rect 53206 34192 53346 34206
rect 53496 34192 54304 34206
rect 54454 34192 54594 34206
rect 54744 34192 55552 34206
rect 55702 34192 55842 34206
rect 55992 34192 56800 34206
rect 56950 34192 57090 34206
rect 57240 34192 58048 34206
rect 58198 34192 58338 34206
rect 58488 34192 58934 34206
rect 16898 34144 16980 34158
rect 17188 34144 17270 34158
rect 18146 34144 18228 34158
rect 18436 34144 18518 34158
rect 19394 34144 19476 34158
rect 19684 34144 19766 34158
rect 20642 34144 20724 34158
rect 20932 34144 21014 34158
rect 21890 34144 21972 34158
rect 22180 34144 22262 34158
rect 23138 34144 23220 34158
rect 23428 34144 23510 34158
rect 24386 34144 24468 34158
rect 24676 34144 24758 34158
rect 25634 34144 25716 34158
rect 25924 34144 26006 34158
rect 26882 34144 26964 34158
rect 27172 34144 27254 34158
rect 28130 34144 28212 34158
rect 28420 34144 28502 34158
rect 29378 34144 29460 34158
rect 29668 34144 29750 34158
rect 30626 34144 30708 34158
rect 30916 34144 30998 34158
rect 31874 34144 31956 34158
rect 32164 34144 32246 34158
rect 33122 34144 33204 34158
rect 33412 34144 33494 34158
rect 34370 34144 34452 34158
rect 34660 34144 34742 34158
rect 35618 34144 35700 34158
rect 35908 34144 35990 34158
rect 36866 34144 36948 34158
rect 37156 34144 37238 34158
rect 38114 34144 38196 34158
rect 38404 34144 38486 34158
rect 39362 34144 39444 34158
rect 39652 34144 39734 34158
rect 40610 34144 40692 34158
rect 40900 34144 40982 34158
rect 41858 34144 41940 34158
rect 42148 34144 42230 34158
rect 43106 34144 43188 34158
rect 43396 34144 43478 34158
rect 44354 34144 44436 34158
rect 44644 34144 44726 34158
rect 45602 34144 45684 34158
rect 45892 34144 45974 34158
rect 46850 34144 46932 34158
rect 47140 34144 47222 34158
rect 48098 34144 48180 34158
rect 48388 34144 48470 34158
rect 49346 34144 49428 34158
rect 49636 34144 49718 34158
rect 50594 34144 50676 34158
rect 50884 34144 50966 34158
rect 51842 34144 51924 34158
rect 52132 34144 52214 34158
rect 53090 34144 53172 34158
rect 53380 34144 53462 34158
rect 54338 34144 54420 34158
rect 54628 34144 54710 34158
rect 55586 34144 55668 34158
rect 55876 34144 55958 34158
rect 56834 34144 56916 34158
rect 57124 34144 57206 34158
rect 58082 34144 58164 34158
rect 58372 34144 58454 34158
rect 16418 34096 58934 34144
rect 16418 33938 58934 34048
rect 16418 33842 58934 33890
rect 16898 33828 16980 33842
rect 17188 33828 17270 33842
rect 18146 33828 18228 33842
rect 18436 33828 18518 33842
rect 19394 33828 19476 33842
rect 19684 33828 19766 33842
rect 20642 33828 20724 33842
rect 20932 33828 21014 33842
rect 21890 33828 21972 33842
rect 22180 33828 22262 33842
rect 23138 33828 23220 33842
rect 23428 33828 23510 33842
rect 24386 33828 24468 33842
rect 24676 33828 24758 33842
rect 25634 33828 25716 33842
rect 25924 33828 26006 33842
rect 26882 33828 26964 33842
rect 27172 33828 27254 33842
rect 28130 33828 28212 33842
rect 28420 33828 28502 33842
rect 29378 33828 29460 33842
rect 29668 33828 29750 33842
rect 30626 33828 30708 33842
rect 30916 33828 30998 33842
rect 31874 33828 31956 33842
rect 32164 33828 32246 33842
rect 33122 33828 33204 33842
rect 33412 33828 33494 33842
rect 34370 33828 34452 33842
rect 34660 33828 34742 33842
rect 35618 33828 35700 33842
rect 35908 33828 35990 33842
rect 36866 33828 36948 33842
rect 37156 33828 37238 33842
rect 38114 33828 38196 33842
rect 38404 33828 38486 33842
rect 39362 33828 39444 33842
rect 39652 33828 39734 33842
rect 40610 33828 40692 33842
rect 40900 33828 40982 33842
rect 41858 33828 41940 33842
rect 42148 33828 42230 33842
rect 43106 33828 43188 33842
rect 43396 33828 43478 33842
rect 44354 33828 44436 33842
rect 44644 33828 44726 33842
rect 45602 33828 45684 33842
rect 45892 33828 45974 33842
rect 46850 33828 46932 33842
rect 47140 33828 47222 33842
rect 48098 33828 48180 33842
rect 48388 33828 48470 33842
rect 49346 33828 49428 33842
rect 49636 33828 49718 33842
rect 50594 33828 50676 33842
rect 50884 33828 50966 33842
rect 51842 33828 51924 33842
rect 52132 33828 52214 33842
rect 53090 33828 53172 33842
rect 53380 33828 53462 33842
rect 54338 33828 54420 33842
rect 54628 33828 54710 33842
rect 55586 33828 55668 33842
rect 55876 33828 55958 33842
rect 56834 33828 56916 33842
rect 57124 33828 57206 33842
rect 58082 33828 58164 33842
rect 58372 33828 58454 33842
rect 16418 33780 16864 33794
rect 17014 33780 17154 33794
rect 17304 33780 18112 33794
rect 18262 33780 18402 33794
rect 18552 33780 19360 33794
rect 19510 33780 19650 33794
rect 19800 33780 20608 33794
rect 20758 33780 20898 33794
rect 21048 33780 21856 33794
rect 22006 33780 22146 33794
rect 22296 33780 23104 33794
rect 23254 33780 23394 33794
rect 23544 33780 24352 33794
rect 24502 33780 24642 33794
rect 24792 33780 25600 33794
rect 25750 33780 25890 33794
rect 26040 33780 26848 33794
rect 26998 33780 27138 33794
rect 27288 33780 28096 33794
rect 28246 33780 28386 33794
rect 28536 33780 29344 33794
rect 29494 33780 29634 33794
rect 29784 33780 30592 33794
rect 30742 33780 30882 33794
rect 31032 33780 31840 33794
rect 31990 33780 32130 33794
rect 32280 33780 33088 33794
rect 33238 33780 33378 33794
rect 33528 33780 34336 33794
rect 34486 33780 34626 33794
rect 34776 33780 35584 33794
rect 35734 33780 35874 33794
rect 36024 33780 36832 33794
rect 36982 33780 37122 33794
rect 37272 33780 38080 33794
rect 38230 33780 38370 33794
rect 38520 33780 39328 33794
rect 39478 33780 39618 33794
rect 39768 33780 40576 33794
rect 40726 33780 40866 33794
rect 41016 33780 41824 33794
rect 41974 33780 42114 33794
rect 42264 33780 43072 33794
rect 43222 33780 43362 33794
rect 43512 33780 44320 33794
rect 44470 33780 44610 33794
rect 44760 33780 45568 33794
rect 45718 33780 45858 33794
rect 46008 33780 46816 33794
rect 46966 33780 47106 33794
rect 47256 33780 48064 33794
rect 48214 33780 48354 33794
rect 48504 33780 49312 33794
rect 49462 33780 49602 33794
rect 49752 33780 50560 33794
rect 50710 33780 50850 33794
rect 51000 33780 51808 33794
rect 51958 33780 52098 33794
rect 52248 33780 53056 33794
rect 53206 33780 53346 33794
rect 53496 33780 54304 33794
rect 54454 33780 54594 33794
rect 54744 33780 55552 33794
rect 55702 33780 55842 33794
rect 55992 33780 56800 33794
rect 56950 33780 57090 33794
rect 57240 33780 58048 33794
rect 58198 33780 58338 33794
rect 58488 33780 58934 33794
rect 16418 33732 58934 33780
rect 16418 33718 16864 33732
rect 17014 33718 17154 33732
rect 17304 33718 18112 33732
rect 18262 33718 18402 33732
rect 18552 33718 19360 33732
rect 19510 33718 19650 33732
rect 19800 33718 20608 33732
rect 20758 33718 20898 33732
rect 21048 33718 21856 33732
rect 22006 33718 22146 33732
rect 22296 33718 23104 33732
rect 23254 33718 23394 33732
rect 23544 33718 24352 33732
rect 24502 33718 24642 33732
rect 24792 33718 25600 33732
rect 25750 33718 25890 33732
rect 26040 33718 26848 33732
rect 26998 33718 27138 33732
rect 27288 33718 28096 33732
rect 28246 33718 28386 33732
rect 28536 33718 29344 33732
rect 29494 33718 29634 33732
rect 29784 33718 30592 33732
rect 30742 33718 30882 33732
rect 31032 33718 31840 33732
rect 31990 33718 32130 33732
rect 32280 33718 33088 33732
rect 33238 33718 33378 33732
rect 33528 33718 34336 33732
rect 34486 33718 34626 33732
rect 34776 33718 35584 33732
rect 35734 33718 35874 33732
rect 36024 33718 36832 33732
rect 36982 33718 37122 33732
rect 37272 33718 38080 33732
rect 38230 33718 38370 33732
rect 38520 33718 39328 33732
rect 39478 33718 39618 33732
rect 39768 33718 40576 33732
rect 40726 33718 40866 33732
rect 41016 33718 41824 33732
rect 41974 33718 42114 33732
rect 42264 33718 43072 33732
rect 43222 33718 43362 33732
rect 43512 33718 44320 33732
rect 44470 33718 44610 33732
rect 44760 33718 45568 33732
rect 45718 33718 45858 33732
rect 46008 33718 46816 33732
rect 46966 33718 47106 33732
rect 47256 33718 48064 33732
rect 48214 33718 48354 33732
rect 48504 33718 49312 33732
rect 49462 33718 49602 33732
rect 49752 33718 50560 33732
rect 50710 33718 50850 33732
rect 51000 33718 51808 33732
rect 51958 33718 52098 33732
rect 52248 33718 53056 33732
rect 53206 33718 53346 33732
rect 53496 33718 54304 33732
rect 54454 33718 54594 33732
rect 54744 33718 55552 33732
rect 55702 33718 55842 33732
rect 55992 33718 56800 33732
rect 56950 33718 57090 33732
rect 57240 33718 58048 33732
rect 58198 33718 58338 33732
rect 58488 33718 58934 33732
rect 16898 33670 16980 33684
rect 17188 33670 17270 33684
rect 18146 33670 18228 33684
rect 18436 33670 18518 33684
rect 19394 33670 19476 33684
rect 19684 33670 19766 33684
rect 20642 33670 20724 33684
rect 20932 33670 21014 33684
rect 21890 33670 21972 33684
rect 22180 33670 22262 33684
rect 23138 33670 23220 33684
rect 23428 33670 23510 33684
rect 24386 33670 24468 33684
rect 24676 33670 24758 33684
rect 25634 33670 25716 33684
rect 25924 33670 26006 33684
rect 26882 33670 26964 33684
rect 27172 33670 27254 33684
rect 28130 33670 28212 33684
rect 28420 33670 28502 33684
rect 29378 33670 29460 33684
rect 29668 33670 29750 33684
rect 30626 33670 30708 33684
rect 30916 33670 30998 33684
rect 31874 33670 31956 33684
rect 32164 33670 32246 33684
rect 33122 33670 33204 33684
rect 33412 33670 33494 33684
rect 34370 33670 34452 33684
rect 34660 33670 34742 33684
rect 35618 33670 35700 33684
rect 35908 33670 35990 33684
rect 36866 33670 36948 33684
rect 37156 33670 37238 33684
rect 38114 33670 38196 33684
rect 38404 33670 38486 33684
rect 39362 33670 39444 33684
rect 39652 33670 39734 33684
rect 40610 33670 40692 33684
rect 40900 33670 40982 33684
rect 41858 33670 41940 33684
rect 42148 33670 42230 33684
rect 43106 33670 43188 33684
rect 43396 33670 43478 33684
rect 44354 33670 44436 33684
rect 44644 33670 44726 33684
rect 45602 33670 45684 33684
rect 45892 33670 45974 33684
rect 46850 33670 46932 33684
rect 47140 33670 47222 33684
rect 48098 33670 48180 33684
rect 48388 33670 48470 33684
rect 49346 33670 49428 33684
rect 49636 33670 49718 33684
rect 50594 33670 50676 33684
rect 50884 33670 50966 33684
rect 51842 33670 51924 33684
rect 52132 33670 52214 33684
rect 53090 33670 53172 33684
rect 53380 33670 53462 33684
rect 54338 33670 54420 33684
rect 54628 33670 54710 33684
rect 55586 33670 55668 33684
rect 55876 33670 55958 33684
rect 56834 33670 56916 33684
rect 57124 33670 57206 33684
rect 58082 33670 58164 33684
rect 58372 33670 58454 33684
rect 16418 33622 58934 33670
rect 16418 33526 58934 33574
rect 16898 33512 16980 33526
rect 17188 33512 17270 33526
rect 18146 33512 18228 33526
rect 18436 33512 18518 33526
rect 19394 33512 19476 33526
rect 19684 33512 19766 33526
rect 20642 33512 20724 33526
rect 20932 33512 21014 33526
rect 21890 33512 21972 33526
rect 22180 33512 22262 33526
rect 23138 33512 23220 33526
rect 23428 33512 23510 33526
rect 24386 33512 24468 33526
rect 24676 33512 24758 33526
rect 25634 33512 25716 33526
rect 25924 33512 26006 33526
rect 26882 33512 26964 33526
rect 27172 33512 27254 33526
rect 28130 33512 28212 33526
rect 28420 33512 28502 33526
rect 29378 33512 29460 33526
rect 29668 33512 29750 33526
rect 30626 33512 30708 33526
rect 30916 33512 30998 33526
rect 31874 33512 31956 33526
rect 32164 33512 32246 33526
rect 33122 33512 33204 33526
rect 33412 33512 33494 33526
rect 34370 33512 34452 33526
rect 34660 33512 34742 33526
rect 35618 33512 35700 33526
rect 35908 33512 35990 33526
rect 36866 33512 36948 33526
rect 37156 33512 37238 33526
rect 38114 33512 38196 33526
rect 38404 33512 38486 33526
rect 39362 33512 39444 33526
rect 39652 33512 39734 33526
rect 40610 33512 40692 33526
rect 40900 33512 40982 33526
rect 41858 33512 41940 33526
rect 42148 33512 42230 33526
rect 43106 33512 43188 33526
rect 43396 33512 43478 33526
rect 44354 33512 44436 33526
rect 44644 33512 44726 33526
rect 45602 33512 45684 33526
rect 45892 33512 45974 33526
rect 46850 33512 46932 33526
rect 47140 33512 47222 33526
rect 48098 33512 48180 33526
rect 48388 33512 48470 33526
rect 49346 33512 49428 33526
rect 49636 33512 49718 33526
rect 50594 33512 50676 33526
rect 50884 33512 50966 33526
rect 51842 33512 51924 33526
rect 52132 33512 52214 33526
rect 53090 33512 53172 33526
rect 53380 33512 53462 33526
rect 54338 33512 54420 33526
rect 54628 33512 54710 33526
rect 55586 33512 55668 33526
rect 55876 33512 55958 33526
rect 56834 33512 56916 33526
rect 57124 33512 57206 33526
rect 58082 33512 58164 33526
rect 58372 33512 58454 33526
rect 16418 33464 16864 33478
rect 17014 33464 17154 33478
rect 17304 33464 18112 33478
rect 18262 33464 18402 33478
rect 18552 33464 19360 33478
rect 19510 33464 19650 33478
rect 19800 33464 20608 33478
rect 20758 33464 20898 33478
rect 21048 33464 21856 33478
rect 22006 33464 22146 33478
rect 22296 33464 23104 33478
rect 23254 33464 23394 33478
rect 23544 33464 24352 33478
rect 24502 33464 24642 33478
rect 24792 33464 25600 33478
rect 25750 33464 25890 33478
rect 26040 33464 26848 33478
rect 26998 33464 27138 33478
rect 27288 33464 28096 33478
rect 28246 33464 28386 33478
rect 28536 33464 29344 33478
rect 29494 33464 29634 33478
rect 29784 33464 30592 33478
rect 30742 33464 30882 33478
rect 31032 33464 31840 33478
rect 31990 33464 32130 33478
rect 32280 33464 33088 33478
rect 33238 33464 33378 33478
rect 33528 33464 34336 33478
rect 34486 33464 34626 33478
rect 34776 33464 35584 33478
rect 35734 33464 35874 33478
rect 36024 33464 36832 33478
rect 36982 33464 37122 33478
rect 37272 33464 38080 33478
rect 38230 33464 38370 33478
rect 38520 33464 39328 33478
rect 39478 33464 39618 33478
rect 39768 33464 40576 33478
rect 40726 33464 40866 33478
rect 41016 33464 41824 33478
rect 41974 33464 42114 33478
rect 42264 33464 43072 33478
rect 43222 33464 43362 33478
rect 43512 33464 44320 33478
rect 44470 33464 44610 33478
rect 44760 33464 45568 33478
rect 45718 33464 45858 33478
rect 46008 33464 46816 33478
rect 46966 33464 47106 33478
rect 47256 33464 48064 33478
rect 48214 33464 48354 33478
rect 48504 33464 49312 33478
rect 49462 33464 49602 33478
rect 49752 33464 50560 33478
rect 50710 33464 50850 33478
rect 51000 33464 51808 33478
rect 51958 33464 52098 33478
rect 52248 33464 53056 33478
rect 53206 33464 53346 33478
rect 53496 33464 54304 33478
rect 54454 33464 54594 33478
rect 54744 33464 55552 33478
rect 55702 33464 55842 33478
rect 55992 33464 56800 33478
rect 56950 33464 57090 33478
rect 57240 33464 58048 33478
rect 58198 33464 58338 33478
rect 58488 33464 58934 33478
rect 16418 33416 58934 33464
rect 16418 33402 16864 33416
rect 17014 33402 17154 33416
rect 17304 33402 18112 33416
rect 18262 33402 18402 33416
rect 18552 33402 19360 33416
rect 19510 33402 19650 33416
rect 19800 33402 20608 33416
rect 20758 33402 20898 33416
rect 21048 33402 21856 33416
rect 22006 33402 22146 33416
rect 22296 33402 23104 33416
rect 23254 33402 23394 33416
rect 23544 33402 24352 33416
rect 24502 33402 24642 33416
rect 24792 33402 25600 33416
rect 25750 33402 25890 33416
rect 26040 33402 26848 33416
rect 26998 33402 27138 33416
rect 27288 33402 28096 33416
rect 28246 33402 28386 33416
rect 28536 33402 29344 33416
rect 29494 33402 29634 33416
rect 29784 33402 30592 33416
rect 30742 33402 30882 33416
rect 31032 33402 31840 33416
rect 31990 33402 32130 33416
rect 32280 33402 33088 33416
rect 33238 33402 33378 33416
rect 33528 33402 34336 33416
rect 34486 33402 34626 33416
rect 34776 33402 35584 33416
rect 35734 33402 35874 33416
rect 36024 33402 36832 33416
rect 36982 33402 37122 33416
rect 37272 33402 38080 33416
rect 38230 33402 38370 33416
rect 38520 33402 39328 33416
rect 39478 33402 39618 33416
rect 39768 33402 40576 33416
rect 40726 33402 40866 33416
rect 41016 33402 41824 33416
rect 41974 33402 42114 33416
rect 42264 33402 43072 33416
rect 43222 33402 43362 33416
rect 43512 33402 44320 33416
rect 44470 33402 44610 33416
rect 44760 33402 45568 33416
rect 45718 33402 45858 33416
rect 46008 33402 46816 33416
rect 46966 33402 47106 33416
rect 47256 33402 48064 33416
rect 48214 33402 48354 33416
rect 48504 33402 49312 33416
rect 49462 33402 49602 33416
rect 49752 33402 50560 33416
rect 50710 33402 50850 33416
rect 51000 33402 51808 33416
rect 51958 33402 52098 33416
rect 52248 33402 53056 33416
rect 53206 33402 53346 33416
rect 53496 33402 54304 33416
rect 54454 33402 54594 33416
rect 54744 33402 55552 33416
rect 55702 33402 55842 33416
rect 55992 33402 56800 33416
rect 56950 33402 57090 33416
rect 57240 33402 58048 33416
rect 58198 33402 58338 33416
rect 58488 33402 58934 33416
rect 16898 33354 16980 33368
rect 17188 33354 17270 33368
rect 18146 33354 18228 33368
rect 18436 33354 18518 33368
rect 19394 33354 19476 33368
rect 19684 33354 19766 33368
rect 20642 33354 20724 33368
rect 20932 33354 21014 33368
rect 21890 33354 21972 33368
rect 22180 33354 22262 33368
rect 23138 33354 23220 33368
rect 23428 33354 23510 33368
rect 24386 33354 24468 33368
rect 24676 33354 24758 33368
rect 25634 33354 25716 33368
rect 25924 33354 26006 33368
rect 26882 33354 26964 33368
rect 27172 33354 27254 33368
rect 28130 33354 28212 33368
rect 28420 33354 28502 33368
rect 29378 33354 29460 33368
rect 29668 33354 29750 33368
rect 30626 33354 30708 33368
rect 30916 33354 30998 33368
rect 31874 33354 31956 33368
rect 32164 33354 32246 33368
rect 33122 33354 33204 33368
rect 33412 33354 33494 33368
rect 34370 33354 34452 33368
rect 34660 33354 34742 33368
rect 35618 33354 35700 33368
rect 35908 33354 35990 33368
rect 36866 33354 36948 33368
rect 37156 33354 37238 33368
rect 38114 33354 38196 33368
rect 38404 33354 38486 33368
rect 39362 33354 39444 33368
rect 39652 33354 39734 33368
rect 40610 33354 40692 33368
rect 40900 33354 40982 33368
rect 41858 33354 41940 33368
rect 42148 33354 42230 33368
rect 43106 33354 43188 33368
rect 43396 33354 43478 33368
rect 44354 33354 44436 33368
rect 44644 33354 44726 33368
rect 45602 33354 45684 33368
rect 45892 33354 45974 33368
rect 46850 33354 46932 33368
rect 47140 33354 47222 33368
rect 48098 33354 48180 33368
rect 48388 33354 48470 33368
rect 49346 33354 49428 33368
rect 49636 33354 49718 33368
rect 50594 33354 50676 33368
rect 50884 33354 50966 33368
rect 51842 33354 51924 33368
rect 52132 33354 52214 33368
rect 53090 33354 53172 33368
rect 53380 33354 53462 33368
rect 54338 33354 54420 33368
rect 54628 33354 54710 33368
rect 55586 33354 55668 33368
rect 55876 33354 55958 33368
rect 56834 33354 56916 33368
rect 57124 33354 57206 33368
rect 58082 33354 58164 33368
rect 58372 33354 58454 33368
rect 16418 33306 58934 33354
rect 16418 33148 58934 33258
rect 16418 33052 58934 33100
rect 16898 33038 16980 33052
rect 17188 33038 17270 33052
rect 18146 33038 18228 33052
rect 18436 33038 18518 33052
rect 19394 33038 19476 33052
rect 19684 33038 19766 33052
rect 20642 33038 20724 33052
rect 20932 33038 21014 33052
rect 21890 33038 21972 33052
rect 22180 33038 22262 33052
rect 23138 33038 23220 33052
rect 23428 33038 23510 33052
rect 24386 33038 24468 33052
rect 24676 33038 24758 33052
rect 25634 33038 25716 33052
rect 25924 33038 26006 33052
rect 26882 33038 26964 33052
rect 27172 33038 27254 33052
rect 28130 33038 28212 33052
rect 28420 33038 28502 33052
rect 29378 33038 29460 33052
rect 29668 33038 29750 33052
rect 30626 33038 30708 33052
rect 30916 33038 30998 33052
rect 31874 33038 31956 33052
rect 32164 33038 32246 33052
rect 33122 33038 33204 33052
rect 33412 33038 33494 33052
rect 34370 33038 34452 33052
rect 34660 33038 34742 33052
rect 35618 33038 35700 33052
rect 35908 33038 35990 33052
rect 36866 33038 36948 33052
rect 37156 33038 37238 33052
rect 38114 33038 38196 33052
rect 38404 33038 38486 33052
rect 39362 33038 39444 33052
rect 39652 33038 39734 33052
rect 40610 33038 40692 33052
rect 40900 33038 40982 33052
rect 41858 33038 41940 33052
rect 42148 33038 42230 33052
rect 43106 33038 43188 33052
rect 43396 33038 43478 33052
rect 44354 33038 44436 33052
rect 44644 33038 44726 33052
rect 45602 33038 45684 33052
rect 45892 33038 45974 33052
rect 46850 33038 46932 33052
rect 47140 33038 47222 33052
rect 48098 33038 48180 33052
rect 48388 33038 48470 33052
rect 49346 33038 49428 33052
rect 49636 33038 49718 33052
rect 50594 33038 50676 33052
rect 50884 33038 50966 33052
rect 51842 33038 51924 33052
rect 52132 33038 52214 33052
rect 53090 33038 53172 33052
rect 53380 33038 53462 33052
rect 54338 33038 54420 33052
rect 54628 33038 54710 33052
rect 55586 33038 55668 33052
rect 55876 33038 55958 33052
rect 56834 33038 56916 33052
rect 57124 33038 57206 33052
rect 58082 33038 58164 33052
rect 58372 33038 58454 33052
rect 16418 32990 16864 33004
rect 17014 32990 17154 33004
rect 17304 32990 18112 33004
rect 18262 32990 18402 33004
rect 18552 32990 19360 33004
rect 19510 32990 19650 33004
rect 19800 32990 20608 33004
rect 20758 32990 20898 33004
rect 21048 32990 21856 33004
rect 22006 32990 22146 33004
rect 22296 32990 23104 33004
rect 23254 32990 23394 33004
rect 23544 32990 24352 33004
rect 24502 32990 24642 33004
rect 24792 32990 25600 33004
rect 25750 32990 25890 33004
rect 26040 32990 26848 33004
rect 26998 32990 27138 33004
rect 27288 32990 28096 33004
rect 28246 32990 28386 33004
rect 28536 32990 29344 33004
rect 29494 32990 29634 33004
rect 29784 32990 30592 33004
rect 30742 32990 30882 33004
rect 31032 32990 31840 33004
rect 31990 32990 32130 33004
rect 32280 32990 33088 33004
rect 33238 32990 33378 33004
rect 33528 32990 34336 33004
rect 34486 32990 34626 33004
rect 34776 32990 35584 33004
rect 35734 32990 35874 33004
rect 36024 32990 36832 33004
rect 36982 32990 37122 33004
rect 37272 32990 38080 33004
rect 38230 32990 38370 33004
rect 38520 32990 39328 33004
rect 39478 32990 39618 33004
rect 39768 32990 40576 33004
rect 40726 32990 40866 33004
rect 41016 32990 41824 33004
rect 41974 32990 42114 33004
rect 42264 32990 43072 33004
rect 43222 32990 43362 33004
rect 43512 32990 44320 33004
rect 44470 32990 44610 33004
rect 44760 32990 45568 33004
rect 45718 32990 45858 33004
rect 46008 32990 46816 33004
rect 46966 32990 47106 33004
rect 47256 32990 48064 33004
rect 48214 32990 48354 33004
rect 48504 32990 49312 33004
rect 49462 32990 49602 33004
rect 49752 32990 50560 33004
rect 50710 32990 50850 33004
rect 51000 32990 51808 33004
rect 51958 32990 52098 33004
rect 52248 32990 53056 33004
rect 53206 32990 53346 33004
rect 53496 32990 54304 33004
rect 54454 32990 54594 33004
rect 54744 32990 55552 33004
rect 55702 32990 55842 33004
rect 55992 32990 56800 33004
rect 56950 32990 57090 33004
rect 57240 32990 58048 33004
rect 58198 32990 58338 33004
rect 58488 32990 58934 33004
rect 16418 32942 58934 32990
rect 16418 32928 16864 32942
rect 17014 32928 17154 32942
rect 17304 32928 18112 32942
rect 18262 32928 18402 32942
rect 18552 32928 19360 32942
rect 19510 32928 19650 32942
rect 19800 32928 20608 32942
rect 20758 32928 20898 32942
rect 21048 32928 21856 32942
rect 22006 32928 22146 32942
rect 22296 32928 23104 32942
rect 23254 32928 23394 32942
rect 23544 32928 24352 32942
rect 24502 32928 24642 32942
rect 24792 32928 25600 32942
rect 25750 32928 25890 32942
rect 26040 32928 26848 32942
rect 26998 32928 27138 32942
rect 27288 32928 28096 32942
rect 28246 32928 28386 32942
rect 28536 32928 29344 32942
rect 29494 32928 29634 32942
rect 29784 32928 30592 32942
rect 30742 32928 30882 32942
rect 31032 32928 31840 32942
rect 31990 32928 32130 32942
rect 32280 32928 33088 32942
rect 33238 32928 33378 32942
rect 33528 32928 34336 32942
rect 34486 32928 34626 32942
rect 34776 32928 35584 32942
rect 35734 32928 35874 32942
rect 36024 32928 36832 32942
rect 36982 32928 37122 32942
rect 37272 32928 38080 32942
rect 38230 32928 38370 32942
rect 38520 32928 39328 32942
rect 39478 32928 39618 32942
rect 39768 32928 40576 32942
rect 40726 32928 40866 32942
rect 41016 32928 41824 32942
rect 41974 32928 42114 32942
rect 42264 32928 43072 32942
rect 43222 32928 43362 32942
rect 43512 32928 44320 32942
rect 44470 32928 44610 32942
rect 44760 32928 45568 32942
rect 45718 32928 45858 32942
rect 46008 32928 46816 32942
rect 46966 32928 47106 32942
rect 47256 32928 48064 32942
rect 48214 32928 48354 32942
rect 48504 32928 49312 32942
rect 49462 32928 49602 32942
rect 49752 32928 50560 32942
rect 50710 32928 50850 32942
rect 51000 32928 51808 32942
rect 51958 32928 52098 32942
rect 52248 32928 53056 32942
rect 53206 32928 53346 32942
rect 53496 32928 54304 32942
rect 54454 32928 54594 32942
rect 54744 32928 55552 32942
rect 55702 32928 55842 32942
rect 55992 32928 56800 32942
rect 56950 32928 57090 32942
rect 57240 32928 58048 32942
rect 58198 32928 58338 32942
rect 58488 32928 58934 32942
rect 16898 32880 16980 32894
rect 17188 32880 17270 32894
rect 18146 32880 18228 32894
rect 18436 32880 18518 32894
rect 19394 32880 19476 32894
rect 19684 32880 19766 32894
rect 20642 32880 20724 32894
rect 20932 32880 21014 32894
rect 21890 32880 21972 32894
rect 22180 32880 22262 32894
rect 23138 32880 23220 32894
rect 23428 32880 23510 32894
rect 24386 32880 24468 32894
rect 24676 32880 24758 32894
rect 25634 32880 25716 32894
rect 25924 32880 26006 32894
rect 26882 32880 26964 32894
rect 27172 32880 27254 32894
rect 28130 32880 28212 32894
rect 28420 32880 28502 32894
rect 29378 32880 29460 32894
rect 29668 32880 29750 32894
rect 30626 32880 30708 32894
rect 30916 32880 30998 32894
rect 31874 32880 31956 32894
rect 32164 32880 32246 32894
rect 33122 32880 33204 32894
rect 33412 32880 33494 32894
rect 34370 32880 34452 32894
rect 34660 32880 34742 32894
rect 35618 32880 35700 32894
rect 35908 32880 35990 32894
rect 36866 32880 36948 32894
rect 37156 32880 37238 32894
rect 38114 32880 38196 32894
rect 38404 32880 38486 32894
rect 39362 32880 39444 32894
rect 39652 32880 39734 32894
rect 40610 32880 40692 32894
rect 40900 32880 40982 32894
rect 41858 32880 41940 32894
rect 42148 32880 42230 32894
rect 43106 32880 43188 32894
rect 43396 32880 43478 32894
rect 44354 32880 44436 32894
rect 44644 32880 44726 32894
rect 45602 32880 45684 32894
rect 45892 32880 45974 32894
rect 46850 32880 46932 32894
rect 47140 32880 47222 32894
rect 48098 32880 48180 32894
rect 48388 32880 48470 32894
rect 49346 32880 49428 32894
rect 49636 32880 49718 32894
rect 50594 32880 50676 32894
rect 50884 32880 50966 32894
rect 51842 32880 51924 32894
rect 52132 32880 52214 32894
rect 53090 32880 53172 32894
rect 53380 32880 53462 32894
rect 54338 32880 54420 32894
rect 54628 32880 54710 32894
rect 55586 32880 55668 32894
rect 55876 32880 55958 32894
rect 56834 32880 56916 32894
rect 57124 32880 57206 32894
rect 58082 32880 58164 32894
rect 58372 32880 58454 32894
rect 16418 32832 58934 32880
rect 16418 32736 58934 32784
rect 16898 32722 16980 32736
rect 17188 32722 17270 32736
rect 18146 32722 18228 32736
rect 18436 32722 18518 32736
rect 19394 32722 19476 32736
rect 19684 32722 19766 32736
rect 20642 32722 20724 32736
rect 20932 32722 21014 32736
rect 21890 32722 21972 32736
rect 22180 32722 22262 32736
rect 23138 32722 23220 32736
rect 23428 32722 23510 32736
rect 24386 32722 24468 32736
rect 24676 32722 24758 32736
rect 25634 32722 25716 32736
rect 25924 32722 26006 32736
rect 26882 32722 26964 32736
rect 27172 32722 27254 32736
rect 28130 32722 28212 32736
rect 28420 32722 28502 32736
rect 29378 32722 29460 32736
rect 29668 32722 29750 32736
rect 30626 32722 30708 32736
rect 30916 32722 30998 32736
rect 31874 32722 31956 32736
rect 32164 32722 32246 32736
rect 33122 32722 33204 32736
rect 33412 32722 33494 32736
rect 34370 32722 34452 32736
rect 34660 32722 34742 32736
rect 35618 32722 35700 32736
rect 35908 32722 35990 32736
rect 36866 32722 36948 32736
rect 37156 32722 37238 32736
rect 38114 32722 38196 32736
rect 38404 32722 38486 32736
rect 39362 32722 39444 32736
rect 39652 32722 39734 32736
rect 40610 32722 40692 32736
rect 40900 32722 40982 32736
rect 41858 32722 41940 32736
rect 42148 32722 42230 32736
rect 43106 32722 43188 32736
rect 43396 32722 43478 32736
rect 44354 32722 44436 32736
rect 44644 32722 44726 32736
rect 45602 32722 45684 32736
rect 45892 32722 45974 32736
rect 46850 32722 46932 32736
rect 47140 32722 47222 32736
rect 48098 32722 48180 32736
rect 48388 32722 48470 32736
rect 49346 32722 49428 32736
rect 49636 32722 49718 32736
rect 50594 32722 50676 32736
rect 50884 32722 50966 32736
rect 51842 32722 51924 32736
rect 52132 32722 52214 32736
rect 53090 32722 53172 32736
rect 53380 32722 53462 32736
rect 54338 32722 54420 32736
rect 54628 32722 54710 32736
rect 55586 32722 55668 32736
rect 55876 32722 55958 32736
rect 56834 32722 56916 32736
rect 57124 32722 57206 32736
rect 58082 32722 58164 32736
rect 58372 32722 58454 32736
rect 16418 32674 16864 32688
rect 17014 32674 17154 32688
rect 17304 32674 18112 32688
rect 18262 32674 18402 32688
rect 18552 32674 19360 32688
rect 19510 32674 19650 32688
rect 19800 32674 20608 32688
rect 20758 32674 20898 32688
rect 21048 32674 21856 32688
rect 22006 32674 22146 32688
rect 22296 32674 23104 32688
rect 23254 32674 23394 32688
rect 23544 32674 24352 32688
rect 24502 32674 24642 32688
rect 24792 32674 25600 32688
rect 25750 32674 25890 32688
rect 26040 32674 26848 32688
rect 26998 32674 27138 32688
rect 27288 32674 28096 32688
rect 28246 32674 28386 32688
rect 28536 32674 29344 32688
rect 29494 32674 29634 32688
rect 29784 32674 30592 32688
rect 30742 32674 30882 32688
rect 31032 32674 31840 32688
rect 31990 32674 32130 32688
rect 32280 32674 33088 32688
rect 33238 32674 33378 32688
rect 33528 32674 34336 32688
rect 34486 32674 34626 32688
rect 34776 32674 35584 32688
rect 35734 32674 35874 32688
rect 36024 32674 36832 32688
rect 36982 32674 37122 32688
rect 37272 32674 38080 32688
rect 38230 32674 38370 32688
rect 38520 32674 39328 32688
rect 39478 32674 39618 32688
rect 39768 32674 40576 32688
rect 40726 32674 40866 32688
rect 41016 32674 41824 32688
rect 41974 32674 42114 32688
rect 42264 32674 43072 32688
rect 43222 32674 43362 32688
rect 43512 32674 44320 32688
rect 44470 32674 44610 32688
rect 44760 32674 45568 32688
rect 45718 32674 45858 32688
rect 46008 32674 46816 32688
rect 46966 32674 47106 32688
rect 47256 32674 48064 32688
rect 48214 32674 48354 32688
rect 48504 32674 49312 32688
rect 49462 32674 49602 32688
rect 49752 32674 50560 32688
rect 50710 32674 50850 32688
rect 51000 32674 51808 32688
rect 51958 32674 52098 32688
rect 52248 32674 53056 32688
rect 53206 32674 53346 32688
rect 53496 32674 54304 32688
rect 54454 32674 54594 32688
rect 54744 32674 55552 32688
rect 55702 32674 55842 32688
rect 55992 32674 56800 32688
rect 56950 32674 57090 32688
rect 57240 32674 58048 32688
rect 58198 32674 58338 32688
rect 58488 32674 58934 32688
rect 16418 32626 58934 32674
rect 16418 32612 16864 32626
rect 17014 32612 17154 32626
rect 17304 32612 18112 32626
rect 18262 32612 18402 32626
rect 18552 32612 19360 32626
rect 19510 32612 19650 32626
rect 19800 32612 20608 32626
rect 20758 32612 20898 32626
rect 21048 32612 21856 32626
rect 22006 32612 22146 32626
rect 22296 32612 23104 32626
rect 23254 32612 23394 32626
rect 23544 32612 24352 32626
rect 24502 32612 24642 32626
rect 24792 32612 25600 32626
rect 25750 32612 25890 32626
rect 26040 32612 26848 32626
rect 26998 32612 27138 32626
rect 27288 32612 28096 32626
rect 28246 32612 28386 32626
rect 28536 32612 29344 32626
rect 29494 32612 29634 32626
rect 29784 32612 30592 32626
rect 30742 32612 30882 32626
rect 31032 32612 31840 32626
rect 31990 32612 32130 32626
rect 32280 32612 33088 32626
rect 33238 32612 33378 32626
rect 33528 32612 34336 32626
rect 34486 32612 34626 32626
rect 34776 32612 35584 32626
rect 35734 32612 35874 32626
rect 36024 32612 36832 32626
rect 36982 32612 37122 32626
rect 37272 32612 38080 32626
rect 38230 32612 38370 32626
rect 38520 32612 39328 32626
rect 39478 32612 39618 32626
rect 39768 32612 40576 32626
rect 40726 32612 40866 32626
rect 41016 32612 41824 32626
rect 41974 32612 42114 32626
rect 42264 32612 43072 32626
rect 43222 32612 43362 32626
rect 43512 32612 44320 32626
rect 44470 32612 44610 32626
rect 44760 32612 45568 32626
rect 45718 32612 45858 32626
rect 46008 32612 46816 32626
rect 46966 32612 47106 32626
rect 47256 32612 48064 32626
rect 48214 32612 48354 32626
rect 48504 32612 49312 32626
rect 49462 32612 49602 32626
rect 49752 32612 50560 32626
rect 50710 32612 50850 32626
rect 51000 32612 51808 32626
rect 51958 32612 52098 32626
rect 52248 32612 53056 32626
rect 53206 32612 53346 32626
rect 53496 32612 54304 32626
rect 54454 32612 54594 32626
rect 54744 32612 55552 32626
rect 55702 32612 55842 32626
rect 55992 32612 56800 32626
rect 56950 32612 57090 32626
rect 57240 32612 58048 32626
rect 58198 32612 58338 32626
rect 58488 32612 58934 32626
rect 16898 32564 16980 32578
rect 17188 32564 17270 32578
rect 18146 32564 18228 32578
rect 18436 32564 18518 32578
rect 19394 32564 19476 32578
rect 19684 32564 19766 32578
rect 20642 32564 20724 32578
rect 20932 32564 21014 32578
rect 21890 32564 21972 32578
rect 22180 32564 22262 32578
rect 23138 32564 23220 32578
rect 23428 32564 23510 32578
rect 24386 32564 24468 32578
rect 24676 32564 24758 32578
rect 25634 32564 25716 32578
rect 25924 32564 26006 32578
rect 26882 32564 26964 32578
rect 27172 32564 27254 32578
rect 28130 32564 28212 32578
rect 28420 32564 28502 32578
rect 29378 32564 29460 32578
rect 29668 32564 29750 32578
rect 30626 32564 30708 32578
rect 30916 32564 30998 32578
rect 31874 32564 31956 32578
rect 32164 32564 32246 32578
rect 33122 32564 33204 32578
rect 33412 32564 33494 32578
rect 34370 32564 34452 32578
rect 34660 32564 34742 32578
rect 35618 32564 35700 32578
rect 35908 32564 35990 32578
rect 36866 32564 36948 32578
rect 37156 32564 37238 32578
rect 38114 32564 38196 32578
rect 38404 32564 38486 32578
rect 39362 32564 39444 32578
rect 39652 32564 39734 32578
rect 40610 32564 40692 32578
rect 40900 32564 40982 32578
rect 41858 32564 41940 32578
rect 42148 32564 42230 32578
rect 43106 32564 43188 32578
rect 43396 32564 43478 32578
rect 44354 32564 44436 32578
rect 44644 32564 44726 32578
rect 45602 32564 45684 32578
rect 45892 32564 45974 32578
rect 46850 32564 46932 32578
rect 47140 32564 47222 32578
rect 48098 32564 48180 32578
rect 48388 32564 48470 32578
rect 49346 32564 49428 32578
rect 49636 32564 49718 32578
rect 50594 32564 50676 32578
rect 50884 32564 50966 32578
rect 51842 32564 51924 32578
rect 52132 32564 52214 32578
rect 53090 32564 53172 32578
rect 53380 32564 53462 32578
rect 54338 32564 54420 32578
rect 54628 32564 54710 32578
rect 55586 32564 55668 32578
rect 55876 32564 55958 32578
rect 56834 32564 56916 32578
rect 57124 32564 57206 32578
rect 58082 32564 58164 32578
rect 58372 32564 58454 32578
rect 16418 32516 58934 32564
rect 16418 32358 58934 32468
rect 16418 32262 58934 32310
rect 16898 32248 16980 32262
rect 17188 32248 17270 32262
rect 18146 32248 18228 32262
rect 18436 32248 18518 32262
rect 19394 32248 19476 32262
rect 19684 32248 19766 32262
rect 20642 32248 20724 32262
rect 20932 32248 21014 32262
rect 21890 32248 21972 32262
rect 22180 32248 22262 32262
rect 23138 32248 23220 32262
rect 23428 32248 23510 32262
rect 24386 32248 24468 32262
rect 24676 32248 24758 32262
rect 25634 32248 25716 32262
rect 25924 32248 26006 32262
rect 26882 32248 26964 32262
rect 27172 32248 27254 32262
rect 28130 32248 28212 32262
rect 28420 32248 28502 32262
rect 29378 32248 29460 32262
rect 29668 32248 29750 32262
rect 30626 32248 30708 32262
rect 30916 32248 30998 32262
rect 31874 32248 31956 32262
rect 32164 32248 32246 32262
rect 33122 32248 33204 32262
rect 33412 32248 33494 32262
rect 34370 32248 34452 32262
rect 34660 32248 34742 32262
rect 35618 32248 35700 32262
rect 35908 32248 35990 32262
rect 36866 32248 36948 32262
rect 37156 32248 37238 32262
rect 38114 32248 38196 32262
rect 38404 32248 38486 32262
rect 39362 32248 39444 32262
rect 39652 32248 39734 32262
rect 40610 32248 40692 32262
rect 40900 32248 40982 32262
rect 41858 32248 41940 32262
rect 42148 32248 42230 32262
rect 43106 32248 43188 32262
rect 43396 32248 43478 32262
rect 44354 32248 44436 32262
rect 44644 32248 44726 32262
rect 45602 32248 45684 32262
rect 45892 32248 45974 32262
rect 46850 32248 46932 32262
rect 47140 32248 47222 32262
rect 48098 32248 48180 32262
rect 48388 32248 48470 32262
rect 49346 32248 49428 32262
rect 49636 32248 49718 32262
rect 50594 32248 50676 32262
rect 50884 32248 50966 32262
rect 51842 32248 51924 32262
rect 52132 32248 52214 32262
rect 53090 32248 53172 32262
rect 53380 32248 53462 32262
rect 54338 32248 54420 32262
rect 54628 32248 54710 32262
rect 55586 32248 55668 32262
rect 55876 32248 55958 32262
rect 56834 32248 56916 32262
rect 57124 32248 57206 32262
rect 58082 32248 58164 32262
rect 58372 32248 58454 32262
rect 16418 32200 16864 32214
rect 17014 32200 17154 32214
rect 17304 32200 18112 32214
rect 18262 32200 18402 32214
rect 18552 32200 19360 32214
rect 19510 32200 19650 32214
rect 19800 32200 20608 32214
rect 20758 32200 20898 32214
rect 21048 32200 21856 32214
rect 22006 32200 22146 32214
rect 22296 32200 23104 32214
rect 23254 32200 23394 32214
rect 23544 32200 24352 32214
rect 24502 32200 24642 32214
rect 24792 32200 25600 32214
rect 25750 32200 25890 32214
rect 26040 32200 26848 32214
rect 26998 32200 27138 32214
rect 27288 32200 28096 32214
rect 28246 32200 28386 32214
rect 28536 32200 29344 32214
rect 29494 32200 29634 32214
rect 29784 32200 30592 32214
rect 30742 32200 30882 32214
rect 31032 32200 31840 32214
rect 31990 32200 32130 32214
rect 32280 32200 33088 32214
rect 33238 32200 33378 32214
rect 33528 32200 34336 32214
rect 34486 32200 34626 32214
rect 34776 32200 35584 32214
rect 35734 32200 35874 32214
rect 36024 32200 36832 32214
rect 36982 32200 37122 32214
rect 37272 32200 38080 32214
rect 38230 32200 38370 32214
rect 38520 32200 39328 32214
rect 39478 32200 39618 32214
rect 39768 32200 40576 32214
rect 40726 32200 40866 32214
rect 41016 32200 41824 32214
rect 41974 32200 42114 32214
rect 42264 32200 43072 32214
rect 43222 32200 43362 32214
rect 43512 32200 44320 32214
rect 44470 32200 44610 32214
rect 44760 32200 45568 32214
rect 45718 32200 45858 32214
rect 46008 32200 46816 32214
rect 46966 32200 47106 32214
rect 47256 32200 48064 32214
rect 48214 32200 48354 32214
rect 48504 32200 49312 32214
rect 49462 32200 49602 32214
rect 49752 32200 50560 32214
rect 50710 32200 50850 32214
rect 51000 32200 51808 32214
rect 51958 32200 52098 32214
rect 52248 32200 53056 32214
rect 53206 32200 53346 32214
rect 53496 32200 54304 32214
rect 54454 32200 54594 32214
rect 54744 32200 55552 32214
rect 55702 32200 55842 32214
rect 55992 32200 56800 32214
rect 56950 32200 57090 32214
rect 57240 32200 58048 32214
rect 58198 32200 58338 32214
rect 58488 32200 58934 32214
rect 16418 32152 58934 32200
rect 16418 32138 16864 32152
rect 17014 32138 17154 32152
rect 17304 32138 18112 32152
rect 18262 32138 18402 32152
rect 18552 32138 19360 32152
rect 19510 32138 19650 32152
rect 19800 32138 20608 32152
rect 20758 32138 20898 32152
rect 21048 32138 21856 32152
rect 22006 32138 22146 32152
rect 22296 32138 23104 32152
rect 23254 32138 23394 32152
rect 23544 32138 24352 32152
rect 24502 32138 24642 32152
rect 24792 32138 25600 32152
rect 25750 32138 25890 32152
rect 26040 32138 26848 32152
rect 26998 32138 27138 32152
rect 27288 32138 28096 32152
rect 28246 32138 28386 32152
rect 28536 32138 29344 32152
rect 29494 32138 29634 32152
rect 29784 32138 30592 32152
rect 30742 32138 30882 32152
rect 31032 32138 31840 32152
rect 31990 32138 32130 32152
rect 32280 32138 33088 32152
rect 33238 32138 33378 32152
rect 33528 32138 34336 32152
rect 34486 32138 34626 32152
rect 34776 32138 35584 32152
rect 35734 32138 35874 32152
rect 36024 32138 36832 32152
rect 36982 32138 37122 32152
rect 37272 32138 38080 32152
rect 38230 32138 38370 32152
rect 38520 32138 39328 32152
rect 39478 32138 39618 32152
rect 39768 32138 40576 32152
rect 40726 32138 40866 32152
rect 41016 32138 41824 32152
rect 41974 32138 42114 32152
rect 42264 32138 43072 32152
rect 43222 32138 43362 32152
rect 43512 32138 44320 32152
rect 44470 32138 44610 32152
rect 44760 32138 45568 32152
rect 45718 32138 45858 32152
rect 46008 32138 46816 32152
rect 46966 32138 47106 32152
rect 47256 32138 48064 32152
rect 48214 32138 48354 32152
rect 48504 32138 49312 32152
rect 49462 32138 49602 32152
rect 49752 32138 50560 32152
rect 50710 32138 50850 32152
rect 51000 32138 51808 32152
rect 51958 32138 52098 32152
rect 52248 32138 53056 32152
rect 53206 32138 53346 32152
rect 53496 32138 54304 32152
rect 54454 32138 54594 32152
rect 54744 32138 55552 32152
rect 55702 32138 55842 32152
rect 55992 32138 56800 32152
rect 56950 32138 57090 32152
rect 57240 32138 58048 32152
rect 58198 32138 58338 32152
rect 58488 32138 58934 32152
rect 16898 32090 16980 32104
rect 17188 32090 17270 32104
rect 18146 32090 18228 32104
rect 18436 32090 18518 32104
rect 19394 32090 19476 32104
rect 19684 32090 19766 32104
rect 20642 32090 20724 32104
rect 20932 32090 21014 32104
rect 21890 32090 21972 32104
rect 22180 32090 22262 32104
rect 23138 32090 23220 32104
rect 23428 32090 23510 32104
rect 24386 32090 24468 32104
rect 24676 32090 24758 32104
rect 25634 32090 25716 32104
rect 25924 32090 26006 32104
rect 26882 32090 26964 32104
rect 27172 32090 27254 32104
rect 28130 32090 28212 32104
rect 28420 32090 28502 32104
rect 29378 32090 29460 32104
rect 29668 32090 29750 32104
rect 30626 32090 30708 32104
rect 30916 32090 30998 32104
rect 31874 32090 31956 32104
rect 32164 32090 32246 32104
rect 33122 32090 33204 32104
rect 33412 32090 33494 32104
rect 34370 32090 34452 32104
rect 34660 32090 34742 32104
rect 35618 32090 35700 32104
rect 35908 32090 35990 32104
rect 36866 32090 36948 32104
rect 37156 32090 37238 32104
rect 38114 32090 38196 32104
rect 38404 32090 38486 32104
rect 39362 32090 39444 32104
rect 39652 32090 39734 32104
rect 40610 32090 40692 32104
rect 40900 32090 40982 32104
rect 41858 32090 41940 32104
rect 42148 32090 42230 32104
rect 43106 32090 43188 32104
rect 43396 32090 43478 32104
rect 44354 32090 44436 32104
rect 44644 32090 44726 32104
rect 45602 32090 45684 32104
rect 45892 32090 45974 32104
rect 46850 32090 46932 32104
rect 47140 32090 47222 32104
rect 48098 32090 48180 32104
rect 48388 32090 48470 32104
rect 49346 32090 49428 32104
rect 49636 32090 49718 32104
rect 50594 32090 50676 32104
rect 50884 32090 50966 32104
rect 51842 32090 51924 32104
rect 52132 32090 52214 32104
rect 53090 32090 53172 32104
rect 53380 32090 53462 32104
rect 54338 32090 54420 32104
rect 54628 32090 54710 32104
rect 55586 32090 55668 32104
rect 55876 32090 55958 32104
rect 56834 32090 56916 32104
rect 57124 32090 57206 32104
rect 58082 32090 58164 32104
rect 58372 32090 58454 32104
rect 16418 32042 58934 32090
rect 16418 31946 58934 31994
rect 16898 31932 16980 31946
rect 17188 31932 17270 31946
rect 18146 31932 18228 31946
rect 18436 31932 18518 31946
rect 19394 31932 19476 31946
rect 19684 31932 19766 31946
rect 20642 31932 20724 31946
rect 20932 31932 21014 31946
rect 21890 31932 21972 31946
rect 22180 31932 22262 31946
rect 23138 31932 23220 31946
rect 23428 31932 23510 31946
rect 24386 31932 24468 31946
rect 24676 31932 24758 31946
rect 25634 31932 25716 31946
rect 25924 31932 26006 31946
rect 26882 31932 26964 31946
rect 27172 31932 27254 31946
rect 28130 31932 28212 31946
rect 28420 31932 28502 31946
rect 29378 31932 29460 31946
rect 29668 31932 29750 31946
rect 30626 31932 30708 31946
rect 30916 31932 30998 31946
rect 31874 31932 31956 31946
rect 32164 31932 32246 31946
rect 33122 31932 33204 31946
rect 33412 31932 33494 31946
rect 34370 31932 34452 31946
rect 34660 31932 34742 31946
rect 35618 31932 35700 31946
rect 35908 31932 35990 31946
rect 36866 31932 36948 31946
rect 37156 31932 37238 31946
rect 38114 31932 38196 31946
rect 38404 31932 38486 31946
rect 39362 31932 39444 31946
rect 39652 31932 39734 31946
rect 40610 31932 40692 31946
rect 40900 31932 40982 31946
rect 41858 31932 41940 31946
rect 42148 31932 42230 31946
rect 43106 31932 43188 31946
rect 43396 31932 43478 31946
rect 44354 31932 44436 31946
rect 44644 31932 44726 31946
rect 45602 31932 45684 31946
rect 45892 31932 45974 31946
rect 46850 31932 46932 31946
rect 47140 31932 47222 31946
rect 48098 31932 48180 31946
rect 48388 31932 48470 31946
rect 49346 31932 49428 31946
rect 49636 31932 49718 31946
rect 50594 31932 50676 31946
rect 50884 31932 50966 31946
rect 51842 31932 51924 31946
rect 52132 31932 52214 31946
rect 53090 31932 53172 31946
rect 53380 31932 53462 31946
rect 54338 31932 54420 31946
rect 54628 31932 54710 31946
rect 55586 31932 55668 31946
rect 55876 31932 55958 31946
rect 56834 31932 56916 31946
rect 57124 31932 57206 31946
rect 58082 31932 58164 31946
rect 58372 31932 58454 31946
rect 16418 31884 16864 31898
rect 17014 31884 17154 31898
rect 17304 31884 18112 31898
rect 18262 31884 18402 31898
rect 18552 31884 19360 31898
rect 19510 31884 19650 31898
rect 19800 31884 20608 31898
rect 20758 31884 20898 31898
rect 21048 31884 21856 31898
rect 22006 31884 22146 31898
rect 22296 31884 23104 31898
rect 23254 31884 23394 31898
rect 23544 31884 24352 31898
rect 24502 31884 24642 31898
rect 24792 31884 25600 31898
rect 25750 31884 25890 31898
rect 26040 31884 26848 31898
rect 26998 31884 27138 31898
rect 27288 31884 28096 31898
rect 28246 31884 28386 31898
rect 28536 31884 29344 31898
rect 29494 31884 29634 31898
rect 29784 31884 30592 31898
rect 30742 31884 30882 31898
rect 31032 31884 31840 31898
rect 31990 31884 32130 31898
rect 32280 31884 33088 31898
rect 33238 31884 33378 31898
rect 33528 31884 34336 31898
rect 34486 31884 34626 31898
rect 34776 31884 35584 31898
rect 35734 31884 35874 31898
rect 36024 31884 36832 31898
rect 36982 31884 37122 31898
rect 37272 31884 38080 31898
rect 38230 31884 38370 31898
rect 38520 31884 39328 31898
rect 39478 31884 39618 31898
rect 39768 31884 40576 31898
rect 40726 31884 40866 31898
rect 41016 31884 41824 31898
rect 41974 31884 42114 31898
rect 42264 31884 43072 31898
rect 43222 31884 43362 31898
rect 43512 31884 44320 31898
rect 44470 31884 44610 31898
rect 44760 31884 45568 31898
rect 45718 31884 45858 31898
rect 46008 31884 46816 31898
rect 46966 31884 47106 31898
rect 47256 31884 48064 31898
rect 48214 31884 48354 31898
rect 48504 31884 49312 31898
rect 49462 31884 49602 31898
rect 49752 31884 50560 31898
rect 50710 31884 50850 31898
rect 51000 31884 51808 31898
rect 51958 31884 52098 31898
rect 52248 31884 53056 31898
rect 53206 31884 53346 31898
rect 53496 31884 54304 31898
rect 54454 31884 54594 31898
rect 54744 31884 55552 31898
rect 55702 31884 55842 31898
rect 55992 31884 56800 31898
rect 56950 31884 57090 31898
rect 57240 31884 58048 31898
rect 58198 31884 58338 31898
rect 58488 31884 58934 31898
rect 16418 31836 58934 31884
rect 16418 31822 16864 31836
rect 17014 31822 17154 31836
rect 17304 31822 18112 31836
rect 18262 31822 18402 31836
rect 18552 31822 19360 31836
rect 19510 31822 19650 31836
rect 19800 31822 20608 31836
rect 20758 31822 20898 31836
rect 21048 31822 21856 31836
rect 22006 31822 22146 31836
rect 22296 31822 23104 31836
rect 23254 31822 23394 31836
rect 23544 31822 24352 31836
rect 24502 31822 24642 31836
rect 24792 31822 25600 31836
rect 25750 31822 25890 31836
rect 26040 31822 26848 31836
rect 26998 31822 27138 31836
rect 27288 31822 28096 31836
rect 28246 31822 28386 31836
rect 28536 31822 29344 31836
rect 29494 31822 29634 31836
rect 29784 31822 30592 31836
rect 30742 31822 30882 31836
rect 31032 31822 31840 31836
rect 31990 31822 32130 31836
rect 32280 31822 33088 31836
rect 33238 31822 33378 31836
rect 33528 31822 34336 31836
rect 34486 31822 34626 31836
rect 34776 31822 35584 31836
rect 35734 31822 35874 31836
rect 36024 31822 36832 31836
rect 36982 31822 37122 31836
rect 37272 31822 38080 31836
rect 38230 31822 38370 31836
rect 38520 31822 39328 31836
rect 39478 31822 39618 31836
rect 39768 31822 40576 31836
rect 40726 31822 40866 31836
rect 41016 31822 41824 31836
rect 41974 31822 42114 31836
rect 42264 31822 43072 31836
rect 43222 31822 43362 31836
rect 43512 31822 44320 31836
rect 44470 31822 44610 31836
rect 44760 31822 45568 31836
rect 45718 31822 45858 31836
rect 46008 31822 46816 31836
rect 46966 31822 47106 31836
rect 47256 31822 48064 31836
rect 48214 31822 48354 31836
rect 48504 31822 49312 31836
rect 49462 31822 49602 31836
rect 49752 31822 50560 31836
rect 50710 31822 50850 31836
rect 51000 31822 51808 31836
rect 51958 31822 52098 31836
rect 52248 31822 53056 31836
rect 53206 31822 53346 31836
rect 53496 31822 54304 31836
rect 54454 31822 54594 31836
rect 54744 31822 55552 31836
rect 55702 31822 55842 31836
rect 55992 31822 56800 31836
rect 56950 31822 57090 31836
rect 57240 31822 58048 31836
rect 58198 31822 58338 31836
rect 58488 31822 58934 31836
rect 16898 31774 16980 31788
rect 17188 31774 17270 31788
rect 18146 31774 18228 31788
rect 18436 31774 18518 31788
rect 19394 31774 19476 31788
rect 19684 31774 19766 31788
rect 20642 31774 20724 31788
rect 20932 31774 21014 31788
rect 21890 31774 21972 31788
rect 22180 31774 22262 31788
rect 23138 31774 23220 31788
rect 23428 31774 23510 31788
rect 24386 31774 24468 31788
rect 24676 31774 24758 31788
rect 25634 31774 25716 31788
rect 25924 31774 26006 31788
rect 26882 31774 26964 31788
rect 27172 31774 27254 31788
rect 28130 31774 28212 31788
rect 28420 31774 28502 31788
rect 29378 31774 29460 31788
rect 29668 31774 29750 31788
rect 30626 31774 30708 31788
rect 30916 31774 30998 31788
rect 31874 31774 31956 31788
rect 32164 31774 32246 31788
rect 33122 31774 33204 31788
rect 33412 31774 33494 31788
rect 34370 31774 34452 31788
rect 34660 31774 34742 31788
rect 35618 31774 35700 31788
rect 35908 31774 35990 31788
rect 36866 31774 36948 31788
rect 37156 31774 37238 31788
rect 38114 31774 38196 31788
rect 38404 31774 38486 31788
rect 39362 31774 39444 31788
rect 39652 31774 39734 31788
rect 40610 31774 40692 31788
rect 40900 31774 40982 31788
rect 41858 31774 41940 31788
rect 42148 31774 42230 31788
rect 43106 31774 43188 31788
rect 43396 31774 43478 31788
rect 44354 31774 44436 31788
rect 44644 31774 44726 31788
rect 45602 31774 45684 31788
rect 45892 31774 45974 31788
rect 46850 31774 46932 31788
rect 47140 31774 47222 31788
rect 48098 31774 48180 31788
rect 48388 31774 48470 31788
rect 49346 31774 49428 31788
rect 49636 31774 49718 31788
rect 50594 31774 50676 31788
rect 50884 31774 50966 31788
rect 51842 31774 51924 31788
rect 52132 31774 52214 31788
rect 53090 31774 53172 31788
rect 53380 31774 53462 31788
rect 54338 31774 54420 31788
rect 54628 31774 54710 31788
rect 55586 31774 55668 31788
rect 55876 31774 55958 31788
rect 56834 31774 56916 31788
rect 57124 31774 57206 31788
rect 58082 31774 58164 31788
rect 58372 31774 58454 31788
rect 16418 31726 58934 31774
rect 16418 31568 58934 31678
rect 16418 31472 58934 31520
rect 16898 31458 16980 31472
rect 17188 31458 17270 31472
rect 18146 31458 18228 31472
rect 18436 31458 18518 31472
rect 19394 31458 19476 31472
rect 19684 31458 19766 31472
rect 20642 31458 20724 31472
rect 20932 31458 21014 31472
rect 21890 31458 21972 31472
rect 22180 31458 22262 31472
rect 23138 31458 23220 31472
rect 23428 31458 23510 31472
rect 24386 31458 24468 31472
rect 24676 31458 24758 31472
rect 25634 31458 25716 31472
rect 25924 31458 26006 31472
rect 26882 31458 26964 31472
rect 27172 31458 27254 31472
rect 28130 31458 28212 31472
rect 28420 31458 28502 31472
rect 29378 31458 29460 31472
rect 29668 31458 29750 31472
rect 30626 31458 30708 31472
rect 30916 31458 30998 31472
rect 31874 31458 31956 31472
rect 32164 31458 32246 31472
rect 33122 31458 33204 31472
rect 33412 31458 33494 31472
rect 34370 31458 34452 31472
rect 34660 31458 34742 31472
rect 35618 31458 35700 31472
rect 35908 31458 35990 31472
rect 36866 31458 36948 31472
rect 37156 31458 37238 31472
rect 38114 31458 38196 31472
rect 38404 31458 38486 31472
rect 39362 31458 39444 31472
rect 39652 31458 39734 31472
rect 40610 31458 40692 31472
rect 40900 31458 40982 31472
rect 41858 31458 41940 31472
rect 42148 31458 42230 31472
rect 43106 31458 43188 31472
rect 43396 31458 43478 31472
rect 44354 31458 44436 31472
rect 44644 31458 44726 31472
rect 45602 31458 45684 31472
rect 45892 31458 45974 31472
rect 46850 31458 46932 31472
rect 47140 31458 47222 31472
rect 48098 31458 48180 31472
rect 48388 31458 48470 31472
rect 49346 31458 49428 31472
rect 49636 31458 49718 31472
rect 50594 31458 50676 31472
rect 50884 31458 50966 31472
rect 51842 31458 51924 31472
rect 52132 31458 52214 31472
rect 53090 31458 53172 31472
rect 53380 31458 53462 31472
rect 54338 31458 54420 31472
rect 54628 31458 54710 31472
rect 55586 31458 55668 31472
rect 55876 31458 55958 31472
rect 56834 31458 56916 31472
rect 57124 31458 57206 31472
rect 58082 31458 58164 31472
rect 58372 31458 58454 31472
rect 16418 31410 16864 31424
rect 17014 31410 17154 31424
rect 17304 31410 18112 31424
rect 18262 31410 18402 31424
rect 18552 31410 19360 31424
rect 19510 31410 19650 31424
rect 19800 31410 20608 31424
rect 20758 31410 20898 31424
rect 21048 31410 21856 31424
rect 22006 31410 22146 31424
rect 22296 31410 23104 31424
rect 23254 31410 23394 31424
rect 23544 31410 24352 31424
rect 24502 31410 24642 31424
rect 24792 31410 25600 31424
rect 25750 31410 25890 31424
rect 26040 31410 26848 31424
rect 26998 31410 27138 31424
rect 27288 31410 28096 31424
rect 28246 31410 28386 31424
rect 28536 31410 29344 31424
rect 29494 31410 29634 31424
rect 29784 31410 30592 31424
rect 30742 31410 30882 31424
rect 31032 31410 31840 31424
rect 31990 31410 32130 31424
rect 32280 31410 33088 31424
rect 33238 31410 33378 31424
rect 33528 31410 34336 31424
rect 34486 31410 34626 31424
rect 34776 31410 35584 31424
rect 35734 31410 35874 31424
rect 36024 31410 36832 31424
rect 36982 31410 37122 31424
rect 37272 31410 38080 31424
rect 38230 31410 38370 31424
rect 38520 31410 39328 31424
rect 39478 31410 39618 31424
rect 39768 31410 40576 31424
rect 40726 31410 40866 31424
rect 41016 31410 41824 31424
rect 41974 31410 42114 31424
rect 42264 31410 43072 31424
rect 43222 31410 43362 31424
rect 43512 31410 44320 31424
rect 44470 31410 44610 31424
rect 44760 31410 45568 31424
rect 45718 31410 45858 31424
rect 46008 31410 46816 31424
rect 46966 31410 47106 31424
rect 47256 31410 48064 31424
rect 48214 31410 48354 31424
rect 48504 31410 49312 31424
rect 49462 31410 49602 31424
rect 49752 31410 50560 31424
rect 50710 31410 50850 31424
rect 51000 31410 51808 31424
rect 51958 31410 52098 31424
rect 52248 31410 53056 31424
rect 53206 31410 53346 31424
rect 53496 31410 54304 31424
rect 54454 31410 54594 31424
rect 54744 31410 55552 31424
rect 55702 31410 55842 31424
rect 55992 31410 56800 31424
rect 56950 31410 57090 31424
rect 57240 31410 58048 31424
rect 58198 31410 58338 31424
rect 58488 31410 58934 31424
rect 16418 31362 58934 31410
rect 16418 31348 16864 31362
rect 17014 31348 17154 31362
rect 17304 31348 18112 31362
rect 18262 31348 18402 31362
rect 18552 31348 19360 31362
rect 19510 31348 19650 31362
rect 19800 31348 20608 31362
rect 20758 31348 20898 31362
rect 21048 31348 21856 31362
rect 22006 31348 22146 31362
rect 22296 31348 23104 31362
rect 23254 31348 23394 31362
rect 23544 31348 24352 31362
rect 24502 31348 24642 31362
rect 24792 31348 25600 31362
rect 25750 31348 25890 31362
rect 26040 31348 26848 31362
rect 26998 31348 27138 31362
rect 27288 31348 28096 31362
rect 28246 31348 28386 31362
rect 28536 31348 29344 31362
rect 29494 31348 29634 31362
rect 29784 31348 30592 31362
rect 30742 31348 30882 31362
rect 31032 31348 31840 31362
rect 31990 31348 32130 31362
rect 32280 31348 33088 31362
rect 33238 31348 33378 31362
rect 33528 31348 34336 31362
rect 34486 31348 34626 31362
rect 34776 31348 35584 31362
rect 35734 31348 35874 31362
rect 36024 31348 36832 31362
rect 36982 31348 37122 31362
rect 37272 31348 38080 31362
rect 38230 31348 38370 31362
rect 38520 31348 39328 31362
rect 39478 31348 39618 31362
rect 39768 31348 40576 31362
rect 40726 31348 40866 31362
rect 41016 31348 41824 31362
rect 41974 31348 42114 31362
rect 42264 31348 43072 31362
rect 43222 31348 43362 31362
rect 43512 31348 44320 31362
rect 44470 31348 44610 31362
rect 44760 31348 45568 31362
rect 45718 31348 45858 31362
rect 46008 31348 46816 31362
rect 46966 31348 47106 31362
rect 47256 31348 48064 31362
rect 48214 31348 48354 31362
rect 48504 31348 49312 31362
rect 49462 31348 49602 31362
rect 49752 31348 50560 31362
rect 50710 31348 50850 31362
rect 51000 31348 51808 31362
rect 51958 31348 52098 31362
rect 52248 31348 53056 31362
rect 53206 31348 53346 31362
rect 53496 31348 54304 31362
rect 54454 31348 54594 31362
rect 54744 31348 55552 31362
rect 55702 31348 55842 31362
rect 55992 31348 56800 31362
rect 56950 31348 57090 31362
rect 57240 31348 58048 31362
rect 58198 31348 58338 31362
rect 58488 31348 58934 31362
rect 16898 31300 16980 31314
rect 17188 31300 17270 31314
rect 18146 31300 18228 31314
rect 18436 31300 18518 31314
rect 19394 31300 19476 31314
rect 19684 31300 19766 31314
rect 20642 31300 20724 31314
rect 20932 31300 21014 31314
rect 21890 31300 21972 31314
rect 22180 31300 22262 31314
rect 23138 31300 23220 31314
rect 23428 31300 23510 31314
rect 24386 31300 24468 31314
rect 24676 31300 24758 31314
rect 25634 31300 25716 31314
rect 25924 31300 26006 31314
rect 26882 31300 26964 31314
rect 27172 31300 27254 31314
rect 28130 31300 28212 31314
rect 28420 31300 28502 31314
rect 29378 31300 29460 31314
rect 29668 31300 29750 31314
rect 30626 31300 30708 31314
rect 30916 31300 30998 31314
rect 31874 31300 31956 31314
rect 32164 31300 32246 31314
rect 33122 31300 33204 31314
rect 33412 31300 33494 31314
rect 34370 31300 34452 31314
rect 34660 31300 34742 31314
rect 35618 31300 35700 31314
rect 35908 31300 35990 31314
rect 36866 31300 36948 31314
rect 37156 31300 37238 31314
rect 38114 31300 38196 31314
rect 38404 31300 38486 31314
rect 39362 31300 39444 31314
rect 39652 31300 39734 31314
rect 40610 31300 40692 31314
rect 40900 31300 40982 31314
rect 41858 31300 41940 31314
rect 42148 31300 42230 31314
rect 43106 31300 43188 31314
rect 43396 31300 43478 31314
rect 44354 31300 44436 31314
rect 44644 31300 44726 31314
rect 45602 31300 45684 31314
rect 45892 31300 45974 31314
rect 46850 31300 46932 31314
rect 47140 31300 47222 31314
rect 48098 31300 48180 31314
rect 48388 31300 48470 31314
rect 49346 31300 49428 31314
rect 49636 31300 49718 31314
rect 50594 31300 50676 31314
rect 50884 31300 50966 31314
rect 51842 31300 51924 31314
rect 52132 31300 52214 31314
rect 53090 31300 53172 31314
rect 53380 31300 53462 31314
rect 54338 31300 54420 31314
rect 54628 31300 54710 31314
rect 55586 31300 55668 31314
rect 55876 31300 55958 31314
rect 56834 31300 56916 31314
rect 57124 31300 57206 31314
rect 58082 31300 58164 31314
rect 58372 31300 58454 31314
rect 16418 31252 58934 31300
rect 16418 31156 58934 31204
rect 16898 31142 16980 31156
rect 17188 31142 17270 31156
rect 18146 31142 18228 31156
rect 18436 31142 18518 31156
rect 19394 31142 19476 31156
rect 19684 31142 19766 31156
rect 20642 31142 20724 31156
rect 20932 31142 21014 31156
rect 21890 31142 21972 31156
rect 22180 31142 22262 31156
rect 23138 31142 23220 31156
rect 23428 31142 23510 31156
rect 24386 31142 24468 31156
rect 24676 31142 24758 31156
rect 25634 31142 25716 31156
rect 25924 31142 26006 31156
rect 26882 31142 26964 31156
rect 27172 31142 27254 31156
rect 28130 31142 28212 31156
rect 28420 31142 28502 31156
rect 29378 31142 29460 31156
rect 29668 31142 29750 31156
rect 30626 31142 30708 31156
rect 30916 31142 30998 31156
rect 31874 31142 31956 31156
rect 32164 31142 32246 31156
rect 33122 31142 33204 31156
rect 33412 31142 33494 31156
rect 34370 31142 34452 31156
rect 34660 31142 34742 31156
rect 35618 31142 35700 31156
rect 35908 31142 35990 31156
rect 36866 31142 36948 31156
rect 37156 31142 37238 31156
rect 38114 31142 38196 31156
rect 38404 31142 38486 31156
rect 39362 31142 39444 31156
rect 39652 31142 39734 31156
rect 40610 31142 40692 31156
rect 40900 31142 40982 31156
rect 41858 31142 41940 31156
rect 42148 31142 42230 31156
rect 43106 31142 43188 31156
rect 43396 31142 43478 31156
rect 44354 31142 44436 31156
rect 44644 31142 44726 31156
rect 45602 31142 45684 31156
rect 45892 31142 45974 31156
rect 46850 31142 46932 31156
rect 47140 31142 47222 31156
rect 48098 31142 48180 31156
rect 48388 31142 48470 31156
rect 49346 31142 49428 31156
rect 49636 31142 49718 31156
rect 50594 31142 50676 31156
rect 50884 31142 50966 31156
rect 51842 31142 51924 31156
rect 52132 31142 52214 31156
rect 53090 31142 53172 31156
rect 53380 31142 53462 31156
rect 54338 31142 54420 31156
rect 54628 31142 54710 31156
rect 55586 31142 55668 31156
rect 55876 31142 55958 31156
rect 56834 31142 56916 31156
rect 57124 31142 57206 31156
rect 58082 31142 58164 31156
rect 58372 31142 58454 31156
rect 16418 31094 16864 31108
rect 17014 31094 17154 31108
rect 17304 31094 18112 31108
rect 18262 31094 18402 31108
rect 18552 31094 19360 31108
rect 19510 31094 19650 31108
rect 19800 31094 20608 31108
rect 20758 31094 20898 31108
rect 21048 31094 21856 31108
rect 22006 31094 22146 31108
rect 22296 31094 23104 31108
rect 23254 31094 23394 31108
rect 23544 31094 24352 31108
rect 24502 31094 24642 31108
rect 24792 31094 25600 31108
rect 25750 31094 25890 31108
rect 26040 31094 26848 31108
rect 26998 31094 27138 31108
rect 27288 31094 28096 31108
rect 28246 31094 28386 31108
rect 28536 31094 29344 31108
rect 29494 31094 29634 31108
rect 29784 31094 30592 31108
rect 30742 31094 30882 31108
rect 31032 31094 31840 31108
rect 31990 31094 32130 31108
rect 32280 31094 33088 31108
rect 33238 31094 33378 31108
rect 33528 31094 34336 31108
rect 34486 31094 34626 31108
rect 34776 31094 35584 31108
rect 35734 31094 35874 31108
rect 36024 31094 36832 31108
rect 36982 31094 37122 31108
rect 37272 31094 38080 31108
rect 38230 31094 38370 31108
rect 38520 31094 39328 31108
rect 39478 31094 39618 31108
rect 39768 31094 40576 31108
rect 40726 31094 40866 31108
rect 41016 31094 41824 31108
rect 41974 31094 42114 31108
rect 42264 31094 43072 31108
rect 43222 31094 43362 31108
rect 43512 31094 44320 31108
rect 44470 31094 44610 31108
rect 44760 31094 45568 31108
rect 45718 31094 45858 31108
rect 46008 31094 46816 31108
rect 46966 31094 47106 31108
rect 47256 31094 48064 31108
rect 48214 31094 48354 31108
rect 48504 31094 49312 31108
rect 49462 31094 49602 31108
rect 49752 31094 50560 31108
rect 50710 31094 50850 31108
rect 51000 31094 51808 31108
rect 51958 31094 52098 31108
rect 52248 31094 53056 31108
rect 53206 31094 53346 31108
rect 53496 31094 54304 31108
rect 54454 31094 54594 31108
rect 54744 31094 55552 31108
rect 55702 31094 55842 31108
rect 55992 31094 56800 31108
rect 56950 31094 57090 31108
rect 57240 31094 58048 31108
rect 58198 31094 58338 31108
rect 58488 31094 58934 31108
rect 16418 31046 58934 31094
rect 16418 31032 16864 31046
rect 17014 31032 17154 31046
rect 17304 31032 18112 31046
rect 18262 31032 18402 31046
rect 18552 31032 19360 31046
rect 19510 31032 19650 31046
rect 19800 31032 20608 31046
rect 20758 31032 20898 31046
rect 21048 31032 21856 31046
rect 22006 31032 22146 31046
rect 22296 31032 23104 31046
rect 23254 31032 23394 31046
rect 23544 31032 24352 31046
rect 24502 31032 24642 31046
rect 24792 31032 25600 31046
rect 25750 31032 25890 31046
rect 26040 31032 26848 31046
rect 26998 31032 27138 31046
rect 27288 31032 28096 31046
rect 28246 31032 28386 31046
rect 28536 31032 29344 31046
rect 29494 31032 29634 31046
rect 29784 31032 30592 31046
rect 30742 31032 30882 31046
rect 31032 31032 31840 31046
rect 31990 31032 32130 31046
rect 32280 31032 33088 31046
rect 33238 31032 33378 31046
rect 33528 31032 34336 31046
rect 34486 31032 34626 31046
rect 34776 31032 35584 31046
rect 35734 31032 35874 31046
rect 36024 31032 36832 31046
rect 36982 31032 37122 31046
rect 37272 31032 38080 31046
rect 38230 31032 38370 31046
rect 38520 31032 39328 31046
rect 39478 31032 39618 31046
rect 39768 31032 40576 31046
rect 40726 31032 40866 31046
rect 41016 31032 41824 31046
rect 41974 31032 42114 31046
rect 42264 31032 43072 31046
rect 43222 31032 43362 31046
rect 43512 31032 44320 31046
rect 44470 31032 44610 31046
rect 44760 31032 45568 31046
rect 45718 31032 45858 31046
rect 46008 31032 46816 31046
rect 46966 31032 47106 31046
rect 47256 31032 48064 31046
rect 48214 31032 48354 31046
rect 48504 31032 49312 31046
rect 49462 31032 49602 31046
rect 49752 31032 50560 31046
rect 50710 31032 50850 31046
rect 51000 31032 51808 31046
rect 51958 31032 52098 31046
rect 52248 31032 53056 31046
rect 53206 31032 53346 31046
rect 53496 31032 54304 31046
rect 54454 31032 54594 31046
rect 54744 31032 55552 31046
rect 55702 31032 55842 31046
rect 55992 31032 56800 31046
rect 56950 31032 57090 31046
rect 57240 31032 58048 31046
rect 58198 31032 58338 31046
rect 58488 31032 58934 31046
rect 16898 30984 16980 30998
rect 17188 30984 17270 30998
rect 18146 30984 18228 30998
rect 18436 30984 18518 30998
rect 19394 30984 19476 30998
rect 19684 30984 19766 30998
rect 20642 30984 20724 30998
rect 20932 30984 21014 30998
rect 21890 30984 21972 30998
rect 22180 30984 22262 30998
rect 23138 30984 23220 30998
rect 23428 30984 23510 30998
rect 24386 30984 24468 30998
rect 24676 30984 24758 30998
rect 25634 30984 25716 30998
rect 25924 30984 26006 30998
rect 26882 30984 26964 30998
rect 27172 30984 27254 30998
rect 28130 30984 28212 30998
rect 28420 30984 28502 30998
rect 29378 30984 29460 30998
rect 29668 30984 29750 30998
rect 30626 30984 30708 30998
rect 30916 30984 30998 30998
rect 31874 30984 31956 30998
rect 32164 30984 32246 30998
rect 33122 30984 33204 30998
rect 33412 30984 33494 30998
rect 34370 30984 34452 30998
rect 34660 30984 34742 30998
rect 35618 30984 35700 30998
rect 35908 30984 35990 30998
rect 36866 30984 36948 30998
rect 37156 30984 37238 30998
rect 38114 30984 38196 30998
rect 38404 30984 38486 30998
rect 39362 30984 39444 30998
rect 39652 30984 39734 30998
rect 40610 30984 40692 30998
rect 40900 30984 40982 30998
rect 41858 30984 41940 30998
rect 42148 30984 42230 30998
rect 43106 30984 43188 30998
rect 43396 30984 43478 30998
rect 44354 30984 44436 30998
rect 44644 30984 44726 30998
rect 45602 30984 45684 30998
rect 45892 30984 45974 30998
rect 46850 30984 46932 30998
rect 47140 30984 47222 30998
rect 48098 30984 48180 30998
rect 48388 30984 48470 30998
rect 49346 30984 49428 30998
rect 49636 30984 49718 30998
rect 50594 30984 50676 30998
rect 50884 30984 50966 30998
rect 51842 30984 51924 30998
rect 52132 30984 52214 30998
rect 53090 30984 53172 30998
rect 53380 30984 53462 30998
rect 54338 30984 54420 30998
rect 54628 30984 54710 30998
rect 55586 30984 55668 30998
rect 55876 30984 55958 30998
rect 56834 30984 56916 30998
rect 57124 30984 57206 30998
rect 58082 30984 58164 30998
rect 58372 30984 58454 30998
rect 16418 30936 58934 30984
rect 16418 30778 58934 30888
rect 16418 30682 58934 30730
rect 16898 30668 16980 30682
rect 17188 30668 17270 30682
rect 18146 30668 18228 30682
rect 18436 30668 18518 30682
rect 19394 30668 19476 30682
rect 19684 30668 19766 30682
rect 20642 30668 20724 30682
rect 20932 30668 21014 30682
rect 21890 30668 21972 30682
rect 22180 30668 22262 30682
rect 23138 30668 23220 30682
rect 23428 30668 23510 30682
rect 24386 30668 24468 30682
rect 24676 30668 24758 30682
rect 25634 30668 25716 30682
rect 25924 30668 26006 30682
rect 26882 30668 26964 30682
rect 27172 30668 27254 30682
rect 28130 30668 28212 30682
rect 28420 30668 28502 30682
rect 29378 30668 29460 30682
rect 29668 30668 29750 30682
rect 30626 30668 30708 30682
rect 30916 30668 30998 30682
rect 31874 30668 31956 30682
rect 32164 30668 32246 30682
rect 33122 30668 33204 30682
rect 33412 30668 33494 30682
rect 34370 30668 34452 30682
rect 34660 30668 34742 30682
rect 35618 30668 35700 30682
rect 35908 30668 35990 30682
rect 36866 30668 36948 30682
rect 37156 30668 37238 30682
rect 38114 30668 38196 30682
rect 38404 30668 38486 30682
rect 39362 30668 39444 30682
rect 39652 30668 39734 30682
rect 40610 30668 40692 30682
rect 40900 30668 40982 30682
rect 41858 30668 41940 30682
rect 42148 30668 42230 30682
rect 43106 30668 43188 30682
rect 43396 30668 43478 30682
rect 44354 30668 44436 30682
rect 44644 30668 44726 30682
rect 45602 30668 45684 30682
rect 45892 30668 45974 30682
rect 46850 30668 46932 30682
rect 47140 30668 47222 30682
rect 48098 30668 48180 30682
rect 48388 30668 48470 30682
rect 49346 30668 49428 30682
rect 49636 30668 49718 30682
rect 50594 30668 50676 30682
rect 50884 30668 50966 30682
rect 51842 30668 51924 30682
rect 52132 30668 52214 30682
rect 53090 30668 53172 30682
rect 53380 30668 53462 30682
rect 54338 30668 54420 30682
rect 54628 30668 54710 30682
rect 55586 30668 55668 30682
rect 55876 30668 55958 30682
rect 56834 30668 56916 30682
rect 57124 30668 57206 30682
rect 58082 30668 58164 30682
rect 58372 30668 58454 30682
rect 16418 30620 16864 30634
rect 17014 30620 17154 30634
rect 17304 30620 18112 30634
rect 18262 30620 18402 30634
rect 18552 30620 19360 30634
rect 19510 30620 19650 30634
rect 19800 30620 20608 30634
rect 20758 30620 20898 30634
rect 21048 30620 21856 30634
rect 22006 30620 22146 30634
rect 22296 30620 23104 30634
rect 23254 30620 23394 30634
rect 23544 30620 24352 30634
rect 24502 30620 24642 30634
rect 24792 30620 25600 30634
rect 25750 30620 25890 30634
rect 26040 30620 26848 30634
rect 26998 30620 27138 30634
rect 27288 30620 28096 30634
rect 28246 30620 28386 30634
rect 28536 30620 29344 30634
rect 29494 30620 29634 30634
rect 29784 30620 30592 30634
rect 30742 30620 30882 30634
rect 31032 30620 31840 30634
rect 31990 30620 32130 30634
rect 32280 30620 33088 30634
rect 33238 30620 33378 30634
rect 33528 30620 34336 30634
rect 34486 30620 34626 30634
rect 34776 30620 35584 30634
rect 35734 30620 35874 30634
rect 36024 30620 36832 30634
rect 36982 30620 37122 30634
rect 37272 30620 38080 30634
rect 38230 30620 38370 30634
rect 38520 30620 39328 30634
rect 39478 30620 39618 30634
rect 39768 30620 40576 30634
rect 40726 30620 40866 30634
rect 41016 30620 41824 30634
rect 41974 30620 42114 30634
rect 42264 30620 43072 30634
rect 43222 30620 43362 30634
rect 43512 30620 44320 30634
rect 44470 30620 44610 30634
rect 44760 30620 45568 30634
rect 45718 30620 45858 30634
rect 46008 30620 46816 30634
rect 46966 30620 47106 30634
rect 47256 30620 48064 30634
rect 48214 30620 48354 30634
rect 48504 30620 49312 30634
rect 49462 30620 49602 30634
rect 49752 30620 50560 30634
rect 50710 30620 50850 30634
rect 51000 30620 51808 30634
rect 51958 30620 52098 30634
rect 52248 30620 53056 30634
rect 53206 30620 53346 30634
rect 53496 30620 54304 30634
rect 54454 30620 54594 30634
rect 54744 30620 55552 30634
rect 55702 30620 55842 30634
rect 55992 30620 56800 30634
rect 56950 30620 57090 30634
rect 57240 30620 58048 30634
rect 58198 30620 58338 30634
rect 58488 30620 58934 30634
rect 16418 30572 58934 30620
rect 16418 30558 16864 30572
rect 17014 30558 17154 30572
rect 17304 30558 18112 30572
rect 18262 30558 18402 30572
rect 18552 30558 19360 30572
rect 19510 30558 19650 30572
rect 19800 30558 20608 30572
rect 20758 30558 20898 30572
rect 21048 30558 21856 30572
rect 22006 30558 22146 30572
rect 22296 30558 23104 30572
rect 23254 30558 23394 30572
rect 23544 30558 24352 30572
rect 24502 30558 24642 30572
rect 24792 30558 25600 30572
rect 25750 30558 25890 30572
rect 26040 30558 26848 30572
rect 26998 30558 27138 30572
rect 27288 30558 28096 30572
rect 28246 30558 28386 30572
rect 28536 30558 29344 30572
rect 29494 30558 29634 30572
rect 29784 30558 30592 30572
rect 30742 30558 30882 30572
rect 31032 30558 31840 30572
rect 31990 30558 32130 30572
rect 32280 30558 33088 30572
rect 33238 30558 33378 30572
rect 33528 30558 34336 30572
rect 34486 30558 34626 30572
rect 34776 30558 35584 30572
rect 35734 30558 35874 30572
rect 36024 30558 36832 30572
rect 36982 30558 37122 30572
rect 37272 30558 38080 30572
rect 38230 30558 38370 30572
rect 38520 30558 39328 30572
rect 39478 30558 39618 30572
rect 39768 30558 40576 30572
rect 40726 30558 40866 30572
rect 41016 30558 41824 30572
rect 41974 30558 42114 30572
rect 42264 30558 43072 30572
rect 43222 30558 43362 30572
rect 43512 30558 44320 30572
rect 44470 30558 44610 30572
rect 44760 30558 45568 30572
rect 45718 30558 45858 30572
rect 46008 30558 46816 30572
rect 46966 30558 47106 30572
rect 47256 30558 48064 30572
rect 48214 30558 48354 30572
rect 48504 30558 49312 30572
rect 49462 30558 49602 30572
rect 49752 30558 50560 30572
rect 50710 30558 50850 30572
rect 51000 30558 51808 30572
rect 51958 30558 52098 30572
rect 52248 30558 53056 30572
rect 53206 30558 53346 30572
rect 53496 30558 54304 30572
rect 54454 30558 54594 30572
rect 54744 30558 55552 30572
rect 55702 30558 55842 30572
rect 55992 30558 56800 30572
rect 56950 30558 57090 30572
rect 57240 30558 58048 30572
rect 58198 30558 58338 30572
rect 58488 30558 58934 30572
rect 16898 30510 16980 30524
rect 17188 30510 17270 30524
rect 18146 30510 18228 30524
rect 18436 30510 18518 30524
rect 19394 30510 19476 30524
rect 19684 30510 19766 30524
rect 20642 30510 20724 30524
rect 20932 30510 21014 30524
rect 21890 30510 21972 30524
rect 22180 30510 22262 30524
rect 23138 30510 23220 30524
rect 23428 30510 23510 30524
rect 24386 30510 24468 30524
rect 24676 30510 24758 30524
rect 25634 30510 25716 30524
rect 25924 30510 26006 30524
rect 26882 30510 26964 30524
rect 27172 30510 27254 30524
rect 28130 30510 28212 30524
rect 28420 30510 28502 30524
rect 29378 30510 29460 30524
rect 29668 30510 29750 30524
rect 30626 30510 30708 30524
rect 30916 30510 30998 30524
rect 31874 30510 31956 30524
rect 32164 30510 32246 30524
rect 33122 30510 33204 30524
rect 33412 30510 33494 30524
rect 34370 30510 34452 30524
rect 34660 30510 34742 30524
rect 35618 30510 35700 30524
rect 35908 30510 35990 30524
rect 36866 30510 36948 30524
rect 37156 30510 37238 30524
rect 38114 30510 38196 30524
rect 38404 30510 38486 30524
rect 39362 30510 39444 30524
rect 39652 30510 39734 30524
rect 40610 30510 40692 30524
rect 40900 30510 40982 30524
rect 41858 30510 41940 30524
rect 42148 30510 42230 30524
rect 43106 30510 43188 30524
rect 43396 30510 43478 30524
rect 44354 30510 44436 30524
rect 44644 30510 44726 30524
rect 45602 30510 45684 30524
rect 45892 30510 45974 30524
rect 46850 30510 46932 30524
rect 47140 30510 47222 30524
rect 48098 30510 48180 30524
rect 48388 30510 48470 30524
rect 49346 30510 49428 30524
rect 49636 30510 49718 30524
rect 50594 30510 50676 30524
rect 50884 30510 50966 30524
rect 51842 30510 51924 30524
rect 52132 30510 52214 30524
rect 53090 30510 53172 30524
rect 53380 30510 53462 30524
rect 54338 30510 54420 30524
rect 54628 30510 54710 30524
rect 55586 30510 55668 30524
rect 55876 30510 55958 30524
rect 56834 30510 56916 30524
rect 57124 30510 57206 30524
rect 58082 30510 58164 30524
rect 58372 30510 58454 30524
rect 16418 30462 58934 30510
rect 16418 30366 58934 30414
rect 16898 30352 16980 30366
rect 17188 30352 17270 30366
rect 18146 30352 18228 30366
rect 18436 30352 18518 30366
rect 19394 30352 19476 30366
rect 19684 30352 19766 30366
rect 20642 30352 20724 30366
rect 20932 30352 21014 30366
rect 21890 30352 21972 30366
rect 22180 30352 22262 30366
rect 23138 30352 23220 30366
rect 23428 30352 23510 30366
rect 24386 30352 24468 30366
rect 24676 30352 24758 30366
rect 25634 30352 25716 30366
rect 25924 30352 26006 30366
rect 26882 30352 26964 30366
rect 27172 30352 27254 30366
rect 28130 30352 28212 30366
rect 28420 30352 28502 30366
rect 29378 30352 29460 30366
rect 29668 30352 29750 30366
rect 30626 30352 30708 30366
rect 30916 30352 30998 30366
rect 31874 30352 31956 30366
rect 32164 30352 32246 30366
rect 33122 30352 33204 30366
rect 33412 30352 33494 30366
rect 34370 30352 34452 30366
rect 34660 30352 34742 30366
rect 35618 30352 35700 30366
rect 35908 30352 35990 30366
rect 36866 30352 36948 30366
rect 37156 30352 37238 30366
rect 38114 30352 38196 30366
rect 38404 30352 38486 30366
rect 39362 30352 39444 30366
rect 39652 30352 39734 30366
rect 40610 30352 40692 30366
rect 40900 30352 40982 30366
rect 41858 30352 41940 30366
rect 42148 30352 42230 30366
rect 43106 30352 43188 30366
rect 43396 30352 43478 30366
rect 44354 30352 44436 30366
rect 44644 30352 44726 30366
rect 45602 30352 45684 30366
rect 45892 30352 45974 30366
rect 46850 30352 46932 30366
rect 47140 30352 47222 30366
rect 48098 30352 48180 30366
rect 48388 30352 48470 30366
rect 49346 30352 49428 30366
rect 49636 30352 49718 30366
rect 50594 30352 50676 30366
rect 50884 30352 50966 30366
rect 51842 30352 51924 30366
rect 52132 30352 52214 30366
rect 53090 30352 53172 30366
rect 53380 30352 53462 30366
rect 54338 30352 54420 30366
rect 54628 30352 54710 30366
rect 55586 30352 55668 30366
rect 55876 30352 55958 30366
rect 56834 30352 56916 30366
rect 57124 30352 57206 30366
rect 58082 30352 58164 30366
rect 58372 30352 58454 30366
rect 16418 30304 16864 30318
rect 17014 30304 17154 30318
rect 17304 30304 18112 30318
rect 18262 30304 18402 30318
rect 18552 30304 19360 30318
rect 19510 30304 19650 30318
rect 19800 30304 20608 30318
rect 20758 30304 20898 30318
rect 21048 30304 21856 30318
rect 22006 30304 22146 30318
rect 22296 30304 23104 30318
rect 23254 30304 23394 30318
rect 23544 30304 24352 30318
rect 24502 30304 24642 30318
rect 24792 30304 25600 30318
rect 25750 30304 25890 30318
rect 26040 30304 26848 30318
rect 26998 30304 27138 30318
rect 27288 30304 28096 30318
rect 28246 30304 28386 30318
rect 28536 30304 29344 30318
rect 29494 30304 29634 30318
rect 29784 30304 30592 30318
rect 30742 30304 30882 30318
rect 31032 30304 31840 30318
rect 31990 30304 32130 30318
rect 32280 30304 33088 30318
rect 33238 30304 33378 30318
rect 33528 30304 34336 30318
rect 34486 30304 34626 30318
rect 34776 30304 35584 30318
rect 35734 30304 35874 30318
rect 36024 30304 36832 30318
rect 36982 30304 37122 30318
rect 37272 30304 38080 30318
rect 38230 30304 38370 30318
rect 38520 30304 39328 30318
rect 39478 30304 39618 30318
rect 39768 30304 40576 30318
rect 40726 30304 40866 30318
rect 41016 30304 41824 30318
rect 41974 30304 42114 30318
rect 42264 30304 43072 30318
rect 43222 30304 43362 30318
rect 43512 30304 44320 30318
rect 44470 30304 44610 30318
rect 44760 30304 45568 30318
rect 45718 30304 45858 30318
rect 46008 30304 46816 30318
rect 46966 30304 47106 30318
rect 47256 30304 48064 30318
rect 48214 30304 48354 30318
rect 48504 30304 49312 30318
rect 49462 30304 49602 30318
rect 49752 30304 50560 30318
rect 50710 30304 50850 30318
rect 51000 30304 51808 30318
rect 51958 30304 52098 30318
rect 52248 30304 53056 30318
rect 53206 30304 53346 30318
rect 53496 30304 54304 30318
rect 54454 30304 54594 30318
rect 54744 30304 55552 30318
rect 55702 30304 55842 30318
rect 55992 30304 56800 30318
rect 56950 30304 57090 30318
rect 57240 30304 58048 30318
rect 58198 30304 58338 30318
rect 58488 30304 58934 30318
rect 16418 30256 58934 30304
rect 16418 30242 16864 30256
rect 17014 30242 17154 30256
rect 17304 30242 18112 30256
rect 18262 30242 18402 30256
rect 18552 30242 19360 30256
rect 19510 30242 19650 30256
rect 19800 30242 20608 30256
rect 20758 30242 20898 30256
rect 21048 30242 21856 30256
rect 22006 30242 22146 30256
rect 22296 30242 23104 30256
rect 23254 30242 23394 30256
rect 23544 30242 24352 30256
rect 24502 30242 24642 30256
rect 24792 30242 25600 30256
rect 25750 30242 25890 30256
rect 26040 30242 26848 30256
rect 26998 30242 27138 30256
rect 27288 30242 28096 30256
rect 28246 30242 28386 30256
rect 28536 30242 29344 30256
rect 29494 30242 29634 30256
rect 29784 30242 30592 30256
rect 30742 30242 30882 30256
rect 31032 30242 31840 30256
rect 31990 30242 32130 30256
rect 32280 30242 33088 30256
rect 33238 30242 33378 30256
rect 33528 30242 34336 30256
rect 34486 30242 34626 30256
rect 34776 30242 35584 30256
rect 35734 30242 35874 30256
rect 36024 30242 36832 30256
rect 36982 30242 37122 30256
rect 37272 30242 38080 30256
rect 38230 30242 38370 30256
rect 38520 30242 39328 30256
rect 39478 30242 39618 30256
rect 39768 30242 40576 30256
rect 40726 30242 40866 30256
rect 41016 30242 41824 30256
rect 41974 30242 42114 30256
rect 42264 30242 43072 30256
rect 43222 30242 43362 30256
rect 43512 30242 44320 30256
rect 44470 30242 44610 30256
rect 44760 30242 45568 30256
rect 45718 30242 45858 30256
rect 46008 30242 46816 30256
rect 46966 30242 47106 30256
rect 47256 30242 48064 30256
rect 48214 30242 48354 30256
rect 48504 30242 49312 30256
rect 49462 30242 49602 30256
rect 49752 30242 50560 30256
rect 50710 30242 50850 30256
rect 51000 30242 51808 30256
rect 51958 30242 52098 30256
rect 52248 30242 53056 30256
rect 53206 30242 53346 30256
rect 53496 30242 54304 30256
rect 54454 30242 54594 30256
rect 54744 30242 55552 30256
rect 55702 30242 55842 30256
rect 55992 30242 56800 30256
rect 56950 30242 57090 30256
rect 57240 30242 58048 30256
rect 58198 30242 58338 30256
rect 58488 30242 58934 30256
rect 16898 30194 16980 30208
rect 17188 30194 17270 30208
rect 18146 30194 18228 30208
rect 18436 30194 18518 30208
rect 19394 30194 19476 30208
rect 19684 30194 19766 30208
rect 20642 30194 20724 30208
rect 20932 30194 21014 30208
rect 21890 30194 21972 30208
rect 22180 30194 22262 30208
rect 23138 30194 23220 30208
rect 23428 30194 23510 30208
rect 24386 30194 24468 30208
rect 24676 30194 24758 30208
rect 25634 30194 25716 30208
rect 25924 30194 26006 30208
rect 26882 30194 26964 30208
rect 27172 30194 27254 30208
rect 28130 30194 28212 30208
rect 28420 30194 28502 30208
rect 29378 30194 29460 30208
rect 29668 30194 29750 30208
rect 30626 30194 30708 30208
rect 30916 30194 30998 30208
rect 31874 30194 31956 30208
rect 32164 30194 32246 30208
rect 33122 30194 33204 30208
rect 33412 30194 33494 30208
rect 34370 30194 34452 30208
rect 34660 30194 34742 30208
rect 35618 30194 35700 30208
rect 35908 30194 35990 30208
rect 36866 30194 36948 30208
rect 37156 30194 37238 30208
rect 38114 30194 38196 30208
rect 38404 30194 38486 30208
rect 39362 30194 39444 30208
rect 39652 30194 39734 30208
rect 40610 30194 40692 30208
rect 40900 30194 40982 30208
rect 41858 30194 41940 30208
rect 42148 30194 42230 30208
rect 43106 30194 43188 30208
rect 43396 30194 43478 30208
rect 44354 30194 44436 30208
rect 44644 30194 44726 30208
rect 45602 30194 45684 30208
rect 45892 30194 45974 30208
rect 46850 30194 46932 30208
rect 47140 30194 47222 30208
rect 48098 30194 48180 30208
rect 48388 30194 48470 30208
rect 49346 30194 49428 30208
rect 49636 30194 49718 30208
rect 50594 30194 50676 30208
rect 50884 30194 50966 30208
rect 51842 30194 51924 30208
rect 52132 30194 52214 30208
rect 53090 30194 53172 30208
rect 53380 30194 53462 30208
rect 54338 30194 54420 30208
rect 54628 30194 54710 30208
rect 55586 30194 55668 30208
rect 55876 30194 55958 30208
rect 56834 30194 56916 30208
rect 57124 30194 57206 30208
rect 58082 30194 58164 30208
rect 58372 30194 58454 30208
rect 16418 30146 58934 30194
rect 16418 29988 58934 30098
rect 16418 29892 58934 29940
rect 16898 29878 16980 29892
rect 17188 29878 17270 29892
rect 18146 29878 18228 29892
rect 18436 29878 18518 29892
rect 19394 29878 19476 29892
rect 19684 29878 19766 29892
rect 20642 29878 20724 29892
rect 20932 29878 21014 29892
rect 21890 29878 21972 29892
rect 22180 29878 22262 29892
rect 23138 29878 23220 29892
rect 23428 29878 23510 29892
rect 24386 29878 24468 29892
rect 24676 29878 24758 29892
rect 25634 29878 25716 29892
rect 25924 29878 26006 29892
rect 26882 29878 26964 29892
rect 27172 29878 27254 29892
rect 28130 29878 28212 29892
rect 28420 29878 28502 29892
rect 29378 29878 29460 29892
rect 29668 29878 29750 29892
rect 30626 29878 30708 29892
rect 30916 29878 30998 29892
rect 31874 29878 31956 29892
rect 32164 29878 32246 29892
rect 33122 29878 33204 29892
rect 33412 29878 33494 29892
rect 34370 29878 34452 29892
rect 34660 29878 34742 29892
rect 35618 29878 35700 29892
rect 35908 29878 35990 29892
rect 36866 29878 36948 29892
rect 37156 29878 37238 29892
rect 38114 29878 38196 29892
rect 38404 29878 38486 29892
rect 39362 29878 39444 29892
rect 39652 29878 39734 29892
rect 40610 29878 40692 29892
rect 40900 29878 40982 29892
rect 41858 29878 41940 29892
rect 42148 29878 42230 29892
rect 43106 29878 43188 29892
rect 43396 29878 43478 29892
rect 44354 29878 44436 29892
rect 44644 29878 44726 29892
rect 45602 29878 45684 29892
rect 45892 29878 45974 29892
rect 46850 29878 46932 29892
rect 47140 29878 47222 29892
rect 48098 29878 48180 29892
rect 48388 29878 48470 29892
rect 49346 29878 49428 29892
rect 49636 29878 49718 29892
rect 50594 29878 50676 29892
rect 50884 29878 50966 29892
rect 51842 29878 51924 29892
rect 52132 29878 52214 29892
rect 53090 29878 53172 29892
rect 53380 29878 53462 29892
rect 54338 29878 54420 29892
rect 54628 29878 54710 29892
rect 55586 29878 55668 29892
rect 55876 29878 55958 29892
rect 56834 29878 56916 29892
rect 57124 29878 57206 29892
rect 58082 29878 58164 29892
rect 58372 29878 58454 29892
rect 16418 29830 16864 29844
rect 17014 29830 17154 29844
rect 17304 29830 18112 29844
rect 18262 29830 18402 29844
rect 18552 29830 19360 29844
rect 19510 29830 19650 29844
rect 19800 29830 20608 29844
rect 20758 29830 20898 29844
rect 21048 29830 21856 29844
rect 22006 29830 22146 29844
rect 22296 29830 23104 29844
rect 23254 29830 23394 29844
rect 23544 29830 24352 29844
rect 24502 29830 24642 29844
rect 24792 29830 25600 29844
rect 25750 29830 25890 29844
rect 26040 29830 26848 29844
rect 26998 29830 27138 29844
rect 27288 29830 28096 29844
rect 28246 29830 28386 29844
rect 28536 29830 29344 29844
rect 29494 29830 29634 29844
rect 29784 29830 30592 29844
rect 30742 29830 30882 29844
rect 31032 29830 31840 29844
rect 31990 29830 32130 29844
rect 32280 29830 33088 29844
rect 33238 29830 33378 29844
rect 33528 29830 34336 29844
rect 34486 29830 34626 29844
rect 34776 29830 35584 29844
rect 35734 29830 35874 29844
rect 36024 29830 36832 29844
rect 36982 29830 37122 29844
rect 37272 29830 38080 29844
rect 38230 29830 38370 29844
rect 38520 29830 39328 29844
rect 39478 29830 39618 29844
rect 39768 29830 40576 29844
rect 40726 29830 40866 29844
rect 41016 29830 41824 29844
rect 41974 29830 42114 29844
rect 42264 29830 43072 29844
rect 43222 29830 43362 29844
rect 43512 29830 44320 29844
rect 44470 29830 44610 29844
rect 44760 29830 45568 29844
rect 45718 29830 45858 29844
rect 46008 29830 46816 29844
rect 46966 29830 47106 29844
rect 47256 29830 48064 29844
rect 48214 29830 48354 29844
rect 48504 29830 49312 29844
rect 49462 29830 49602 29844
rect 49752 29830 50560 29844
rect 50710 29830 50850 29844
rect 51000 29830 51808 29844
rect 51958 29830 52098 29844
rect 52248 29830 53056 29844
rect 53206 29830 53346 29844
rect 53496 29830 54304 29844
rect 54454 29830 54594 29844
rect 54744 29830 55552 29844
rect 55702 29830 55842 29844
rect 55992 29830 56800 29844
rect 56950 29830 57090 29844
rect 57240 29830 58048 29844
rect 58198 29830 58338 29844
rect 58488 29830 58934 29844
rect 16418 29782 58934 29830
rect 16418 29768 16864 29782
rect 17014 29768 17154 29782
rect 17304 29768 18112 29782
rect 18262 29768 18402 29782
rect 18552 29768 19360 29782
rect 19510 29768 19650 29782
rect 19800 29768 20608 29782
rect 20758 29768 20898 29782
rect 21048 29768 21856 29782
rect 22006 29768 22146 29782
rect 22296 29768 23104 29782
rect 23254 29768 23394 29782
rect 23544 29768 24352 29782
rect 24502 29768 24642 29782
rect 24792 29768 25600 29782
rect 25750 29768 25890 29782
rect 26040 29768 26848 29782
rect 26998 29768 27138 29782
rect 27288 29768 28096 29782
rect 28246 29768 28386 29782
rect 28536 29768 29344 29782
rect 29494 29768 29634 29782
rect 29784 29768 30592 29782
rect 30742 29768 30882 29782
rect 31032 29768 31840 29782
rect 31990 29768 32130 29782
rect 32280 29768 33088 29782
rect 33238 29768 33378 29782
rect 33528 29768 34336 29782
rect 34486 29768 34626 29782
rect 34776 29768 35584 29782
rect 35734 29768 35874 29782
rect 36024 29768 36832 29782
rect 36982 29768 37122 29782
rect 37272 29768 38080 29782
rect 38230 29768 38370 29782
rect 38520 29768 39328 29782
rect 39478 29768 39618 29782
rect 39768 29768 40576 29782
rect 40726 29768 40866 29782
rect 41016 29768 41824 29782
rect 41974 29768 42114 29782
rect 42264 29768 43072 29782
rect 43222 29768 43362 29782
rect 43512 29768 44320 29782
rect 44470 29768 44610 29782
rect 44760 29768 45568 29782
rect 45718 29768 45858 29782
rect 46008 29768 46816 29782
rect 46966 29768 47106 29782
rect 47256 29768 48064 29782
rect 48214 29768 48354 29782
rect 48504 29768 49312 29782
rect 49462 29768 49602 29782
rect 49752 29768 50560 29782
rect 50710 29768 50850 29782
rect 51000 29768 51808 29782
rect 51958 29768 52098 29782
rect 52248 29768 53056 29782
rect 53206 29768 53346 29782
rect 53496 29768 54304 29782
rect 54454 29768 54594 29782
rect 54744 29768 55552 29782
rect 55702 29768 55842 29782
rect 55992 29768 56800 29782
rect 56950 29768 57090 29782
rect 57240 29768 58048 29782
rect 58198 29768 58338 29782
rect 58488 29768 58934 29782
rect 16898 29720 16980 29734
rect 17188 29720 17270 29734
rect 18146 29720 18228 29734
rect 18436 29720 18518 29734
rect 19394 29720 19476 29734
rect 19684 29720 19766 29734
rect 20642 29720 20724 29734
rect 20932 29720 21014 29734
rect 21890 29720 21972 29734
rect 22180 29720 22262 29734
rect 23138 29720 23220 29734
rect 23428 29720 23510 29734
rect 24386 29720 24468 29734
rect 24676 29720 24758 29734
rect 25634 29720 25716 29734
rect 25924 29720 26006 29734
rect 26882 29720 26964 29734
rect 27172 29720 27254 29734
rect 28130 29720 28212 29734
rect 28420 29720 28502 29734
rect 29378 29720 29460 29734
rect 29668 29720 29750 29734
rect 30626 29720 30708 29734
rect 30916 29720 30998 29734
rect 31874 29720 31956 29734
rect 32164 29720 32246 29734
rect 33122 29720 33204 29734
rect 33412 29720 33494 29734
rect 34370 29720 34452 29734
rect 34660 29720 34742 29734
rect 35618 29720 35700 29734
rect 35908 29720 35990 29734
rect 36866 29720 36948 29734
rect 37156 29720 37238 29734
rect 38114 29720 38196 29734
rect 38404 29720 38486 29734
rect 39362 29720 39444 29734
rect 39652 29720 39734 29734
rect 40610 29720 40692 29734
rect 40900 29720 40982 29734
rect 41858 29720 41940 29734
rect 42148 29720 42230 29734
rect 43106 29720 43188 29734
rect 43396 29720 43478 29734
rect 44354 29720 44436 29734
rect 44644 29720 44726 29734
rect 45602 29720 45684 29734
rect 45892 29720 45974 29734
rect 46850 29720 46932 29734
rect 47140 29720 47222 29734
rect 48098 29720 48180 29734
rect 48388 29720 48470 29734
rect 49346 29720 49428 29734
rect 49636 29720 49718 29734
rect 50594 29720 50676 29734
rect 50884 29720 50966 29734
rect 51842 29720 51924 29734
rect 52132 29720 52214 29734
rect 53090 29720 53172 29734
rect 53380 29720 53462 29734
rect 54338 29720 54420 29734
rect 54628 29720 54710 29734
rect 55586 29720 55668 29734
rect 55876 29720 55958 29734
rect 56834 29720 56916 29734
rect 57124 29720 57206 29734
rect 58082 29720 58164 29734
rect 58372 29720 58454 29734
rect 16418 29672 58934 29720
rect 16418 29576 58934 29624
rect 16898 29562 16980 29576
rect 17188 29562 17270 29576
rect 18146 29562 18228 29576
rect 18436 29562 18518 29576
rect 19394 29562 19476 29576
rect 19684 29562 19766 29576
rect 20642 29562 20724 29576
rect 20932 29562 21014 29576
rect 21890 29562 21972 29576
rect 22180 29562 22262 29576
rect 23138 29562 23220 29576
rect 23428 29562 23510 29576
rect 24386 29562 24468 29576
rect 24676 29562 24758 29576
rect 25634 29562 25716 29576
rect 25924 29562 26006 29576
rect 26882 29562 26964 29576
rect 27172 29562 27254 29576
rect 28130 29562 28212 29576
rect 28420 29562 28502 29576
rect 29378 29562 29460 29576
rect 29668 29562 29750 29576
rect 30626 29562 30708 29576
rect 30916 29562 30998 29576
rect 31874 29562 31956 29576
rect 32164 29562 32246 29576
rect 33122 29562 33204 29576
rect 33412 29562 33494 29576
rect 34370 29562 34452 29576
rect 34660 29562 34742 29576
rect 35618 29562 35700 29576
rect 35908 29562 35990 29576
rect 36866 29562 36948 29576
rect 37156 29562 37238 29576
rect 38114 29562 38196 29576
rect 38404 29562 38486 29576
rect 39362 29562 39444 29576
rect 39652 29562 39734 29576
rect 40610 29562 40692 29576
rect 40900 29562 40982 29576
rect 41858 29562 41940 29576
rect 42148 29562 42230 29576
rect 43106 29562 43188 29576
rect 43396 29562 43478 29576
rect 44354 29562 44436 29576
rect 44644 29562 44726 29576
rect 45602 29562 45684 29576
rect 45892 29562 45974 29576
rect 46850 29562 46932 29576
rect 47140 29562 47222 29576
rect 48098 29562 48180 29576
rect 48388 29562 48470 29576
rect 49346 29562 49428 29576
rect 49636 29562 49718 29576
rect 50594 29562 50676 29576
rect 50884 29562 50966 29576
rect 51842 29562 51924 29576
rect 52132 29562 52214 29576
rect 53090 29562 53172 29576
rect 53380 29562 53462 29576
rect 54338 29562 54420 29576
rect 54628 29562 54710 29576
rect 55586 29562 55668 29576
rect 55876 29562 55958 29576
rect 56834 29562 56916 29576
rect 57124 29562 57206 29576
rect 58082 29562 58164 29576
rect 58372 29562 58454 29576
rect 16418 29514 16864 29528
rect 17014 29514 17154 29528
rect 17304 29514 18112 29528
rect 18262 29514 18402 29528
rect 18552 29514 19360 29528
rect 19510 29514 19650 29528
rect 19800 29514 20608 29528
rect 20758 29514 20898 29528
rect 21048 29514 21856 29528
rect 22006 29514 22146 29528
rect 22296 29514 23104 29528
rect 23254 29514 23394 29528
rect 23544 29514 24352 29528
rect 24502 29514 24642 29528
rect 24792 29514 25600 29528
rect 25750 29514 25890 29528
rect 26040 29514 26848 29528
rect 26998 29514 27138 29528
rect 27288 29514 28096 29528
rect 28246 29514 28386 29528
rect 28536 29514 29344 29528
rect 29494 29514 29634 29528
rect 29784 29514 30592 29528
rect 30742 29514 30882 29528
rect 31032 29514 31840 29528
rect 31990 29514 32130 29528
rect 32280 29514 33088 29528
rect 33238 29514 33378 29528
rect 33528 29514 34336 29528
rect 34486 29514 34626 29528
rect 34776 29514 35584 29528
rect 35734 29514 35874 29528
rect 36024 29514 36832 29528
rect 36982 29514 37122 29528
rect 37272 29514 38080 29528
rect 38230 29514 38370 29528
rect 38520 29514 39328 29528
rect 39478 29514 39618 29528
rect 39768 29514 40576 29528
rect 40726 29514 40866 29528
rect 41016 29514 41824 29528
rect 41974 29514 42114 29528
rect 42264 29514 43072 29528
rect 43222 29514 43362 29528
rect 43512 29514 44320 29528
rect 44470 29514 44610 29528
rect 44760 29514 45568 29528
rect 45718 29514 45858 29528
rect 46008 29514 46816 29528
rect 46966 29514 47106 29528
rect 47256 29514 48064 29528
rect 48214 29514 48354 29528
rect 48504 29514 49312 29528
rect 49462 29514 49602 29528
rect 49752 29514 50560 29528
rect 50710 29514 50850 29528
rect 51000 29514 51808 29528
rect 51958 29514 52098 29528
rect 52248 29514 53056 29528
rect 53206 29514 53346 29528
rect 53496 29514 54304 29528
rect 54454 29514 54594 29528
rect 54744 29514 55552 29528
rect 55702 29514 55842 29528
rect 55992 29514 56800 29528
rect 56950 29514 57090 29528
rect 57240 29514 58048 29528
rect 58198 29514 58338 29528
rect 58488 29514 58934 29528
rect 16418 29466 58934 29514
rect 16418 29452 16864 29466
rect 17014 29452 17154 29466
rect 17304 29452 18112 29466
rect 18262 29452 18402 29466
rect 18552 29452 19360 29466
rect 19510 29452 19650 29466
rect 19800 29452 20608 29466
rect 20758 29452 20898 29466
rect 21048 29452 21856 29466
rect 22006 29452 22146 29466
rect 22296 29452 23104 29466
rect 23254 29452 23394 29466
rect 23544 29452 24352 29466
rect 24502 29452 24642 29466
rect 24792 29452 25600 29466
rect 25750 29452 25890 29466
rect 26040 29452 26848 29466
rect 26998 29452 27138 29466
rect 27288 29452 28096 29466
rect 28246 29452 28386 29466
rect 28536 29452 29344 29466
rect 29494 29452 29634 29466
rect 29784 29452 30592 29466
rect 30742 29452 30882 29466
rect 31032 29452 31840 29466
rect 31990 29452 32130 29466
rect 32280 29452 33088 29466
rect 33238 29452 33378 29466
rect 33528 29452 34336 29466
rect 34486 29452 34626 29466
rect 34776 29452 35584 29466
rect 35734 29452 35874 29466
rect 36024 29452 36832 29466
rect 36982 29452 37122 29466
rect 37272 29452 38080 29466
rect 38230 29452 38370 29466
rect 38520 29452 39328 29466
rect 39478 29452 39618 29466
rect 39768 29452 40576 29466
rect 40726 29452 40866 29466
rect 41016 29452 41824 29466
rect 41974 29452 42114 29466
rect 42264 29452 43072 29466
rect 43222 29452 43362 29466
rect 43512 29452 44320 29466
rect 44470 29452 44610 29466
rect 44760 29452 45568 29466
rect 45718 29452 45858 29466
rect 46008 29452 46816 29466
rect 46966 29452 47106 29466
rect 47256 29452 48064 29466
rect 48214 29452 48354 29466
rect 48504 29452 49312 29466
rect 49462 29452 49602 29466
rect 49752 29452 50560 29466
rect 50710 29452 50850 29466
rect 51000 29452 51808 29466
rect 51958 29452 52098 29466
rect 52248 29452 53056 29466
rect 53206 29452 53346 29466
rect 53496 29452 54304 29466
rect 54454 29452 54594 29466
rect 54744 29452 55552 29466
rect 55702 29452 55842 29466
rect 55992 29452 56800 29466
rect 56950 29452 57090 29466
rect 57240 29452 58048 29466
rect 58198 29452 58338 29466
rect 58488 29452 58934 29466
rect 16898 29404 16980 29418
rect 17188 29404 17270 29418
rect 18146 29404 18228 29418
rect 18436 29404 18518 29418
rect 19394 29404 19476 29418
rect 19684 29404 19766 29418
rect 20642 29404 20724 29418
rect 20932 29404 21014 29418
rect 21890 29404 21972 29418
rect 22180 29404 22262 29418
rect 23138 29404 23220 29418
rect 23428 29404 23510 29418
rect 24386 29404 24468 29418
rect 24676 29404 24758 29418
rect 25634 29404 25716 29418
rect 25924 29404 26006 29418
rect 26882 29404 26964 29418
rect 27172 29404 27254 29418
rect 28130 29404 28212 29418
rect 28420 29404 28502 29418
rect 29378 29404 29460 29418
rect 29668 29404 29750 29418
rect 30626 29404 30708 29418
rect 30916 29404 30998 29418
rect 31874 29404 31956 29418
rect 32164 29404 32246 29418
rect 33122 29404 33204 29418
rect 33412 29404 33494 29418
rect 34370 29404 34452 29418
rect 34660 29404 34742 29418
rect 35618 29404 35700 29418
rect 35908 29404 35990 29418
rect 36866 29404 36948 29418
rect 37156 29404 37238 29418
rect 38114 29404 38196 29418
rect 38404 29404 38486 29418
rect 39362 29404 39444 29418
rect 39652 29404 39734 29418
rect 40610 29404 40692 29418
rect 40900 29404 40982 29418
rect 41858 29404 41940 29418
rect 42148 29404 42230 29418
rect 43106 29404 43188 29418
rect 43396 29404 43478 29418
rect 44354 29404 44436 29418
rect 44644 29404 44726 29418
rect 45602 29404 45684 29418
rect 45892 29404 45974 29418
rect 46850 29404 46932 29418
rect 47140 29404 47222 29418
rect 48098 29404 48180 29418
rect 48388 29404 48470 29418
rect 49346 29404 49428 29418
rect 49636 29404 49718 29418
rect 50594 29404 50676 29418
rect 50884 29404 50966 29418
rect 51842 29404 51924 29418
rect 52132 29404 52214 29418
rect 53090 29404 53172 29418
rect 53380 29404 53462 29418
rect 54338 29404 54420 29418
rect 54628 29404 54710 29418
rect 55586 29404 55668 29418
rect 55876 29404 55958 29418
rect 56834 29404 56916 29418
rect 57124 29404 57206 29418
rect 58082 29404 58164 29418
rect 58372 29404 58454 29418
rect 16418 29356 58934 29404
rect 16418 29198 58934 29308
rect 63080 29253 63108 79813
rect 75079 71121 75107 80603
rect 16418 29102 58934 29150
rect 1804 28463 1832 28985
rect 3426 27582 4494 27610
rect 4300 24754 4494 24782
rect 3426 23340 4494 23368
rect 4348 21926 4494 21954
rect 193 19229 259 19281
rect 425 19127 453 19819
rect 1060 19309 1126 19361
rect 1912 19300 1940 19328
rect 1138 19158 1204 19210
rect 425 19063 479 19127
rect 15840 19078 15868 29093
rect 15964 19078 15992 29093
rect 16088 19078 16116 29093
rect 16212 19078 16240 29093
rect 16898 29088 16980 29102
rect 17188 29088 17270 29102
rect 18146 29088 18228 29102
rect 18436 29088 18518 29102
rect 19394 29088 19476 29102
rect 19684 29088 19766 29102
rect 20642 29088 20724 29102
rect 20932 29088 21014 29102
rect 21890 29088 21972 29102
rect 22180 29088 22262 29102
rect 23138 29088 23220 29102
rect 23428 29088 23510 29102
rect 24386 29088 24468 29102
rect 24676 29088 24758 29102
rect 25634 29088 25716 29102
rect 25924 29088 26006 29102
rect 26882 29088 26964 29102
rect 27172 29088 27254 29102
rect 28130 29088 28212 29102
rect 28420 29088 28502 29102
rect 29378 29088 29460 29102
rect 29668 29088 29750 29102
rect 30626 29088 30708 29102
rect 30916 29088 30998 29102
rect 31874 29088 31956 29102
rect 32164 29088 32246 29102
rect 33122 29088 33204 29102
rect 33412 29088 33494 29102
rect 34370 29088 34452 29102
rect 34660 29088 34742 29102
rect 35618 29088 35700 29102
rect 35908 29088 35990 29102
rect 36866 29088 36948 29102
rect 37156 29088 37238 29102
rect 38114 29088 38196 29102
rect 38404 29088 38486 29102
rect 39362 29088 39444 29102
rect 39652 29088 39734 29102
rect 40610 29088 40692 29102
rect 40900 29088 40982 29102
rect 41858 29088 41940 29102
rect 42148 29088 42230 29102
rect 43106 29088 43188 29102
rect 43396 29088 43478 29102
rect 44354 29088 44436 29102
rect 44644 29088 44726 29102
rect 45602 29088 45684 29102
rect 45892 29088 45974 29102
rect 46850 29088 46932 29102
rect 47140 29088 47222 29102
rect 48098 29088 48180 29102
rect 48388 29088 48470 29102
rect 49346 29088 49428 29102
rect 49636 29088 49718 29102
rect 50594 29088 50676 29102
rect 50884 29088 50966 29102
rect 51842 29088 51924 29102
rect 52132 29088 52214 29102
rect 53090 29088 53172 29102
rect 53380 29088 53462 29102
rect 54338 29088 54420 29102
rect 54628 29088 54710 29102
rect 55586 29088 55668 29102
rect 55876 29088 55958 29102
rect 56834 29088 56916 29102
rect 57124 29088 57206 29102
rect 58082 29088 58164 29102
rect 58372 29088 58454 29102
rect 16418 29040 16864 29054
rect 17014 29040 17154 29054
rect 17304 29040 18112 29054
rect 18262 29040 18402 29054
rect 18552 29040 19360 29054
rect 19510 29040 19650 29054
rect 19800 29040 20608 29054
rect 20758 29040 20898 29054
rect 21048 29040 21856 29054
rect 22006 29040 22146 29054
rect 22296 29040 23104 29054
rect 23254 29040 23394 29054
rect 23544 29040 24352 29054
rect 24502 29040 24642 29054
rect 24792 29040 25600 29054
rect 25750 29040 25890 29054
rect 26040 29040 26848 29054
rect 26998 29040 27138 29054
rect 27288 29040 28096 29054
rect 28246 29040 28386 29054
rect 28536 29040 29344 29054
rect 29494 29040 29634 29054
rect 29784 29040 30592 29054
rect 30742 29040 30882 29054
rect 31032 29040 31840 29054
rect 31990 29040 32130 29054
rect 32280 29040 33088 29054
rect 33238 29040 33378 29054
rect 33528 29040 34336 29054
rect 34486 29040 34626 29054
rect 34776 29040 35584 29054
rect 35734 29040 35874 29054
rect 36024 29040 36832 29054
rect 36982 29040 37122 29054
rect 37272 29040 38080 29054
rect 38230 29040 38370 29054
rect 38520 29040 39328 29054
rect 39478 29040 39618 29054
rect 39768 29040 40576 29054
rect 40726 29040 40866 29054
rect 41016 29040 41824 29054
rect 41974 29040 42114 29054
rect 42264 29040 43072 29054
rect 43222 29040 43362 29054
rect 43512 29040 44320 29054
rect 44470 29040 44610 29054
rect 44760 29040 45568 29054
rect 45718 29040 45858 29054
rect 46008 29040 46816 29054
rect 46966 29040 47106 29054
rect 47256 29040 48064 29054
rect 48214 29040 48354 29054
rect 48504 29040 49312 29054
rect 49462 29040 49602 29054
rect 49752 29040 50560 29054
rect 50710 29040 50850 29054
rect 51000 29040 51808 29054
rect 51958 29040 52098 29054
rect 52248 29040 53056 29054
rect 53206 29040 53346 29054
rect 53496 29040 54304 29054
rect 54454 29040 54594 29054
rect 54744 29040 55552 29054
rect 55702 29040 55842 29054
rect 55992 29040 56800 29054
rect 56950 29040 57090 29054
rect 57240 29040 58048 29054
rect 58198 29040 58338 29054
rect 58488 29040 58934 29054
rect 16418 28992 58934 29040
rect 16418 28978 16864 28992
rect 17014 28978 17154 28992
rect 17304 28978 18112 28992
rect 18262 28978 18402 28992
rect 18552 28978 19360 28992
rect 19510 28978 19650 28992
rect 19800 28978 20608 28992
rect 20758 28978 20898 28992
rect 21048 28978 21856 28992
rect 22006 28978 22146 28992
rect 22296 28978 23104 28992
rect 23254 28978 23394 28992
rect 23544 28978 24352 28992
rect 24502 28978 24642 28992
rect 24792 28978 25600 28992
rect 25750 28978 25890 28992
rect 26040 28978 26848 28992
rect 26998 28978 27138 28992
rect 27288 28978 28096 28992
rect 28246 28978 28386 28992
rect 28536 28978 29344 28992
rect 29494 28978 29634 28992
rect 29784 28978 30592 28992
rect 30742 28978 30882 28992
rect 31032 28978 31840 28992
rect 31990 28978 32130 28992
rect 32280 28978 33088 28992
rect 33238 28978 33378 28992
rect 33528 28978 34336 28992
rect 34486 28978 34626 28992
rect 34776 28978 35584 28992
rect 35734 28978 35874 28992
rect 36024 28978 36832 28992
rect 36982 28978 37122 28992
rect 37272 28978 38080 28992
rect 38230 28978 38370 28992
rect 38520 28978 39328 28992
rect 39478 28978 39618 28992
rect 39768 28978 40576 28992
rect 40726 28978 40866 28992
rect 41016 28978 41824 28992
rect 41974 28978 42114 28992
rect 42264 28978 43072 28992
rect 43222 28978 43362 28992
rect 43512 28978 44320 28992
rect 44470 28978 44610 28992
rect 44760 28978 45568 28992
rect 45718 28978 45858 28992
rect 46008 28978 46816 28992
rect 46966 28978 47106 28992
rect 47256 28978 48064 28992
rect 48214 28978 48354 28992
rect 48504 28978 49312 28992
rect 49462 28978 49602 28992
rect 49752 28978 50560 28992
rect 50710 28978 50850 28992
rect 51000 28978 51808 28992
rect 51958 28978 52098 28992
rect 52248 28978 53056 28992
rect 53206 28978 53346 28992
rect 53496 28978 54304 28992
rect 54454 28978 54594 28992
rect 54744 28978 55552 28992
rect 55702 28978 55842 28992
rect 55992 28978 56800 28992
rect 56950 28978 57090 28992
rect 57240 28978 58048 28992
rect 58198 28978 58338 28992
rect 58488 28978 58934 28992
rect 16898 28930 16980 28944
rect 17188 28930 17270 28944
rect 18146 28930 18228 28944
rect 18436 28930 18518 28944
rect 19394 28930 19476 28944
rect 19684 28930 19766 28944
rect 20642 28930 20724 28944
rect 20932 28930 21014 28944
rect 21890 28930 21972 28944
rect 22180 28930 22262 28944
rect 23138 28930 23220 28944
rect 23428 28930 23510 28944
rect 24386 28930 24468 28944
rect 24676 28930 24758 28944
rect 25634 28930 25716 28944
rect 25924 28930 26006 28944
rect 26882 28930 26964 28944
rect 27172 28930 27254 28944
rect 28130 28930 28212 28944
rect 28420 28930 28502 28944
rect 29378 28930 29460 28944
rect 29668 28930 29750 28944
rect 30626 28930 30708 28944
rect 30916 28930 30998 28944
rect 31874 28930 31956 28944
rect 32164 28930 32246 28944
rect 33122 28930 33204 28944
rect 33412 28930 33494 28944
rect 34370 28930 34452 28944
rect 34660 28930 34742 28944
rect 35618 28930 35700 28944
rect 35908 28930 35990 28944
rect 36866 28930 36948 28944
rect 37156 28930 37238 28944
rect 38114 28930 38196 28944
rect 38404 28930 38486 28944
rect 39362 28930 39444 28944
rect 39652 28930 39734 28944
rect 40610 28930 40692 28944
rect 40900 28930 40982 28944
rect 41858 28930 41940 28944
rect 42148 28930 42230 28944
rect 43106 28930 43188 28944
rect 43396 28930 43478 28944
rect 44354 28930 44436 28944
rect 44644 28930 44726 28944
rect 45602 28930 45684 28944
rect 45892 28930 45974 28944
rect 46850 28930 46932 28944
rect 47140 28930 47222 28944
rect 48098 28930 48180 28944
rect 48388 28930 48470 28944
rect 49346 28930 49428 28944
rect 49636 28930 49718 28944
rect 50594 28930 50676 28944
rect 50884 28930 50966 28944
rect 51842 28930 51924 28944
rect 52132 28930 52214 28944
rect 53090 28930 53172 28944
rect 53380 28930 53462 28944
rect 54338 28930 54420 28944
rect 54628 28930 54710 28944
rect 55586 28930 55668 28944
rect 55876 28930 55958 28944
rect 56834 28930 56916 28944
rect 57124 28930 57206 28944
rect 58082 28930 58164 28944
rect 58372 28930 58454 28944
rect 16418 28882 58934 28930
rect 17084 28637 58268 28747
rect 71040 28466 71106 28518
rect 71907 28386 71973 28438
rect 70962 28315 71028 28367
rect 71687 28220 71741 28284
rect 17084 27468 57644 27496
rect 71687 26840 71741 26904
rect 70962 26757 71028 26809
rect 71907 26686 71973 26738
rect 71040 26606 71106 26658
rect 71040 25638 71106 25690
rect 71907 25558 71973 25610
rect 70962 25487 71028 25539
rect 71687 25392 71741 25456
rect 71687 24012 71741 24076
rect 70962 23929 71028 23981
rect 71907 23858 71973 23910
rect 71040 23778 71106 23830
rect 71040 22810 71106 22862
rect 71907 22730 71973 22782
rect 70962 22659 71028 22711
rect 71687 22564 71741 22628
rect 71687 21184 71741 21248
rect 70962 21101 71028 21153
rect 71907 21030 71973 21082
rect 71040 20950 71106 21002
rect 71040 19982 71106 20034
rect 71907 19902 71973 19954
rect 70962 19831 71028 19883
rect 71687 19736 71741 19800
rect 17694 19334 17722 19362
rect 27678 19334 27706 19362
rect 37662 19334 37690 19362
rect 47646 19334 47674 19362
rect 425 17747 453 19063
rect 1568 18913 1596 18941
rect 1568 17869 1596 17897
rect 425 17683 479 17747
rect 4348 17684 4494 17712
rect 193 17529 259 17581
rect 425 16991 453 17683
rect 1138 17600 1204 17652
rect 2819 17646 2847 17674
rect 1060 17449 1126 17501
rect 1912 17482 1940 17510
rect 6031 788 6085 852
rect 7199 788 7253 852
rect 8367 788 8421 852
rect 9535 788 9589 852
rect 10703 788 10757 852
rect 11871 788 11925 852
rect 13039 788 13093 852
rect 14207 788 14261 852
rect 15375 788 15429 852
rect 16543 788 16597 852
rect 17711 788 17765 852
rect 18879 788 18933 852
rect 20047 788 20101 852
rect 21215 788 21269 852
rect 22383 788 22437 852
rect 23551 788 23605 852
rect 24719 788 24773 852
rect 25887 788 25941 852
rect 27055 788 27109 852
rect 28223 788 28277 852
rect 29391 788 29445 852
rect 30559 788 30613 852
rect 31727 788 31781 852
rect 32895 788 32949 852
rect 34063 788 34117 852
rect 35231 788 35285 852
rect 36399 788 36453 852
rect 37567 788 37621 852
rect 38735 788 38789 852
rect 39903 788 39957 852
rect 41071 788 41125 852
rect 42239 788 42293 852
rect 43407 788 43461 852
rect 44575 788 44629 852
rect 45743 788 45797 852
rect 46911 788 46965 852
rect 48079 788 48133 852
rect 6744 705 6810 757
rect 7912 705 7978 757
rect 9080 705 9146 757
rect 10248 705 10314 757
rect 11416 705 11482 757
rect 12584 705 12650 757
rect 13752 705 13818 757
rect 14920 705 14986 757
rect 16088 705 16154 757
rect 17256 705 17322 757
rect 18424 705 18490 757
rect 19592 705 19658 757
rect 20760 705 20826 757
rect 21928 705 21994 757
rect 23096 705 23162 757
rect 24264 705 24330 757
rect 25432 705 25498 757
rect 26600 705 26666 757
rect 27768 705 27834 757
rect 28936 705 29002 757
rect 30104 705 30170 757
rect 31272 705 31338 757
rect 32440 705 32506 757
rect 33608 705 33674 757
rect 34776 705 34842 757
rect 35944 705 36010 757
rect 37112 705 37178 757
rect 38280 705 38346 757
rect 39448 705 39514 757
rect 40616 705 40682 757
rect 41784 705 41850 757
rect 42952 705 43018 757
rect 44120 705 44186 757
rect 45288 705 45354 757
rect 46456 705 46522 757
rect 47624 705 47690 757
rect 48792 705 48858 757
rect 5799 634 5865 686
rect 6967 634 7033 686
rect 8135 634 8201 686
rect 9303 634 9369 686
rect 10471 634 10537 686
rect 11639 634 11705 686
rect 12807 634 12873 686
rect 13975 634 14041 686
rect 15143 634 15209 686
rect 16311 634 16377 686
rect 17479 634 17545 686
rect 18647 634 18713 686
rect 19815 634 19881 686
rect 20983 634 21049 686
rect 22151 634 22217 686
rect 23319 634 23385 686
rect 24487 634 24553 686
rect 25655 634 25721 686
rect 26823 634 26889 686
rect 27991 634 28057 686
rect 29159 634 29225 686
rect 30327 634 30393 686
rect 31495 634 31561 686
rect 32663 634 32729 686
rect 33831 634 33897 686
rect 34999 634 35065 686
rect 36167 634 36233 686
rect 37335 634 37401 686
rect 38503 634 38569 686
rect 39671 634 39737 686
rect 40839 634 40905 686
rect 42007 634 42073 686
rect 43175 634 43241 686
rect 44343 634 44409 686
rect 45511 634 45577 686
rect 46679 634 46745 686
rect 47847 634 47913 686
rect 6666 554 6732 606
rect 7834 554 7900 606
rect 9002 554 9068 606
rect 10170 554 10236 606
rect 11338 554 11404 606
rect 12506 554 12572 606
rect 13674 554 13740 606
rect 14842 554 14908 606
rect 16010 554 16076 606
rect 17178 554 17244 606
rect 18346 554 18412 606
rect 19514 554 19580 606
rect 20682 554 20748 606
rect 21850 554 21916 606
rect 23018 554 23084 606
rect 24186 554 24252 606
rect 25354 554 25420 606
rect 26522 554 26588 606
rect 27690 554 27756 606
rect 28858 554 28924 606
rect 30026 554 30092 606
rect 31194 554 31260 606
rect 32362 554 32428 606
rect 33530 554 33596 606
rect 34698 554 34764 606
rect 35866 554 35932 606
rect 37034 554 37100 606
rect 38202 554 38268 606
rect 39370 554 39436 606
rect 40538 554 40604 606
rect 41706 554 41772 606
rect 42874 554 42940 606
rect 44042 554 44108 606
rect 45210 554 45276 606
rect 46378 554 46444 606
rect 47546 554 47612 606
rect 48714 554 48780 606
<< metal3 >>
rect 0 89080 70660 89156
rect 73304 89080 75012 89156
rect 0 88944 70796 89020
rect 73304 88944 75284 89020
rect 0 88808 67668 88884
rect 68272 88808 72564 88884
rect 73712 88808 75284 88884
rect 0 88672 72564 88748
rect 75266 88653 75326 88713
rect 0 88536 67124 88612
rect 72896 88536 74876 88612
rect 0 88400 67124 88476
rect 0 88264 67260 88340
rect 68000 88264 72564 88340
rect 0 88128 67260 88204
rect 68000 88128 75284 88204
rect 0 87992 75284 88068
rect 0 87856 70660 87932
rect 0 87784 70977 87796
rect 71400 87856 75012 87932
rect 71075 87784 71476 87796
rect 0 87720 71476 87784
rect 73440 87784 75247 87796
rect 73440 87720 75284 87784
rect 0 87584 71476 87660
rect 73440 87584 75284 87660
rect 0 87462 75284 87524
rect 0 87448 67973 87462
rect 0 87312 67668 87388
rect 68071 87448 75284 87462
rect 68272 87312 75284 87388
rect 0 87176 75284 87252
rect 0 87040 75284 87116
rect 0 86904 71748 86980
rect 73168 86904 75284 86980
rect 0 86768 75284 86844
rect 0 86632 75284 86708
rect 0 86496 3612 86572
rect 4080 86496 75284 86572
rect 0 86388 3861 86436
rect 3959 86388 70660 86436
rect 0 86360 70660 86388
rect 71400 86360 75284 86436
rect 0 86224 17484 86300
rect 56848 86224 75284 86300
rect 0 86088 17484 86164
rect 57120 86088 75284 86164
rect 0 85952 17756 86028
rect 0 85874 18040 85892
rect 18138 85874 19288 85892
rect 19386 85874 20536 85892
rect 20634 85874 21784 85892
rect 21882 85874 23032 85892
rect 23130 85874 24280 85892
rect 24378 85874 25528 85892
rect 25626 85874 26776 85892
rect 26874 85874 28024 85892
rect 28122 85874 29272 85892
rect 29370 85874 30520 85892
rect 30618 85874 31768 85892
rect 31866 85874 33016 85892
rect 33114 85874 34264 85892
rect 34362 85874 35512 85892
rect 35610 85874 36760 85892
rect 36858 85874 38008 85892
rect 38106 85874 39256 85892
rect 39354 85874 40504 85892
rect 40602 85874 41752 85892
rect 41850 85874 43000 85892
rect 43098 85874 44248 85892
rect 44346 85874 45496 85892
rect 45594 85874 46744 85892
rect 46842 85874 47992 85892
rect 48090 85874 49240 85892
rect 49338 85874 50488 85892
rect 50586 85874 51736 85892
rect 51834 85874 52984 85892
rect 53082 85874 54232 85892
rect 54330 85874 55480 85892
rect 55578 85874 56728 85892
rect 57120 85952 75284 86028
rect 56826 85874 71748 85892
rect 0 85816 71748 85874
rect 73440 85816 75284 85892
rect 0 85680 3204 85756
rect 5440 85680 71748 85756
rect 73440 85680 75284 85756
rect 26 85557 86 85617
rect 5440 85544 75284 85620
rect 0 85408 75284 85484
rect 0 85272 63724 85348
rect 64328 85272 75284 85348
rect 0 85136 17756 85212
rect 57120 85150 64029 85212
rect 64127 85150 75284 85212
rect 57120 85136 75284 85150
rect 0 85000 3612 85076
rect 4080 85036 18028 85076
rect 18126 85036 19276 85076
rect 19374 85036 20524 85076
rect 20622 85036 21772 85076
rect 21870 85036 23020 85076
rect 23118 85036 24268 85076
rect 24366 85036 25516 85076
rect 25614 85036 26764 85076
rect 26862 85036 28012 85076
rect 28110 85036 29260 85076
rect 29358 85036 30508 85076
rect 30606 85036 31756 85076
rect 31854 85036 33004 85076
rect 33102 85036 34252 85076
rect 34350 85036 35500 85076
rect 35598 85036 36748 85076
rect 36846 85036 37996 85076
rect 38094 85036 39244 85076
rect 39342 85036 40492 85076
rect 40590 85036 41740 85076
rect 41838 85036 42988 85076
rect 43086 85036 44236 85076
rect 44334 85036 45484 85076
rect 45582 85036 46732 85076
rect 46830 85036 47980 85076
rect 48078 85036 49228 85076
rect 49326 85036 50476 85076
rect 50574 85036 51724 85076
rect 51822 85036 52972 85076
rect 53070 85036 54220 85076
rect 54318 85036 55468 85076
rect 55566 85036 56716 85076
rect 56814 85054 75284 85076
rect 56814 85036 70977 85054
rect 4080 85000 70977 85036
rect 71075 85000 75284 85054
rect 0 84864 70660 84940
rect 71400 84864 75284 84940
rect 0 84728 75284 84804
rect 0 84592 75284 84668
rect 26 84429 86 84489
rect 5440 84456 62908 84532
rect 63920 84456 75284 84532
rect 5440 84360 58692 84396
rect 5440 84320 18110 84360
rect 18208 84320 19358 84360
rect 19456 84320 20606 84360
rect 20704 84320 21854 84360
rect 21952 84320 23102 84360
rect 23200 84320 24350 84360
rect 24448 84320 25598 84360
rect 25696 84320 26846 84360
rect 26944 84320 28094 84360
rect 28192 84320 29342 84360
rect 29440 84320 30590 84360
rect 30688 84320 31838 84360
rect 31936 84320 33086 84360
rect 33184 84320 34334 84360
rect 34432 84320 35582 84360
rect 35680 84320 36830 84360
rect 36928 84320 38078 84360
rect 38176 84320 39326 84360
rect 39424 84320 40574 84360
rect 40672 84320 41822 84360
rect 41920 84320 43070 84360
rect 43168 84320 44318 84360
rect 44416 84320 45566 84360
rect 45664 84320 46814 84360
rect 46912 84320 48062 84360
rect 48160 84320 49310 84360
rect 49408 84320 50558 84360
rect 50656 84320 51806 84360
rect 51904 84320 53054 84360
rect 53152 84320 54302 84360
rect 54400 84320 55550 84360
rect 55648 84320 56798 84360
rect 56896 84320 58692 84360
rect 71264 84320 75284 84396
rect 0 84184 17484 84260
rect 71264 84184 75284 84260
rect 0 84048 17484 84124
rect 59568 84048 75284 84124
rect 0 83912 75284 83988
rect 0 83776 18028 83852
rect 57392 83776 63724 83852
rect 64328 83776 75284 83852
rect 0 83658 17484 83716
rect 0 83640 3861 83658
rect 0 83504 3612 83580
rect 3959 83640 17484 83658
rect 57800 83640 70660 83716
rect 71400 83640 75284 83716
rect 4080 83504 17484 83580
rect 63512 83542 70977 83580
rect 71075 83542 75284 83580
rect 63512 83504 75284 83542
rect 0 83368 17484 83444
rect 63648 83368 75284 83444
rect 0 83232 17484 83308
rect 63648 83232 75284 83308
rect 0 83096 63044 83172
rect 63920 83096 75284 83172
rect 0 82960 58828 83036
rect 71264 82960 75284 83036
rect 5304 82824 58828 82900
rect 71264 82824 75284 82900
rect 26 82729 86 82789
rect 5304 82688 75284 82764
rect 0 82552 18028 82628
rect 0 82489 18283 82492
rect 18381 82489 19531 82492
rect 19629 82489 20779 82492
rect 20877 82489 22027 82492
rect 22125 82489 23275 82492
rect 23373 82489 24523 82492
rect 24621 82489 25771 82492
rect 25869 82489 27019 82492
rect 27117 82489 28267 82492
rect 28365 82489 29515 82492
rect 29613 82489 30763 82492
rect 30861 82489 32011 82492
rect 32109 82489 33259 82492
rect 33357 82489 34507 82492
rect 34605 82489 35755 82492
rect 35853 82489 37003 82492
rect 37101 82489 38251 82492
rect 38349 82489 39499 82492
rect 39597 82489 40747 82492
rect 40845 82489 41995 82492
rect 42093 82489 43243 82492
rect 43341 82489 44491 82492
rect 44589 82489 45739 82492
rect 45837 82489 46987 82492
rect 47085 82489 48235 82492
rect 48333 82489 49483 82492
rect 49581 82489 50731 82492
rect 50829 82489 51979 82492
rect 52077 82489 53227 82492
rect 53325 82489 54475 82492
rect 54573 82489 55723 82492
rect 55821 82489 56971 82492
rect 57392 82552 75284 82628
rect 57069 82489 75284 82492
rect 0 82420 75284 82489
rect 0 82416 64029 82420
rect 0 82280 3612 82356
rect 4080 82280 63724 82356
rect 64127 82416 75284 82420
rect 64328 82280 75284 82356
rect 0 82146 3861 82220
rect 3959 82146 70660 82220
rect 0 82144 70660 82146
rect 71400 82144 75284 82220
rect 0 82008 75284 82084
rect 0 81872 75284 81948
rect 0 81736 57468 81812
rect 26 81601 86 81661
rect 5168 81600 17484 81676
rect 0 81464 3204 81540
rect 5168 81464 17484 81540
rect 71264 81464 75284 81540
rect 0 81328 58964 81404
rect 71264 81328 75284 81404
rect 0 81192 75284 81268
rect 0 81056 17620 81132
rect 58208 81056 75284 81132
rect 0 80920 17852 80996
rect 17950 80920 18714 80996
rect 18812 80920 19100 80996
rect 19198 80920 19962 80996
rect 20060 80920 20348 80996
rect 20446 80920 21210 80996
rect 21308 80920 21596 80996
rect 21694 80920 22458 80996
rect 22556 80920 22844 80996
rect 22942 80920 23706 80996
rect 23804 80920 24092 80996
rect 24190 80920 24954 80996
rect 25052 80920 25340 80996
rect 25438 80920 26202 80996
rect 26300 80920 26588 80996
rect 26686 80920 27450 80996
rect 27548 80920 27836 80996
rect 27934 80920 28698 80996
rect 28796 80920 29084 80996
rect 29182 80920 29946 80996
rect 30044 80920 30332 80996
rect 30430 80920 31194 80996
rect 31292 80920 31580 80996
rect 31678 80920 32442 80996
rect 32540 80920 32828 80996
rect 32926 80920 33690 80996
rect 33788 80920 34076 80996
rect 34174 80920 34938 80996
rect 35036 80920 35324 80996
rect 35422 80920 36186 80996
rect 36284 80920 36572 80996
rect 36670 80920 37434 80996
rect 37532 80920 37820 80996
rect 37918 80920 38682 80996
rect 38780 80920 39068 80996
rect 39166 80920 39930 80996
rect 40028 80920 40316 80996
rect 40414 80920 41178 80996
rect 41276 80920 41564 80996
rect 41662 80920 42426 80996
rect 42524 80920 42812 80996
rect 42910 80920 43674 80996
rect 43772 80920 44060 80996
rect 44158 80920 44922 80996
rect 45020 80920 45308 80996
rect 45406 80920 46170 80996
rect 46268 80920 46556 80996
rect 46654 80920 47418 80996
rect 47516 80920 47804 80996
rect 47902 80920 48666 80996
rect 48764 80920 49052 80996
rect 49150 80920 49914 80996
rect 50012 80920 50300 80996
rect 50398 80920 51162 80996
rect 51260 80920 51548 80996
rect 51646 80920 52410 80996
rect 52508 80920 52796 80996
rect 52894 80920 53658 80996
rect 53756 80920 54044 80996
rect 54142 80920 54906 80996
rect 55004 80920 55292 80996
rect 55390 80920 56154 80996
rect 56252 80920 56540 80996
rect 56638 80920 57402 80996
rect 57500 80920 57788 80996
rect 57886 80920 75284 80996
rect 0 80784 3612 80860
rect 4080 80784 17620 80860
rect 58208 80812 75284 80860
rect 58208 80784 70977 80812
rect 0 80648 70660 80724
rect 71075 80784 75284 80812
rect 71400 80648 73788 80724
rect 0 80554 74063 80588
rect 74161 80554 74799 80588
rect 74897 80554 75284 80588
rect 0 80512 75284 80554
rect 0 80423 73244 80452
rect 0 80376 17347 80423
rect 17445 80376 17971 80423
rect 18069 80376 18595 80423
rect 18693 80376 19219 80423
rect 19317 80376 19843 80423
rect 19941 80376 20467 80423
rect 20565 80376 21091 80423
rect 21189 80376 21715 80423
rect 21813 80376 22339 80423
rect 22437 80376 22963 80423
rect 23061 80376 23587 80423
rect 23685 80376 24211 80423
rect 24309 80376 24835 80423
rect 24933 80376 25459 80423
rect 25557 80376 26083 80423
rect 26181 80376 26707 80423
rect 26805 80376 27331 80423
rect 27429 80376 27955 80423
rect 28053 80376 28579 80423
rect 28677 80376 29203 80423
rect 29301 80376 29827 80423
rect 29925 80376 30451 80423
rect 30549 80376 31075 80423
rect 31173 80376 31699 80423
rect 31797 80376 32323 80423
rect 32421 80376 32947 80423
rect 33045 80376 33571 80423
rect 33669 80376 34195 80423
rect 34293 80376 34819 80423
rect 34917 80376 35443 80423
rect 35541 80376 36067 80423
rect 36165 80376 36691 80423
rect 36789 80376 37315 80423
rect 37413 80376 37939 80423
rect 38037 80376 38563 80423
rect 38661 80376 39187 80423
rect 39285 80376 39811 80423
rect 39909 80376 40435 80423
rect 40533 80376 41059 80423
rect 41157 80376 41683 80423
rect 41781 80376 42307 80423
rect 42405 80376 42931 80423
rect 43029 80376 43555 80423
rect 43653 80376 44179 80423
rect 44277 80376 44803 80423
rect 44901 80376 45427 80423
rect 45525 80376 46051 80423
rect 46149 80376 46675 80423
rect 46773 80376 47299 80423
rect 47397 80376 47923 80423
rect 48021 80376 48547 80423
rect 48645 80376 49171 80423
rect 49269 80376 49795 80423
rect 49893 80376 50419 80423
rect 50517 80376 51043 80423
rect 51141 80376 51667 80423
rect 51765 80376 52291 80423
rect 52389 80376 52915 80423
rect 53013 80376 53539 80423
rect 53637 80376 54163 80423
rect 54261 80376 54787 80423
rect 54885 80376 55411 80423
rect 55509 80376 56035 80423
rect 56133 80376 56659 80423
rect 56757 80376 57283 80423
rect 57381 80376 57907 80423
rect 58005 80376 73244 80423
rect 0 80240 17076 80316
rect 58208 80240 73244 80316
rect 0 80104 16396 80180
rect 17000 80104 58284 80180
rect 59024 80104 73380 80180
rect 5168 80001 16651 80044
rect 16749 80001 58603 80044
rect 58701 80001 73380 80044
rect 5168 79968 73380 80001
rect 26 79901 86 79961
rect 3672 79832 16396 79908
rect 0 79764 16651 79772
rect 17000 79832 58284 79908
rect 16749 79764 58603 79772
rect 59024 79832 75284 79908
rect 58701 79764 75284 79772
rect 0 79696 75284 79764
rect 0 79560 10140 79636
rect 10744 79560 16396 79636
rect 17000 79560 58284 79636
rect 59024 79560 64540 79636
rect 65144 79560 75284 79636
rect 0 79424 10438 79500
rect 10536 79424 10548 79500
rect 0 79288 3612 79364
rect 12376 79424 63044 79500
rect 64736 79424 64816 79500
rect 64914 79424 73788 79500
rect 4080 79288 10140 79364
rect 12104 79288 16396 79364
rect 0 79152 11636 79228
rect 12376 79211 16651 79228
rect 17000 79288 58284 79364
rect 16749 79211 58603 79228
rect 59024 79288 63316 79364
rect 65144 79288 75284 79364
rect 58701 79211 63044 79228
rect 12376 79152 63044 79211
rect 63648 79152 75284 79228
rect 0 79016 10140 79092
rect 12104 79016 16396 79092
rect 17000 79016 58284 79092
rect 59024 79016 63305 79092
rect 65144 79016 75284 79092
rect 3672 78880 10548 78956
rect 12376 78880 63044 78956
rect 64736 78880 73380 78956
rect 26 78773 86 78833
rect 5032 78744 10140 78820
rect 12104 78744 16396 78820
rect 17000 78744 58284 78820
rect 59024 78744 63316 78820
rect 65144 78744 73380 78820
rect 0 78608 4156 78684
rect 5032 78631 10438 78684
rect 10536 78631 10548 78684
rect 5032 78608 10548 78631
rect 12240 78608 63044 78684
rect 64736 78631 64816 78684
rect 64914 78631 75284 78684
rect 64736 78608 75284 78631
rect 0 78472 11364 78548
rect 12104 78472 16396 78548
rect 17000 78472 58284 78548
rect 59024 78472 63316 78548
rect 63920 78472 73788 78548
rect 0 78355 10548 78412
rect 0 78336 10438 78355
rect 0 78200 10140 78276
rect 10536 78336 10548 78355
rect 12376 78336 63044 78412
rect 64736 78355 74063 78412
rect 64736 78336 64816 78355
rect 12104 78200 16396 78276
rect 17000 78200 58284 78276
rect 59024 78213 63305 78276
rect 59024 78200 63316 78213
rect 64914 78336 74063 78355
rect 74161 78336 74799 78412
rect 74897 78336 75284 78412
rect 65144 78200 73788 78276
rect 0 78064 10548 78140
rect 11696 78064 63724 78140
rect 64736 78064 75284 78140
rect 0 78002 10140 78004
rect 0 77928 3861 78002
rect 3959 77928 10140 78002
rect 0 77792 3612 77868
rect 4080 77841 10438 77868
rect 10536 77841 10548 77868
rect 12104 77928 16396 78004
rect 17000 77928 58284 78004
rect 59024 77928 63316 78004
rect 4080 77792 10548 77841
rect 12376 77792 63044 77868
rect 64736 77841 64816 77868
rect 65144 77928 73380 78004
rect 64914 77841 73380 77868
rect 64736 77792 73380 77841
rect 0 77656 16396 77732
rect 17000 77656 58284 77732
rect 59024 77656 75284 77732
rect 0 77565 10548 77596
rect 0 77520 10438 77565
rect 10536 77520 10548 77565
rect 0 77384 10140 77460
rect 12376 77520 63044 77596
rect 64736 77565 75284 77596
rect 12104 77384 16396 77460
rect 17000 77384 58284 77460
rect 59024 77423 63305 77460
rect 64736 77520 64816 77565
rect 59024 77384 63316 77423
rect 64914 77520 75284 77565
rect 65144 77384 75284 77460
rect 0 77248 4156 77324
rect 5032 77255 73788 77324
rect 5032 77248 16651 77255
rect 26 77073 86 77133
rect 5032 77112 10140 77188
rect 3672 77051 10438 77052
rect 10536 77051 10548 77052
rect 3672 76976 10548 77051
rect 12104 77112 16396 77188
rect 16749 77248 58603 77255
rect 17000 77112 58284 77188
rect 58701 77248 73788 77255
rect 59024 77126 63316 77188
rect 59024 77112 63305 77126
rect 12376 76976 63044 77052
rect 64736 77051 64816 77052
rect 65144 77112 75284 77188
rect 64914 77051 75284 77052
rect 64736 76976 75284 77051
rect 0 76840 3068 76916
rect 4896 76840 16396 76916
rect 17000 76840 58284 76916
rect 59024 76840 75284 76916
rect 0 76704 3068 76780
rect 4896 76775 10548 76780
rect 4896 76704 10438 76775
rect 10536 76704 10548 76775
rect 0 76568 3612 76644
rect 0 76490 3861 76508
rect 4080 76568 10140 76644
rect 12376 76704 63044 76780
rect 64736 76775 73380 76780
rect 12104 76568 16396 76644
rect 17000 76568 58284 76644
rect 59024 76633 63305 76644
rect 59024 76568 63316 76633
rect 64736 76704 64816 76775
rect 64914 76704 73380 76775
rect 65144 76568 73380 76644
rect 3959 76490 75284 76508
rect 0 76465 75284 76490
rect 0 76432 16651 76465
rect 0 76296 10140 76372
rect 12104 76296 16396 76372
rect 16749 76432 58603 76465
rect 17000 76296 58284 76372
rect 58701 76432 75284 76465
rect 59024 76336 63316 76372
rect 59024 76296 63305 76336
rect 65144 76296 75284 76372
rect 0 76160 10548 76236
rect 12376 76160 63044 76236
rect 64736 76172 75284 76236
rect 64736 76160 74063 76172
rect 0 76024 10140 76100
rect 10744 76024 16396 76100
rect 17000 76024 58284 76100
rect 59024 76024 64540 76100
rect 65144 76024 73788 76100
rect 74161 76160 74799 76172
rect 74897 76160 75284 76172
rect 0 75888 10438 75964
rect 10536 75888 10548 75964
rect 12376 75912 63044 75964
rect 12376 75888 16651 75912
rect 0 75752 10140 75828
rect 12104 75752 16396 75828
rect 16749 75888 58603 75912
rect 17000 75752 58284 75828
rect 58701 75888 63044 75912
rect 64736 75888 64816 75964
rect 64914 75888 75284 75964
rect 59024 75752 63316 75828
rect 65144 75752 75284 75828
rect 0 75616 10548 75692
rect 11696 75675 63724 75692
rect 11696 75616 16651 75675
rect 16749 75616 58603 75675
rect 58701 75616 63724 75675
rect 64736 75616 73380 75692
rect 0 75480 10140 75556
rect 12104 75480 16396 75556
rect 17000 75480 58284 75556
rect 59024 75546 63316 75556
rect 59024 75480 63305 75546
rect 65144 75480 73380 75556
rect 0 75344 10548 75420
rect 12376 75359 63044 75420
rect 12376 75344 16651 75359
rect 0 75208 10140 75284
rect 12104 75208 16396 75284
rect 16749 75344 58603 75359
rect 17000 75208 58284 75284
rect 58701 75344 63044 75359
rect 64736 75344 75284 75420
rect 59024 75208 63316 75284
rect 65144 75208 75284 75284
rect 0 75097 10438 75148
rect 10536 75097 10548 75148
rect 0 75072 10548 75097
rect 12376 75122 63044 75148
rect 12376 75072 16651 75122
rect 16749 75072 58603 75122
rect 58701 75072 63044 75122
rect 64736 75097 64816 75148
rect 64914 75097 73788 75148
rect 64736 75072 73788 75097
rect 0 74936 11364 75012
rect 12104 74936 16396 75012
rect 17000 74936 58284 75012
rect 59024 74936 63316 75012
rect 63920 74954 74063 75012
rect 74161 74954 74799 75012
rect 74897 74954 75284 75012
rect 63920 74936 75284 74954
rect 0 74800 10548 74876
rect 12376 74800 16651 74876
rect 16749 74800 58603 74876
rect 58701 74800 63044 74876
rect 64736 74800 75284 74876
rect 0 74664 10140 74740
rect 12104 74664 16396 74740
rect 17000 74664 58284 74740
rect 59024 74664 63305 74740
rect 65144 74664 75284 74740
rect 0 74528 11636 74604
rect 12376 74569 63044 74604
rect 12376 74528 16651 74569
rect 16749 74528 58603 74569
rect 58701 74528 63044 74569
rect 63648 74528 75284 74604
rect 0 74392 10140 74468
rect 0 74307 10438 74332
rect 12104 74392 16396 74468
rect 17000 74392 58284 74468
rect 59024 74392 63316 74468
rect 10536 74307 10548 74332
rect 0 74256 10548 74307
rect 12376 74256 16651 74332
rect 16749 74256 58603 74332
rect 58701 74256 63044 74332
rect 64736 74307 64816 74332
rect 65144 74392 73380 74468
rect 64914 74307 73380 74332
rect 64736 74256 73380 74307
rect 0 74120 16396 74196
rect 17000 74120 58284 74196
rect 59024 74120 75284 74196
rect 0 73989 10548 74060
rect 12376 73997 16651 74060
rect 16749 73997 58603 74060
rect 58701 73997 63044 74060
rect 0 73984 10438 73989
rect 0 73848 10140 73924
rect 10536 73984 10548 73989
rect 12376 73984 63044 73997
rect 64736 73989 75284 74060
rect 12104 73868 63305 73924
rect 64736 73984 64816 73989
rect 64914 73984 75284 73989
rect 12104 73848 63316 73868
rect 65144 73848 73788 73924
rect 0 73779 75284 73788
rect 0 73712 16651 73779
rect 16749 73712 58603 73779
rect 58701 73712 75284 73779
rect 0 73576 10140 73652
rect 12104 73576 16396 73652
rect 17000 73576 58284 73652
rect 59024 73576 63316 73652
rect 0 73440 10548 73516
rect 12376 73444 16651 73516
rect 16749 73444 58603 73516
rect 58701 73444 63044 73516
rect 65144 73576 75284 73652
rect 12376 73440 63044 73444
rect 64736 73440 73380 73516
rect 0 73304 16396 73380
rect 0 73199 10548 73244
rect 12376 73207 16651 73244
rect 17000 73304 58284 73380
rect 16749 73207 58603 73244
rect 59024 73304 73380 73380
rect 58701 73207 63044 73244
rect 0 73168 10438 73199
rect 0 73032 10140 73108
rect 10536 73168 10548 73199
rect 12376 73168 63044 73207
rect 64736 73199 75284 73244
rect 12104 73032 16396 73108
rect 17000 73032 58284 73108
rect 59024 73078 63305 73108
rect 64736 73168 64816 73199
rect 64914 73168 75284 73199
rect 59024 73032 63316 73078
rect 65144 73032 75284 73108
rect 0 72896 16651 72972
rect 16749 72896 58603 72972
rect 58701 72896 75284 72972
rect 0 72760 10140 72836
rect 0 72624 10548 72700
rect 12104 72760 16396 72836
rect 17000 72760 58284 72836
rect 59024 72781 63316 72836
rect 59024 72760 63305 72781
rect 12376 72654 16651 72700
rect 16749 72654 58603 72700
rect 58701 72654 63044 72700
rect 65144 72812 75284 72836
rect 65144 72760 74063 72812
rect 74161 72760 74799 72812
rect 74897 72760 75284 72812
rect 12376 72624 63044 72654
rect 64736 72624 73788 72700
rect 0 72488 16396 72564
rect 0 72409 10548 72428
rect 12376 72417 16651 72428
rect 17000 72488 58284 72564
rect 16749 72417 58603 72428
rect 59024 72488 75284 72564
rect 58701 72417 63044 72428
rect 0 72352 10438 72409
rect 10536 72352 10548 72409
rect 0 72216 10140 72292
rect 12376 72352 63044 72417
rect 64736 72409 75284 72428
rect 12104 72216 16396 72292
rect 17000 72216 58284 72292
rect 59024 72288 63305 72292
rect 64736 72352 64816 72409
rect 64914 72352 75284 72409
rect 59024 72216 63316 72288
rect 65144 72216 73380 72292
rect 0 72101 16651 72156
rect 16749 72101 58603 72156
rect 58701 72101 73380 72156
rect 0 72080 73380 72101
rect 0 71944 10140 72020
rect 0 71808 10548 71884
rect 12104 71944 16396 72020
rect 12376 71864 16651 71884
rect 17000 71944 58284 72020
rect 59024 71991 63316 72020
rect 16749 71864 58603 71884
rect 59024 71944 63305 71991
rect 58701 71864 63044 71884
rect 65144 71944 75284 72020
rect 12376 71808 63044 71864
rect 64736 71808 75284 71884
rect 0 71672 10140 71748
rect 10744 71672 16396 71748
rect 17000 71672 58284 71748
rect 59024 71672 64540 71748
rect 65144 71672 73788 71748
rect 0 71536 10438 71612
rect 10536 71536 10548 71612
rect 12376 71536 63044 71612
rect 64736 71536 64816 71612
rect 64914 71594 74063 71612
rect 74161 71594 74799 71612
rect 74897 71594 75284 71612
rect 64914 71536 75284 71594
rect 0 71400 10140 71476
rect 12104 71400 16396 71476
rect 0 71311 16651 71340
rect 17000 71400 58284 71476
rect 16749 71311 58603 71340
rect 59024 71400 63316 71476
rect 65144 71400 75284 71476
rect 58701 71311 75284 71340
rect 0 71264 75284 71311
rect 0 71128 10140 71204
rect 12104 71128 16396 71204
rect 17000 71128 58284 71204
rect 59024 71201 63316 71204
rect 59024 71128 63305 71201
rect 65144 71128 73380 71204
rect 0 70992 10548 71068
rect 12376 70992 63044 71068
rect 64736 70992 73380 71068
rect 0 70856 10140 70932
rect 12104 70856 16396 70932
rect 17000 70856 58284 70932
rect 59024 70856 63316 70932
rect 65144 70856 75284 70932
rect 0 70731 10438 70796
rect 10536 70731 10548 70796
rect 0 70720 10548 70731
rect 12376 70720 63044 70796
rect 64736 70731 64816 70796
rect 64914 70731 75284 70796
rect 64736 70720 75284 70731
rect 0 70584 11364 70660
rect 12104 70584 16396 70660
rect 0 70455 10548 70524
rect 0 70448 10438 70455
rect 0 70312 10140 70388
rect 10536 70448 10548 70455
rect 12376 70521 16651 70524
rect 17000 70584 58284 70660
rect 16749 70521 58603 70524
rect 59024 70584 63316 70660
rect 63920 70584 75284 70660
rect 58701 70521 63044 70524
rect 12376 70448 63044 70521
rect 64736 70455 73788 70524
rect 64736 70448 64816 70455
rect 12104 70312 16396 70388
rect 17000 70312 58284 70388
rect 59024 70313 63305 70388
rect 59024 70312 63316 70313
rect 64914 70448 73788 70455
rect 65144 70312 75284 70388
rect 0 70176 10548 70252
rect 11696 70176 63724 70252
rect 64736 70176 75284 70252
rect 0 70040 10140 70116
rect 12104 70040 16396 70116
rect 17000 70040 58284 70116
rect 59024 70040 63316 70116
rect 65144 70040 75284 70116
rect 0 69941 10438 69980
rect 10536 69941 10548 69980
rect 0 69904 10548 69941
rect 12376 69904 63044 69980
rect 64736 69941 64816 69980
rect 64914 69941 75284 69980
rect 64736 69904 75284 69941
rect 0 69768 16396 69844
rect 17000 69768 58284 69844
rect 59024 69768 75284 69844
rect 0 69665 10548 69708
rect 0 69632 10438 69665
rect 0 69496 10140 69572
rect 10536 69632 10548 69665
rect 12376 69632 63044 69708
rect 64736 69665 75284 69708
rect 64736 69632 64816 69665
rect 12104 69496 16396 69572
rect 17000 69496 58284 69572
rect 59024 69523 63305 69572
rect 59024 69496 63316 69523
rect 64914 69632 75284 69665
rect 65144 69496 75284 69572
rect 0 69360 75284 69436
rect 0 69224 10140 69300
rect 0 69151 10438 69164
rect 10536 69151 10548 69164
rect 0 69088 10548 69151
rect 12104 69224 16396 69300
rect 17000 69224 58284 69300
rect 59024 69226 63316 69300
rect 59024 69224 63305 69226
rect 12376 69088 63044 69164
rect 64736 69151 64816 69164
rect 65144 69224 75284 69300
rect 64914 69151 75284 69164
rect 64736 69088 75284 69151
rect 0 68952 16396 69028
rect 17000 68952 58284 69028
rect 59024 68952 75284 69028
rect 0 68875 10548 68892
rect 0 68816 10438 68875
rect 10536 68816 10548 68875
rect 0 68680 10140 68756
rect 12376 68816 63044 68892
rect 64736 68875 75284 68892
rect 12104 68680 16396 68756
rect 17000 68680 58284 68756
rect 59024 68733 63305 68756
rect 59024 68680 63316 68733
rect 64736 68816 64816 68875
rect 64914 68816 75284 68875
rect 65144 68680 75284 68756
rect 0 68565 75284 68620
rect 0 68544 16651 68565
rect 0 68408 10140 68484
rect 0 68272 10548 68348
rect 12104 68408 16396 68484
rect 16749 68544 58603 68565
rect 17000 68408 58284 68484
rect 58701 68544 75284 68565
rect 59024 68436 63316 68484
rect 59024 68408 63305 68436
rect 12376 68272 63044 68348
rect 65144 68408 75284 68484
rect 64736 68272 75284 68348
rect 0 68136 10140 68212
rect 10744 68136 16396 68212
rect 17000 68136 58284 68212
rect 59024 68136 64540 68212
rect 65144 68136 75284 68212
rect 0 68000 10438 68076
rect 10536 68000 10548 68076
rect 0 67864 10140 67940
rect 12376 68012 63044 68076
rect 12376 68000 16651 68012
rect 12104 67864 16396 67940
rect 16749 68000 58603 68012
rect 17000 67864 58284 67940
rect 58701 68000 63044 68012
rect 59024 67864 63316 67940
rect 64736 68000 64816 68076
rect 64914 68000 75284 68076
rect 65144 67864 75284 67940
rect 0 67728 10548 67804
rect 11696 67775 63724 67804
rect 11696 67728 16651 67775
rect 16749 67728 58603 67775
rect 58701 67728 63724 67775
rect 64736 67728 75284 67804
rect 0 67592 10140 67668
rect 12104 67592 16396 67668
rect 17000 67592 58284 67668
rect 59024 67646 63316 67668
rect 59024 67592 63305 67646
rect 65144 67592 75284 67668
rect 0 67456 10548 67532
rect 12376 67459 63044 67532
rect 12376 67456 16651 67459
rect 0 67320 10140 67396
rect 10744 67320 16396 67396
rect 16749 67456 58603 67459
rect 17000 67320 58284 67396
rect 58701 67456 63044 67459
rect 64736 67456 75284 67532
rect 59024 67320 64540 67396
rect 65144 67320 75284 67396
rect 0 67197 10438 67260
rect 10536 67197 10548 67260
rect 0 67184 10548 67197
rect 12376 67222 63044 67260
rect 12376 67184 16651 67222
rect 16749 67184 58603 67222
rect 58701 67184 63044 67222
rect 64736 67197 64816 67260
rect 64914 67197 75284 67260
rect 64736 67184 75284 67197
rect 0 67048 11364 67124
rect 12104 67048 16396 67124
rect 17000 67048 58284 67124
rect 59024 67048 63316 67124
rect 63920 67048 75284 67124
rect 0 66912 10548 66988
rect 12376 66985 63044 66988
rect 12376 66912 16651 66985
rect 16749 66912 58603 66985
rect 58701 66912 63044 66985
rect 64736 66912 75284 66988
rect 0 66776 10140 66852
rect 12104 66776 16396 66852
rect 17000 66776 58284 66852
rect 59024 66776 63305 66852
rect 65144 66776 75284 66852
rect 0 66640 11636 66716
rect 12376 66669 63044 66716
rect 12376 66640 16651 66669
rect 0 66504 10140 66580
rect 0 66407 10438 66444
rect 12104 66504 16396 66580
rect 16749 66640 58603 66669
rect 17000 66504 58284 66580
rect 58701 66640 63044 66669
rect 63648 66640 75284 66716
rect 59024 66504 63316 66580
rect 10536 66407 10548 66444
rect 0 66368 10548 66407
rect 12376 66432 63044 66444
rect 12376 66368 16651 66432
rect 16749 66368 58603 66432
rect 58701 66368 63044 66432
rect 64736 66407 64816 66444
rect 65144 66504 75284 66580
rect 64914 66407 75284 66444
rect 64736 66368 75284 66407
rect 0 66232 11364 66308
rect 12104 66232 16396 66308
rect 17000 66232 58284 66308
rect 59024 66232 63316 66308
rect 63920 66232 75284 66308
rect 0 66096 10548 66172
rect 12376 66097 16651 66172
rect 16749 66097 58603 66172
rect 58701 66097 63044 66172
rect 12376 66096 63044 66097
rect 64736 66096 75284 66172
rect 0 65960 10140 66036
rect 12104 65968 63305 66036
rect 12104 65960 63316 65968
rect 65144 65960 75284 66036
rect 0 65879 75284 65900
rect 0 65824 16651 65879
rect 16749 65824 58603 65879
rect 58701 65824 75284 65879
rect 0 65688 10140 65764
rect 0 65617 10438 65628
rect 12104 65688 16396 65764
rect 17000 65688 58284 65764
rect 59024 65688 63316 65764
rect 10536 65617 10548 65628
rect 0 65552 10548 65617
rect 12376 65552 16651 65628
rect 16749 65552 58603 65628
rect 58701 65552 63044 65628
rect 64736 65617 64816 65628
rect 65144 65688 75284 65764
rect 64914 65617 75284 65628
rect 64736 65552 75284 65617
rect 0 65416 16396 65492
rect 17000 65416 58284 65492
rect 59024 65416 75284 65492
rect 0 65299 10548 65356
rect 12376 65307 16651 65356
rect 16749 65307 58603 65356
rect 58701 65307 63044 65356
rect 0 65280 10438 65299
rect 0 65144 10140 65220
rect 10536 65280 10548 65299
rect 12376 65280 63044 65307
rect 64736 65299 75284 65356
rect 12104 65144 16396 65220
rect 17000 65144 58284 65220
rect 59024 65178 63305 65220
rect 64736 65280 64816 65299
rect 64914 65280 75284 65299
rect 59024 65144 63316 65178
rect 65144 65144 75284 65220
rect 0 65008 16651 65084
rect 16749 65008 58603 65084
rect 58701 65008 75284 65084
rect 0 64872 10140 64948
rect 0 64736 10548 64812
rect 12104 64872 16396 64948
rect 17000 64872 58284 64948
rect 59024 64881 63316 64948
rect 59024 64872 63305 64881
rect 12376 64754 16651 64812
rect 16749 64754 58603 64812
rect 58701 64754 63044 64812
rect 65144 64872 75284 64948
rect 12376 64736 63044 64754
rect 64736 64736 75284 64812
rect 0 64600 16396 64676
rect 0 64509 10548 64540
rect 12376 64517 16651 64540
rect 17000 64600 58284 64676
rect 16749 64517 58603 64540
rect 59024 64600 75284 64676
rect 58701 64517 63044 64540
rect 0 64464 10438 64509
rect 10536 64464 10548 64509
rect 0 64328 10140 64404
rect 12376 64464 63044 64517
rect 64736 64509 75284 64540
rect 12104 64328 16396 64404
rect 17000 64328 58284 64404
rect 59024 64388 63305 64404
rect 64736 64464 64816 64509
rect 64914 64464 75284 64509
rect 59024 64328 63316 64388
rect 65144 64328 75284 64404
rect 0 64201 16651 64268
rect 16749 64201 58603 64268
rect 58701 64201 75284 64268
rect 0 64192 75284 64201
rect 0 64056 10140 64132
rect 0 63920 10548 63996
rect 12104 64056 16396 64132
rect 12376 63964 16651 63996
rect 17000 64056 58284 64132
rect 59024 64091 63316 64132
rect 16749 63964 58603 63996
rect 59024 64056 63305 64091
rect 58701 63964 63044 63996
rect 65144 64056 75284 64132
rect 12376 63920 63044 63964
rect 64736 63920 75284 63996
rect 0 63784 16396 63860
rect 17000 63784 58284 63860
rect 59024 63784 75284 63860
rect 0 63719 10548 63724
rect 0 63648 10438 63719
rect 10536 63648 10548 63719
rect 12376 63648 63044 63724
rect 64736 63719 75284 63724
rect 64736 63648 64816 63719
rect 64914 63648 75284 63719
rect 0 63512 10140 63588
rect 12104 63512 16396 63588
rect 17000 63512 58284 63588
rect 59024 63512 63316 63588
rect 65144 63512 75284 63588
rect 0 63411 16651 63452
rect 16749 63411 58603 63452
rect 58701 63411 75284 63452
rect 0 63376 75284 63411
rect 0 63240 10140 63316
rect 12104 63240 16396 63316
rect 0 63104 10548 63180
rect 12376 63174 16651 63180
rect 17000 63240 58284 63316
rect 59024 63301 63316 63316
rect 16749 63174 58603 63180
rect 59024 63240 63305 63301
rect 65144 63240 75284 63316
rect 58701 63174 63044 63180
rect 12376 63104 63044 63174
rect 64736 63104 75284 63180
rect 0 62968 10140 63044
rect 10744 62968 16396 63044
rect 17000 62968 58284 63044
rect 59024 62968 64540 63044
rect 65144 62968 75284 63044
rect 0 62832 10438 62908
rect 10536 62832 10548 62908
rect 12376 62832 63044 62908
rect 64736 62832 64816 62908
rect 64914 62832 75284 62908
rect 0 62696 10140 62772
rect 12104 62696 16396 62772
rect 0 62560 11636 62636
rect 12376 62621 16651 62636
rect 17000 62696 58284 62772
rect 16749 62621 58603 62636
rect 59024 62696 63316 62772
rect 65144 62696 75284 62772
rect 58701 62621 63044 62636
rect 12376 62560 63044 62621
rect 63648 62560 75284 62636
rect 0 62424 10140 62500
rect 12104 62424 16396 62500
rect 17000 62424 58284 62500
rect 59024 62424 63305 62500
rect 65144 62424 75284 62500
rect 0 62288 10548 62364
rect 12376 62288 63044 62364
rect 64736 62288 75284 62364
rect 0 62152 10140 62228
rect 12104 62152 16396 62228
rect 17000 62152 58284 62228
rect 59024 62152 63316 62228
rect 65144 62152 75284 62228
rect 0 62041 10438 62092
rect 10536 62041 10548 62092
rect 0 62016 10548 62041
rect 12376 62016 63044 62092
rect 64736 62041 64816 62092
rect 64914 62041 75284 62092
rect 64736 62016 75284 62041
rect 0 61880 16396 61956
rect 17000 61880 58284 61956
rect 59024 61880 75284 61956
rect 0 61765 10548 61820
rect 0 61744 10438 61765
rect 0 61608 10140 61684
rect 10536 61744 10548 61765
rect 12376 61744 63044 61820
rect 64736 61765 75284 61820
rect 64736 61744 64816 61765
rect 12104 61608 16396 61684
rect 17000 61608 58284 61684
rect 59024 61623 63305 61684
rect 59024 61608 63316 61623
rect 64914 61744 75284 61765
rect 65144 61608 75284 61684
rect 0 61472 75284 61548
rect 0 61336 10140 61412
rect 0 61251 10438 61276
rect 10536 61251 10548 61276
rect 12104 61336 16396 61412
rect 17000 61336 58284 61412
rect 59024 61336 63316 61412
rect 0 61200 10548 61251
rect 12376 61200 63044 61276
rect 64736 61251 64816 61276
rect 65144 61336 75284 61412
rect 64914 61251 75284 61276
rect 64736 61200 75284 61251
rect 0 61064 16396 61140
rect 17000 61064 58284 61140
rect 59024 61064 75284 61140
rect 0 60975 10548 61004
rect 0 60928 10438 60975
rect 10536 60928 10548 60975
rect 0 60792 10140 60868
rect 12376 60928 63044 61004
rect 64736 60975 75284 61004
rect 12104 60792 16396 60868
rect 17000 60792 58284 60868
rect 59024 60833 63305 60868
rect 64736 60928 64816 60975
rect 59024 60792 63316 60833
rect 64914 60928 75284 60975
rect 65144 60792 75284 60868
rect 0 60665 75284 60732
rect 0 60656 16651 60665
rect 0 60520 10140 60596
rect 0 60384 10548 60460
rect 12104 60520 16396 60596
rect 16749 60656 58603 60665
rect 17000 60520 58284 60596
rect 58701 60656 75284 60665
rect 59024 60536 63316 60596
rect 59024 60520 63305 60536
rect 12376 60384 63044 60460
rect 65144 60520 75284 60596
rect 64736 60384 75284 60460
rect 0 60248 16396 60324
rect 17000 60248 58284 60324
rect 59024 60248 75284 60324
rect 0 60185 10548 60188
rect 0 60112 10438 60185
rect 10536 60112 10548 60185
rect 0 59976 10140 60052
rect 12376 60112 63044 60188
rect 64736 60185 75284 60188
rect 12104 59976 16396 60052
rect 17000 59976 58284 60052
rect 59024 60043 63305 60052
rect 59024 59976 63316 60043
rect 64736 60112 64816 60185
rect 64914 60112 75284 60185
rect 65144 59976 75284 60052
rect 0 59875 75284 59916
rect 0 59840 16651 59875
rect 0 59704 10140 59780
rect 12104 59704 16396 59780
rect 16749 59840 58603 59875
rect 17000 59704 58284 59780
rect 58701 59840 75284 59875
rect 59024 59746 63316 59780
rect 59024 59704 63305 59746
rect 65144 59704 75284 59780
rect 0 59568 10548 59644
rect 12376 59568 63044 59644
rect 64736 59568 75284 59644
rect 0 59432 10140 59508
rect 10744 59432 16396 59508
rect 17000 59432 58284 59508
rect 59024 59432 64540 59508
rect 65144 59432 75284 59508
rect 0 59297 10438 59372
rect 10536 59297 10548 59372
rect 0 59296 10548 59297
rect 12376 59322 63044 59372
rect 12376 59296 16651 59322
rect 0 59160 11364 59236
rect 12104 59160 16396 59236
rect 16749 59296 58603 59322
rect 17000 59160 58284 59236
rect 58701 59296 63044 59322
rect 64736 59297 64816 59372
rect 64914 59297 75284 59372
rect 64736 59296 75284 59297
rect 59024 59160 63316 59236
rect 63920 59160 75284 59236
rect 0 59024 10548 59100
rect 11696 59085 63724 59100
rect 11696 59024 16651 59085
rect 16749 59024 58603 59085
rect 58701 59024 63724 59085
rect 64736 59024 75284 59100
rect 0 58888 10140 58964
rect 12104 58888 16396 58964
rect 17000 58888 58284 58964
rect 59024 58956 63316 58964
rect 59024 58888 63305 58956
rect 65144 58888 75284 58964
rect 0 58752 10548 58828
rect 12376 58769 63044 58828
rect 12376 58752 16651 58769
rect 0 58616 10140 58692
rect 12104 58616 16396 58692
rect 16749 58752 58603 58769
rect 17000 58616 58284 58692
rect 58701 58752 63044 58769
rect 64736 58752 75284 58828
rect 59024 58616 63316 58692
rect 65144 58616 75284 58692
rect 0 58507 10438 58556
rect 10536 58507 10548 58556
rect 0 58480 10548 58507
rect 12376 58532 63044 58556
rect 12376 58480 16651 58532
rect 16749 58480 58603 58532
rect 58701 58480 63044 58532
rect 64736 58507 64816 58556
rect 64914 58507 75284 58556
rect 64736 58480 75284 58507
rect 0 58344 11364 58420
rect 12104 58344 16396 58420
rect 17000 58344 58284 58420
rect 59024 58344 63316 58420
rect 63920 58344 75284 58420
rect 0 58208 10548 58284
rect 12376 58208 16651 58284
rect 16749 58208 58603 58284
rect 58701 58208 63044 58284
rect 64736 58208 75284 58284
rect 0 58072 10140 58148
rect 12104 58072 16396 58148
rect 17000 58072 58284 58148
rect 59024 58072 63305 58148
rect 65144 58072 75284 58148
rect 0 57936 11636 58012
rect 12376 57979 63044 58012
rect 12376 57936 16651 57979
rect 16749 57936 58603 57979
rect 58701 57936 63044 57979
rect 63648 57936 75284 58012
rect 0 57800 10140 57876
rect 0 57717 10438 57740
rect 12104 57800 16396 57876
rect 17000 57800 58284 57876
rect 59024 57800 63316 57876
rect 10536 57717 10548 57740
rect 0 57664 10548 57717
rect 12376 57664 16651 57740
rect 16749 57664 58603 57740
rect 58701 57664 63044 57740
rect 64736 57717 64816 57740
rect 65144 57800 75284 57876
rect 64914 57717 75284 57740
rect 64736 57664 75284 57717
rect 0 57528 16396 57604
rect 17000 57528 58284 57604
rect 59024 57528 75284 57604
rect 0 57399 10548 57468
rect 12376 57407 16651 57468
rect 16749 57407 58603 57468
rect 58701 57407 63044 57468
rect 0 57392 10438 57399
rect 0 57256 10140 57332
rect 10536 57392 10548 57399
rect 12376 57392 63044 57407
rect 64736 57399 75284 57468
rect 12104 57278 63305 57332
rect 64736 57392 64816 57399
rect 64914 57392 75284 57399
rect 12104 57256 63316 57278
rect 65144 57256 75284 57332
rect 0 57189 75284 57196
rect 0 57120 16651 57189
rect 16749 57120 58603 57189
rect 58701 57120 75284 57189
rect 0 56984 10140 57060
rect 12104 56984 16396 57060
rect 17000 56984 58284 57060
rect 59024 56984 63316 57060
rect 0 56848 10548 56924
rect 12376 56854 16651 56924
rect 16749 56854 58603 56924
rect 58701 56854 63044 56924
rect 65144 56984 75284 57060
rect 12376 56848 63044 56854
rect 64736 56848 75284 56924
rect 0 56712 16396 56788
rect 0 56609 10548 56652
rect 12376 56617 16651 56652
rect 17000 56712 58284 56788
rect 16749 56617 58603 56652
rect 59024 56712 75284 56788
rect 58701 56617 63044 56652
rect 0 56576 10438 56609
rect 0 56440 10140 56516
rect 10536 56576 10548 56609
rect 12376 56576 63044 56617
rect 64736 56609 75284 56652
rect 12104 56440 16396 56516
rect 17000 56440 58284 56516
rect 59024 56488 63305 56516
rect 64736 56576 64816 56609
rect 64914 56576 75284 56609
rect 59024 56440 63316 56488
rect 65144 56440 75284 56516
rect 0 56304 16651 56380
rect 16749 56304 58603 56380
rect 58701 56304 75284 56380
rect 0 56168 10140 56244
rect 0 56032 10548 56108
rect 12104 56168 16396 56244
rect 17000 56168 58284 56244
rect 59024 56191 63316 56244
rect 59024 56168 63305 56191
rect 12376 56064 16651 56108
rect 16749 56064 58603 56108
rect 58701 56064 63044 56108
rect 65144 56168 75284 56244
rect 12376 56032 63044 56064
rect 64736 56032 75284 56108
rect 0 55896 16396 55972
rect 0 55819 10548 55836
rect 12376 55827 16651 55836
rect 17000 55896 58284 55972
rect 16749 55827 58603 55836
rect 59024 55896 75284 55972
rect 58701 55827 63044 55836
rect 0 55760 10438 55819
rect 10536 55760 10548 55819
rect 0 55624 10140 55700
rect 12376 55760 63044 55827
rect 64736 55819 75284 55836
rect 12104 55624 16396 55700
rect 17000 55624 58284 55700
rect 59024 55698 63305 55700
rect 64736 55760 64816 55819
rect 64914 55760 75284 55819
rect 59024 55624 63316 55698
rect 65144 55624 75284 55700
rect 0 55511 16651 55564
rect 16749 55511 58603 55564
rect 58701 55511 75284 55564
rect 0 55488 75284 55511
rect 0 55352 10140 55428
rect 0 55216 10548 55292
rect 12104 55352 16396 55428
rect 12376 55274 16651 55292
rect 17000 55352 58284 55428
rect 59024 55401 63316 55428
rect 16749 55274 58603 55292
rect 59024 55352 63305 55401
rect 58701 55274 63044 55292
rect 65144 55352 75284 55428
rect 12376 55216 63044 55274
rect 64736 55216 75284 55292
rect 0 55080 10140 55156
rect 10744 55080 16396 55156
rect 17000 55080 58284 55156
rect 59024 55080 64540 55156
rect 65144 55080 75284 55156
rect 0 54944 10438 55020
rect 10536 54944 10548 55020
rect 12376 54944 63044 55020
rect 64736 54944 64816 55020
rect 64914 54944 75284 55020
rect 0 54808 10140 54884
rect 12104 54808 16396 54884
rect 0 54721 16651 54748
rect 17000 54808 58284 54884
rect 16749 54721 58603 54748
rect 59024 54808 63316 54884
rect 65144 54808 75284 54884
rect 58701 54721 75284 54748
rect 0 54672 75284 54721
rect 0 54536 10140 54612
rect 14280 54582 16396 54612
rect 0 54400 10548 54476
rect 14280 54536 15387 54582
rect 15485 54536 16396 54582
rect 17000 54536 58284 54612
rect 59024 54582 61140 54612
rect 59024 54536 59867 54582
rect 59965 54536 61140 54582
rect 13192 54400 15172 54476
rect 15776 54400 59644 54476
rect 60248 54400 62228 54476
rect 65144 54536 75284 54612
rect 64736 54400 75284 54476
rect 0 54264 10140 54340
rect 12104 54264 16396 54340
rect 17000 54264 58284 54340
rect 59024 54264 63316 54340
rect 65144 54264 75284 54340
rect 0 54141 10438 54204
rect 10536 54141 10548 54204
rect 0 54128 10548 54141
rect 12376 54128 63044 54204
rect 64736 54141 64816 54204
rect 64914 54141 75284 54204
rect 64736 54128 75284 54141
rect 0 53992 11364 54068
rect 12104 53992 16396 54068
rect 0 53865 10548 53932
rect 0 53856 10438 53865
rect 0 53720 10140 53796
rect 10536 53856 10548 53865
rect 12376 53931 16651 53932
rect 17000 53992 58284 54068
rect 16749 53931 58603 53932
rect 59024 53992 63316 54068
rect 63920 53992 75284 54068
rect 58701 53931 63044 53932
rect 12376 53856 63044 53931
rect 64736 53865 75284 53932
rect 64736 53856 64816 53865
rect 12104 53720 16396 53796
rect 17000 53720 58284 53796
rect 59024 53723 63305 53796
rect 59024 53720 63316 53723
rect 64914 53856 75284 53865
rect 65144 53720 75284 53796
rect 0 53584 10548 53660
rect 11696 53584 63724 53660
rect 64736 53584 75284 53660
rect 0 53448 10140 53524
rect 0 53351 10438 53388
rect 10536 53351 10548 53388
rect 12104 53448 16396 53524
rect 17000 53448 58284 53524
rect 59024 53448 63316 53524
rect 0 53312 10548 53351
rect 12376 53312 63044 53388
rect 64736 53351 64816 53388
rect 65144 53448 75284 53524
rect 64914 53351 75284 53388
rect 64736 53312 75284 53351
rect 0 53176 16396 53252
rect 17000 53176 58284 53252
rect 59024 53176 75284 53252
rect 0 53075 10548 53116
rect 0 53040 10438 53075
rect 0 52904 10140 52980
rect 10536 53040 10548 53075
rect 12376 53040 63044 53116
rect 64736 53075 75284 53116
rect 64736 53040 64816 53075
rect 12104 52904 16396 52980
rect 17000 52904 58420 52980
rect 58888 52933 63305 52980
rect 58888 52904 63316 52933
rect 64914 53040 75284 53075
rect 65144 52904 75284 52980
rect 0 52768 75284 52844
rect 0 52632 10140 52708
rect 0 52561 10438 52572
rect 10536 52561 10548 52572
rect 0 52496 10548 52561
rect 12104 52632 16396 52708
rect 17000 52632 58284 52708
rect 59024 52636 63316 52708
rect 59024 52632 63305 52636
rect 12376 52496 63044 52572
rect 64736 52561 64816 52572
rect 65144 52632 75284 52708
rect 64914 52561 75284 52572
rect 64736 52496 75284 52561
rect 0 52360 16396 52436
rect 17000 52360 58284 52436
rect 59024 52360 75284 52436
rect 0 52285 10548 52300
rect 0 52224 10438 52285
rect 10536 52224 10548 52285
rect 0 52088 10140 52164
rect 12376 52224 63044 52300
rect 64736 52285 75284 52300
rect 12104 52088 16396 52164
rect 17000 52088 58284 52164
rect 59024 52143 63305 52164
rect 59024 52088 63316 52143
rect 64736 52224 64816 52285
rect 64914 52224 75284 52285
rect 65144 52088 75284 52164
rect 0 51975 75284 52028
rect 0 51952 16651 51975
rect 0 51816 10140 51892
rect 0 51680 10548 51756
rect 12104 51816 16396 51892
rect 16749 51952 58603 51975
rect 17000 51816 58284 51892
rect 58701 51952 75284 51975
rect 59024 51846 63316 51892
rect 59024 51816 63305 51846
rect 12376 51680 63044 51756
rect 65144 51816 75284 51892
rect 64736 51680 75284 51756
rect 0 51544 10140 51620
rect 10744 51544 16396 51620
rect 17000 51544 58284 51620
rect 59024 51544 64540 51620
rect 65144 51544 75284 51620
rect 0 51408 10438 51484
rect 10536 51408 10548 51484
rect 0 51272 10140 51348
rect 12376 51422 63044 51484
rect 12376 51408 16651 51422
rect 12104 51272 16396 51348
rect 16749 51408 58603 51422
rect 17000 51272 58284 51348
rect 58701 51408 63044 51422
rect 59024 51272 63316 51348
rect 64736 51408 64816 51484
rect 64914 51408 75284 51484
rect 65144 51272 75284 51348
rect 0 51136 10548 51212
rect 11696 51185 63724 51212
rect 11696 51136 16651 51185
rect 16749 51136 58603 51185
rect 58701 51136 63724 51185
rect 64736 51136 75284 51212
rect 0 51000 10140 51076
rect 12104 51000 16396 51076
rect 17000 51000 58284 51076
rect 59024 51056 63316 51076
rect 59024 51000 63305 51056
rect 65144 51000 75284 51076
rect 0 50864 10548 50940
rect 12376 50869 63044 50940
rect 12376 50864 16651 50869
rect 0 50728 10140 50804
rect 10744 50728 16396 50804
rect 16749 50864 58603 50869
rect 17000 50728 58284 50804
rect 58701 50864 63044 50869
rect 64736 50864 75284 50940
rect 59024 50728 64540 50804
rect 65144 50728 75284 50804
rect 0 50607 10438 50668
rect 10536 50607 10548 50668
rect 0 50592 10548 50607
rect 12376 50632 63044 50668
rect 12376 50592 16651 50632
rect 16749 50592 58603 50632
rect 58701 50592 63044 50632
rect 64736 50607 64816 50668
rect 64914 50607 75284 50668
rect 64736 50592 75284 50607
rect 0 50456 11364 50532
rect 12104 50456 16396 50532
rect 17000 50456 58284 50532
rect 59024 50456 63316 50532
rect 63920 50456 75284 50532
rect 0 50320 10548 50396
rect 12376 50395 63044 50396
rect 12376 50320 16651 50395
rect 16749 50320 58603 50395
rect 58701 50320 63044 50395
rect 64736 50320 75284 50396
rect 0 50184 10140 50260
rect 12104 50184 16396 50260
rect 17000 50184 58284 50260
rect 59024 50184 63305 50260
rect 65144 50184 75284 50260
rect 0 50048 11636 50124
rect 12376 50079 63044 50124
rect 12376 50048 16651 50079
rect 0 49912 10140 49988
rect 0 49817 10438 49852
rect 12104 49912 16396 49988
rect 16749 50048 58603 50079
rect 17000 49912 58284 49988
rect 58701 50048 63044 50079
rect 63648 50048 75284 50124
rect 59024 49912 63316 49988
rect 10536 49817 10548 49852
rect 0 49776 10548 49817
rect 12376 49842 63044 49852
rect 12376 49776 16651 49842
rect 16749 49776 58603 49842
rect 58701 49776 63044 49842
rect 64736 49817 64816 49852
rect 65144 49912 75284 49988
rect 64914 49817 75284 49852
rect 64736 49776 75284 49817
rect 0 49640 11364 49716
rect 12104 49640 16396 49716
rect 17000 49640 58284 49716
rect 59024 49640 63316 49716
rect 63920 49640 75284 49716
rect 0 49504 10548 49580
rect 12376 49507 16651 49580
rect 16749 49507 58603 49580
rect 58701 49507 63044 49580
rect 12376 49504 63044 49507
rect 64736 49504 75284 49580
rect 0 49368 10140 49444
rect 12104 49378 63305 49444
rect 12104 49368 63316 49378
rect 65144 49368 75284 49444
rect 0 49289 75284 49308
rect 0 49232 16651 49289
rect 16749 49232 58603 49289
rect 58701 49232 75284 49289
rect 0 49096 10140 49172
rect 0 49027 10438 49036
rect 12104 49096 16396 49172
rect 17000 49096 58284 49172
rect 59024 49096 63316 49172
rect 10536 49027 10548 49036
rect 0 48960 10548 49027
rect 12376 48960 16651 49036
rect 16749 48960 58603 49036
rect 58701 48960 63044 49036
rect 64736 49027 64816 49036
rect 65144 49096 75284 49172
rect 64914 49027 75284 49036
rect 64736 48960 75284 49027
rect 0 48824 16396 48900
rect 17000 48824 58284 48900
rect 59024 48824 75284 48900
rect 0 48709 10548 48764
rect 12376 48717 16651 48764
rect 16749 48717 58603 48764
rect 58701 48717 63044 48764
rect 0 48688 10438 48709
rect 0 48552 10140 48628
rect 10536 48688 10548 48709
rect 12376 48688 63044 48717
rect 64736 48709 75284 48764
rect 12104 48552 16396 48628
rect 17000 48552 58284 48628
rect 59024 48588 63305 48628
rect 64736 48688 64816 48709
rect 64914 48688 75284 48709
rect 59024 48552 63316 48588
rect 65144 48552 75284 48628
rect 0 48416 16651 48492
rect 16749 48416 58603 48492
rect 58701 48416 75284 48492
rect 0 48280 10140 48356
rect 0 48144 10548 48220
rect 12104 48280 16396 48356
rect 17000 48280 58284 48356
rect 59024 48291 63316 48356
rect 59024 48280 63305 48291
rect 12376 48164 16651 48220
rect 16749 48164 58603 48220
rect 58701 48164 63044 48220
rect 65144 48280 75284 48356
rect 12376 48144 63044 48164
rect 64736 48144 75284 48220
rect 0 48008 16396 48084
rect 0 47919 10548 47948
rect 12376 47927 16651 47948
rect 17000 48008 58284 48084
rect 16749 47927 58603 47948
rect 59024 48008 75284 48084
rect 58701 47927 63044 47948
rect 0 47872 10438 47919
rect 10536 47872 10548 47919
rect 0 47736 10140 47812
rect 12376 47872 63044 47927
rect 64736 47919 75284 47948
rect 12104 47736 16396 47812
rect 17000 47736 58284 47812
rect 59024 47798 63305 47812
rect 64736 47872 64816 47919
rect 64914 47872 75284 47919
rect 59024 47736 63316 47798
rect 65144 47736 75284 47812
rect 0 47611 16651 47676
rect 16749 47611 58603 47676
rect 58701 47611 75284 47676
rect 0 47600 75284 47611
rect 0 47464 10140 47540
rect 0 47328 10548 47404
rect 12104 47464 16396 47540
rect 12376 47374 16651 47404
rect 17000 47464 58284 47540
rect 59024 47501 63316 47540
rect 16749 47374 58603 47404
rect 59024 47464 63305 47501
rect 58701 47374 63044 47404
rect 65144 47464 75284 47540
rect 12376 47328 63044 47374
rect 64736 47328 75284 47404
rect 0 47192 16396 47268
rect 17000 47192 58284 47268
rect 59024 47192 75284 47268
rect 0 47129 10548 47132
rect 0 47056 10438 47129
rect 10536 47056 10548 47129
rect 12376 47056 63044 47132
rect 64736 47129 75284 47132
rect 64736 47056 64816 47129
rect 64914 47056 75284 47129
rect 0 46920 10140 46996
rect 12104 46920 16396 46996
rect 17000 46920 58284 46996
rect 59024 46920 63316 46996
rect 65144 46920 75284 46996
rect 0 46821 16651 46860
rect 16749 46821 58603 46860
rect 58701 46821 75284 46860
rect 0 46784 75284 46821
rect 0 46648 10140 46724
rect 12104 46648 16396 46724
rect 0 46512 10548 46588
rect 12376 46584 16651 46588
rect 17000 46648 58284 46724
rect 59024 46711 63316 46724
rect 16749 46584 58603 46588
rect 59024 46648 63305 46711
rect 65144 46648 75284 46724
rect 58701 46584 63044 46588
rect 12376 46512 63044 46584
rect 64736 46512 75284 46588
rect 0 46376 10140 46452
rect 12104 46376 16396 46452
rect 17000 46376 58284 46452
rect 59024 46376 63316 46452
rect 65144 46376 75284 46452
rect 0 46241 10438 46316
rect 10536 46241 10548 46316
rect 0 46240 10548 46241
rect 12240 46240 63044 46316
rect 64736 46241 64816 46316
rect 64914 46241 75284 46316
rect 64736 46240 75284 46241
rect 0 46104 11364 46180
rect 12104 46104 16396 46180
rect 0 45968 11636 46044
rect 12376 46031 16651 46044
rect 17000 46104 58284 46180
rect 16749 46031 58603 46044
rect 59024 46104 63316 46180
rect 63920 46104 75284 46180
rect 58701 46031 63044 46044
rect 12376 45968 63044 46031
rect 63648 45968 75284 46044
rect 0 45832 10140 45908
rect 12104 45832 16396 45908
rect 17000 45832 58284 45908
rect 59024 45832 63305 45908
rect 65144 45832 75284 45908
rect 0 45696 10548 45772
rect 12376 45696 63044 45772
rect 64736 45696 75284 45772
rect 0 45560 10140 45636
rect 12104 45560 16396 45636
rect 17000 45560 58284 45636
rect 59024 45560 63316 45636
rect 65144 45560 75284 45636
rect 0 45451 10438 45500
rect 10536 45451 10548 45500
rect 0 45424 10548 45451
rect 12376 45424 63044 45500
rect 64736 45451 64816 45500
rect 64914 45451 75284 45500
rect 64736 45424 75284 45451
rect 0 45288 16396 45364
rect 17000 45288 58284 45364
rect 59024 45288 75284 45364
rect 0 45175 10548 45228
rect 0 45152 10438 45175
rect 0 45016 10140 45092
rect 10536 45152 10548 45175
rect 12376 45152 63044 45228
rect 64736 45175 75284 45228
rect 64736 45152 64816 45175
rect 12104 45016 16396 45092
rect 17000 45016 58284 45092
rect 59024 45033 63305 45092
rect 59024 45016 63316 45033
rect 64914 45152 75284 45175
rect 65144 45016 75284 45092
rect 0 44880 75284 44956
rect 0 44744 10140 44820
rect 0 44661 10438 44684
rect 10536 44661 10548 44684
rect 12104 44744 16396 44820
rect 17000 44744 58284 44820
rect 59024 44744 63316 44820
rect 0 44608 10548 44661
rect 12376 44608 63044 44684
rect 64736 44661 64816 44684
rect 65144 44744 75284 44820
rect 64914 44661 75284 44684
rect 64736 44608 75284 44661
rect 0 44472 16396 44548
rect 17000 44472 58284 44548
rect 59024 44472 75284 44548
rect 0 44385 10548 44412
rect 0 44336 10438 44385
rect 10536 44336 10548 44385
rect 0 44200 10140 44276
rect 12376 44336 63044 44412
rect 64736 44385 75284 44412
rect 12104 44200 16396 44276
rect 17000 44200 58284 44276
rect 59024 44243 63305 44276
rect 64736 44336 64816 44385
rect 59024 44200 63316 44243
rect 64914 44336 75284 44385
rect 65144 44200 75284 44276
rect 0 44075 75284 44140
rect 0 44064 16651 44075
rect 0 43928 10140 44004
rect 0 43792 10548 43868
rect 12104 43928 16396 44004
rect 16749 44064 58603 44075
rect 17000 43928 58284 44004
rect 58701 44064 75284 44075
rect 59024 43946 63316 44004
rect 59024 43928 63305 43946
rect 12376 43792 63044 43868
rect 65144 43928 75284 44004
rect 64736 43792 75284 43868
rect 0 43656 16396 43732
rect 17000 43656 58284 43732
rect 59024 43656 75284 43732
rect 0 43595 10548 43596
rect 0 43520 10438 43595
rect 10536 43520 10548 43595
rect 0 43384 10140 43460
rect 12376 43522 63044 43596
rect 64736 43595 75284 43596
rect 12376 43520 16651 43522
rect 12104 43384 16396 43460
rect 16749 43520 58603 43522
rect 17000 43384 58284 43460
rect 58701 43520 63044 43522
rect 59024 43453 63305 43460
rect 59024 43384 63316 43453
rect 64736 43520 64816 43595
rect 64914 43520 75284 43595
rect 65144 43384 75284 43460
rect 0 43285 75284 43324
rect 0 43248 16651 43285
rect 0 43112 10140 43188
rect 12104 43112 16396 43188
rect 16749 43248 58603 43285
rect 17000 43112 58284 43188
rect 58701 43248 75284 43285
rect 59024 43156 63316 43188
rect 59024 43112 63305 43156
rect 65144 43112 75284 43188
rect 0 42976 10548 43052
rect 12376 42976 63044 43052
rect 64736 42976 75284 43052
rect 0 42840 10140 42916
rect 10744 42840 16396 42916
rect 17000 42840 58284 42916
rect 59024 42840 64540 42916
rect 65144 42840 75284 42916
rect 0 42707 10438 42780
rect 10536 42707 10548 42780
rect 0 42704 10548 42707
rect 12376 42732 63044 42780
rect 12376 42704 16651 42732
rect 0 42568 11364 42644
rect 12104 42568 16396 42644
rect 16749 42704 58603 42732
rect 17000 42568 58284 42644
rect 58701 42704 63044 42732
rect 64736 42707 64816 42780
rect 64914 42707 75284 42780
rect 64736 42704 75284 42707
rect 59024 42568 63316 42644
rect 63920 42568 75284 42644
rect 0 42432 10548 42508
rect 11696 42495 63724 42508
rect 11696 42432 16651 42495
rect 16749 42432 58603 42495
rect 58701 42432 63724 42495
rect 64736 42432 75284 42508
rect 0 42296 10140 42372
rect 12104 42296 16396 42372
rect 17000 42296 58284 42372
rect 59024 42366 63316 42372
rect 59024 42296 63305 42366
rect 65144 42296 75284 42372
rect 0 42160 10548 42236
rect 12376 42179 63044 42236
rect 12376 42160 16651 42179
rect 0 42024 10140 42100
rect 12104 42024 16396 42100
rect 16749 42160 58603 42179
rect 17000 42024 58284 42100
rect 58701 42160 63044 42179
rect 64736 42160 75284 42236
rect 59024 42024 63316 42100
rect 65144 42024 75284 42100
rect 0 41917 10438 41964
rect 10536 41917 10548 41964
rect 0 41888 10548 41917
rect 12376 41942 63044 41964
rect 12376 41888 16651 41942
rect 16749 41888 58603 41942
rect 58701 41888 63044 41942
rect 64736 41917 64816 41964
rect 64914 41917 75284 41964
rect 64736 41888 75284 41917
rect 0 41752 11364 41828
rect 12104 41752 16396 41828
rect 17000 41752 58284 41828
rect 59024 41752 63316 41828
rect 63920 41752 75284 41828
rect 0 41616 10548 41692
rect 12376 41616 16651 41692
rect 16749 41616 58603 41692
rect 58701 41616 63044 41692
rect 64736 41616 75284 41692
rect 0 41480 10140 41556
rect 12104 41480 16396 41556
rect 17000 41480 58284 41556
rect 59024 41480 63305 41556
rect 65144 41480 75284 41556
rect 0 41344 11636 41420
rect 12376 41389 63044 41420
rect 12376 41344 16651 41389
rect 16749 41344 58603 41389
rect 58701 41344 63044 41389
rect 63648 41344 75284 41420
rect 0 41208 10140 41284
rect 0 41127 10438 41148
rect 12104 41208 16396 41284
rect 17000 41208 58284 41284
rect 59024 41208 63316 41284
rect 10536 41127 10548 41148
rect 0 41072 10548 41127
rect 12376 41072 16651 41148
rect 16749 41072 58603 41148
rect 58701 41072 63044 41148
rect 64736 41127 64816 41148
rect 65144 41208 75284 41284
rect 64914 41127 75284 41148
rect 64736 41072 75284 41127
rect 0 40936 16396 41012
rect 17000 40936 58284 41012
rect 59024 40936 75284 41012
rect 0 40809 10548 40876
rect 12376 40817 16651 40876
rect 16749 40817 58603 40876
rect 58701 40817 63044 40876
rect 0 40800 10438 40809
rect 0 40664 10140 40740
rect 10536 40800 10548 40809
rect 12376 40800 63044 40817
rect 64736 40809 75284 40876
rect 12104 40688 63305 40740
rect 64736 40800 64816 40809
rect 64914 40800 75284 40809
rect 12104 40664 63316 40688
rect 65144 40664 75284 40740
rect 0 40599 75284 40604
rect 0 40528 16651 40599
rect 16749 40528 58603 40599
rect 58701 40528 75284 40599
rect 0 40392 10140 40468
rect 12104 40392 16396 40468
rect 17000 40392 58284 40468
rect 59024 40392 63316 40468
rect 0 40256 10548 40332
rect 12376 40264 16651 40332
rect 16749 40264 58603 40332
rect 58701 40264 63044 40332
rect 65144 40392 75284 40468
rect 12376 40256 63044 40264
rect 64736 40256 75284 40332
rect 0 40120 16396 40196
rect 0 40019 10548 40060
rect 12376 40027 16651 40060
rect 17000 40120 58284 40196
rect 16749 40027 58603 40060
rect 59024 40120 75284 40196
rect 58701 40027 63044 40060
rect 0 39984 10438 40019
rect 0 39848 10140 39924
rect 10536 39984 10548 40019
rect 12376 39984 63044 40027
rect 64736 40019 75284 40060
rect 12104 39848 16396 39924
rect 17000 39848 58284 39924
rect 59024 39898 63305 39924
rect 64736 39984 64816 40019
rect 64914 39984 75284 40019
rect 59024 39848 63316 39898
rect 65144 39848 75284 39924
rect 0 39712 16651 39788
rect 16749 39712 58603 39788
rect 58701 39712 75284 39788
rect 0 39576 10140 39652
rect 0 39440 10548 39516
rect 12104 39576 16396 39652
rect 17000 39576 58284 39652
rect 59024 39601 63316 39652
rect 59024 39576 63305 39601
rect 12376 39474 16651 39516
rect 16749 39474 58603 39516
rect 58701 39474 63044 39516
rect 65144 39576 75284 39652
rect 12376 39440 63044 39474
rect 64736 39440 75284 39516
rect 0 39304 16396 39380
rect 0 39229 10548 39244
rect 12376 39237 16651 39244
rect 17000 39304 58284 39380
rect 16749 39237 58603 39244
rect 59024 39304 75284 39380
rect 58701 39237 63044 39244
rect 0 39168 10438 39229
rect 10536 39168 10548 39229
rect 12376 39168 63044 39237
rect 64736 39229 75284 39244
rect 64736 39168 64816 39229
rect 64914 39168 75284 39229
rect 0 39032 10140 39108
rect 12104 39032 16396 39108
rect 17000 39032 58284 39108
rect 59024 39032 63316 39108
rect 65144 39032 75284 39108
rect 0 38921 16651 38972
rect 16749 38921 58603 38972
rect 58701 38921 75284 38972
rect 0 38896 75284 38921
rect 0 38760 10140 38836
rect 1360 38624 10548 38700
rect 12104 38760 16396 38836
rect 12376 38684 16651 38700
rect 17000 38760 58284 38836
rect 59024 38811 63316 38836
rect 16749 38684 58603 38700
rect 59024 38760 63305 38811
rect 58701 38684 63044 38700
rect 65144 38760 75284 38836
rect 12376 38624 63044 38684
rect 64736 38624 75284 38700
rect 0 38494 455 38564
rect 553 38494 1191 38564
rect 1289 38494 10140 38564
rect 0 38488 10140 38494
rect 10744 38488 16396 38564
rect 17000 38488 58284 38564
rect 59024 38488 64540 38564
rect 65144 38488 75284 38564
rect 0 38352 10438 38428
rect 10536 38352 10548 38428
rect 12376 38352 63044 38428
rect 64736 38352 64816 38428
rect 64914 38352 75284 38428
rect 0 38216 10140 38292
rect 12104 38216 16396 38292
rect 0 38080 11636 38156
rect 12376 38131 16651 38156
rect 17000 38216 58284 38292
rect 16749 38131 58603 38156
rect 59024 38216 63316 38292
rect 65144 38216 75284 38292
rect 58701 38131 63044 38156
rect 12376 38080 63044 38131
rect 63648 38080 75284 38156
rect 1904 37944 10140 38020
rect 12104 37944 16396 38020
rect 17000 37944 58284 38020
rect 59024 37944 63305 38020
rect 65144 37944 75284 38020
rect 1904 37808 10548 37884
rect 12376 37808 63044 37884
rect 64736 37808 75284 37884
rect 0 37672 10140 37748
rect 12104 37672 16396 37748
rect 17000 37672 58284 37748
rect 59024 37672 63316 37748
rect 65144 37672 75284 37748
rect 0 37551 10438 37612
rect 10536 37551 10548 37612
rect 0 37536 10548 37551
rect 12376 37536 63044 37612
rect 64736 37551 64816 37612
rect 64914 37551 75284 37612
rect 64736 37536 75284 37551
rect 1360 37400 11364 37476
rect 12104 37400 16396 37476
rect 17000 37400 58284 37476
rect 59024 37400 63316 37476
rect 63920 37400 75284 37476
rect 0 37275 10548 37340
rect 0 37264 10438 37275
rect 0 37128 10140 37204
rect 10536 37264 10548 37275
rect 12376 37264 63044 37340
rect 64736 37275 75284 37340
rect 64736 37264 64816 37275
rect 12104 37128 16396 37204
rect 17000 37128 58284 37204
rect 59024 37133 63305 37204
rect 59024 37128 63316 37133
rect 64914 37264 75284 37275
rect 65144 37128 75284 37204
rect 1904 36992 10548 37068
rect 11696 36992 63724 37068
rect 64736 36992 75284 37068
rect 1904 36856 6876 36932
rect 0 36761 7148 36796
rect 7246 36761 7284 36796
rect 0 36720 7284 36761
rect 8976 36761 10438 36796
rect 10536 36761 10548 36796
rect 12104 36856 16396 36932
rect 17000 36856 58284 36932
rect 59024 36856 63316 36932
rect 8976 36720 10548 36761
rect 12376 36720 63044 36796
rect 64736 36761 64816 36796
rect 64914 36761 66308 36796
rect 64736 36720 66308 36761
rect 68000 36761 68106 36796
rect 68408 36856 75284 36932
rect 68204 36761 75284 36796
rect 68000 36720 75284 36761
rect 0 36584 16396 36660
rect 17000 36584 58284 36660
rect 59024 36584 75284 36660
rect 0 36485 10548 36524
rect 0 36448 10438 36485
rect 0 36352 10140 36388
rect 10536 36448 10548 36485
rect 12376 36448 63044 36524
rect 64736 36485 75284 36524
rect 64736 36448 64816 36485
rect 0 36312 455 36352
rect 553 36312 1191 36352
rect 1289 36312 10140 36352
rect 12104 36312 16396 36388
rect 17000 36312 58284 36388
rect 59024 36343 63305 36388
rect 59024 36312 63316 36343
rect 64914 36448 75284 36485
rect 65144 36312 75284 36388
rect 1360 36176 75284 36252
rect 0 36040 6876 36116
rect 0 35971 7148 35980
rect 7246 35971 7284 35980
rect 0 35904 7284 35971
rect 8976 35971 10438 35980
rect 10536 35971 10548 35980
rect 8976 35904 10548 35971
rect 12104 36040 16396 36116
rect 17000 36040 58284 36116
rect 59024 36046 63316 36116
rect 59024 36040 63305 36046
rect 12376 35904 63044 35980
rect 64736 35971 64816 35980
rect 64914 35971 66308 35980
rect 64736 35904 66308 35971
rect 68000 35971 68106 35980
rect 68408 36040 75284 36116
rect 68204 35971 75284 35980
rect 68000 35904 75284 35971
rect 1904 35768 16396 35844
rect 17000 35768 58284 35844
rect 59024 35768 75284 35844
rect 1904 35695 10548 35708
rect 1904 35632 10438 35695
rect 10536 35632 10548 35695
rect 0 35496 10140 35572
rect 12376 35632 63044 35708
rect 64736 35695 75284 35708
rect 12104 35496 16396 35572
rect 17000 35496 58284 35572
rect 59024 35553 63305 35572
rect 59024 35496 63316 35553
rect 64736 35632 64816 35695
rect 64914 35632 75284 35695
rect 65144 35496 75284 35572
rect 0 35385 75284 35436
rect 0 35360 16651 35385
rect 0 35134 455 35164
rect 553 35134 1191 35164
rect 1360 35224 6876 35300
rect 1289 35134 7284 35164
rect 0 35088 7284 35134
rect 8976 35088 10548 35164
rect 12104 35224 16396 35300
rect 16749 35360 58603 35385
rect 17000 35224 58284 35300
rect 58701 35360 75284 35385
rect 59024 35256 63316 35300
rect 59024 35224 63305 35256
rect 12376 35088 63044 35164
rect 64736 35088 66308 35164
rect 68408 35224 75284 35300
rect 68000 35088 75284 35164
rect 0 34952 10140 35028
rect 10744 34952 16396 35028
rect 17000 34952 58284 35028
rect 59024 34952 64540 35028
rect 65144 34952 75284 35028
rect 0 34816 10438 34892
rect 10536 34816 10548 34892
rect 1904 34680 10140 34756
rect 12376 34832 63044 34892
rect 12376 34816 16651 34832
rect 12104 34680 16396 34756
rect 16749 34816 58603 34832
rect 17000 34680 58284 34756
rect 58701 34816 63044 34832
rect 59024 34680 63316 34756
rect 64736 34816 64816 34892
rect 64914 34816 75284 34892
rect 65144 34680 75284 34756
rect 1904 34544 7284 34620
rect 8432 34544 10548 34620
rect 11696 34595 63724 34620
rect 11696 34544 16651 34595
rect 16749 34544 58603 34595
rect 58701 34544 63724 34595
rect 64736 34544 66988 34620
rect 68000 34544 75284 34620
rect 0 34408 5516 34484
rect 12104 34408 16396 34484
rect 17000 34408 58284 34484
rect 59024 34466 63316 34484
rect 59024 34408 63305 34466
rect 69768 34408 75284 34484
rect 0 34272 5788 34348
rect 8976 34272 10548 34348
rect 12376 34279 63044 34348
rect 12376 34272 16651 34279
rect 0 34136 10140 34212
rect 10744 34136 16396 34212
rect 16749 34272 58603 34279
rect 17000 34136 58284 34212
rect 58701 34272 63044 34279
rect 64736 34272 66308 34348
rect 69496 34272 75284 34348
rect 59024 34136 64540 34212
rect 65144 34136 75284 34212
rect 1360 34017 10438 34076
rect 10536 34017 10548 34076
rect 1360 34000 10548 34017
rect 12376 34042 63044 34076
rect 12376 34000 16651 34042
rect 16749 34000 58603 34042
rect 58701 34000 63044 34042
rect 64736 34017 64816 34076
rect 64914 34017 75284 34076
rect 64736 34000 75284 34017
rect 0 33864 11364 33940
rect 12104 33864 16396 33940
rect 17000 33864 58284 33940
rect 59024 33864 63316 33940
rect 63920 33864 75284 33940
rect 0 33728 10548 33804
rect 12376 33728 16651 33804
rect 16749 33728 58603 33804
rect 58701 33728 63044 33804
rect 64736 33728 75284 33804
rect 0 33592 10140 33668
rect 12104 33592 16396 33668
rect 17000 33592 58284 33668
rect 59024 33592 63305 33668
rect 65144 33592 75284 33668
rect 1904 33456 11636 33532
rect 12376 33489 63044 33532
rect 12376 33456 16651 33489
rect 1904 33320 10140 33396
rect 0 33227 10438 33260
rect 12104 33320 16396 33396
rect 16749 33456 58603 33489
rect 17000 33320 58284 33396
rect 58701 33456 63044 33489
rect 63648 33456 75284 33532
rect 59024 33320 63316 33396
rect 10536 33227 10548 33260
rect 0 33184 10548 33227
rect 12376 33252 63044 33260
rect 12376 33184 16651 33252
rect 16749 33184 58603 33252
rect 58701 33184 63044 33252
rect 64736 33227 64816 33260
rect 65144 33320 75284 33396
rect 64914 33227 75284 33260
rect 64736 33184 75284 33227
rect 1360 33048 11364 33124
rect 12104 33048 16396 33124
rect 17000 33048 58284 33124
rect 59024 33048 63316 33124
rect 63920 33048 75284 33124
rect 0 32912 455 32988
rect 553 32912 1191 32988
rect 1289 32912 7692 32988
rect 8976 32912 10548 32988
rect 12376 32917 16651 32988
rect 16749 32917 58603 32988
rect 58701 32917 63044 32988
rect 12376 32912 63044 32917
rect 64736 32912 66308 32988
rect 67592 32912 75284 32988
rect 1360 32776 7284 32852
rect 12104 32788 63305 32852
rect 12104 32776 63316 32788
rect 68000 32776 75284 32852
rect 0 32699 75284 32716
rect 0 32640 16651 32699
rect 16749 32640 58603 32699
rect 58701 32640 75284 32699
rect 1904 32504 10140 32580
rect 1904 32437 10438 32444
rect 12104 32504 16396 32580
rect 17000 32504 58284 32580
rect 59024 32504 63316 32580
rect 10536 32437 10548 32444
rect 1904 32368 10548 32437
rect 12376 32368 16651 32444
rect 16749 32368 58603 32444
rect 58701 32368 63044 32444
rect 64736 32437 64816 32444
rect 65144 32504 75284 32580
rect 64914 32437 75284 32444
rect 64736 32368 75284 32437
rect 0 32232 16396 32308
rect 17000 32232 58284 32308
rect 59024 32232 75284 32308
rect 0 32096 6468 32172
rect 8976 32119 10548 32172
rect 12376 32127 16651 32172
rect 16749 32127 58603 32172
rect 58701 32127 63044 32172
rect 0 31960 6196 32036
rect 8976 32096 10438 32119
rect 10536 32096 10548 32119
rect 12376 32096 63044 32127
rect 64736 32119 66308 32172
rect 12104 31960 16396 32036
rect 17000 31960 58284 32036
rect 59024 31998 63305 32036
rect 64736 32096 64816 32119
rect 64914 32096 66308 32119
rect 68952 32096 75284 32172
rect 59024 31960 63316 31998
rect 69224 31960 75284 32036
rect 1360 31824 16651 31900
rect 16749 31824 58603 31900
rect 58701 31824 75284 31900
rect 0 31688 10140 31764
rect 0 31552 10548 31628
rect 12104 31688 16396 31764
rect 17000 31688 58284 31764
rect 59024 31701 63316 31764
rect 59024 31688 63305 31701
rect 12376 31574 16651 31628
rect 16749 31574 58603 31628
rect 58701 31574 63044 31628
rect 65144 31688 75284 31764
rect 12376 31552 63044 31574
rect 64736 31552 75284 31628
rect 0 31416 16396 31492
rect 1904 31329 10548 31356
rect 12376 31337 16651 31356
rect 17000 31416 58284 31492
rect 16749 31337 58603 31356
rect 59024 31416 75284 31492
rect 58701 31337 63044 31356
rect 1904 31280 10438 31329
rect 10536 31280 10548 31329
rect 1904 31144 10140 31220
rect 12376 31280 63044 31337
rect 64736 31329 75284 31356
rect 12104 31144 16396 31220
rect 17000 31144 58284 31220
rect 59024 31208 63305 31220
rect 64736 31280 64816 31329
rect 64914 31280 75284 31329
rect 59024 31144 63316 31208
rect 65144 31144 75284 31220
rect 0 31021 16651 31084
rect 16749 31021 58603 31084
rect 58701 31021 75284 31084
rect 0 31008 75284 31021
rect 0 30872 10140 30948
rect 0 30752 10548 30812
rect 12104 30872 16396 30948
rect 0 30736 455 30752
rect 553 30736 1191 30752
rect 1289 30736 10548 30752
rect 12376 30784 16651 30812
rect 17000 30872 58284 30948
rect 59024 30911 63316 30948
rect 16749 30784 58603 30812
rect 59024 30872 63305 30911
rect 58701 30784 63044 30812
rect 65144 30872 75284 30948
rect 12376 30736 63044 30784
rect 64736 30736 75284 30812
rect 1360 30600 16396 30676
rect 17000 30600 58284 30676
rect 59024 30600 75284 30676
rect 0 30523 7692 30540
rect 8976 30539 10548 30540
rect 0 30464 7583 30523
rect 7681 30464 7692 30523
rect 8976 30464 10438 30539
rect 10536 30464 10548 30539
rect 12376 30464 63044 30540
rect 64736 30539 66308 30540
rect 64736 30464 64816 30539
rect 64914 30464 66308 30539
rect 67592 30523 75284 30540
rect 67592 30464 67671 30523
rect 67769 30464 75284 30523
rect 0 30328 7284 30404
rect 12104 30328 16396 30404
rect 1904 30231 16651 30268
rect 17000 30328 58284 30404
rect 16749 30231 58603 30268
rect 59024 30328 63316 30404
rect 68000 30328 75284 30404
rect 58701 30231 75284 30268
rect 1904 30192 75284 30231
rect 1904 30056 10140 30132
rect 12104 30056 16396 30132
rect 0 29920 10548 29996
rect 12376 29994 16651 29996
rect 17000 30056 58284 30132
rect 59024 30121 63316 30132
rect 16749 29994 58603 29996
rect 59024 30056 63305 30121
rect 65144 30056 75284 30132
rect 58701 29994 63044 29996
rect 12376 29920 63044 29994
rect 64736 29920 75284 29996
rect 0 29784 6196 29860
rect 12104 29784 16396 29860
rect 17000 29784 58284 29860
rect 59024 29784 63316 29860
rect 69224 29784 75284 29860
rect 1360 29648 6413 29724
rect 0 29534 455 29588
rect 553 29534 1191 29588
rect 8976 29651 10438 29724
rect 10536 29651 10548 29724
rect 8976 29648 10548 29651
rect 12376 29648 63044 29724
rect 64736 29651 64816 29724
rect 64914 29651 66308 29724
rect 64736 29648 66308 29651
rect 68952 29648 75284 29724
rect 1289 29534 6196 29588
rect 0 29512 6196 29534
rect 8704 29512 11364 29588
rect 12104 29512 16396 29588
rect 0 29441 16651 29452
rect 17000 29512 58284 29588
rect 16749 29441 58603 29452
rect 59024 29512 63316 29588
rect 63920 29512 66580 29588
rect 69224 29512 75284 29588
rect 58701 29441 75284 29452
rect 0 29376 75284 29441
rect 0 29240 16396 29316
rect 17000 29240 58284 29316
rect 59024 29240 75284 29316
rect 0 29104 75284 29180
rect 1904 28968 16396 29044
rect 17000 28968 58284 29044
rect 59024 28968 71204 29044
rect 71808 28968 75284 29044
rect 1904 28832 75284 28908
rect 2040 28741 70524 28772
rect 2040 28696 17347 28741
rect 17445 28696 17971 28741
rect 18069 28696 18595 28741
rect 18693 28696 19219 28741
rect 19317 28696 19843 28741
rect 19941 28696 20467 28741
rect 20565 28696 21091 28741
rect 21189 28696 21715 28741
rect 21813 28696 22339 28741
rect 22437 28696 22963 28741
rect 23061 28696 23587 28741
rect 23685 28696 24211 28741
rect 24309 28696 24835 28741
rect 24933 28696 25459 28741
rect 25557 28696 26083 28741
rect 26181 28696 26707 28741
rect 26805 28696 27331 28741
rect 27429 28696 27955 28741
rect 28053 28696 28579 28741
rect 28677 28696 29203 28741
rect 29301 28696 29827 28741
rect 29925 28696 30451 28741
rect 30549 28696 31075 28741
rect 31173 28696 31699 28741
rect 31797 28696 32323 28741
rect 32421 28696 32947 28741
rect 33045 28696 33571 28741
rect 33669 28696 34195 28741
rect 34293 28696 34819 28741
rect 34917 28696 35443 28741
rect 35541 28696 36067 28741
rect 36165 28696 36691 28741
rect 36789 28696 37315 28741
rect 37413 28696 37939 28741
rect 38037 28696 38563 28741
rect 38661 28696 39187 28741
rect 39285 28696 39811 28741
rect 39909 28696 40435 28741
rect 40533 28696 41059 28741
rect 41157 28696 41683 28741
rect 41781 28696 42307 28741
rect 42405 28696 42931 28741
rect 43029 28696 43555 28741
rect 43653 28696 44179 28741
rect 44277 28696 44803 28741
rect 44901 28696 45427 28741
rect 45525 28696 46051 28741
rect 46149 28696 46675 28741
rect 46773 28696 47299 28741
rect 47397 28696 47923 28741
rect 48021 28696 48547 28741
rect 48645 28696 49171 28741
rect 49269 28696 49795 28741
rect 49893 28696 50419 28741
rect 50517 28696 51043 28741
rect 51141 28696 51667 28741
rect 51765 28696 52291 28741
rect 52389 28696 52915 28741
rect 53013 28696 53539 28741
rect 53637 28696 54163 28741
rect 54261 28696 54787 28741
rect 54885 28696 55411 28741
rect 55509 28696 56035 28741
rect 56133 28696 56659 28741
rect 56757 28696 57283 28741
rect 57381 28696 57907 28741
rect 58005 28696 70524 28741
rect 72352 28696 75284 28772
rect 2040 28560 17076 28636
rect 58208 28560 70524 28636
rect 72352 28560 75284 28636
rect 1360 28424 70388 28500
rect 75266 28382 75326 28442
rect 0 28352 70388 28364
rect 0 28288 4361 28352
rect 4459 28288 70388 28352
rect 0 28152 4156 28228
rect 4624 28152 75284 28228
rect 0 28016 17212 28092
rect 57800 28016 75284 28092
rect 0 27880 75284 27956
rect 0 27744 75284 27820
rect 0 27608 4156 27684
rect 16184 27611 75284 27684
rect 16184 27608 71477 27611
rect 0 27472 4156 27548
rect 57936 27472 71204 27548
rect 71575 27608 75284 27611
rect 71808 27472 75284 27548
rect 0 27336 1572 27412
rect 57936 27336 75284 27412
rect 0 27200 1572 27276
rect 17952 27200 75284 27276
rect 0 27064 75284 27140
rect 0 26928 4156 27004
rect 0 26840 4361 26868
rect 4624 26928 75284 27004
rect 4459 26840 10820 26868
rect 0 26792 10820 26840
rect 11424 26792 70252 26868
rect 0 26656 11101 26732
rect 11199 26656 70252 26732
rect 75266 26682 75326 26742
rect 0 26520 10820 26596
rect 11424 26520 18028 26596
rect 57392 26520 75284 26596
rect 0 26384 75284 26460
rect 0 26248 71204 26324
rect 71808 26248 75284 26324
rect 0 26112 71477 26188
rect 71575 26112 75284 26188
rect 0 25976 11228 26052
rect 12240 25976 71204 26052
rect 71808 25976 75284 26052
rect 0 25840 11228 25916
rect 12240 25840 18300 25916
rect 57664 25840 75284 25916
rect 0 25704 11500 25780
rect 57936 25704 75284 25780
rect 0 25568 1708 25644
rect 3128 25568 11500 25644
rect 57936 25568 70252 25644
rect 75266 25554 75326 25614
rect 0 25432 1708 25508
rect 4624 25432 17484 25508
rect 57800 25432 70252 25508
rect 0 25296 10820 25372
rect 0 25232 11101 25236
rect 11424 25296 18028 25372
rect 57392 25296 75284 25372
rect 11199 25232 75284 25236
rect 0 25160 75284 25232
rect 0 25024 75284 25100
rect 0 24888 15580 24964
rect 57936 24888 75284 24964
rect 0 24752 4156 24828
rect 57936 24752 71204 24828
rect 0 24616 4156 24692
rect 57120 24685 71477 24692
rect 71808 24752 75284 24828
rect 71575 24685 75284 24692
rect 57120 24616 75284 24685
rect 0 24480 10276 24556
rect 12104 24480 75284 24556
rect 0 24344 75284 24420
rect 0 24208 75284 24284
rect 0 24110 75284 24148
rect 0 24072 4361 24110
rect 4459 24072 75284 24110
rect 0 23936 4156 24012
rect 4624 23936 17756 24012
rect 57120 23936 70116 24012
rect 0 23800 10820 23876
rect 11424 23800 70116 23876
rect 75266 23854 75326 23914
rect 0 23664 75284 23740
rect 0 23528 75284 23604
rect 0 23392 4156 23468
rect 16320 23392 75284 23468
rect 0 23256 4156 23332
rect 16320 23256 71204 23332
rect 71808 23256 75284 23332
rect 0 23120 17756 23196
rect 57120 23120 75284 23196
rect 0 22984 75284 23060
rect 0 22870 71612 22924
rect 0 22848 18040 22870
rect 0 22712 4156 22788
rect 4624 22712 17484 22788
rect 18138 22848 19288 22870
rect 19386 22848 20536 22870
rect 20634 22848 21784 22870
rect 21882 22848 23032 22870
rect 23130 22848 24280 22870
rect 24378 22848 25528 22870
rect 25626 22848 26776 22870
rect 26874 22848 28024 22870
rect 28122 22848 29272 22870
rect 29370 22848 30520 22870
rect 30618 22848 31768 22870
rect 31866 22848 33016 22870
rect 33114 22848 34264 22870
rect 34362 22848 35512 22870
rect 35610 22848 36760 22870
rect 36858 22848 38008 22870
rect 38106 22848 39256 22870
rect 39354 22848 40504 22870
rect 40602 22848 41752 22870
rect 41850 22848 43000 22870
rect 43098 22848 44248 22870
rect 44346 22848 45496 22870
rect 45594 22848 46744 22870
rect 46842 22848 47992 22870
rect 48090 22848 49240 22870
rect 49338 22848 50488 22870
rect 50586 22848 51736 22870
rect 51834 22848 52984 22870
rect 53082 22848 54232 22870
rect 54330 22848 55480 22870
rect 55578 22848 56728 22870
rect 56826 22848 71612 22870
rect 72216 22848 75284 22924
rect 57120 22712 69980 22788
rect 75266 22726 75326 22786
rect 0 22598 4361 22652
rect 4459 22598 17484 22652
rect 0 22576 17484 22598
rect 56848 22576 69980 22652
rect 71264 22576 75284 22652
rect 0 22440 75284 22516
rect 0 22304 75284 22380
rect 0 22168 75284 22244
rect 0 22032 4156 22108
rect 4624 22032 15988 22108
rect 16456 22077 75284 22108
rect 16456 22032 17926 22077
rect 18024 22032 19174 22077
rect 19272 22032 20422 22077
rect 20520 22032 21670 22077
rect 21768 22032 22918 22077
rect 23016 22032 24166 22077
rect 24264 22032 25414 22077
rect 25512 22032 26662 22077
rect 26760 22032 27910 22077
rect 28008 22032 29158 22077
rect 29256 22032 30406 22077
rect 30504 22032 31654 22077
rect 31752 22032 32902 22077
rect 33000 22032 34150 22077
rect 34248 22032 35398 22077
rect 35496 22032 36646 22077
rect 36744 22032 37894 22077
rect 37992 22032 39142 22077
rect 39240 22032 40390 22077
rect 40488 22032 41638 22077
rect 41736 22032 42886 22077
rect 42984 22032 44134 22077
rect 44232 22032 45382 22077
rect 45480 22032 46630 22077
rect 46728 22032 47878 22077
rect 47976 22032 49126 22077
rect 49224 22032 50374 22077
rect 50472 22032 51622 22077
rect 51720 22032 52870 22077
rect 52968 22032 54118 22077
rect 54216 22032 55366 22077
rect 55464 22032 56614 22077
rect 56712 22032 75284 22077
rect 0 21896 4156 21972
rect 56984 21955 75284 21972
rect 56984 21896 71477 21955
rect 71575 21896 75284 21955
rect 0 21760 71204 21836
rect 71808 21760 75284 21836
rect 0 21640 75284 21700
rect 0 21624 17915 21640
rect 0 21488 17620 21564
rect 18013 21624 19163 21640
rect 19261 21624 20411 21640
rect 20509 21624 21659 21640
rect 21757 21624 22907 21640
rect 23005 21624 24155 21640
rect 24253 21624 25403 21640
rect 25501 21624 26651 21640
rect 26749 21624 27899 21640
rect 27997 21624 29147 21640
rect 29245 21624 30395 21640
rect 30493 21624 31643 21640
rect 31741 21624 32891 21640
rect 32989 21624 34139 21640
rect 34237 21624 35387 21640
rect 35485 21624 36635 21640
rect 36733 21624 37883 21640
rect 37981 21624 39131 21640
rect 39229 21624 40379 21640
rect 40477 21624 41627 21640
rect 41725 21624 42875 21640
rect 42973 21624 44123 21640
rect 44221 21624 45371 21640
rect 45469 21624 46619 21640
rect 46717 21624 47867 21640
rect 47965 21624 49115 21640
rect 49213 21624 50363 21640
rect 50461 21624 51611 21640
rect 51709 21624 52859 21640
rect 52957 21624 54107 21640
rect 54205 21624 55355 21640
rect 55453 21624 56603 21640
rect 56701 21624 75284 21640
rect 56984 21488 75284 21564
rect 0 21352 17756 21428
rect 57120 21352 75284 21428
rect 0 21216 4156 21292
rect 4624 21216 18036 21292
rect 18134 21216 19284 21292
rect 19382 21216 20532 21292
rect 20630 21216 21780 21292
rect 21878 21216 23028 21292
rect 23126 21216 24276 21292
rect 24374 21216 25524 21292
rect 25622 21216 26772 21292
rect 26870 21216 28020 21292
rect 28118 21216 29268 21292
rect 29366 21216 30516 21292
rect 30614 21216 31764 21292
rect 31862 21216 33012 21292
rect 33110 21216 34260 21292
rect 34358 21216 35508 21292
rect 35606 21216 36756 21292
rect 36854 21216 38004 21292
rect 38102 21216 39252 21292
rect 39350 21216 40500 21292
rect 40598 21216 41748 21292
rect 41846 21216 42996 21292
rect 43094 21216 44244 21292
rect 44342 21216 45492 21292
rect 45590 21216 46740 21292
rect 46838 21216 47988 21292
rect 48086 21216 49236 21292
rect 49334 21216 50484 21292
rect 50582 21216 51732 21292
rect 51830 21216 52980 21292
rect 53078 21216 54228 21292
rect 54326 21216 55476 21292
rect 55574 21216 56724 21292
rect 56822 21216 69980 21292
rect 71264 21216 75284 21292
rect 0 21080 17620 21156
rect 0 21008 17921 21020
rect 18019 21008 19169 21020
rect 19267 21008 20417 21020
rect 20515 21008 21665 21020
rect 21763 21008 22913 21020
rect 23011 21008 24161 21020
rect 24259 21008 25409 21020
rect 25507 21008 26657 21020
rect 26755 21008 27905 21020
rect 28003 21008 29153 21020
rect 29251 21008 30401 21020
rect 30499 21008 31649 21020
rect 31747 21008 32897 21020
rect 32995 21008 34145 21020
rect 34243 21008 35393 21020
rect 35491 21008 36641 21020
rect 36739 21008 37889 21020
rect 37987 21008 39137 21020
rect 39235 21008 40385 21020
rect 40483 21008 41633 21020
rect 41731 21008 42881 21020
rect 42979 21008 44129 21020
rect 44227 21008 45377 21020
rect 45475 21008 46625 21020
rect 46723 21008 47873 21020
rect 47971 21008 49121 21020
rect 49219 21008 50369 21020
rect 50467 21008 51617 21020
rect 51715 21008 52865 21020
rect 52963 21008 54113 21020
rect 54211 21008 55361 21020
rect 55459 21008 56609 21020
rect 57120 21080 69980 21156
rect 75266 21026 75326 21086
rect 56707 21008 71612 21020
rect 0 20944 71612 21008
rect 0 20808 75284 20884
rect 0 20672 17620 20748
rect 0 20536 1980 20612
rect 3536 20536 17620 20612
rect 56984 20672 75284 20748
rect 56984 20536 71204 20612
rect 0 20400 1980 20476
rect 3536 20400 17620 20476
rect 56984 20443 71477 20476
rect 71808 20536 75284 20612
rect 71575 20443 75284 20476
rect 56984 20400 75284 20443
rect 0 20264 75284 20340
rect 0 20128 17756 20204
rect 18360 20128 27684 20204
rect 28424 20128 37748 20204
rect 38352 20128 47676 20204
rect 48280 20128 75284 20204
rect 0 19992 71612 20068
rect 0 19870 69844 19932
rect 75266 19898 75326 19958
rect 0 19856 7 19870
rect 105 19868 69844 19870
rect 105 19856 4361 19868
rect 272 19720 4156 19796
rect 4459 19856 69844 19868
rect 4624 19720 69844 19796
rect 71264 19720 75284 19796
rect 0 19584 15716 19660
rect 57936 19584 75284 19660
rect 0 19448 15716 19524
rect 57936 19448 75284 19524
rect 3536 19312 17348 19388
rect 18088 19312 27412 19388
rect 28016 19312 37340 19388
rect 38080 19312 47268 19388
rect 48008 19312 75284 19388
rect 26 19225 86 19285
rect 3536 19176 17348 19252
rect 18360 19176 27412 19252
rect 28424 19176 37340 19252
rect 38352 19176 47268 19252
rect 48280 19176 75284 19252
rect 0 19040 18032 19116
rect 18130 19040 28016 19116
rect 28114 19040 38000 19116
rect 38098 19040 47984 19116
rect 48082 19040 71204 19116
rect 71808 19040 75284 19116
rect 2448 18904 17756 18980
rect 18360 18904 27684 18980
rect 28424 18904 37748 18980
rect 38352 18904 47676 18980
rect 48280 18904 75284 18980
rect 2448 18768 75284 18844
rect 0 18632 1844 18708
rect 3808 18632 75284 18708
rect 272 18496 1844 18572
rect 4624 18496 75284 18572
rect 0 18360 7 18436
rect 105 18360 4361 18436
rect 4459 18360 75284 18436
rect 272 18224 4156 18300
rect 4624 18224 39516 18300
rect 48144 18224 75284 18300
rect 0 18088 25508 18164
rect 33048 18088 75284 18164
rect 2720 17952 25508 18028
rect 33048 17952 75284 18028
rect 2720 17816 19660 17892
rect 26928 17816 75284 17892
rect 0 17680 2524 17756
rect 2992 17680 19660 17756
rect 26928 17680 75284 17756
rect 26 17525 86 17585
rect 408 17544 2524 17620
rect 2992 17544 20476 17620
rect 27064 17544 75284 17620
rect 408 17408 20476 17484
rect 27064 17408 75284 17484
rect 0 17272 26324 17348
rect 33320 17272 75284 17348
rect 0 17136 2252 17212
rect 4488 17136 26324 17212
rect 33320 17136 75284 17212
rect 272 17000 2252 17076
rect 4624 17000 32580 17076
rect 40664 17000 75284 17076
rect 0 16864 33396 16940
rect 40800 16864 75284 16940
rect 0 16728 33396 16804
rect 40800 16728 75284 16804
rect 0 16592 40332 16668
rect 48280 16592 75284 16668
rect 0 16456 40332 16532
rect 48280 16456 75284 16532
rect 0 16320 47676 16396
rect 56848 16320 75284 16396
rect 0 16184 47676 16260
rect 56848 16184 75284 16260
rect 0 16048 38292 16124
rect 46784 16048 75284 16124
rect 0 15912 38292 15988
rect 47056 15912 75284 15988
rect 0 15776 39244 15852
rect 47056 15776 75284 15852
rect 0 15640 46588 15716
rect 55624 15640 75284 15716
rect 0 15504 46588 15580
rect 55624 15504 75284 15580
rect 0 15368 23196 15444
rect 30600 15368 75284 15444
rect 0 15232 23196 15308
rect 30600 15232 75284 15308
rect 0 15096 11500 15172
rect 18088 15096 75284 15172
rect 0 14960 11500 15036
rect 18088 14960 75284 15036
rect 0 14824 7692 14900
rect 17952 14824 75284 14900
rect 0 14688 7692 14764
rect 24344 14688 75284 14764
rect 0 14552 17348 14628
rect 24344 14552 75284 14628
rect 0 14416 18164 14492
rect 24480 14416 75284 14492
rect 0 14280 18164 14356
rect 24480 14280 75284 14356
rect 0 14144 24012 14220
rect 30736 14144 75284 14220
rect 0 14008 24012 14084
rect 30736 14008 75284 14084
rect 0 13872 30132 13948
rect 38080 13872 75284 13948
rect 0 13736 30132 13812
rect 38080 13736 75284 13812
rect 0 13600 10004 13676
rect 37944 13600 75284 13676
rect 0 13464 10004 13540
rect 45560 13464 75284 13540
rect 0 13328 37204 13404
rect 45560 13328 75284 13404
rect 0 13192 38020 13268
rect 45696 13192 75284 13268
rect 0 13056 38020 13132
rect 45696 13056 75284 13132
rect 0 12920 45364 12996
rect 54264 12920 75284 12996
rect 0 12784 45364 12860
rect 54264 12784 75284 12860
rect 0 12648 44140 12724
rect 53040 12648 75284 12724
rect 0 12512 44140 12588
rect 53040 12512 75284 12588
rect 0 12376 43052 12452
rect 51816 12376 75284 12452
rect 0 12240 41828 12316
rect 51816 12240 75284 12316
rect 0 12104 41828 12180
rect 50592 12104 75284 12180
rect 0 11968 40740 12044
rect 49368 11968 75284 12044
rect 0 11832 40740 11908
rect 49368 11832 75284 11908
rect 0 11696 21972 11772
rect 29376 11696 75284 11772
rect 0 11560 21972 11636
rect 29376 11560 75284 11636
rect 0 11424 16124 11500
rect 23120 11424 75284 11500
rect 0 11288 16124 11364
rect 23120 11288 75284 11364
rect 0 11152 16940 11228
rect 23256 11152 75284 11228
rect 0 11016 22788 11092
rect 29512 11016 75284 11092
rect 0 10880 22788 10956
rect 29512 10880 75284 10956
rect 0 10744 29044 10820
rect 36856 10744 75284 10820
rect 0 10608 29044 10684
rect 36856 10608 75284 10684
rect 0 10472 35980 10548
rect 44336 10472 75284 10548
rect 0 10336 35980 10412
rect 44336 10336 75284 10412
rect 0 10200 20884 10276
rect 28152 10200 75284 10276
rect 0 10064 20884 10140
rect 28152 10064 75284 10140
rect 0 9928 15036 10004
rect 21896 9928 75284 10004
rect 0 9792 15852 9868
rect 22032 9792 75284 9868
rect 0 9656 15852 9732
rect 22032 9656 75284 9732
rect 0 9520 21700 9596
rect 28288 9520 75284 9596
rect 0 9384 21700 9460
rect 28288 9384 75284 9460
rect 0 9248 27820 9324
rect 35632 9248 75284 9324
rect 0 9112 27820 9188
rect 35632 9112 75284 9188
rect 0 8976 34892 9052
rect 43112 8976 75284 9052
rect 0 8840 34892 8916
rect 43112 8840 75284 8916
rect 0 8704 26732 8780
rect 34408 8704 75284 8780
rect 0 8568 8780 8644
rect 28016 8568 75284 8644
rect 0 8432 8780 8508
rect 28016 8432 75284 8508
rect 0 8296 27548 8372
rect 34544 8296 75284 8372
rect 0 8160 27548 8236
rect 34544 8160 75284 8236
rect 0 8024 33668 8100
rect 41888 8024 75284 8100
rect 0 7888 33668 7964
rect 41888 7888 75284 7964
rect 0 7752 24284 7828
rect 31824 7752 75284 7828
rect 0 7616 18436 7692
rect 19040 7616 24284 7692
rect 31824 7616 75284 7692
rect 0 7480 18436 7556
rect 25568 7480 75284 7556
rect 0 7344 19388 7420
rect 25840 7344 75284 7420
rect 0 7208 19388 7284
rect 25840 7208 75284 7284
rect 0 7072 25100 7148
rect 31960 7072 75284 7148
rect 0 6936 25100 7012
rect 31960 6936 75284 7012
rect 0 6800 31356 6876
rect 39304 6800 75284 6876
rect 0 6664 31356 6740
rect 39304 6664 75284 6740
rect 0 6528 13812 6604
rect 20672 6528 75284 6604
rect 0 6392 12724 6468
rect 20672 6392 75284 6468
rect 0 6256 12724 6332
rect 19448 6256 75284 6332
rect 0 6120 48492 6196
rect 56984 6120 75284 6196
rect 0 5984 48492 6060
rect 56984 5984 75284 6060
rect 0 5848 11092 5924
rect 48008 5848 75284 5924
rect 0 5712 11092 5788
rect 48008 5712 75284 5788
rect 0 5576 47404 5652
rect 55760 5576 75284 5652
rect 0 5440 47404 5516
rect 55760 5440 75284 5516
rect 0 5304 46180 5380
rect 54536 5304 75284 5380
rect 0 5168 44956 5244
rect 54536 5168 75284 5244
rect 0 5032 44956 5108
rect 53176 5032 75284 5108
rect 0 4896 36796 4972
rect 44472 4896 75284 4972
rect 0 4760 36796 4836
rect 44472 4760 75284 4836
rect 0 4624 43868 4700
rect 51952 4624 75284 4700
rect 0 4488 43868 4564
rect 51952 4488 75284 4564
rect 0 4352 35708 4428
rect 43248 4352 75284 4428
rect 0 4216 35708 4292
rect 43248 4216 75284 4292
rect 0 4080 42644 4156
rect 50728 4080 75284 4156
rect 0 3944 34484 4020
rect 50728 3944 75284 4020
rect 0 3808 34484 3884
rect 42024 3808 75284 3884
rect 0 3672 41556 3748
rect 49504 3672 75284 3748
rect 0 3536 41556 3612
rect 49504 3536 75284 3612
rect 0 3400 32172 3476
rect 39576 3400 75284 3476
rect 0 3264 32172 3340
rect 39576 3264 75284 3340
rect 0 3128 30948 3204
rect 38216 3128 75284 3204
rect 0 2992 30948 3068
rect 38216 2992 75284 3068
rect 0 2856 29860 2932
rect 36992 2856 75284 2932
rect 0 2720 28636 2796
rect 35768 2720 75284 2796
rect 0 2584 28636 2660
rect 35768 2584 75284 2660
rect 0 2448 14628 2524
rect 20808 2448 75284 2524
rect 0 2312 14628 2388
rect 20808 2312 75284 2388
rect 0 2176 13540 2252
rect 19584 2176 75284 2252
rect 0 2040 13540 2116
rect 19584 2040 75284 2116
rect 0 1904 12316 1980
rect 18360 1904 75284 1980
rect 0 1768 12316 1844
rect 18360 1768 75284 1844
rect 0 1632 6468 1708
rect 11016 1632 75284 1708
rect 0 1559 75284 1572
rect 0 1496 6197 1559
rect 6295 1496 7365 1559
rect 7463 1496 8533 1559
rect 8631 1496 9701 1559
rect 9799 1496 10869 1559
rect 10967 1496 12037 1559
rect 12135 1496 13205 1559
rect 13303 1496 14373 1559
rect 14471 1496 15541 1559
rect 15639 1496 16709 1559
rect 16807 1496 17877 1559
rect 17975 1496 19045 1559
rect 19143 1496 20213 1559
rect 20311 1496 21381 1559
rect 21479 1496 22549 1559
rect 22647 1496 23717 1559
rect 23815 1496 24885 1559
rect 24983 1496 26053 1559
rect 26151 1496 27221 1559
rect 27319 1496 28389 1559
rect 28487 1496 29557 1559
rect 29655 1496 30725 1559
rect 30823 1496 31893 1559
rect 31991 1496 33061 1559
rect 33159 1496 34229 1559
rect 34327 1496 35397 1559
rect 35495 1496 36565 1559
rect 36663 1496 37733 1559
rect 37831 1496 38901 1559
rect 38999 1496 40069 1559
rect 40167 1496 41237 1559
rect 41335 1496 42405 1559
rect 42503 1496 43573 1559
rect 43671 1496 44741 1559
rect 44839 1496 45909 1559
rect 46007 1496 47077 1559
rect 47175 1496 48245 1559
rect 48343 1496 75284 1559
rect 0 1360 5924 1436
rect 48552 1360 75284 1436
rect 0 1224 75284 1300
rect 0 1088 75284 1164
rect 0 952 75284 1028
rect 0 816 6468 892
rect 49232 816 75284 892
rect 0 680 5516 756
rect 49232 680 75284 756
rect 0 544 5516 620
rect 48280 544 75284 620
rect 0 408 4292 484
rect 49096 408 75284 484
rect 0 272 4292 348
rect 49096 272 75284 348
rect 0 136 5924 212
rect 0 47 6197 76
rect 6295 47 7365 76
rect 7463 47 8533 76
rect 8631 47 9701 76
rect 9799 47 10869 76
rect 10967 47 12037 76
rect 12135 47 13205 76
rect 13303 47 14373 76
rect 14471 47 15541 76
rect 15639 47 16709 76
rect 16807 47 17877 76
rect 17975 47 19045 76
rect 19143 47 20213 76
rect 20311 47 21381 76
rect 21479 47 22549 76
rect 22647 47 23717 76
rect 23815 47 24885 76
rect 24983 47 26053 76
rect 26151 47 27221 76
rect 27319 47 28389 76
rect 28487 47 29557 76
rect 29655 47 30725 76
rect 30823 47 31893 76
rect 31991 47 33061 76
rect 33159 47 34229 76
rect 34327 47 35397 76
rect 35495 47 36565 76
rect 36663 47 37733 76
rect 37831 47 38901 76
rect 38999 47 40069 76
rect 40167 47 41237 76
rect 41335 47 42405 76
rect 42503 47 43573 76
rect 43671 47 44741 76
rect 44839 47 45909 76
rect 46007 47 47077 76
rect 47175 47 48245 76
rect 48552 136 75284 212
rect 48343 47 75284 76
rect 0 0 75284 47
<< obsm3 >>
rect 70977 89198 71075 89296
rect 75247 89200 75345 89298
rect 67973 88778 68071 88876
rect 67438 88489 68606 88549
rect 70977 87784 71075 87882
rect 75247 87784 75345 87882
rect 67973 87364 68071 87462
rect 3861 86388 3959 86486
rect 70977 86370 71075 86468
rect 18040 86196 18138 86294
rect 19288 86196 19386 86294
rect 20536 86196 20634 86294
rect 21784 86196 21882 86294
rect 23032 86196 23130 86294
rect 24280 86196 24378 86294
rect 25528 86196 25626 86294
rect 26776 86196 26874 86294
rect 28024 86196 28122 86294
rect 29272 86196 29370 86294
rect 30520 86196 30618 86294
rect 31768 86196 31866 86294
rect 33016 86196 33114 86294
rect 34264 86196 34362 86294
rect 35512 86196 35610 86294
rect 36760 86196 36858 86294
rect 38008 86196 38106 86294
rect 39256 86196 39354 86294
rect 40504 86196 40602 86294
rect 41752 86196 41850 86294
rect 43000 86196 43098 86294
rect 44248 86196 44346 86294
rect 45496 86196 45594 86294
rect 46744 86196 46842 86294
rect 47992 86196 48090 86294
rect 49240 86196 49338 86294
rect 50488 86196 50586 86294
rect 51736 86196 51834 86294
rect 52984 86196 53082 86294
rect 54232 86196 54330 86294
rect 55480 86196 55578 86294
rect 56728 86196 56826 86294
rect 18040 85874 18138 85972
rect 19288 85874 19386 85972
rect 20536 85874 20634 85972
rect 21784 85874 21882 85972
rect 23032 85874 23130 85972
rect 24280 85874 24378 85972
rect 25528 85874 25626 85972
rect 26776 85874 26874 85972
rect 28024 85874 28122 85972
rect 29272 85874 29370 85972
rect 30520 85874 30618 85972
rect 31768 85874 31866 85972
rect 33016 85874 33114 85972
rect 34264 85874 34362 85972
rect 35512 85874 35610 85972
rect 36760 85874 36858 85972
rect 38008 85874 38106 85972
rect 39256 85874 39354 85972
rect 40504 85874 40602 85972
rect 41752 85874 41850 85972
rect 43000 85874 43098 85972
rect 44248 85874 44346 85972
rect 45496 85874 45594 85972
rect 46744 85874 46842 85972
rect 47992 85874 48090 85972
rect 49240 85874 49338 85972
rect 50488 85874 50586 85972
rect 51736 85874 51834 85972
rect 52984 85874 53082 85972
rect 54232 85874 54330 85972
rect 55480 85874 55578 85972
rect 56728 85874 56826 85972
rect 64029 85150 64127 85248
rect 3861 84974 3959 85072
rect 18028 85036 18126 85134
rect 19276 85036 19374 85134
rect 20524 85036 20622 85134
rect 21772 85036 21870 85134
rect 23020 85036 23118 85134
rect 24268 85036 24366 85134
rect 25516 85036 25614 85134
rect 26764 85036 26862 85134
rect 28012 85036 28110 85134
rect 29260 85036 29358 85134
rect 30508 85036 30606 85134
rect 31756 85036 31854 85134
rect 33004 85036 33102 85134
rect 34252 85036 34350 85134
rect 35500 85036 35598 85134
rect 36748 85036 36846 85134
rect 37996 85036 38094 85134
rect 39244 85036 39342 85134
rect 40492 85036 40590 85134
rect 41740 85036 41838 85134
rect 42988 85036 43086 85134
rect 44236 85036 44334 85134
rect 45484 85036 45582 85134
rect 46732 85036 46830 85134
rect 47980 85036 48078 85134
rect 49228 85036 49326 85134
rect 50476 85036 50574 85134
rect 51724 85036 51822 85134
rect 52972 85036 53070 85134
rect 54220 85036 54318 85134
rect 55468 85036 55566 85134
rect 56716 85036 56814 85134
rect 70977 84956 71075 85054
rect 18110 84262 18208 84360
rect 19358 84262 19456 84360
rect 20606 84262 20704 84360
rect 21854 84262 21952 84360
rect 23102 84262 23200 84360
rect 24350 84262 24448 84360
rect 25598 84262 25696 84360
rect 26846 84262 26944 84360
rect 28094 84262 28192 84360
rect 29342 84262 29440 84360
rect 30590 84262 30688 84360
rect 31838 84262 31936 84360
rect 33086 84262 33184 84360
rect 34334 84262 34432 84360
rect 35582 84262 35680 84360
rect 36830 84262 36928 84360
rect 38078 84262 38176 84360
rect 39326 84262 39424 84360
rect 40574 84262 40672 84360
rect 41822 84262 41920 84360
rect 43070 84262 43168 84360
rect 44318 84262 44416 84360
rect 45566 84262 45664 84360
rect 46814 84262 46912 84360
rect 48062 84262 48160 84360
rect 49310 84262 49408 84360
rect 50558 84262 50656 84360
rect 51806 84262 51904 84360
rect 53054 84262 53152 84360
rect 54302 84262 54400 84360
rect 55550 84262 55648 84360
rect 56798 84262 56896 84360
rect 17708 84129 57644 84189
rect 64029 83736 64127 83834
rect 3861 83560 3959 83658
rect 70977 83542 71075 83640
rect 17708 83413 57644 83473
rect 17708 83289 57644 83349
rect 18283 82489 18381 82587
rect 19531 82489 19629 82587
rect 20779 82489 20877 82587
rect 22027 82489 22125 82587
rect 23275 82489 23373 82587
rect 24523 82489 24621 82587
rect 25771 82489 25869 82587
rect 27019 82489 27117 82587
rect 28267 82489 28365 82587
rect 29515 82489 29613 82587
rect 30763 82489 30861 82587
rect 32011 82489 32109 82587
rect 33259 82489 33357 82587
rect 34507 82489 34605 82587
rect 35755 82489 35853 82587
rect 37003 82489 37101 82587
rect 38251 82489 38349 82587
rect 39499 82489 39597 82587
rect 40747 82489 40845 82587
rect 41995 82489 42093 82587
rect 43243 82489 43341 82587
rect 44491 82489 44589 82587
rect 45739 82489 45837 82587
rect 46987 82489 47085 82587
rect 48235 82489 48333 82587
rect 49483 82489 49581 82587
rect 50731 82489 50829 82587
rect 51979 82489 52077 82587
rect 53227 82489 53325 82587
rect 54475 82489 54573 82587
rect 55723 82489 55821 82587
rect 56971 82489 57069 82587
rect 64029 82322 64127 82420
rect 3861 82146 3959 82244
rect 70977 82128 71075 82226
rect 17708 81554 58268 81614
rect 17852 80916 17950 81014
rect 18714 80916 18812 81014
rect 19100 80916 19198 81014
rect 19962 80916 20060 81014
rect 20348 80916 20446 81014
rect 21210 80916 21308 81014
rect 21596 80916 21694 81014
rect 22458 80916 22556 81014
rect 22844 80916 22942 81014
rect 23706 80916 23804 81014
rect 24092 80916 24190 81014
rect 24954 80916 25052 81014
rect 25340 80916 25438 81014
rect 26202 80916 26300 81014
rect 26588 80916 26686 81014
rect 27450 80916 27548 81014
rect 27836 80916 27934 81014
rect 28698 80916 28796 81014
rect 29084 80916 29182 81014
rect 29946 80916 30044 81014
rect 30332 80916 30430 81014
rect 31194 80916 31292 81014
rect 31580 80916 31678 81014
rect 32442 80916 32540 81014
rect 32828 80916 32926 81014
rect 33690 80916 33788 81014
rect 34076 80916 34174 81014
rect 34938 80916 35036 81014
rect 35324 80916 35422 81014
rect 36186 80916 36284 81014
rect 36572 80916 36670 81014
rect 37434 80916 37532 81014
rect 37820 80916 37918 81014
rect 38682 80916 38780 81014
rect 39068 80916 39166 81014
rect 39930 80916 40028 81014
rect 40316 80916 40414 81014
rect 41178 80916 41276 81014
rect 41564 80916 41662 81014
rect 42426 80916 42524 81014
rect 42812 80916 42910 81014
rect 43674 80916 43772 81014
rect 44060 80916 44158 81014
rect 44922 80916 45020 81014
rect 45308 80916 45406 81014
rect 46170 80916 46268 81014
rect 46556 80916 46654 81014
rect 47418 80916 47516 81014
rect 47804 80916 47902 81014
rect 48666 80916 48764 81014
rect 49052 80916 49150 81014
rect 49914 80916 50012 81014
rect 50300 80916 50398 81014
rect 51162 80916 51260 81014
rect 51548 80916 51646 81014
rect 52410 80916 52508 81014
rect 52796 80916 52894 81014
rect 53658 80916 53756 81014
rect 54044 80916 54142 81014
rect 54906 80916 55004 81014
rect 55292 80916 55390 81014
rect 56154 80916 56252 81014
rect 56540 80916 56638 81014
rect 57402 80916 57500 81014
rect 57788 80916 57886 81014
rect 3861 80732 3959 80830
rect 70977 80714 71075 80812
rect 74063 80554 74161 80652
rect 74799 80554 74897 80652
rect 17347 80325 17445 80423
rect 17971 80325 18069 80423
rect 18595 80325 18693 80423
rect 19219 80325 19317 80423
rect 19843 80325 19941 80423
rect 20467 80325 20565 80423
rect 21091 80325 21189 80423
rect 21715 80325 21813 80423
rect 22339 80325 22437 80423
rect 22963 80325 23061 80423
rect 23587 80325 23685 80423
rect 24211 80325 24309 80423
rect 24835 80325 24933 80423
rect 25459 80325 25557 80423
rect 26083 80325 26181 80423
rect 26707 80325 26805 80423
rect 27331 80325 27429 80423
rect 27955 80325 28053 80423
rect 28579 80325 28677 80423
rect 29203 80325 29301 80423
rect 29827 80325 29925 80423
rect 30451 80325 30549 80423
rect 31075 80325 31173 80423
rect 31699 80325 31797 80423
rect 32323 80325 32421 80423
rect 32947 80325 33045 80423
rect 33571 80325 33669 80423
rect 34195 80325 34293 80423
rect 34819 80325 34917 80423
rect 35443 80325 35541 80423
rect 36067 80325 36165 80423
rect 36691 80325 36789 80423
rect 37315 80325 37413 80423
rect 37939 80325 38037 80423
rect 38563 80325 38661 80423
rect 39187 80325 39285 80423
rect 39811 80325 39909 80423
rect 40435 80325 40533 80423
rect 41059 80325 41157 80423
rect 41683 80325 41781 80423
rect 42307 80325 42405 80423
rect 42931 80325 43029 80423
rect 43555 80325 43653 80423
rect 44179 80325 44277 80423
rect 44803 80325 44901 80423
rect 45427 80325 45525 80423
rect 46051 80325 46149 80423
rect 46675 80325 46773 80423
rect 47299 80325 47397 80423
rect 47923 80325 48021 80423
rect 48547 80325 48645 80423
rect 49171 80325 49269 80423
rect 49795 80325 49893 80423
rect 50419 80325 50517 80423
rect 51043 80325 51141 80423
rect 51667 80325 51765 80423
rect 52291 80325 52389 80423
rect 52915 80325 53013 80423
rect 53539 80325 53637 80423
rect 54163 80325 54261 80423
rect 54787 80325 54885 80423
rect 55411 80325 55509 80423
rect 56035 80325 56133 80423
rect 56659 80325 56757 80423
rect 57283 80325 57381 80423
rect 57907 80325 58005 80423
rect 16651 80001 16749 80099
rect 58603 80001 58701 80099
rect 16651 79764 16749 79862
rect 58603 79764 58701 79862
rect 16651 79527 16749 79625
rect 58603 79527 58701 79625
rect 10438 79421 10536 79519
rect 10863 79421 10961 79519
rect 11295 79421 11393 79519
rect 3861 79318 3959 79416
rect 11677 79398 11775 79496
rect 11949 79398 12047 79496
rect 63305 79398 63403 79496
rect 63577 79398 63675 79496
rect 63959 79421 64057 79519
rect 64391 79421 64489 79519
rect 64816 79421 64914 79519
rect 74063 79434 74161 79532
rect 74799 79434 74897 79532
rect 16651 79211 16749 79309
rect 58603 79211 58701 79309
rect 10438 79047 10536 79145
rect 10863 78989 10961 79087
rect 11295 78989 11393 79087
rect 11677 79003 11775 79101
rect 11949 79003 12047 79101
rect 16651 78974 16749 79072
rect 58603 78974 58701 79072
rect 63305 79003 63403 79101
rect 63577 79003 63675 79101
rect 63959 78989 64057 79087
rect 64391 78989 64489 79087
rect 64816 79047 64914 79145
rect 16651 78737 16749 78835
rect 58603 78737 58701 78835
rect 10438 78631 10536 78729
rect 10863 78631 10961 78729
rect 11295 78631 11393 78729
rect 11677 78608 11775 78706
rect 11949 78608 12047 78706
rect 63305 78608 63403 78706
rect 63577 78608 63675 78706
rect 63959 78631 64057 78729
rect 64391 78631 64489 78729
rect 64816 78631 64914 78729
rect 16651 78421 16749 78519
rect 58603 78421 58701 78519
rect 10438 78257 10536 78355
rect 10863 78199 10961 78297
rect 11295 78199 11393 78297
rect 11677 78213 11775 78311
rect 11949 78213 12047 78311
rect 16651 78184 16749 78282
rect 58603 78184 58701 78282
rect 63305 78213 63403 78311
rect 63577 78213 63675 78311
rect 63959 78199 64057 78297
rect 64391 78199 64489 78297
rect 64816 78257 64914 78355
rect 74063 78314 74161 78412
rect 74799 78314 74897 78412
rect 3861 77904 3959 78002
rect 10438 77841 10536 77939
rect 10863 77841 10961 77939
rect 11295 77841 11393 77939
rect 16651 77947 16749 78045
rect 58603 77947 58701 78045
rect 11677 77818 11775 77916
rect 11949 77818 12047 77916
rect 63305 77818 63403 77916
rect 63577 77818 63675 77916
rect 63959 77841 64057 77939
rect 64391 77841 64489 77939
rect 64816 77841 64914 77939
rect 16651 77631 16749 77729
rect 58603 77631 58701 77729
rect 10438 77467 10536 77565
rect 10863 77409 10961 77507
rect 11295 77409 11393 77507
rect 11677 77423 11775 77521
rect 11949 77423 12047 77521
rect 16651 77394 16749 77492
rect 58603 77394 58701 77492
rect 63305 77423 63403 77521
rect 63577 77423 63675 77521
rect 63959 77409 64057 77507
rect 64391 77409 64489 77507
rect 64816 77467 64914 77565
rect 10438 77051 10536 77149
rect 10863 77051 10961 77149
rect 11295 77051 11393 77149
rect 11677 77028 11775 77126
rect 11949 77028 12047 77126
rect 16651 77157 16749 77255
rect 58603 77157 58701 77255
rect 74063 77194 74161 77292
rect 74799 77194 74897 77292
rect 63305 77028 63403 77126
rect 63577 77028 63675 77126
rect 63959 77051 64057 77149
rect 64391 77051 64489 77149
rect 64816 77051 64914 77149
rect 3326 76817 4494 76877
rect 16651 76841 16749 76939
rect 58603 76841 58701 76939
rect 10438 76677 10536 76775
rect 3861 76490 3959 76588
rect 10863 76619 10961 76717
rect 11295 76619 11393 76717
rect 11677 76633 11775 76731
rect 11949 76633 12047 76731
rect 16651 76604 16749 76702
rect 58603 76604 58701 76702
rect 63305 76633 63403 76731
rect 63577 76633 63675 76731
rect 63959 76619 64057 76717
rect 64391 76619 64489 76717
rect 64816 76677 64914 76775
rect 10438 76261 10536 76359
rect 10863 76261 10961 76359
rect 11295 76261 11393 76359
rect 11677 76238 11775 76336
rect 11949 76238 12047 76336
rect 16651 76367 16749 76465
rect 58603 76367 58701 76465
rect 63305 76238 63403 76336
rect 63577 76238 63675 76336
rect 63959 76261 64057 76359
rect 64391 76261 64489 76359
rect 64816 76261 64914 76359
rect 16651 76051 16749 76149
rect 58603 76051 58701 76149
rect 74063 76074 74161 76172
rect 74799 76074 74897 76172
rect 10438 75887 10536 75985
rect 10863 75829 10961 75927
rect 11295 75829 11393 75927
rect 11677 75843 11775 75941
rect 11949 75843 12047 75941
rect 16651 75814 16749 75912
rect 58603 75814 58701 75912
rect 63305 75843 63403 75941
rect 63577 75843 63675 75941
rect 63959 75829 64057 75927
rect 64391 75829 64489 75927
rect 64816 75887 64914 75985
rect 16651 75577 16749 75675
rect 58603 75577 58701 75675
rect 10438 75471 10536 75569
rect 10863 75471 10961 75569
rect 11295 75471 11393 75569
rect 11677 75448 11775 75546
rect 11949 75448 12047 75546
rect 63305 75448 63403 75546
rect 63577 75448 63675 75546
rect 63959 75471 64057 75569
rect 64391 75471 64489 75569
rect 64816 75471 64914 75569
rect 16651 75261 16749 75359
rect 58603 75261 58701 75359
rect 10438 75097 10536 75195
rect 10863 75039 10961 75137
rect 11295 75039 11393 75137
rect 11677 75053 11775 75151
rect 11949 75053 12047 75151
rect 16651 75024 16749 75122
rect 58603 75024 58701 75122
rect 63305 75053 63403 75151
rect 63577 75053 63675 75151
rect 63959 75039 64057 75137
rect 64391 75039 64489 75137
rect 64816 75097 64914 75195
rect 74063 74954 74161 75052
rect 74799 74954 74897 75052
rect 16651 74787 16749 74885
rect 58603 74787 58701 74885
rect 10438 74681 10536 74779
rect 10863 74681 10961 74779
rect 11295 74681 11393 74779
rect 11677 74658 11775 74756
rect 11949 74658 12047 74756
rect 63305 74658 63403 74756
rect 63577 74658 63675 74756
rect 63959 74681 64057 74779
rect 64391 74681 64489 74779
rect 64816 74681 64914 74779
rect 16651 74471 16749 74569
rect 58603 74471 58701 74569
rect 10438 74307 10536 74405
rect 10863 74249 10961 74347
rect 11295 74249 11393 74347
rect 11677 74263 11775 74361
rect 11949 74263 12047 74361
rect 16651 74234 16749 74332
rect 58603 74234 58701 74332
rect 63305 74263 63403 74361
rect 63577 74263 63675 74361
rect 63959 74249 64057 74347
rect 64391 74249 64489 74347
rect 64816 74307 64914 74405
rect 16651 73997 16749 74095
rect 58603 73997 58701 74095
rect 10438 73891 10536 73989
rect 10863 73891 10961 73989
rect 11295 73891 11393 73989
rect 11677 73868 11775 73966
rect 11949 73868 12047 73966
rect 63305 73868 63403 73966
rect 63577 73868 63675 73966
rect 63959 73891 64057 73989
rect 64391 73891 64489 73989
rect 64816 73891 64914 73989
rect 74063 73834 74161 73932
rect 74799 73834 74897 73932
rect 16651 73681 16749 73779
rect 58603 73681 58701 73779
rect 10438 73517 10536 73615
rect 10863 73459 10961 73557
rect 11295 73459 11393 73557
rect 11677 73473 11775 73571
rect 11949 73473 12047 73571
rect 16651 73444 16749 73542
rect 58603 73444 58701 73542
rect 63305 73473 63403 73571
rect 63577 73473 63675 73571
rect 63959 73459 64057 73557
rect 64391 73459 64489 73557
rect 64816 73517 64914 73615
rect 16651 73207 16749 73305
rect 58603 73207 58701 73305
rect 10438 73101 10536 73199
rect 10863 73101 10961 73199
rect 11295 73101 11393 73199
rect 11677 73078 11775 73176
rect 11949 73078 12047 73176
rect 63305 73078 63403 73176
rect 63577 73078 63675 73176
rect 63959 73101 64057 73199
rect 64391 73101 64489 73199
rect 64816 73101 64914 73199
rect 16651 72891 16749 72989
rect 58603 72891 58701 72989
rect 10438 72727 10536 72825
rect 10863 72669 10961 72767
rect 11295 72669 11393 72767
rect 11677 72683 11775 72781
rect 11949 72683 12047 72781
rect 16651 72654 16749 72752
rect 58603 72654 58701 72752
rect 63305 72683 63403 72781
rect 63577 72683 63675 72781
rect 63959 72669 64057 72767
rect 64391 72669 64489 72767
rect 64816 72727 64914 72825
rect 74063 72714 74161 72812
rect 74799 72714 74897 72812
rect 16651 72417 16749 72515
rect 58603 72417 58701 72515
rect 10438 72311 10536 72409
rect 10863 72311 10961 72409
rect 11295 72311 11393 72409
rect 11677 72288 11775 72386
rect 11949 72288 12047 72386
rect 63305 72288 63403 72386
rect 63577 72288 63675 72386
rect 63959 72311 64057 72409
rect 64391 72311 64489 72409
rect 64816 72311 64914 72409
rect 16651 72101 16749 72199
rect 58603 72101 58701 72199
rect 10438 71937 10536 72035
rect 10863 71879 10961 71977
rect 11295 71879 11393 71977
rect 11677 71893 11775 71991
rect 11949 71893 12047 71991
rect 16651 71864 16749 71962
rect 58603 71864 58701 71962
rect 63305 71893 63403 71991
rect 63577 71893 63675 71991
rect 63959 71879 64057 71977
rect 64391 71879 64489 71977
rect 64816 71937 64914 72035
rect 16651 71627 16749 71725
rect 58603 71627 58701 71725
rect 10438 71521 10536 71619
rect 10863 71521 10961 71619
rect 11295 71521 11393 71619
rect 11677 71498 11775 71596
rect 11949 71498 12047 71596
rect 63305 71498 63403 71596
rect 63577 71498 63675 71596
rect 63959 71521 64057 71619
rect 64391 71521 64489 71619
rect 64816 71521 64914 71619
rect 74063 71594 74161 71692
rect 74799 71594 74897 71692
rect 16651 71311 16749 71409
rect 58603 71311 58701 71409
rect 10438 71147 10536 71245
rect 10863 71089 10961 71187
rect 11295 71089 11393 71187
rect 11677 71103 11775 71201
rect 11949 71103 12047 71201
rect 16651 71074 16749 71172
rect 58603 71074 58701 71172
rect 63305 71103 63403 71201
rect 63577 71103 63675 71201
rect 63959 71089 64057 71187
rect 64391 71089 64489 71187
rect 64816 71147 64914 71245
rect 16651 70837 16749 70935
rect 58603 70837 58701 70935
rect 10438 70731 10536 70829
rect 10863 70731 10961 70829
rect 11295 70731 11393 70829
rect 11677 70708 11775 70806
rect 11949 70708 12047 70806
rect 63305 70708 63403 70806
rect 63577 70708 63675 70806
rect 63959 70731 64057 70829
rect 64391 70731 64489 70829
rect 64816 70731 64914 70829
rect 10438 70357 10536 70455
rect 16651 70521 16749 70619
rect 58603 70521 58701 70619
rect 74063 70474 74161 70572
rect 74799 70474 74897 70572
rect 10863 70299 10961 70397
rect 11295 70299 11393 70397
rect 11677 70313 11775 70411
rect 11949 70313 12047 70411
rect 16651 70284 16749 70382
rect 58603 70284 58701 70382
rect 63305 70313 63403 70411
rect 63577 70313 63675 70411
rect 63959 70299 64057 70397
rect 64391 70299 64489 70397
rect 64816 70357 64914 70455
rect 16651 70047 16749 70145
rect 58603 70047 58701 70145
rect 10438 69941 10536 70039
rect 10863 69941 10961 70039
rect 11295 69941 11393 70039
rect 11677 69918 11775 70016
rect 11949 69918 12047 70016
rect 63305 69918 63403 70016
rect 63577 69918 63675 70016
rect 63959 69941 64057 70039
rect 64391 69941 64489 70039
rect 64816 69941 64914 70039
rect 16651 69731 16749 69829
rect 58603 69731 58701 69829
rect 10438 69567 10536 69665
rect 10863 69509 10961 69607
rect 11295 69509 11393 69607
rect 11677 69523 11775 69621
rect 11949 69523 12047 69621
rect 16651 69494 16749 69592
rect 58603 69494 58701 69592
rect 63305 69523 63403 69621
rect 63577 69523 63675 69621
rect 63959 69509 64057 69607
rect 64391 69509 64489 69607
rect 64816 69567 64914 69665
rect 10438 69151 10536 69249
rect 10863 69151 10961 69249
rect 11295 69151 11393 69249
rect 11677 69128 11775 69226
rect 11949 69128 12047 69226
rect 16651 69257 16749 69355
rect 58603 69257 58701 69355
rect 63305 69128 63403 69226
rect 63577 69128 63675 69226
rect 63959 69151 64057 69249
rect 64391 69151 64489 69249
rect 64816 69151 64914 69249
rect 16651 68941 16749 69039
rect 58603 68941 58701 69039
rect 10438 68777 10536 68875
rect 10863 68719 10961 68817
rect 11295 68719 11393 68817
rect 11677 68733 11775 68831
rect 11949 68733 12047 68831
rect 16651 68704 16749 68802
rect 58603 68704 58701 68802
rect 63305 68733 63403 68831
rect 63577 68733 63675 68831
rect 63959 68719 64057 68817
rect 64391 68719 64489 68817
rect 64816 68777 64914 68875
rect 10438 68361 10536 68459
rect 10863 68361 10961 68459
rect 11295 68361 11393 68459
rect 11677 68338 11775 68436
rect 11949 68338 12047 68436
rect 16651 68467 16749 68565
rect 58603 68467 58701 68565
rect 63305 68338 63403 68436
rect 63577 68338 63675 68436
rect 63959 68361 64057 68459
rect 64391 68361 64489 68459
rect 64816 68361 64914 68459
rect 16651 68151 16749 68249
rect 58603 68151 58701 68249
rect 10438 67987 10536 68085
rect 10863 67929 10961 68027
rect 11295 67929 11393 68027
rect 11677 67943 11775 68041
rect 11949 67943 12047 68041
rect 16651 67914 16749 68012
rect 58603 67914 58701 68012
rect 63305 67943 63403 68041
rect 63577 67943 63675 68041
rect 63959 67929 64057 68027
rect 64391 67929 64489 68027
rect 64816 67987 64914 68085
rect 16651 67677 16749 67775
rect 58603 67677 58701 67775
rect 10438 67571 10536 67669
rect 10863 67571 10961 67669
rect 11295 67571 11393 67669
rect 11677 67548 11775 67646
rect 11949 67548 12047 67646
rect 63305 67548 63403 67646
rect 63577 67548 63675 67646
rect 63959 67571 64057 67669
rect 64391 67571 64489 67669
rect 64816 67571 64914 67669
rect 16651 67361 16749 67459
rect 58603 67361 58701 67459
rect 10438 67197 10536 67295
rect 10863 67139 10961 67237
rect 11295 67139 11393 67237
rect 11677 67153 11775 67251
rect 11949 67153 12047 67251
rect 16651 67124 16749 67222
rect 58603 67124 58701 67222
rect 63305 67153 63403 67251
rect 63577 67153 63675 67251
rect 63959 67139 64057 67237
rect 64391 67139 64489 67237
rect 64816 67197 64914 67295
rect 16651 66887 16749 66985
rect 58603 66887 58701 66985
rect 10438 66781 10536 66879
rect 10863 66781 10961 66879
rect 11295 66781 11393 66879
rect 11677 66758 11775 66856
rect 11949 66758 12047 66856
rect 63305 66758 63403 66856
rect 63577 66758 63675 66856
rect 63959 66781 64057 66879
rect 64391 66781 64489 66879
rect 64816 66781 64914 66879
rect 10438 66407 10536 66505
rect 16651 66571 16749 66669
rect 58603 66571 58701 66669
rect 10863 66349 10961 66447
rect 11295 66349 11393 66447
rect 11677 66363 11775 66461
rect 11949 66363 12047 66461
rect 16651 66334 16749 66432
rect 58603 66334 58701 66432
rect 63305 66363 63403 66461
rect 63577 66363 63675 66461
rect 63959 66349 64057 66447
rect 64391 66349 64489 66447
rect 64816 66407 64914 66505
rect 16651 66097 16749 66195
rect 58603 66097 58701 66195
rect 10438 65991 10536 66089
rect 10863 65991 10961 66089
rect 11295 65991 11393 66089
rect 11677 65968 11775 66066
rect 11949 65968 12047 66066
rect 63305 65968 63403 66066
rect 63577 65968 63675 66066
rect 63959 65991 64057 66089
rect 64391 65991 64489 66089
rect 64816 65991 64914 66089
rect 16651 65781 16749 65879
rect 58603 65781 58701 65879
rect 10438 65617 10536 65715
rect 10863 65559 10961 65657
rect 11295 65559 11393 65657
rect 11677 65573 11775 65671
rect 11949 65573 12047 65671
rect 16651 65544 16749 65642
rect 58603 65544 58701 65642
rect 63305 65573 63403 65671
rect 63577 65573 63675 65671
rect 63959 65559 64057 65657
rect 64391 65559 64489 65657
rect 64816 65617 64914 65715
rect 16651 65307 16749 65405
rect 58603 65307 58701 65405
rect 10438 65201 10536 65299
rect 10863 65201 10961 65299
rect 11295 65201 11393 65299
rect 11677 65178 11775 65276
rect 11949 65178 12047 65276
rect 63305 65178 63403 65276
rect 63577 65178 63675 65276
rect 63959 65201 64057 65299
rect 64391 65201 64489 65299
rect 64816 65201 64914 65299
rect 16651 64991 16749 65089
rect 58603 64991 58701 65089
rect 10438 64827 10536 64925
rect 10863 64769 10961 64867
rect 11295 64769 11393 64867
rect 11677 64783 11775 64881
rect 11949 64783 12047 64881
rect 16651 64754 16749 64852
rect 58603 64754 58701 64852
rect 63305 64783 63403 64881
rect 63577 64783 63675 64881
rect 63959 64769 64057 64867
rect 64391 64769 64489 64867
rect 64816 64827 64914 64925
rect 16651 64517 16749 64615
rect 58603 64517 58701 64615
rect 10438 64411 10536 64509
rect 10863 64411 10961 64509
rect 11295 64411 11393 64509
rect 11677 64388 11775 64486
rect 11949 64388 12047 64486
rect 63305 64388 63403 64486
rect 63577 64388 63675 64486
rect 63959 64411 64057 64509
rect 64391 64411 64489 64509
rect 64816 64411 64914 64509
rect 16651 64201 16749 64299
rect 58603 64201 58701 64299
rect 10438 64037 10536 64135
rect 10863 63979 10961 64077
rect 11295 63979 11393 64077
rect 11677 63993 11775 64091
rect 11949 63993 12047 64091
rect 16651 63964 16749 64062
rect 58603 63964 58701 64062
rect 63305 63993 63403 64091
rect 63577 63993 63675 64091
rect 63959 63979 64057 64077
rect 64391 63979 64489 64077
rect 64816 64037 64914 64135
rect 16651 63727 16749 63825
rect 58603 63727 58701 63825
rect 10438 63621 10536 63719
rect 10863 63621 10961 63719
rect 11295 63621 11393 63719
rect 11677 63598 11775 63696
rect 11949 63598 12047 63696
rect 63305 63598 63403 63696
rect 63577 63598 63675 63696
rect 63959 63621 64057 63719
rect 64391 63621 64489 63719
rect 64816 63621 64914 63719
rect 16651 63411 16749 63509
rect 58603 63411 58701 63509
rect 10438 63247 10536 63345
rect 10863 63189 10961 63287
rect 11295 63189 11393 63287
rect 11677 63203 11775 63301
rect 11949 63203 12047 63301
rect 16651 63174 16749 63272
rect 58603 63174 58701 63272
rect 63305 63203 63403 63301
rect 63577 63203 63675 63301
rect 63959 63189 64057 63287
rect 64391 63189 64489 63287
rect 64816 63247 64914 63345
rect 16651 62937 16749 63035
rect 58603 62937 58701 63035
rect 10438 62831 10536 62929
rect 10863 62831 10961 62929
rect 11295 62831 11393 62929
rect 11677 62808 11775 62906
rect 11949 62808 12047 62906
rect 63305 62808 63403 62906
rect 63577 62808 63675 62906
rect 63959 62831 64057 62929
rect 64391 62831 64489 62929
rect 64816 62831 64914 62929
rect 16651 62621 16749 62719
rect 58603 62621 58701 62719
rect 10438 62457 10536 62555
rect 10863 62399 10961 62497
rect 11295 62399 11393 62497
rect 11677 62413 11775 62511
rect 11949 62413 12047 62511
rect 16651 62384 16749 62482
rect 58603 62384 58701 62482
rect 63305 62413 63403 62511
rect 63577 62413 63675 62511
rect 63959 62399 64057 62497
rect 64391 62399 64489 62497
rect 64816 62457 64914 62555
rect 16651 62147 16749 62245
rect 58603 62147 58701 62245
rect 10438 62041 10536 62139
rect 10863 62041 10961 62139
rect 11295 62041 11393 62139
rect 11677 62018 11775 62116
rect 11949 62018 12047 62116
rect 63305 62018 63403 62116
rect 63577 62018 63675 62116
rect 63959 62041 64057 62139
rect 64391 62041 64489 62139
rect 64816 62041 64914 62139
rect 16651 61831 16749 61929
rect 58603 61831 58701 61929
rect 10438 61667 10536 61765
rect 10863 61609 10961 61707
rect 11295 61609 11393 61707
rect 11677 61623 11775 61721
rect 11949 61623 12047 61721
rect 16651 61594 16749 61692
rect 58603 61594 58701 61692
rect 63305 61623 63403 61721
rect 63577 61623 63675 61721
rect 63959 61609 64057 61707
rect 64391 61609 64489 61707
rect 64816 61667 64914 61765
rect 10438 61251 10536 61349
rect 10863 61251 10961 61349
rect 11295 61251 11393 61349
rect 16651 61357 16749 61455
rect 58603 61357 58701 61455
rect 11677 61228 11775 61326
rect 11949 61228 12047 61326
rect 63305 61228 63403 61326
rect 63577 61228 63675 61326
rect 63959 61251 64057 61349
rect 64391 61251 64489 61349
rect 64816 61251 64914 61349
rect 16651 61041 16749 61139
rect 58603 61041 58701 61139
rect 10438 60877 10536 60975
rect 10863 60819 10961 60917
rect 11295 60819 11393 60917
rect 11677 60833 11775 60931
rect 11949 60833 12047 60931
rect 16651 60804 16749 60902
rect 58603 60804 58701 60902
rect 63305 60833 63403 60931
rect 63577 60833 63675 60931
rect 63959 60819 64057 60917
rect 64391 60819 64489 60917
rect 64816 60877 64914 60975
rect 10438 60461 10536 60559
rect 10863 60461 10961 60559
rect 11295 60461 11393 60559
rect 11677 60438 11775 60536
rect 11949 60438 12047 60536
rect 16651 60567 16749 60665
rect 58603 60567 58701 60665
rect 63305 60438 63403 60536
rect 63577 60438 63675 60536
rect 63959 60461 64057 60559
rect 64391 60461 64489 60559
rect 64816 60461 64914 60559
rect 16651 60251 16749 60349
rect 58603 60251 58701 60349
rect 10438 60087 10536 60185
rect 10863 60029 10961 60127
rect 11295 60029 11393 60127
rect 11677 60043 11775 60141
rect 11949 60043 12047 60141
rect 16651 60014 16749 60112
rect 58603 60014 58701 60112
rect 63305 60043 63403 60141
rect 63577 60043 63675 60141
rect 63959 60029 64057 60127
rect 64391 60029 64489 60127
rect 64816 60087 64914 60185
rect 10438 59671 10536 59769
rect 10863 59671 10961 59769
rect 11295 59671 11393 59769
rect 11677 59648 11775 59746
rect 11949 59648 12047 59746
rect 16651 59777 16749 59875
rect 58603 59777 58701 59875
rect 63305 59648 63403 59746
rect 63577 59648 63675 59746
rect 63959 59671 64057 59769
rect 64391 59671 64489 59769
rect 64816 59671 64914 59769
rect 16651 59461 16749 59559
rect 58603 59461 58701 59559
rect 10438 59297 10536 59395
rect 10863 59239 10961 59337
rect 11295 59239 11393 59337
rect 11677 59253 11775 59351
rect 11949 59253 12047 59351
rect 16651 59224 16749 59322
rect 58603 59224 58701 59322
rect 63305 59253 63403 59351
rect 63577 59253 63675 59351
rect 63959 59239 64057 59337
rect 64391 59239 64489 59337
rect 64816 59297 64914 59395
rect 16651 58987 16749 59085
rect 58603 58987 58701 59085
rect 10438 58881 10536 58979
rect 10863 58881 10961 58979
rect 11295 58881 11393 58979
rect 11677 58858 11775 58956
rect 11949 58858 12047 58956
rect 63305 58858 63403 58956
rect 63577 58858 63675 58956
rect 63959 58881 64057 58979
rect 64391 58881 64489 58979
rect 64816 58881 64914 58979
rect 16651 58671 16749 58769
rect 58603 58671 58701 58769
rect 10438 58507 10536 58605
rect 10863 58449 10961 58547
rect 11295 58449 11393 58547
rect 11677 58463 11775 58561
rect 11949 58463 12047 58561
rect 16651 58434 16749 58532
rect 58603 58434 58701 58532
rect 63305 58463 63403 58561
rect 63577 58463 63675 58561
rect 63959 58449 64057 58547
rect 64391 58449 64489 58547
rect 64816 58507 64914 58605
rect 16651 58197 16749 58295
rect 58603 58197 58701 58295
rect 10438 58091 10536 58189
rect 10863 58091 10961 58189
rect 11295 58091 11393 58189
rect 11677 58068 11775 58166
rect 11949 58068 12047 58166
rect 63305 58068 63403 58166
rect 63577 58068 63675 58166
rect 63959 58091 64057 58189
rect 64391 58091 64489 58189
rect 64816 58091 64914 58189
rect 16651 57881 16749 57979
rect 58603 57881 58701 57979
rect 10438 57717 10536 57815
rect 10863 57659 10961 57757
rect 11295 57659 11393 57757
rect 11677 57673 11775 57771
rect 11949 57673 12047 57771
rect 16651 57644 16749 57742
rect 58603 57644 58701 57742
rect 63305 57673 63403 57771
rect 63577 57673 63675 57771
rect 63959 57659 64057 57757
rect 64391 57659 64489 57757
rect 64816 57717 64914 57815
rect 16651 57407 16749 57505
rect 58603 57407 58701 57505
rect 10438 57301 10536 57399
rect 10863 57301 10961 57399
rect 11295 57301 11393 57399
rect 11677 57278 11775 57376
rect 11949 57278 12047 57376
rect 63305 57278 63403 57376
rect 63577 57278 63675 57376
rect 63959 57301 64057 57399
rect 64391 57301 64489 57399
rect 64816 57301 64914 57399
rect 16651 57091 16749 57189
rect 58603 57091 58701 57189
rect 10438 56927 10536 57025
rect 10863 56869 10961 56967
rect 11295 56869 11393 56967
rect 11677 56883 11775 56981
rect 11949 56883 12047 56981
rect 16651 56854 16749 56952
rect 58603 56854 58701 56952
rect 63305 56883 63403 56981
rect 63577 56883 63675 56981
rect 63959 56869 64057 56967
rect 64391 56869 64489 56967
rect 64816 56927 64914 57025
rect 16651 56617 16749 56715
rect 58603 56617 58701 56715
rect 10438 56511 10536 56609
rect 10863 56511 10961 56609
rect 11295 56511 11393 56609
rect 11677 56488 11775 56586
rect 11949 56488 12047 56586
rect 63305 56488 63403 56586
rect 63577 56488 63675 56586
rect 63959 56511 64057 56609
rect 64391 56511 64489 56609
rect 64816 56511 64914 56609
rect 16651 56301 16749 56399
rect 58603 56301 58701 56399
rect 10438 56137 10536 56235
rect 10863 56079 10961 56177
rect 11295 56079 11393 56177
rect 11677 56093 11775 56191
rect 11949 56093 12047 56191
rect 16651 56064 16749 56162
rect 58603 56064 58701 56162
rect 63305 56093 63403 56191
rect 63577 56093 63675 56191
rect 63959 56079 64057 56177
rect 64391 56079 64489 56177
rect 64816 56137 64914 56235
rect 16651 55827 16749 55925
rect 58603 55827 58701 55925
rect 10438 55721 10536 55819
rect 10863 55721 10961 55819
rect 11295 55721 11393 55819
rect 11677 55698 11775 55796
rect 11949 55698 12047 55796
rect 63305 55698 63403 55796
rect 63577 55698 63675 55796
rect 63959 55721 64057 55819
rect 64391 55721 64489 55819
rect 64816 55721 64914 55819
rect 16651 55511 16749 55609
rect 58603 55511 58701 55609
rect 10438 55347 10536 55445
rect 10863 55289 10961 55387
rect 11295 55289 11393 55387
rect 11677 55303 11775 55401
rect 11949 55303 12047 55401
rect 16651 55274 16749 55372
rect 58603 55274 58701 55372
rect 63305 55303 63403 55401
rect 63577 55303 63675 55401
rect 63959 55289 64057 55387
rect 64391 55289 64489 55387
rect 64816 55347 64914 55445
rect 16651 55037 16749 55135
rect 58603 55037 58701 55135
rect 10438 54931 10536 55029
rect 10863 54931 10961 55029
rect 11295 54931 11393 55029
rect 11677 54908 11775 55006
rect 11949 54908 12047 55006
rect 63305 54908 63403 55006
rect 63577 54908 63675 55006
rect 63959 54931 64057 55029
rect 64391 54931 64489 55029
rect 64816 54931 64914 55029
rect 16651 54721 16749 54819
rect 58603 54721 58701 54819
rect 10438 54557 10536 54655
rect 10863 54499 10961 54597
rect 11295 54499 11393 54597
rect 11677 54513 11775 54611
rect 11949 54513 12047 54611
rect 12395 54469 12493 54567
rect 12820 54468 12918 54566
rect 13863 54484 13961 54582
rect 15387 54484 15485 54582
rect 16651 54484 16749 54582
rect 58603 54484 58701 54582
rect 59867 54484 59965 54582
rect 61391 54484 61489 54582
rect 62434 54468 62532 54566
rect 62859 54469 62957 54567
rect 63305 54513 63403 54611
rect 63577 54513 63675 54611
rect 63959 54499 64057 54597
rect 64391 54499 64489 54597
rect 64816 54557 64914 54655
rect 16651 54247 16749 54345
rect 58603 54247 58701 54345
rect 10438 54141 10536 54239
rect 10863 54141 10961 54239
rect 11295 54141 11393 54239
rect 11677 54118 11775 54216
rect 11949 54118 12047 54216
rect 63305 54118 63403 54216
rect 63577 54118 63675 54216
rect 63959 54141 64057 54239
rect 64391 54141 64489 54239
rect 64816 54141 64914 54239
rect 10438 53767 10536 53865
rect 16651 53931 16749 54029
rect 58603 53931 58701 54029
rect 10863 53709 10961 53807
rect 11295 53709 11393 53807
rect 11677 53723 11775 53821
rect 11949 53723 12047 53821
rect 16651 53694 16749 53792
rect 58603 53694 58701 53792
rect 63305 53723 63403 53821
rect 63577 53723 63675 53821
rect 63959 53709 64057 53807
rect 64391 53709 64489 53807
rect 64816 53767 64914 53865
rect 10438 53351 10536 53449
rect 10863 53351 10961 53449
rect 11295 53351 11393 53449
rect 16651 53457 16749 53555
rect 58603 53457 58701 53555
rect 11677 53328 11775 53426
rect 11949 53328 12047 53426
rect 63305 53328 63403 53426
rect 63577 53328 63675 53426
rect 63959 53351 64057 53449
rect 64391 53351 64489 53449
rect 64816 53351 64914 53449
rect 16651 53141 16749 53239
rect 58603 53141 58701 53239
rect 10438 52977 10536 53075
rect 10863 52919 10961 53017
rect 11295 52919 11393 53017
rect 11677 52933 11775 53031
rect 11949 52933 12047 53031
rect 16651 52904 16749 53002
rect 58603 52904 58701 53002
rect 63305 52933 63403 53031
rect 63577 52933 63675 53031
rect 63959 52919 64057 53017
rect 64391 52919 64489 53017
rect 64816 52977 64914 53075
rect 10438 52561 10536 52659
rect 10863 52561 10961 52659
rect 11295 52561 11393 52659
rect 11677 52538 11775 52636
rect 11949 52538 12047 52636
rect 16651 52667 16749 52765
rect 58603 52667 58701 52765
rect 63305 52538 63403 52636
rect 63577 52538 63675 52636
rect 63959 52561 64057 52659
rect 64391 52561 64489 52659
rect 64816 52561 64914 52659
rect 16651 52351 16749 52449
rect 58603 52351 58701 52449
rect 10438 52187 10536 52285
rect 10863 52129 10961 52227
rect 11295 52129 11393 52227
rect 11677 52143 11775 52241
rect 11949 52143 12047 52241
rect 16651 52114 16749 52212
rect 58603 52114 58701 52212
rect 63305 52143 63403 52241
rect 63577 52143 63675 52241
rect 63959 52129 64057 52227
rect 64391 52129 64489 52227
rect 64816 52187 64914 52285
rect 10438 51771 10536 51869
rect 10863 51771 10961 51869
rect 11295 51771 11393 51869
rect 11677 51748 11775 51846
rect 11949 51748 12047 51846
rect 16651 51877 16749 51975
rect 58603 51877 58701 51975
rect 63305 51748 63403 51846
rect 63577 51748 63675 51846
rect 63959 51771 64057 51869
rect 64391 51771 64489 51869
rect 64816 51771 64914 51869
rect 16651 51561 16749 51659
rect 58603 51561 58701 51659
rect 10438 51397 10536 51495
rect 10863 51339 10961 51437
rect 11295 51339 11393 51437
rect 11677 51353 11775 51451
rect 11949 51353 12047 51451
rect 16651 51324 16749 51422
rect 58603 51324 58701 51422
rect 63305 51353 63403 51451
rect 63577 51353 63675 51451
rect 63959 51339 64057 51437
rect 64391 51339 64489 51437
rect 64816 51397 64914 51495
rect 16651 51087 16749 51185
rect 58603 51087 58701 51185
rect 10438 50981 10536 51079
rect 10863 50981 10961 51079
rect 11295 50981 11393 51079
rect 11677 50958 11775 51056
rect 11949 50958 12047 51056
rect 63305 50958 63403 51056
rect 63577 50958 63675 51056
rect 63959 50981 64057 51079
rect 64391 50981 64489 51079
rect 64816 50981 64914 51079
rect 16651 50771 16749 50869
rect 58603 50771 58701 50869
rect 10438 50607 10536 50705
rect 10863 50549 10961 50647
rect 11295 50549 11393 50647
rect 11677 50563 11775 50661
rect 11949 50563 12047 50661
rect 16651 50534 16749 50632
rect 58603 50534 58701 50632
rect 63305 50563 63403 50661
rect 63577 50563 63675 50661
rect 63959 50549 64057 50647
rect 64391 50549 64489 50647
rect 64816 50607 64914 50705
rect 16651 50297 16749 50395
rect 58603 50297 58701 50395
rect 10438 50191 10536 50289
rect 10863 50191 10961 50289
rect 11295 50191 11393 50289
rect 11677 50168 11775 50266
rect 11949 50168 12047 50266
rect 63305 50168 63403 50266
rect 63577 50168 63675 50266
rect 63959 50191 64057 50289
rect 64391 50191 64489 50289
rect 64816 50191 64914 50289
rect 10438 49817 10536 49915
rect 16651 49981 16749 50079
rect 58603 49981 58701 50079
rect 10863 49759 10961 49857
rect 11295 49759 11393 49857
rect 11677 49773 11775 49871
rect 11949 49773 12047 49871
rect 16651 49744 16749 49842
rect 58603 49744 58701 49842
rect 63305 49773 63403 49871
rect 63577 49773 63675 49871
rect 63959 49759 64057 49857
rect 64391 49759 64489 49857
rect 64816 49817 64914 49915
rect 16651 49507 16749 49605
rect 58603 49507 58701 49605
rect 10438 49401 10536 49499
rect 10863 49401 10961 49499
rect 11295 49401 11393 49499
rect 11677 49378 11775 49476
rect 11949 49378 12047 49476
rect 63305 49378 63403 49476
rect 63577 49378 63675 49476
rect 63959 49401 64057 49499
rect 64391 49401 64489 49499
rect 64816 49401 64914 49499
rect 16651 49191 16749 49289
rect 58603 49191 58701 49289
rect 10438 49027 10536 49125
rect 10863 48969 10961 49067
rect 11295 48969 11393 49067
rect 11677 48983 11775 49081
rect 11949 48983 12047 49081
rect 16651 48954 16749 49052
rect 58603 48954 58701 49052
rect 63305 48983 63403 49081
rect 63577 48983 63675 49081
rect 63959 48969 64057 49067
rect 64391 48969 64489 49067
rect 64816 49027 64914 49125
rect 16651 48717 16749 48815
rect 58603 48717 58701 48815
rect 10438 48611 10536 48709
rect 10863 48611 10961 48709
rect 11295 48611 11393 48709
rect 11677 48588 11775 48686
rect 11949 48588 12047 48686
rect 63305 48588 63403 48686
rect 63577 48588 63675 48686
rect 63959 48611 64057 48709
rect 64391 48611 64489 48709
rect 64816 48611 64914 48709
rect 16651 48401 16749 48499
rect 58603 48401 58701 48499
rect 10438 48237 10536 48335
rect 10863 48179 10961 48277
rect 11295 48179 11393 48277
rect 11677 48193 11775 48291
rect 11949 48193 12047 48291
rect 16651 48164 16749 48262
rect 58603 48164 58701 48262
rect 63305 48193 63403 48291
rect 63577 48193 63675 48291
rect 63959 48179 64057 48277
rect 64391 48179 64489 48277
rect 64816 48237 64914 48335
rect 16651 47927 16749 48025
rect 58603 47927 58701 48025
rect 10438 47821 10536 47919
rect 10863 47821 10961 47919
rect 11295 47821 11393 47919
rect 11677 47798 11775 47896
rect 11949 47798 12047 47896
rect 63305 47798 63403 47896
rect 63577 47798 63675 47896
rect 63959 47821 64057 47919
rect 64391 47821 64489 47919
rect 64816 47821 64914 47919
rect 16651 47611 16749 47709
rect 58603 47611 58701 47709
rect 10438 47447 10536 47545
rect 10863 47389 10961 47487
rect 11295 47389 11393 47487
rect 11677 47403 11775 47501
rect 11949 47403 12047 47501
rect 16651 47374 16749 47472
rect 58603 47374 58701 47472
rect 63305 47403 63403 47501
rect 63577 47403 63675 47501
rect 63959 47389 64057 47487
rect 64391 47389 64489 47487
rect 64816 47447 64914 47545
rect 16651 47137 16749 47235
rect 58603 47137 58701 47235
rect 10438 47031 10536 47129
rect 10863 47031 10961 47129
rect 11295 47031 11393 47129
rect 11677 47008 11775 47106
rect 11949 47008 12047 47106
rect 63305 47008 63403 47106
rect 63577 47008 63675 47106
rect 63959 47031 64057 47129
rect 64391 47031 64489 47129
rect 64816 47031 64914 47129
rect 16651 46821 16749 46919
rect 58603 46821 58701 46919
rect 10438 46657 10536 46755
rect 10863 46599 10961 46697
rect 11295 46599 11393 46697
rect 11677 46613 11775 46711
rect 11949 46613 12047 46711
rect 16651 46584 16749 46682
rect 58603 46584 58701 46682
rect 63305 46613 63403 46711
rect 63577 46613 63675 46711
rect 63959 46599 64057 46697
rect 64391 46599 64489 46697
rect 64816 46657 64914 46755
rect 16651 46347 16749 46445
rect 58603 46347 58701 46445
rect 10438 46241 10536 46339
rect 10863 46241 10961 46339
rect 11295 46241 11393 46339
rect 11677 46218 11775 46316
rect 11949 46218 12047 46316
rect 63305 46218 63403 46316
rect 63577 46218 63675 46316
rect 63959 46241 64057 46339
rect 64391 46241 64489 46339
rect 64816 46241 64914 46339
rect 16651 46031 16749 46129
rect 58603 46031 58701 46129
rect 10438 45867 10536 45965
rect 10863 45809 10961 45907
rect 11295 45809 11393 45907
rect 11677 45823 11775 45921
rect 11949 45823 12047 45921
rect 16651 45794 16749 45892
rect 58603 45794 58701 45892
rect 63305 45823 63403 45921
rect 63577 45823 63675 45921
rect 63959 45809 64057 45907
rect 64391 45809 64489 45907
rect 64816 45867 64914 45965
rect 16651 45557 16749 45655
rect 58603 45557 58701 45655
rect 10438 45451 10536 45549
rect 10863 45451 10961 45549
rect 11295 45451 11393 45549
rect 11677 45428 11775 45526
rect 11949 45428 12047 45526
rect 63305 45428 63403 45526
rect 63577 45428 63675 45526
rect 63959 45451 64057 45549
rect 64391 45451 64489 45549
rect 64816 45451 64914 45549
rect 16651 45241 16749 45339
rect 58603 45241 58701 45339
rect 10438 45077 10536 45175
rect 10863 45019 10961 45117
rect 11295 45019 11393 45117
rect 11677 45033 11775 45131
rect 11949 45033 12047 45131
rect 16651 45004 16749 45102
rect 58603 45004 58701 45102
rect 63305 45033 63403 45131
rect 63577 45033 63675 45131
rect 63959 45019 64057 45117
rect 64391 45019 64489 45117
rect 64816 45077 64914 45175
rect 10438 44661 10536 44759
rect 10863 44661 10961 44759
rect 11295 44661 11393 44759
rect 16651 44767 16749 44865
rect 58603 44767 58701 44865
rect 11677 44638 11775 44736
rect 11949 44638 12047 44736
rect 63305 44638 63403 44736
rect 63577 44638 63675 44736
rect 63959 44661 64057 44759
rect 64391 44661 64489 44759
rect 64816 44661 64914 44759
rect 16651 44451 16749 44549
rect 58603 44451 58701 44549
rect 10438 44287 10536 44385
rect 10863 44229 10961 44327
rect 11295 44229 11393 44327
rect 11677 44243 11775 44341
rect 11949 44243 12047 44341
rect 16651 44214 16749 44312
rect 58603 44214 58701 44312
rect 63305 44243 63403 44341
rect 63577 44243 63675 44341
rect 63959 44229 64057 44327
rect 64391 44229 64489 44327
rect 64816 44287 64914 44385
rect 10438 43871 10536 43969
rect 10863 43871 10961 43969
rect 11295 43871 11393 43969
rect 11677 43848 11775 43946
rect 11949 43848 12047 43946
rect 16651 43977 16749 44075
rect 58603 43977 58701 44075
rect 63305 43848 63403 43946
rect 63577 43848 63675 43946
rect 63959 43871 64057 43969
rect 64391 43871 64489 43969
rect 64816 43871 64914 43969
rect 16651 43661 16749 43759
rect 58603 43661 58701 43759
rect 10438 43497 10536 43595
rect 10863 43439 10961 43537
rect 11295 43439 11393 43537
rect 11677 43453 11775 43551
rect 11949 43453 12047 43551
rect 16651 43424 16749 43522
rect 58603 43424 58701 43522
rect 63305 43453 63403 43551
rect 63577 43453 63675 43551
rect 63959 43439 64057 43537
rect 64391 43439 64489 43537
rect 64816 43497 64914 43595
rect 10438 43081 10536 43179
rect 10863 43081 10961 43179
rect 11295 43081 11393 43179
rect 11677 43058 11775 43156
rect 11949 43058 12047 43156
rect 16651 43187 16749 43285
rect 58603 43187 58701 43285
rect 63305 43058 63403 43156
rect 63577 43058 63675 43156
rect 63959 43081 64057 43179
rect 64391 43081 64489 43179
rect 64816 43081 64914 43179
rect 16651 42871 16749 42969
rect 58603 42871 58701 42969
rect 10438 42707 10536 42805
rect 10863 42649 10961 42747
rect 11295 42649 11393 42747
rect 11677 42663 11775 42761
rect 11949 42663 12047 42761
rect 16651 42634 16749 42732
rect 58603 42634 58701 42732
rect 63305 42663 63403 42761
rect 63577 42663 63675 42761
rect 63959 42649 64057 42747
rect 64391 42649 64489 42747
rect 64816 42707 64914 42805
rect 16651 42397 16749 42495
rect 58603 42397 58701 42495
rect 10438 42291 10536 42389
rect 10863 42291 10961 42389
rect 11295 42291 11393 42389
rect 11677 42268 11775 42366
rect 11949 42268 12047 42366
rect 63305 42268 63403 42366
rect 63577 42268 63675 42366
rect 63959 42291 64057 42389
rect 64391 42291 64489 42389
rect 64816 42291 64914 42389
rect 16651 42081 16749 42179
rect 58603 42081 58701 42179
rect 10438 41917 10536 42015
rect 10863 41859 10961 41957
rect 11295 41859 11393 41957
rect 11677 41873 11775 41971
rect 11949 41873 12047 41971
rect 16651 41844 16749 41942
rect 58603 41844 58701 41942
rect 63305 41873 63403 41971
rect 63577 41873 63675 41971
rect 63959 41859 64057 41957
rect 64391 41859 64489 41957
rect 64816 41917 64914 42015
rect 16651 41607 16749 41705
rect 58603 41607 58701 41705
rect 10438 41501 10536 41599
rect 10863 41501 10961 41599
rect 11295 41501 11393 41599
rect 11677 41478 11775 41576
rect 11949 41478 12047 41576
rect 63305 41478 63403 41576
rect 63577 41478 63675 41576
rect 63959 41501 64057 41599
rect 64391 41501 64489 41599
rect 64816 41501 64914 41599
rect 16651 41291 16749 41389
rect 58603 41291 58701 41389
rect 10438 41127 10536 41225
rect 10863 41069 10961 41167
rect 11295 41069 11393 41167
rect 11677 41083 11775 41181
rect 11949 41083 12047 41181
rect 16651 41054 16749 41152
rect 58603 41054 58701 41152
rect 63305 41083 63403 41181
rect 63577 41083 63675 41181
rect 63959 41069 64057 41167
rect 64391 41069 64489 41167
rect 64816 41127 64914 41225
rect 16651 40817 16749 40915
rect 58603 40817 58701 40915
rect 10438 40711 10536 40809
rect 10863 40711 10961 40809
rect 11295 40711 11393 40809
rect 11677 40688 11775 40786
rect 11949 40688 12047 40786
rect 63305 40688 63403 40786
rect 63577 40688 63675 40786
rect 63959 40711 64057 40809
rect 64391 40711 64489 40809
rect 64816 40711 64914 40809
rect 16651 40501 16749 40599
rect 58603 40501 58701 40599
rect 10438 40337 10536 40435
rect 10863 40279 10961 40377
rect 11295 40279 11393 40377
rect 11677 40293 11775 40391
rect 11949 40293 12047 40391
rect 16651 40264 16749 40362
rect 58603 40264 58701 40362
rect 63305 40293 63403 40391
rect 63577 40293 63675 40391
rect 63959 40279 64057 40377
rect 64391 40279 64489 40377
rect 64816 40337 64914 40435
rect 16651 40027 16749 40125
rect 58603 40027 58701 40125
rect 10438 39921 10536 40019
rect 10863 39921 10961 40019
rect 11295 39921 11393 40019
rect 11677 39898 11775 39996
rect 11949 39898 12047 39996
rect 63305 39898 63403 39996
rect 63577 39898 63675 39996
rect 63959 39921 64057 40019
rect 64391 39921 64489 40019
rect 64816 39921 64914 40019
rect 16651 39711 16749 39809
rect 58603 39711 58701 39809
rect 10438 39547 10536 39645
rect 10863 39489 10961 39587
rect 11295 39489 11393 39587
rect 11677 39503 11775 39601
rect 11949 39503 12047 39601
rect 16651 39474 16749 39572
rect 58603 39474 58701 39572
rect 63305 39503 63403 39601
rect 63577 39503 63675 39601
rect 63959 39489 64057 39587
rect 64391 39489 64489 39587
rect 64816 39547 64914 39645
rect 16651 39237 16749 39335
rect 58603 39237 58701 39335
rect 10438 39131 10536 39229
rect 10863 39131 10961 39229
rect 11295 39131 11393 39229
rect 11677 39108 11775 39206
rect 11949 39108 12047 39206
rect 63305 39108 63403 39206
rect 63577 39108 63675 39206
rect 63959 39131 64057 39229
rect 64391 39131 64489 39229
rect 64816 39131 64914 39229
rect 16651 38921 16749 39019
rect 58603 38921 58701 39019
rect 10438 38757 10536 38855
rect 10863 38699 10961 38797
rect 11295 38699 11393 38797
rect 11677 38713 11775 38811
rect 11949 38713 12047 38811
rect 16651 38684 16749 38782
rect 58603 38684 58701 38782
rect 63305 38713 63403 38811
rect 63577 38713 63675 38811
rect 63959 38699 64057 38797
rect 64391 38699 64489 38797
rect 64816 38757 64914 38855
rect 455 38494 553 38592
rect 1191 38494 1289 38592
rect 16651 38447 16749 38545
rect 58603 38447 58701 38545
rect 10438 38341 10536 38439
rect 10863 38341 10961 38439
rect 11295 38341 11393 38439
rect 11677 38318 11775 38416
rect 11949 38318 12047 38416
rect 63305 38318 63403 38416
rect 63577 38318 63675 38416
rect 63959 38341 64057 38439
rect 64391 38341 64489 38439
rect 64816 38341 64914 38439
rect 16651 38131 16749 38229
rect 58603 38131 58701 38229
rect 10438 37967 10536 38065
rect 10863 37909 10961 38007
rect 11295 37909 11393 38007
rect 11677 37923 11775 38021
rect 11949 37923 12047 38021
rect 16651 37894 16749 37992
rect 58603 37894 58701 37992
rect 63305 37923 63403 38021
rect 63577 37923 63675 38021
rect 63959 37909 64057 38007
rect 64391 37909 64489 38007
rect 64816 37967 64914 38065
rect 16651 37657 16749 37755
rect 58603 37657 58701 37755
rect 10438 37551 10536 37649
rect 10863 37551 10961 37649
rect 11295 37551 11393 37649
rect 11677 37528 11775 37626
rect 11949 37528 12047 37626
rect 63305 37528 63403 37626
rect 63577 37528 63675 37626
rect 63959 37551 64057 37649
rect 64391 37551 64489 37649
rect 64816 37551 64914 37649
rect 455 37374 553 37472
rect 1191 37374 1289 37472
rect 16651 37341 16749 37439
rect 58603 37341 58701 37439
rect 10438 37177 10536 37275
rect 10863 37119 10961 37217
rect 11295 37119 11393 37217
rect 11677 37133 11775 37231
rect 11949 37133 12047 37231
rect 16651 37104 16749 37202
rect 58603 37104 58701 37202
rect 63305 37133 63403 37231
rect 63577 37133 63675 37231
rect 63959 37119 64057 37217
rect 64391 37119 64489 37217
rect 64816 37177 64914 37275
rect 7148 36761 7246 36859
rect 7573 36761 7671 36859
rect 8005 36761 8103 36859
rect 8387 36738 8485 36836
rect 8659 36738 8757 36836
rect 10438 36761 10536 36859
rect 10863 36761 10961 36859
rect 11295 36761 11393 36859
rect 16651 36867 16749 36965
rect 58603 36867 58701 36965
rect 11677 36738 11775 36836
rect 11949 36738 12047 36836
rect 63305 36738 63403 36836
rect 63577 36738 63675 36836
rect 63959 36761 64057 36859
rect 64391 36761 64489 36859
rect 64816 36761 64914 36859
rect 66595 36738 66693 36836
rect 66867 36738 66965 36836
rect 67249 36761 67347 36859
rect 67681 36761 67779 36859
rect 68106 36761 68204 36859
rect 16651 36551 16749 36649
rect 58603 36551 58701 36649
rect 10438 36387 10536 36485
rect 455 36254 553 36352
rect 1191 36254 1289 36352
rect 10863 36329 10961 36427
rect 11295 36329 11393 36427
rect 11677 36343 11775 36441
rect 11949 36343 12047 36441
rect 16651 36314 16749 36412
rect 58603 36314 58701 36412
rect 63305 36343 63403 36441
rect 63577 36343 63675 36441
rect 63959 36329 64057 36427
rect 64391 36329 64489 36427
rect 64816 36387 64914 36485
rect 7148 35971 7246 36069
rect 7573 35971 7671 36069
rect 8005 35971 8103 36069
rect 8387 35948 8485 36046
rect 8659 35948 8757 36046
rect 10438 35971 10536 36069
rect 10863 35971 10961 36069
rect 11295 35971 11393 36069
rect 11677 35948 11775 36046
rect 11949 35948 12047 36046
rect 16651 36077 16749 36175
rect 58603 36077 58701 36175
rect 63305 35948 63403 36046
rect 63577 35948 63675 36046
rect 63959 35971 64057 36069
rect 64391 35971 64489 36069
rect 64816 35971 64914 36069
rect 66595 35948 66693 36046
rect 66867 35948 66965 36046
rect 67249 35971 67347 36069
rect 67681 35971 67779 36069
rect 68106 35971 68204 36069
rect 16651 35761 16749 35859
rect 58603 35761 58701 35859
rect 10438 35597 10536 35695
rect 10863 35539 10961 35637
rect 11295 35539 11393 35637
rect 11677 35553 11775 35651
rect 11949 35553 12047 35651
rect 16651 35524 16749 35622
rect 58603 35524 58701 35622
rect 63305 35553 63403 35651
rect 63577 35553 63675 35651
rect 63959 35539 64057 35637
rect 64391 35539 64489 35637
rect 64816 35597 64914 35695
rect 455 35134 553 35232
rect 1191 35134 1289 35232
rect 7148 35181 7246 35279
rect 7573 35181 7671 35279
rect 8005 35181 8103 35279
rect 8387 35158 8485 35256
rect 8659 35158 8757 35256
rect 10438 35181 10536 35279
rect 10863 35181 10961 35279
rect 11295 35181 11393 35279
rect 11677 35158 11775 35256
rect 11949 35158 12047 35256
rect 16651 35287 16749 35385
rect 58603 35287 58701 35385
rect 63305 35158 63403 35256
rect 63577 35158 63675 35256
rect 63959 35181 64057 35279
rect 64391 35181 64489 35279
rect 64816 35181 64914 35279
rect 66595 35158 66693 35256
rect 66867 35158 66965 35256
rect 67249 35181 67347 35279
rect 67681 35181 67779 35279
rect 68106 35181 68204 35279
rect 16651 34971 16749 35069
rect 58603 34971 58701 35069
rect 10438 34807 10536 34905
rect 10863 34749 10961 34847
rect 11295 34749 11393 34847
rect 11677 34763 11775 34861
rect 11949 34763 12047 34861
rect 16651 34734 16749 34832
rect 58603 34734 58701 34832
rect 63305 34763 63403 34861
rect 63577 34763 63675 34861
rect 63959 34749 64057 34847
rect 64391 34749 64489 34847
rect 64816 34807 64914 34905
rect 16651 34497 16749 34595
rect 58603 34497 58701 34595
rect 5817 34368 5915 34466
rect 6089 34368 6187 34466
rect 7148 34391 7246 34489
rect 7573 34391 7671 34489
rect 8005 34391 8103 34489
rect 8387 34368 8485 34466
rect 8659 34368 8757 34466
rect 10438 34391 10536 34489
rect 10863 34391 10961 34489
rect 11295 34391 11393 34489
rect 11677 34368 11775 34466
rect 11949 34368 12047 34466
rect 63305 34368 63403 34466
rect 63577 34368 63675 34466
rect 63959 34391 64057 34489
rect 64391 34391 64489 34489
rect 64816 34391 64914 34489
rect 66595 34368 66693 34466
rect 66867 34368 66965 34466
rect 67249 34391 67347 34489
rect 67681 34391 67779 34489
rect 68106 34391 68204 34489
rect 69165 34368 69263 34466
rect 69437 34368 69535 34466
rect 16651 34181 16749 34279
rect 58603 34181 58701 34279
rect 455 34014 553 34112
rect 1191 34014 1289 34112
rect 10438 34017 10536 34115
rect 10863 33959 10961 34057
rect 11295 33959 11393 34057
rect 11677 33973 11775 34071
rect 11949 33973 12047 34071
rect 16651 33944 16749 34042
rect 58603 33944 58701 34042
rect 63305 33973 63403 34071
rect 63577 33973 63675 34071
rect 63959 33959 64057 34057
rect 64391 33959 64489 34057
rect 64816 34017 64914 34115
rect 16651 33707 16749 33805
rect 58603 33707 58701 33805
rect 10438 33601 10536 33699
rect 10863 33601 10961 33699
rect 11295 33601 11393 33699
rect 11677 33578 11775 33676
rect 11949 33578 12047 33676
rect 63305 33578 63403 33676
rect 63577 33578 63675 33676
rect 63959 33601 64057 33699
rect 64391 33601 64489 33699
rect 64816 33601 64914 33699
rect 10438 33227 10536 33325
rect 16651 33391 16749 33489
rect 58603 33391 58701 33489
rect 10863 33169 10961 33267
rect 11295 33169 11393 33267
rect 11677 33183 11775 33281
rect 11949 33183 12047 33281
rect 16651 33154 16749 33252
rect 58603 33154 58701 33252
rect 63305 33183 63403 33281
rect 63577 33183 63675 33281
rect 63959 33169 64057 33267
rect 64391 33169 64489 33267
rect 64816 33227 64914 33325
rect 455 32894 553 32992
rect 1191 32894 1289 32992
rect 16651 32917 16749 33015
rect 58603 32917 58701 33015
rect 7583 32795 7681 32893
rect 8008 32795 8106 32893
rect 8387 32788 8485 32886
rect 8659 32788 8757 32886
rect 10438 32811 10536 32909
rect 10863 32811 10961 32909
rect 11295 32811 11393 32909
rect 11677 32788 11775 32886
rect 11949 32788 12047 32886
rect 63305 32788 63403 32886
rect 63577 32788 63675 32886
rect 63959 32811 64057 32909
rect 64391 32811 64489 32909
rect 64816 32811 64914 32909
rect 66595 32788 66693 32886
rect 66867 32788 66965 32886
rect 67246 32795 67344 32893
rect 67671 32795 67769 32893
rect 16651 32601 16749 32699
rect 58603 32601 58701 32699
rect 10438 32437 10536 32535
rect 10863 32379 10961 32477
rect 11295 32379 11393 32477
rect 11677 32393 11775 32491
rect 11949 32393 12047 32491
rect 16651 32364 16749 32462
rect 58603 32364 58701 32462
rect 63305 32393 63403 32491
rect 63577 32393 63675 32491
rect 63959 32379 64057 32477
rect 64391 32379 64489 32477
rect 64816 32437 64914 32535
rect 16651 32127 16749 32225
rect 58603 32127 58701 32225
rect 6413 31998 6511 32096
rect 6685 31998 6783 32096
rect 7583 32005 7681 32103
rect 8008 32005 8106 32103
rect 8387 31998 8485 32096
rect 8659 31998 8757 32096
rect 10438 32021 10536 32119
rect 10863 32021 10961 32119
rect 11295 32021 11393 32119
rect 11677 31998 11775 32096
rect 11949 31998 12047 32096
rect 63305 31998 63403 32096
rect 63577 31998 63675 32096
rect 63959 32021 64057 32119
rect 64391 32021 64489 32119
rect 64816 32021 64914 32119
rect 66595 31998 66693 32096
rect 66867 31998 66965 32096
rect 67246 32005 67344 32103
rect 67671 32005 67769 32103
rect 68569 31998 68667 32096
rect 68841 31998 68939 32096
rect 455 31774 553 31872
rect 1191 31774 1289 31872
rect 16651 31811 16749 31909
rect 58603 31811 58701 31909
rect 10438 31647 10536 31745
rect 10863 31589 10961 31687
rect 11295 31589 11393 31687
rect 11677 31603 11775 31701
rect 11949 31603 12047 31701
rect 16651 31574 16749 31672
rect 58603 31574 58701 31672
rect 63305 31603 63403 31701
rect 63577 31603 63675 31701
rect 63959 31589 64057 31687
rect 64391 31589 64489 31687
rect 64816 31647 64914 31745
rect 16651 31337 16749 31435
rect 58603 31337 58701 31435
rect 10438 31231 10536 31329
rect 10863 31231 10961 31329
rect 11295 31231 11393 31329
rect 11677 31208 11775 31306
rect 11949 31208 12047 31306
rect 63305 31208 63403 31306
rect 63577 31208 63675 31306
rect 63959 31231 64057 31329
rect 64391 31231 64489 31329
rect 64816 31231 64914 31329
rect 16651 31021 16749 31119
rect 58603 31021 58701 31119
rect 10438 30857 10536 30955
rect 10863 30799 10961 30897
rect 11295 30799 11393 30897
rect 11677 30813 11775 30911
rect 11949 30813 12047 30911
rect 455 30654 553 30752
rect 1191 30654 1289 30752
rect 16651 30784 16749 30882
rect 58603 30784 58701 30882
rect 63305 30813 63403 30911
rect 63577 30813 63675 30911
rect 63959 30799 64057 30897
rect 64391 30799 64489 30897
rect 64816 30857 64914 30955
rect 16651 30547 16749 30645
rect 58603 30547 58701 30645
rect 7583 30425 7681 30523
rect 8008 30425 8106 30523
rect 8387 30418 8485 30516
rect 8659 30418 8757 30516
rect 10438 30441 10536 30539
rect 10863 30441 10961 30539
rect 11295 30441 11393 30539
rect 11677 30418 11775 30516
rect 11949 30418 12047 30516
rect 63305 30418 63403 30516
rect 63577 30418 63675 30516
rect 63959 30441 64057 30539
rect 64391 30441 64489 30539
rect 64816 30441 64914 30539
rect 66595 30418 66693 30516
rect 66867 30418 66965 30516
rect 67246 30425 67344 30523
rect 67671 30425 67769 30523
rect 16651 30231 16749 30329
rect 58603 30231 58701 30329
rect 10438 30067 10536 30165
rect 10863 30009 10961 30107
rect 11295 30009 11393 30107
rect 11677 30023 11775 30121
rect 11949 30023 12047 30121
rect 16651 29994 16749 30092
rect 58603 29994 58701 30092
rect 63305 30023 63403 30121
rect 63577 30023 63675 30121
rect 63959 30009 64057 30107
rect 64391 30009 64489 30107
rect 64816 30067 64914 30165
rect 16651 29757 16749 29855
rect 58603 29757 58701 29855
rect 455 29534 553 29632
rect 1191 29534 1289 29632
rect 6413 29628 6511 29726
rect 6685 29628 6783 29726
rect 7583 29635 7681 29733
rect 8008 29635 8106 29733
rect 8387 29628 8485 29726
rect 8659 29628 8757 29726
rect 10438 29651 10536 29749
rect 10863 29651 10961 29749
rect 11295 29651 11393 29749
rect 11677 29628 11775 29726
rect 11949 29628 12047 29726
rect 63305 29628 63403 29726
rect 63577 29628 63675 29726
rect 63959 29651 64057 29749
rect 64391 29651 64489 29749
rect 64816 29651 64914 29749
rect 66595 29628 66693 29726
rect 66867 29628 66965 29726
rect 67246 29635 67344 29733
rect 67671 29635 67769 29733
rect 68569 29628 68667 29726
rect 68841 29628 68939 29726
rect 16651 29441 16749 29539
rect 58603 29441 58701 29539
rect 16651 29204 16749 29302
rect 58603 29204 58701 29302
rect 16651 28967 16749 29065
rect 58603 28967 58701 29065
rect 71477 28927 71575 29025
rect 17347 28643 17445 28741
rect 17971 28643 18069 28741
rect 18595 28643 18693 28741
rect 19219 28643 19317 28741
rect 19843 28643 19941 28741
rect 20467 28643 20565 28741
rect 21091 28643 21189 28741
rect 21715 28643 21813 28741
rect 22339 28643 22437 28741
rect 22963 28643 23061 28741
rect 23587 28643 23685 28741
rect 24211 28643 24309 28741
rect 24835 28643 24933 28741
rect 25459 28643 25557 28741
rect 26083 28643 26181 28741
rect 26707 28643 26805 28741
rect 27331 28643 27429 28741
rect 27955 28643 28053 28741
rect 28579 28643 28677 28741
rect 29203 28643 29301 28741
rect 29827 28643 29925 28741
rect 30451 28643 30549 28741
rect 31075 28643 31173 28741
rect 31699 28643 31797 28741
rect 32323 28643 32421 28741
rect 32947 28643 33045 28741
rect 33571 28643 33669 28741
rect 34195 28643 34293 28741
rect 34819 28643 34917 28741
rect 35443 28643 35541 28741
rect 36067 28643 36165 28741
rect 36691 28643 36789 28741
rect 37315 28643 37413 28741
rect 37939 28643 38037 28741
rect 38563 28643 38661 28741
rect 39187 28643 39285 28741
rect 39811 28643 39909 28741
rect 40435 28643 40533 28741
rect 41059 28643 41157 28741
rect 41683 28643 41781 28741
rect 42307 28643 42405 28741
rect 42931 28643 43029 28741
rect 43555 28643 43653 28741
rect 44179 28643 44277 28741
rect 44803 28643 44901 28741
rect 45427 28643 45525 28741
rect 46051 28643 46149 28741
rect 46675 28643 46773 28741
rect 47299 28643 47397 28741
rect 47923 28643 48021 28741
rect 48547 28643 48645 28741
rect 49171 28643 49269 28741
rect 49795 28643 49893 28741
rect 50419 28643 50517 28741
rect 51043 28643 51141 28741
rect 51667 28643 51765 28741
rect 52291 28643 52389 28741
rect 52915 28643 53013 28741
rect 53539 28643 53637 28741
rect 54163 28643 54261 28741
rect 54787 28643 54885 28741
rect 55411 28643 55509 28741
rect 56035 28643 56133 28741
rect 56659 28643 56757 28741
rect 57283 28643 57381 28741
rect 57907 28643 58005 28741
rect 70942 28638 72110 28698
rect 455 28414 553 28512
rect 1191 28414 1289 28512
rect 4361 28254 4459 28352
rect 17466 28052 17564 28150
rect 17852 28052 17950 28150
rect 18714 28052 18812 28150
rect 19100 28052 19198 28150
rect 19962 28052 20060 28150
rect 20348 28052 20446 28150
rect 21210 28052 21308 28150
rect 21596 28052 21694 28150
rect 22458 28052 22556 28150
rect 22844 28052 22942 28150
rect 23706 28052 23804 28150
rect 24092 28052 24190 28150
rect 24954 28052 25052 28150
rect 25340 28052 25438 28150
rect 26202 28052 26300 28150
rect 26588 28052 26686 28150
rect 27450 28052 27548 28150
rect 27836 28052 27934 28150
rect 28698 28052 28796 28150
rect 29084 28052 29182 28150
rect 29946 28052 30044 28150
rect 30332 28052 30430 28150
rect 31194 28052 31292 28150
rect 31580 28052 31678 28150
rect 32442 28052 32540 28150
rect 32828 28052 32926 28150
rect 33690 28052 33788 28150
rect 34076 28052 34174 28150
rect 34938 28052 35036 28150
rect 35324 28052 35422 28150
rect 36186 28052 36284 28150
rect 36572 28052 36670 28150
rect 37434 28052 37532 28150
rect 37820 28052 37918 28150
rect 38682 28052 38780 28150
rect 39068 28052 39166 28150
rect 39930 28052 40028 28150
rect 40316 28052 40414 28150
rect 41178 28052 41276 28150
rect 41564 28052 41662 28150
rect 42426 28052 42524 28150
rect 42812 28052 42910 28150
rect 43674 28052 43772 28150
rect 44060 28052 44158 28150
rect 44922 28052 45020 28150
rect 45308 28052 45406 28150
rect 46170 28052 46268 28150
rect 46556 28052 46654 28150
rect 47418 28052 47516 28150
rect 47804 28052 47902 28150
rect 48666 28052 48764 28150
rect 49052 28052 49150 28150
rect 49914 28052 50012 28150
rect 50300 28052 50398 28150
rect 51162 28052 51260 28150
rect 51548 28052 51646 28150
rect 52410 28052 52508 28150
rect 52796 28052 52894 28150
rect 53658 28052 53756 28150
rect 54044 28052 54142 28150
rect 54906 28052 55004 28150
rect 55292 28052 55390 28150
rect 56154 28052 56252 28150
rect 56540 28052 56638 28150
rect 57402 28052 57500 28150
rect 17084 27452 57644 27512
rect 71477 27513 71575 27611
rect 4361 26840 4459 26938
rect 11101 26646 11199 26744
rect 18283 26479 18381 26577
rect 19531 26479 19629 26577
rect 20779 26479 20877 26577
rect 22027 26479 22125 26577
rect 23275 26479 23373 26577
rect 24523 26479 24621 26577
rect 25771 26479 25869 26577
rect 27019 26479 27117 26577
rect 28267 26479 28365 26577
rect 29515 26479 29613 26577
rect 30763 26479 30861 26577
rect 32011 26479 32109 26577
rect 33259 26479 33357 26577
rect 34507 26479 34605 26577
rect 35755 26479 35853 26577
rect 37003 26479 37101 26577
rect 38251 26479 38349 26577
rect 39499 26479 39597 26577
rect 40747 26479 40845 26577
rect 41995 26479 42093 26577
rect 43243 26479 43341 26577
rect 44491 26479 44589 26577
rect 45739 26479 45837 26577
rect 46987 26479 47085 26577
rect 48235 26479 48333 26577
rect 49483 26479 49581 26577
rect 50731 26479 50829 26577
rect 51979 26479 52077 26577
rect 53227 26479 53325 26577
rect 54475 26479 54573 26577
rect 55723 26479 55821 26577
rect 56971 26479 57069 26577
rect 71477 26099 71575 26197
rect 17708 25717 57644 25777
rect 17708 25593 57644 25653
rect 4361 25426 4459 25524
rect 11101 25232 11199 25330
rect 17708 24877 57644 24937
rect 18110 24706 18208 24804
rect 19358 24706 19456 24804
rect 20606 24706 20704 24804
rect 21854 24706 21952 24804
rect 23102 24706 23200 24804
rect 24350 24706 24448 24804
rect 25598 24706 25696 24804
rect 26846 24706 26944 24804
rect 28094 24706 28192 24804
rect 29342 24706 29440 24804
rect 30590 24706 30688 24804
rect 31838 24706 31936 24804
rect 33086 24706 33184 24804
rect 34334 24706 34432 24804
rect 35582 24706 35680 24804
rect 36830 24706 36928 24804
rect 38078 24706 38176 24804
rect 39326 24706 39424 24804
rect 40574 24706 40672 24804
rect 41822 24706 41920 24804
rect 43070 24706 43168 24804
rect 44318 24706 44416 24804
rect 45566 24706 45664 24804
rect 46814 24706 46912 24804
rect 48062 24706 48160 24804
rect 49310 24706 49408 24804
rect 50558 24706 50656 24804
rect 51806 24706 51904 24804
rect 53054 24706 53152 24804
rect 54302 24706 54400 24804
rect 55550 24706 55648 24804
rect 56798 24706 56896 24804
rect 71477 24685 71575 24783
rect 4361 24012 4459 24110
rect 18028 23932 18126 24030
rect 19276 23932 19374 24030
rect 20524 23932 20622 24030
rect 21772 23932 21870 24030
rect 23020 23932 23118 24030
rect 24268 23932 24366 24030
rect 25516 23932 25614 24030
rect 26764 23932 26862 24030
rect 28012 23932 28110 24030
rect 29260 23932 29358 24030
rect 30508 23932 30606 24030
rect 31756 23932 31854 24030
rect 33004 23932 33102 24030
rect 34252 23932 34350 24030
rect 35500 23932 35598 24030
rect 36748 23932 36846 24030
rect 37996 23932 38094 24030
rect 39244 23932 39342 24030
rect 40492 23932 40590 24030
rect 41740 23932 41838 24030
rect 42988 23932 43086 24030
rect 44236 23932 44334 24030
rect 45484 23932 45582 24030
rect 46732 23932 46830 24030
rect 47980 23932 48078 24030
rect 49228 23932 49326 24030
rect 50476 23932 50574 24030
rect 51724 23932 51822 24030
rect 52972 23932 53070 24030
rect 54220 23932 54318 24030
rect 55468 23932 55566 24030
rect 56716 23932 56814 24030
rect 11101 23818 11199 23916
rect 71477 23271 71575 23369
rect 18040 23094 18138 23192
rect 19288 23094 19386 23192
rect 20536 23094 20634 23192
rect 21784 23094 21882 23192
rect 23032 23094 23130 23192
rect 24280 23094 24378 23192
rect 25528 23094 25626 23192
rect 26776 23094 26874 23192
rect 28024 23094 28122 23192
rect 29272 23094 29370 23192
rect 30520 23094 30618 23192
rect 31768 23094 31866 23192
rect 33016 23094 33114 23192
rect 34264 23094 34362 23192
rect 35512 23094 35610 23192
rect 36760 23094 36858 23192
rect 38008 23094 38106 23192
rect 39256 23094 39354 23192
rect 40504 23094 40602 23192
rect 41752 23094 41850 23192
rect 43000 23094 43098 23192
rect 44248 23094 44346 23192
rect 45496 23094 45594 23192
rect 46744 23094 46842 23192
rect 47992 23094 48090 23192
rect 49240 23094 49338 23192
rect 50488 23094 50586 23192
rect 51736 23094 51834 23192
rect 52984 23094 53082 23192
rect 54232 23094 54330 23192
rect 55480 23094 55578 23192
rect 56728 23094 56826 23192
rect 18040 22772 18138 22870
rect 19288 22772 19386 22870
rect 20536 22772 20634 22870
rect 21784 22772 21882 22870
rect 23032 22772 23130 22870
rect 24280 22772 24378 22870
rect 25528 22772 25626 22870
rect 26776 22772 26874 22870
rect 28024 22772 28122 22870
rect 29272 22772 29370 22870
rect 30520 22772 30618 22870
rect 31768 22772 31866 22870
rect 33016 22772 33114 22870
rect 34264 22772 34362 22870
rect 35512 22772 35610 22870
rect 36760 22772 36858 22870
rect 38008 22772 38106 22870
rect 39256 22772 39354 22870
rect 40504 22772 40602 22870
rect 41752 22772 41850 22870
rect 43000 22772 43098 22870
rect 44248 22772 44346 22870
rect 45496 22772 45594 22870
rect 46744 22772 46842 22870
rect 47992 22772 48090 22870
rect 49240 22772 49338 22870
rect 50488 22772 50586 22870
rect 51736 22772 51834 22870
rect 52984 22772 53082 22870
rect 54232 22772 54330 22870
rect 55480 22772 55578 22870
rect 56728 22772 56826 22870
rect 4361 22598 4459 22696
rect 17926 21979 18024 22077
rect 19174 21979 19272 22077
rect 20422 21979 20520 22077
rect 21670 21979 21768 22077
rect 22918 21979 23016 22077
rect 24166 21979 24264 22077
rect 25414 21979 25512 22077
rect 26662 21979 26760 22077
rect 27910 21979 28008 22077
rect 29158 21979 29256 22077
rect 30406 21979 30504 22077
rect 31654 21979 31752 22077
rect 32902 21979 33000 22077
rect 34150 21979 34248 22077
rect 35398 21979 35496 22077
rect 36646 21979 36744 22077
rect 37894 21979 37992 22077
rect 39142 21979 39240 22077
rect 40390 21979 40488 22077
rect 41638 21979 41736 22077
rect 42886 21979 42984 22077
rect 44134 21979 44232 22077
rect 45382 21979 45480 22077
rect 46630 21979 46728 22077
rect 47878 21979 47976 22077
rect 49126 21979 49224 22077
rect 50374 21979 50472 22077
rect 51622 21979 51720 22077
rect 52870 21979 52968 22077
rect 54118 21979 54216 22077
rect 55366 21979 55464 22077
rect 56614 21979 56712 22077
rect 71477 21857 71575 21955
rect 17915 21542 18013 21640
rect 19163 21542 19261 21640
rect 20411 21542 20509 21640
rect 21659 21542 21757 21640
rect 22907 21542 23005 21640
rect 24155 21542 24253 21640
rect 25403 21542 25501 21640
rect 26651 21542 26749 21640
rect 27899 21542 27997 21640
rect 29147 21542 29245 21640
rect 30395 21542 30493 21640
rect 31643 21542 31741 21640
rect 32891 21542 32989 21640
rect 34139 21542 34237 21640
rect 35387 21542 35485 21640
rect 36635 21542 36733 21640
rect 37883 21542 37981 21640
rect 39131 21542 39229 21640
rect 40379 21542 40477 21640
rect 41627 21542 41725 21640
rect 42875 21542 42973 21640
rect 44123 21542 44221 21640
rect 45371 21542 45469 21640
rect 46619 21542 46717 21640
rect 47867 21542 47965 21640
rect 49115 21542 49213 21640
rect 50363 21542 50461 21640
rect 51611 21542 51709 21640
rect 52859 21542 52957 21640
rect 54107 21542 54205 21640
rect 55355 21542 55453 21640
rect 56603 21542 56701 21640
rect 4361 21184 4459 21282
rect 18036 21210 18134 21308
rect 19284 21210 19382 21308
rect 20532 21210 20630 21308
rect 21780 21210 21878 21308
rect 23028 21210 23126 21308
rect 24276 21210 24374 21308
rect 25524 21210 25622 21308
rect 26772 21210 26870 21308
rect 28020 21210 28118 21308
rect 29268 21210 29366 21308
rect 30516 21210 30614 21308
rect 31764 21210 31862 21308
rect 33012 21210 33110 21308
rect 34260 21210 34358 21308
rect 35508 21210 35606 21308
rect 36756 21210 36854 21308
rect 38004 21210 38102 21308
rect 39252 21210 39350 21308
rect 40500 21210 40598 21308
rect 41748 21210 41846 21308
rect 42996 21210 43094 21308
rect 44244 21210 44342 21308
rect 45492 21210 45590 21308
rect 46740 21210 46838 21308
rect 47988 21210 48086 21308
rect 49236 21210 49334 21308
rect 50484 21210 50582 21308
rect 51732 21210 51830 21308
rect 52980 21210 53078 21308
rect 54228 21210 54326 21308
rect 55476 21210 55574 21308
rect 56724 21210 56822 21308
rect 17921 21008 18019 21106
rect 19169 21008 19267 21106
rect 20417 21008 20515 21106
rect 21665 21008 21763 21106
rect 22913 21008 23011 21106
rect 24161 21008 24259 21106
rect 25409 21008 25507 21106
rect 26657 21008 26755 21106
rect 27905 21008 28003 21106
rect 29153 21008 29251 21106
rect 30401 21008 30499 21106
rect 31649 21008 31747 21106
rect 32897 21008 32995 21106
rect 34145 21008 34243 21106
rect 35393 21008 35491 21106
rect 36641 21008 36739 21106
rect 37889 21008 37987 21106
rect 39137 21008 39235 21106
rect 40385 21008 40483 21106
rect 41633 21008 41731 21106
rect 42881 21008 42979 21106
rect 44129 21008 44227 21106
rect 45377 21008 45475 21106
rect 46625 21008 46723 21106
rect 47873 21008 47971 21106
rect 49121 21008 49219 21106
rect 50369 21008 50467 21106
rect 51617 21008 51715 21106
rect 52865 21008 52963 21106
rect 54113 21008 54211 21106
rect 55361 21008 55459 21106
rect 56609 21008 56707 21106
rect 17935 20592 18033 20690
rect 19183 20592 19281 20690
rect 20431 20592 20529 20690
rect 21679 20592 21777 20690
rect 22927 20592 23025 20690
rect 24175 20592 24273 20690
rect 25423 20592 25521 20690
rect 26671 20592 26769 20690
rect 27919 20592 28017 20690
rect 29167 20592 29265 20690
rect 30415 20592 30513 20690
rect 31663 20592 31761 20690
rect 32911 20592 33009 20690
rect 34159 20592 34257 20690
rect 35407 20592 35505 20690
rect 36655 20592 36753 20690
rect 37903 20592 38001 20690
rect 39151 20592 39249 20690
rect 40399 20592 40497 20690
rect 41647 20592 41745 20690
rect 42895 20592 42993 20690
rect 44143 20592 44241 20690
rect 45391 20592 45489 20690
rect 46639 20592 46737 20690
rect 47887 20592 47985 20690
rect 49135 20592 49233 20690
rect 50383 20592 50481 20690
rect 51631 20592 51729 20690
rect 52879 20592 52977 20690
rect 54127 20592 54225 20690
rect 55375 20592 55473 20690
rect 56623 20592 56721 20690
rect 71477 20443 71575 20541
rect 18032 20149 18130 20247
rect 28016 20149 28114 20247
rect 38000 20149 38098 20247
rect 47984 20149 48082 20247
rect 7 19772 105 19870
rect 4361 19770 4459 19868
rect 17708 19566 57644 19626
rect 18032 19029 18130 19127
rect 28016 19029 28114 19127
rect 38000 19029 38098 19127
rect 47984 19029 48082 19127
rect 71477 19029 71575 19127
rect 7 18356 105 18454
rect 4361 18356 4459 18454
rect 7 16940 105 17038
rect 4361 16942 4459 17040
rect 6197 1461 6295 1559
rect 7365 1461 7463 1559
rect 8533 1461 8631 1559
rect 9701 1461 9799 1559
rect 10869 1461 10967 1559
rect 12037 1461 12135 1559
rect 13205 1461 13303 1559
rect 14373 1461 14471 1559
rect 15541 1461 15639 1559
rect 16709 1461 16807 1559
rect 17877 1461 17975 1559
rect 19045 1461 19143 1559
rect 20213 1461 20311 1559
rect 21381 1461 21479 1559
rect 22549 1461 22647 1559
rect 23717 1461 23815 1559
rect 24885 1461 24983 1559
rect 26053 1461 26151 1559
rect 27221 1461 27319 1559
rect 28389 1461 28487 1559
rect 29557 1461 29655 1559
rect 30725 1461 30823 1559
rect 31893 1461 31991 1559
rect 33061 1461 33159 1559
rect 34229 1461 34327 1559
rect 35397 1461 35495 1559
rect 36565 1461 36663 1559
rect 37733 1461 37831 1559
rect 38901 1461 38999 1559
rect 40069 1461 40167 1559
rect 41237 1461 41335 1559
rect 42405 1461 42503 1559
rect 43573 1461 43671 1559
rect 44741 1461 44839 1559
rect 45909 1461 46007 1559
rect 47077 1461 47175 1559
rect 48245 1461 48343 1559
rect 5662 374 48878 434
rect 6197 47 6295 145
rect 7365 47 7463 145
rect 8533 47 8631 145
rect 9701 47 9799 145
rect 10869 47 10967 145
rect 12037 47 12135 145
rect 13205 47 13303 145
rect 14373 47 14471 145
rect 15541 47 15639 145
rect 16709 47 16807 145
rect 17877 47 17975 145
rect 19045 47 19143 145
rect 20213 47 20311 145
rect 21381 47 21479 145
rect 22549 47 22647 145
rect 23717 47 23815 145
rect 24885 47 24983 145
rect 26053 47 26151 145
rect 27221 47 27319 145
rect 28389 47 28487 145
rect 29557 47 29655 145
rect 30725 47 30823 145
rect 31893 47 31991 145
rect 33061 47 33159 145
rect 34229 47 34327 145
rect 35397 47 35495 145
rect 36565 47 36663 145
rect 37733 47 37831 145
rect 38901 47 38999 145
rect 40069 47 40167 145
rect 41237 47 41335 145
rect 42405 47 42503 145
rect 43573 47 43671 145
rect 44741 47 44839 145
rect 45909 47 46007 145
rect 47077 47 47175 145
rect 48245 47 48343 145
<< metal4 >>
rect 17805 89217 17865 89277
rect 19053 89217 19113 89277
rect 20301 89217 20361 89277
rect 21549 89217 21609 89277
rect 22797 89217 22857 89277
rect 24045 89217 24105 89277
rect 25293 89217 25353 89277
rect 26541 89217 26601 89277
rect 27789 89217 27849 89277
rect 29037 89217 29097 89277
rect 30285 89217 30345 89277
rect 31533 89217 31593 89277
rect 32781 89217 32841 89277
rect 34029 89217 34089 89277
rect 35277 89217 35337 89277
rect 36525 89217 36585 89277
rect 37773 89217 37833 89277
rect 39021 89217 39081 89277
rect 40269 89217 40329 89277
rect 41517 89217 41577 89277
rect 42765 89217 42825 89277
rect 44013 89217 44073 89277
rect 45261 89217 45321 89277
rect 46509 89217 46569 89277
rect 47757 89217 47817 89277
rect 49005 89217 49065 89277
rect 50253 89217 50313 89277
rect 51501 89217 51561 89277
rect 52749 89217 52809 89277
rect 53997 89217 54057 89277
rect 55245 89217 55305 89277
rect 56493 89217 56553 89277
rect 67578 89217 67638 89277
rect 72573 89217 72633 89277
rect 0 0 76 89156
rect 136 0 212 89156
rect 272 0 348 89156
rect 408 0 484 89156
rect 544 0 620 89156
rect 680 0 756 89156
rect 816 0 892 89156
rect 952 0 1028 89156
rect 1088 0 1164 89156
rect 1224 0 1300 89156
rect 1360 0 1436 89156
rect 1496 0 1572 89156
rect 1632 0 1708 89156
rect 1768 0 1844 89156
rect 1904 0 1980 89156
rect 2040 0 2116 89156
rect 2176 0 2252 89156
rect 2312 0 2388 89156
rect 2448 0 2524 89156
rect 2584 0 2660 89156
rect 2720 17816 2796 89156
rect 2856 17816 2932 89156
rect 2803 66 2863 126
rect 2992 0 3068 89156
rect 3128 0 3204 89156
rect 3264 0 3340 89156
rect 3400 0 3476 89156
rect 3536 0 3612 89156
rect 3672 0 3748 89156
rect 3808 0 3884 89156
rect 3944 0 4020 89156
rect 4080 0 4156 89156
rect 4216 0 4292 89156
rect 4352 0 4428 89156
rect 4488 0 4564 89156
rect 4624 0 4700 89156
rect 4760 0 4836 89156
rect 4896 0 4972 89156
rect 5032 0 5108 89156
rect 5168 0 5244 89156
rect 5304 0 5380 89156
rect 5440 0 5516 89156
rect 5576 0 5652 89156
rect 5712 816 5788 89156
rect 5848 816 5924 89156
rect 5802 66 5862 126
rect 5984 0 6060 89156
rect 6120 0 6196 89156
rect 6256 0 6332 89156
rect 6392 0 6468 89156
rect 6528 0 6604 89156
rect 6664 1768 6740 89156
rect 6800 1768 6876 89156
rect 6936 816 7012 89156
rect 7072 816 7148 89156
rect 6970 66 7030 126
rect 7208 0 7284 89156
rect 7344 0 7420 89156
rect 7480 0 7556 89156
rect 7616 0 7692 89156
rect 7752 0 7828 89156
rect 7888 14960 7964 89156
rect 8024 14960 8100 89156
rect 8160 816 8236 89156
rect 8138 66 8198 126
rect 8296 0 8372 89156
rect 8432 0 8508 89156
rect 8568 0 8644 89156
rect 8704 0 8780 89156
rect 8840 0 8916 89156
rect 8976 8704 9052 89156
rect 9112 8704 9188 89156
rect 9248 816 9324 89156
rect 9384 816 9460 89156
rect 9306 66 9366 126
rect 9520 0 9596 89156
rect 9656 0 9732 89156
rect 9792 0 9868 89156
rect 9928 0 10004 89156
rect 10064 0 10140 89156
rect 10200 13736 10276 89156
rect 10336 13736 10412 89156
rect 10472 816 10548 89156
rect 10608 24752 10684 89156
rect 10744 24752 10820 89156
rect 10474 66 10534 126
rect 10880 0 10956 89156
rect 11016 0 11092 89156
rect 11152 0 11228 89156
rect 11288 5984 11364 89156
rect 11424 5984 11500 89156
rect 11560 816 11636 89156
rect 11696 15232 11772 89156
rect 11832 15232 11908 89156
rect 11642 66 11702 126
rect 11766 66 11826 126
rect 11968 0 12044 89156
rect 12104 0 12180 89156
rect 12240 0 12316 89156
rect 12376 0 12452 89156
rect 12512 2040 12588 89156
rect 12648 2040 12724 89156
rect 12784 816 12860 89156
rect 12920 6528 12996 89156
rect 13056 6528 13132 89156
rect 12810 66 12870 126
rect 12934 66 12994 126
rect 13056 0 13132 6060
rect 13192 0 13268 89156
rect 13328 0 13404 89156
rect 13464 0 13540 89156
rect 13600 0 13676 89156
rect 13736 2312 13812 89156
rect 13872 2312 13948 89156
rect 14008 6664 14084 89156
rect 14144 6664 14220 89156
rect 13978 66 14038 126
rect 14102 66 14162 126
rect 14280 0 14356 89156
rect 14416 0 14492 89156
rect 14552 0 14628 89156
rect 14688 0 14764 89156
rect 14824 2584 14900 89156
rect 14960 2584 15036 89156
rect 15096 816 15172 89156
rect 15232 10064 15308 89156
rect 15368 10064 15444 89156
rect 15146 66 15206 126
rect 15270 66 15330 126
rect 15504 0 15580 89156
rect 15640 0 15716 89156
rect 15776 0 15852 89156
rect 15912 0 15988 89156
rect 16048 9928 16124 89156
rect 16184 9928 16260 89156
rect 16320 11560 16396 89156
rect 16456 11560 16532 89156
rect 16314 66 16374 126
rect 16438 66 16498 126
rect 16592 0 16668 89156
rect 16728 0 16804 89156
rect 16864 0 16940 89156
rect 17000 0 17076 89156
rect 17136 11288 17212 89156
rect 17272 11288 17348 89156
rect 17408 816 17484 89156
rect 17544 19584 17620 89156
rect 17680 22984 17756 85892
rect 17816 22984 17892 85892
rect 17952 20808 18028 89156
rect 17482 66 17542 126
rect 17606 66 17666 126
rect 17816 0 17892 14764
rect 17952 0 18028 1572
rect 18088 0 18164 89156
rect 18224 0 18300 89156
rect 18360 14552 18436 89156
rect 18496 14552 18572 89156
rect 18632 816 18708 89156
rect 18768 7752 18844 89156
rect 18650 66 18710 126
rect 18774 66 18834 126
rect 18904 0 18980 89156
rect 19176 86496 19252 89156
rect 19040 22984 19116 85892
rect 19176 22984 19252 85892
rect 19176 20808 19252 22380
rect 19312 20808 19388 89156
rect 19040 0 19116 6060
rect 19176 0 19252 1844
rect 19312 0 19388 1844
rect 19448 0 19524 89156
rect 19584 7480 19660 89156
rect 19720 816 19796 89156
rect 19856 17952 19932 89156
rect 19992 17952 20068 89156
rect 19818 66 19878 126
rect 19942 66 20002 126
rect 20128 0 20204 89156
rect 20264 22984 20340 85892
rect 20400 22984 20476 85892
rect 20536 20808 20612 89156
rect 20672 17680 20748 89156
rect 20808 17680 20884 89156
rect 20264 0 20340 6196
rect 20400 0 20476 2116
rect 20536 0 20612 2116
rect 20944 816 21020 89156
rect 21080 10336 21156 89156
rect 21216 10336 21292 89156
rect 20986 66 21046 126
rect 21110 66 21170 126
rect 21352 0 21428 89156
rect 21488 22984 21564 85892
rect 21624 22984 21700 85892
rect 21760 20808 21836 89156
rect 21488 0 21564 9732
rect 21896 9656 21972 89156
rect 22032 9656 22108 89156
rect 22168 11832 22244 89156
rect 22304 11832 22380 89156
rect 21624 0 21700 9460
rect 21760 0 21836 9460
rect 22154 66 22214 126
rect 22278 66 22338 126
rect 22440 0 22516 89156
rect 22576 0 22652 89156
rect 22712 22984 22788 85892
rect 22848 22984 22924 85892
rect 22984 20808 23060 89156
rect 23120 11152 23196 89156
rect 22712 0 22788 11092
rect 22848 0 22924 10956
rect 23256 816 23332 89156
rect 23392 15504 23468 89156
rect 23528 15504 23604 89156
rect 23322 66 23382 126
rect 23446 66 23506 126
rect 23664 0 23740 89156
rect 23800 0 23876 89156
rect 23936 22984 24012 85892
rect 24072 22984 24148 85892
rect 24208 20808 24284 89156
rect 23936 0 24012 14356
rect 24344 14280 24420 89156
rect 24072 0 24148 14084
rect 24480 7888 24556 89156
rect 24616 7888 24692 89156
rect 24490 66 24550 126
rect 24614 66 24674 126
rect 24752 0 24828 89156
rect 24888 0 24964 89156
rect 25024 0 25100 89156
rect 25160 22984 25236 85892
rect 25296 22984 25372 85892
rect 25432 20808 25508 89156
rect 25568 20808 25644 89156
rect 25704 18224 25780 89156
rect 25840 18224 25916 89156
rect 25160 0 25236 7284
rect 25296 0 25372 7284
rect 25568 816 25644 7012
rect 25658 66 25718 126
rect 25782 66 25842 126
rect 25976 0 26052 89156
rect 26112 0 26188 89156
rect 26248 0 26324 89156
rect 26384 0 26460 89156
rect 26520 22984 26596 85892
rect 26656 22984 26732 85892
rect 26792 20808 26868 89156
rect 26792 816 26868 17212
rect 26928 8840 27004 89156
rect 27064 8840 27140 89156
rect 26826 66 26886 126
rect 26950 66 27010 126
rect 27200 0 27276 89156
rect 27336 0 27412 89156
rect 27472 0 27548 89156
rect 27608 19584 27684 89156
rect 27744 22984 27820 85892
rect 27880 22984 27956 85892
rect 28016 20808 28092 89156
rect 28152 9384 28228 89156
rect 27608 0 27684 8236
rect 27994 66 28054 126
rect 28118 66 28178 126
rect 28288 0 28364 89156
rect 28424 0 28500 89156
rect 28560 0 28636 89156
rect 28696 0 28772 89156
rect 28832 2856 28908 89156
rect 28968 22984 29044 85892
rect 29104 22984 29180 85892
rect 29240 20808 29316 89156
rect 28968 2856 29044 11364
rect 29376 10880 29452 89156
rect 29104 816 29180 10684
rect 29162 66 29222 126
rect 29286 66 29346 126
rect 29512 0 29588 89156
rect 29648 0 29724 89156
rect 29784 0 29860 89156
rect 29920 0 29996 89156
rect 30056 2992 30132 89156
rect 30192 22984 30268 85892
rect 30328 22984 30404 85892
rect 30464 20808 30540 89156
rect 30192 2992 30268 15036
rect 30330 66 30390 126
rect 30454 66 30514 126
rect 30600 0 30676 89156
rect 30736 0 30812 89156
rect 30872 0 30948 89156
rect 31008 0 31084 89156
rect 31144 3264 31220 89156
rect 31280 3264 31356 89156
rect 31416 22984 31492 85892
rect 31552 22984 31628 85892
rect 31688 20808 31764 89156
rect 31416 816 31492 7420
rect 31498 66 31558 126
rect 31622 66 31682 126
rect 31824 0 31900 89156
rect 31960 0 32036 89156
rect 32096 0 32172 89156
rect 32232 0 32308 89156
rect 32368 3536 32444 89156
rect 32504 3536 32580 89156
rect 32640 816 32716 89156
rect 32776 22984 32852 85892
rect 32912 20808 32988 89156
rect 33048 20808 33124 89156
rect 32666 66 32726 126
rect 32790 66 32850 126
rect 32912 0 32988 16804
rect 33048 0 33124 16940
rect 33184 0 33260 89156
rect 33320 0 33396 89156
rect 33456 0 33532 89156
rect 33592 17000 33668 89156
rect 33728 17000 33804 89156
rect 33864 8160 33940 89156
rect 34000 22984 34076 85892
rect 34136 22984 34212 85892
rect 34272 20808 34348 89156
rect 33834 66 33894 126
rect 33958 66 34018 126
rect 34136 0 34212 7964
rect 34272 0 34348 7964
rect 34408 0 34484 89156
rect 34544 0 34620 89156
rect 34680 4080 34756 89156
rect 34816 4080 34892 89156
rect 34952 816 35028 89156
rect 35088 9112 35164 89156
rect 35224 22984 35300 85892
rect 35360 22984 35436 85892
rect 35496 20808 35572 89156
rect 35002 66 35062 126
rect 35126 66 35186 126
rect 35360 0 35436 2388
rect 35496 0 35572 2388
rect 35632 0 35708 89156
rect 35768 0 35844 89156
rect 35904 4488 35980 89156
rect 36040 4488 36116 89156
rect 36176 10608 36252 89156
rect 36312 10608 36388 89156
rect 36448 22984 36524 85892
rect 36584 22984 36660 85892
rect 36720 20808 36796 89156
rect 36170 66 36230 126
rect 36294 66 36354 126
rect 36448 0 36524 10412
rect 36584 0 36660 2660
rect 36720 0 36796 2660
rect 36856 0 36932 89156
rect 36992 5032 37068 89156
rect 37128 5032 37204 89156
rect 37264 816 37340 89156
rect 37400 13600 37476 89156
rect 37536 19584 37612 89156
rect 37672 22984 37748 85892
rect 37808 22984 37884 85892
rect 37944 20808 38020 89156
rect 37338 66 37398 126
rect 37462 66 37522 126
rect 37672 0 37748 13268
rect 37808 0 37884 2796
rect 37944 0 38020 2796
rect 38080 0 38156 89156
rect 38216 13328 38292 89156
rect 38352 13328 38428 89156
rect 38488 816 38564 89156
rect 38624 16184 38700 89156
rect 38506 66 38566 126
rect 38630 66 38690 126
rect 38760 0 38836 89156
rect 38896 22984 38972 85892
rect 39032 22984 39108 85892
rect 39168 20808 39244 89156
rect 38896 0 38972 6468
rect 39032 0 39108 6468
rect 39168 0 39244 3068
rect 39304 0 39380 89156
rect 39440 16048 39516 89156
rect 39576 816 39652 89156
rect 39712 18360 39788 89156
rect 39848 18360 39924 89156
rect 39674 66 39734 126
rect 39798 66 39858 126
rect 39984 0 40060 89156
rect 40120 0 40196 89156
rect 40256 22984 40332 85892
rect 40392 20808 40468 89156
rect 40528 20808 40604 89156
rect 40256 0 40332 16804
rect 40664 16728 40740 89156
rect 40392 0 40468 16532
rect 40800 816 40876 89156
rect 40936 12104 41012 89156
rect 41072 12104 41148 89156
rect 40842 66 40902 126
rect 40966 66 41026 126
rect 41208 0 41284 89156
rect 41344 0 41420 89156
rect 41480 22984 41556 85892
rect 41616 22984 41692 85892
rect 41752 20808 41828 89156
rect 41480 0 41556 7692
rect 41888 3808 41964 89156
rect 42024 12376 42100 89156
rect 42160 12376 42236 89156
rect 41616 0 41692 3612
rect 42010 66 42070 126
rect 42134 66 42194 126
rect 42296 0 42372 89156
rect 42432 0 42508 89156
rect 42568 0 42644 89156
rect 42704 22984 42780 85892
rect 42840 22984 42916 85892
rect 42976 20808 43052 89156
rect 42704 0 42780 8644
rect 43112 816 43188 89156
rect 43248 12512 43324 89156
rect 43384 12512 43460 89156
rect 43178 66 43238 126
rect 43302 66 43362 126
rect 43520 0 43596 89156
rect 43656 0 43732 89156
rect 43792 0 43868 89156
rect 43928 22984 44004 85892
rect 44064 22984 44140 85892
rect 44200 20808 44276 89156
rect 44336 12784 44412 89156
rect 44472 12784 44548 89156
rect 43928 0 44004 10140
rect 44346 66 44406 126
rect 44470 66 44530 126
rect 44608 0 44684 89156
rect 44744 0 44820 89156
rect 44880 0 44956 89156
rect 45016 0 45092 89156
rect 45152 22984 45228 85892
rect 45288 22984 45364 85892
rect 45424 20808 45500 89156
rect 45152 0 45228 13132
rect 45560 13056 45636 89156
rect 45696 13056 45772 89156
rect 45288 5304 45364 12860
rect 45424 816 45500 12860
rect 45514 66 45574 126
rect 45638 66 45698 126
rect 45832 0 45908 89156
rect 45968 0 46044 89156
rect 46104 0 46180 89156
rect 46240 0 46316 89156
rect 46376 22984 46452 85892
rect 46512 22984 46588 85892
rect 46648 20808 46724 89156
rect 46784 20808 46860 89156
rect 46920 15776 46996 89156
rect 46376 5440 46452 15716
rect 46512 5440 46588 15716
rect 46648 816 46724 15580
rect 46682 66 46742 126
rect 46806 66 46866 126
rect 47056 0 47132 89156
rect 47192 0 47268 89156
rect 47328 0 47404 89156
rect 47464 0 47540 89156
rect 47600 19584 47676 89156
rect 47736 22984 47812 85892
rect 47872 22984 47948 85892
rect 48008 20808 48084 89156
rect 47850 66 47910 126
rect 47974 66 48034 126
rect 48144 0 48220 89156
rect 48280 0 48356 89156
rect 48416 0 48492 89156
rect 48552 0 48628 89156
rect 48688 6256 48764 89156
rect 48824 6256 48900 89156
rect 48960 22984 49036 85892
rect 49096 22984 49172 85892
rect 49232 20808 49308 89156
rect 48960 0 49036 11636
rect 49096 0 49172 3340
rect 49232 0 49308 3340
rect 49368 0 49444 89156
rect 49504 0 49580 89156
rect 49640 0 49716 89156
rect 49776 0 49852 89156
rect 49912 0 49988 89156
rect 50048 0 50124 89156
rect 50184 22984 50260 85892
rect 50320 22984 50396 85892
rect 50456 20808 50532 89156
rect 50184 0 50260 11908
rect 50320 0 50396 3748
rect 50456 0 50532 3748
rect 50592 0 50668 89156
rect 50728 0 50804 89156
rect 50864 0 50940 89156
rect 51000 0 51076 89156
rect 51136 0 51212 89156
rect 51272 0 51348 89156
rect 51408 22984 51484 85892
rect 51544 22984 51620 85892
rect 51680 20808 51756 89156
rect 51408 0 51484 12044
rect 51544 0 51620 4292
rect 51680 0 51756 4292
rect 51816 0 51892 89156
rect 51952 0 52028 89156
rect 52088 0 52164 89156
rect 52224 0 52300 89156
rect 52360 0 52436 89156
rect 52496 0 52572 89156
rect 52632 22984 52708 85892
rect 52768 22984 52844 85892
rect 52904 20808 52980 89156
rect 52632 0 52708 12316
rect 52768 0 52844 12316
rect 52904 0 52980 4836
rect 53040 0 53116 89156
rect 53176 0 53252 89156
rect 53312 0 53388 89156
rect 53448 0 53524 89156
rect 53584 0 53660 89156
rect 53720 0 53796 89156
rect 53856 0 53932 89156
rect 53992 22984 54068 85892
rect 54128 20808 54204 89156
rect 54264 20808 54340 89156
rect 53992 0 54068 12588
rect 54128 0 54204 4972
rect 54264 0 54340 4972
rect 54400 0 54476 89156
rect 54536 0 54612 89156
rect 54672 0 54748 89156
rect 54808 0 54884 89156
rect 54944 0 55020 89156
rect 55080 0 55156 89156
rect 55216 22984 55292 85892
rect 55352 22984 55428 85892
rect 55488 20808 55564 89156
rect 55216 0 55292 15308
rect 55352 0 55428 5244
rect 55488 0 55564 5244
rect 55624 0 55700 89156
rect 55760 0 55836 89156
rect 55896 0 55972 89156
rect 56032 0 56108 89156
rect 56168 0 56244 89156
rect 56304 0 56380 89156
rect 56440 22984 56516 85892
rect 56576 22984 56652 85892
rect 56712 20808 56788 89156
rect 56440 0 56516 15988
rect 56576 0 56652 5788
rect 56712 0 56788 5788
rect 56848 0 56924 89156
rect 56984 0 57060 89156
rect 57120 0 57196 89156
rect 57256 0 57332 89156
rect 57392 0 57468 89156
rect 57528 0 57604 89156
rect 57664 0 57740 89156
rect 57800 0 57876 89156
rect 57936 0 58012 89156
rect 58072 0 58148 89156
rect 58208 0 58284 89156
rect 58344 0 58420 89156
rect 58480 0 58556 89156
rect 58616 0 58692 89156
rect 58752 0 58828 89156
rect 58888 0 58964 89156
rect 59024 0 59100 89156
rect 59160 0 59236 89156
rect 59296 0 59372 89156
rect 59432 0 59508 89156
rect 59568 0 59644 89156
rect 59704 0 59780 89156
rect 59840 0 59916 89156
rect 59976 0 60052 89156
rect 60112 0 60188 89156
rect 60248 0 60324 89156
rect 60384 0 60460 89156
rect 60520 0 60596 89156
rect 60656 0 60732 89156
rect 60792 0 60868 89156
rect 60928 0 61004 89156
rect 61064 0 61140 89156
rect 61200 0 61276 89156
rect 61336 0 61412 89156
rect 61472 0 61548 89156
rect 61608 0 61684 89156
rect 61744 0 61820 89156
rect 61880 0 61956 89156
rect 62016 0 62092 89156
rect 62152 0 62228 89156
rect 62288 0 62364 89156
rect 62424 0 62500 89156
rect 62560 0 62636 89156
rect 62696 0 62772 89156
rect 62832 0 62908 89156
rect 62968 0 63044 89156
rect 63104 0 63180 89156
rect 63240 0 63316 89156
rect 63376 0 63452 89156
rect 63512 0 63588 89156
rect 63648 0 63724 89156
rect 63784 0 63860 89156
rect 63920 0 63996 89156
rect 64056 0 64132 89156
rect 64192 0 64268 89156
rect 64328 0 64404 89156
rect 64464 0 64540 89156
rect 64600 0 64676 89156
rect 64736 0 64812 89156
rect 64872 0 64948 89156
rect 65008 0 65084 89156
rect 65144 0 65220 89156
rect 65280 0 65356 89156
rect 65416 0 65492 89156
rect 65552 0 65628 89156
rect 65688 0 65764 89156
rect 65824 0 65900 89156
rect 65960 0 66036 89156
rect 66096 0 66172 89156
rect 66232 0 66308 89156
rect 66368 0 66444 89156
rect 66504 0 66580 89156
rect 66640 0 66716 89156
rect 66776 0 66852 89156
rect 66912 0 66988 89156
rect 67048 0 67124 89156
rect 67184 0 67260 89156
rect 67320 0 67396 89156
rect 67456 0 67532 87932
rect 67592 0 67668 87932
rect 67728 0 67804 89156
rect 67864 0 67940 89156
rect 68000 0 68076 89156
rect 68136 0 68212 89156
rect 68272 0 68348 89156
rect 68408 0 68484 89156
rect 68544 0 68620 89156
rect 68680 0 68756 89156
rect 68816 0 68892 89156
rect 68952 0 69028 89156
rect 69088 0 69164 89156
rect 69224 0 69300 89156
rect 69360 0 69436 89156
rect 69496 0 69572 89156
rect 69632 0 69708 89156
rect 69768 0 69844 89156
rect 69904 0 69980 89156
rect 70040 0 70116 89156
rect 70176 0 70252 89156
rect 70312 0 70388 89156
rect 70448 0 70524 89156
rect 70584 0 70660 89156
rect 70720 0 70796 89156
rect 70856 0 70932 89156
rect 70992 0 71068 89156
rect 71128 0 71204 89156
rect 71264 0 71340 89156
rect 71400 0 71476 89156
rect 71536 0 71612 89156
rect 71672 0 71748 89156
rect 71808 0 71884 89156
rect 71944 0 72020 89156
rect 72080 0 72156 89156
rect 72216 0 72292 89156
rect 72352 0 72428 89156
rect 72488 0 72564 88340
rect 72624 0 72700 88340
rect 72760 0 72836 89156
rect 72896 0 72972 89156
rect 73032 0 73108 89156
rect 73168 0 73244 89156
rect 73304 0 73380 89156
rect 73440 0 73516 89156
rect 73576 0 73652 89156
rect 73712 0 73788 89156
rect 73848 0 73924 89156
rect 73984 0 74060 89156
rect 74120 0 74196 89156
rect 74256 0 74332 89156
rect 74392 0 74468 89156
rect 74528 0 74604 89156
rect 74664 0 74740 89156
rect 74800 0 74876 89156
rect 74936 0 75012 89156
rect 75072 0 75148 89156
rect 75208 0 75284 89156
<< labels >>
rlabel metal4 s 11642 66 11702 126 6 din0[0]
port 32 nsew default input
rlabel metal4 s 12810 66 12870 126 6 din0[1]
port 31 nsew default input
rlabel metal4 s 13978 66 14038 126 6 din0[2]
port 30 nsew default input
rlabel metal4 s 15146 66 15206 126 6 din0[3]
port 29 nsew default input
rlabel metal4 s 16314 66 16374 126 6 din0[4]
port 28 nsew default input
rlabel metal4 s 17482 66 17542 126 6 din0[5]
port 27 nsew default input
rlabel metal4 s 18650 66 18710 126 6 din0[6]
port 26 nsew default input
rlabel metal4 s 19818 66 19878 126 6 din0[7]
port 25 nsew default input
rlabel metal4 s 20986 66 21046 126 6 din0[8]
port 24 nsew default input
rlabel metal4 s 22154 66 22214 126 6 din0[9]
port 23 nsew default input
rlabel metal4 s 23322 66 23382 126 6 din0[10]
port 22 nsew default input
rlabel metal4 s 24490 66 24550 126 6 din0[11]
port 21 nsew default input
rlabel metal4 s 25658 66 25718 126 6 din0[12]
port 20 nsew default input
rlabel metal4 s 26826 66 26886 126 6 din0[13]
port 19 nsew default input
rlabel metal4 s 27994 66 28054 126 6 din0[14]
port 18 nsew default input
rlabel metal4 s 29162 66 29222 126 6 din0[15]
port 17 nsew default input
rlabel metal4 s 30330 66 30390 126 6 din0[16]
port 16 nsew default input
rlabel metal4 s 31498 66 31558 126 6 din0[17]
port 15 nsew default input
rlabel metal4 s 32666 66 32726 126 6 din0[18]
port 14 nsew default input
rlabel metal4 s 33834 66 33894 126 6 din0[19]
port 13 nsew default input
rlabel metal4 s 35002 66 35062 126 6 din0[20]
port 12 nsew default input
rlabel metal4 s 36170 66 36230 126 6 din0[21]
port 11 nsew default input
rlabel metal4 s 37338 66 37398 126 6 din0[22]
port 10 nsew default input
rlabel metal4 s 38506 66 38566 126 6 din0[23]
port 9 nsew default input
rlabel metal4 s 39674 66 39734 126 6 din0[24]
port 8 nsew default input
rlabel metal4 s 40842 66 40902 126 6 din0[25]
port 7 nsew default input
rlabel metal4 s 42010 66 42070 126 6 din0[26]
port 6 nsew default input
rlabel metal4 s 43178 66 43238 126 6 din0[27]
port 5 nsew default input
rlabel metal4 s 44346 66 44406 126 6 din0[28]
port 4 nsew default input
rlabel metal4 s 45514 66 45574 126 6 din0[29]
port 3 nsew default input
rlabel metal4 s 46682 66 46742 126 6 din0[30]
port 2 nsew default input
rlabel metal4 s 47850 66 47910 126 6 din0[31]
port 1 nsew default input
rlabel metal4 s 5802 66 5862 126 6 addr0[0]
port 40 nsew default input
rlabel metal3 s 26 77073 86 77133 6 addr0[1]
port 39 nsew default input
rlabel metal3 s 26 78773 86 78833 6 addr0[2]
port 38 nsew default input
rlabel metal3 s 26 79901 86 79961 6 addr0[3]
port 37 nsew default input
rlabel metal3 s 26 81601 86 81661 6 addr0[4]
port 36 nsew default input
rlabel metal3 s 26 82729 86 82789 6 addr0[5]
port 35 nsew default input
rlabel metal3 s 26 84429 86 84489 6 addr0[6]
port 34 nsew default input
rlabel metal3 s 26 85557 86 85617 6 addr0[7]
port 33 nsew default input
rlabel metal4 s 67578 89217 67638 89277 6 addr1[0]
port 48 nsew default input
rlabel metal3 s 75266 28382 75326 28442 6 addr1[1]
port 47 nsew default input
rlabel metal3 s 75266 26682 75326 26742 6 addr1[2]
port 46 nsew default input
rlabel metal3 s 75266 25554 75326 25614 6 addr1[3]
port 45 nsew default input
rlabel metal3 s 75266 23854 75326 23914 6 addr1[4]
port 44 nsew default input
rlabel metal3 s 75266 22726 75326 22786 6 addr1[5]
port 43 nsew default input
rlabel metal3 s 75266 21026 75326 21086 6 addr1[6]
port 42 nsew default input
rlabel metal3 s 75266 19898 75326 19958 6 addr1[7]
port 41 nsew default input
rlabel metal3 s 26 17525 86 17585 6 csb0
port 49 nsew default input
rlabel metal3 s 75266 88653 75326 88713 6 csb1
port 50 nsew default input
rlabel metal3 s 26 19225 86 19285 6 web0
port 51 nsew default input
rlabel metal4 s 2803 66 2863 126 6 clk0
port 52 nsew default input
rlabel metal4 s 72573 89217 72633 89277 6 clk1
port 53 nsew default input
rlabel metal4 s 6970 66 7030 126 6 wmask0[0]
port 57 nsew default input
rlabel metal4 s 8138 66 8198 126 6 wmask0[1]
port 56 nsew default input
rlabel metal4 s 9306 66 9366 126 6 wmask0[2]
port 55 nsew default input
rlabel metal4 s 10474 66 10534 126 6 wmask0[3]
port 54 nsew default input
rlabel metal4 s 11766 66 11826 126 6 dout0[0]
port 89 nsew default output
rlabel metal4 s 12934 66 12994 126 6 dout0[1]
port 88 nsew default output
rlabel metal4 s 14102 66 14162 126 6 dout0[2]
port 87 nsew default output
rlabel metal4 s 15270 66 15330 126 6 dout0[3]
port 86 nsew default output
rlabel metal4 s 16438 66 16498 126 6 dout0[4]
port 85 nsew default output
rlabel metal4 s 17606 66 17666 126 6 dout0[5]
port 84 nsew default output
rlabel metal4 s 18774 66 18834 126 6 dout0[6]
port 83 nsew default output
rlabel metal4 s 19942 66 20002 126 6 dout0[7]
port 82 nsew default output
rlabel metal4 s 21110 66 21170 126 6 dout0[8]
port 81 nsew default output
rlabel metal4 s 22278 66 22338 126 6 dout0[9]
port 80 nsew default output
rlabel metal4 s 23446 66 23506 126 6 dout0[10]
port 79 nsew default output
rlabel metal4 s 24614 66 24674 126 6 dout0[11]
port 78 nsew default output
rlabel metal4 s 25782 66 25842 126 6 dout0[12]
port 77 nsew default output
rlabel metal4 s 26950 66 27010 126 6 dout0[13]
port 76 nsew default output
rlabel metal4 s 28118 66 28178 126 6 dout0[14]
port 75 nsew default output
rlabel metal4 s 29286 66 29346 126 6 dout0[15]
port 74 nsew default output
rlabel metal4 s 30454 66 30514 126 6 dout0[16]
port 73 nsew default output
rlabel metal4 s 31622 66 31682 126 6 dout0[17]
port 72 nsew default output
rlabel metal4 s 32790 66 32850 126 6 dout0[18]
port 71 nsew default output
rlabel metal4 s 33958 66 34018 126 6 dout0[19]
port 70 nsew default output
rlabel metal4 s 35126 66 35186 126 6 dout0[20]
port 69 nsew default output
rlabel metal4 s 36294 66 36354 126 6 dout0[21]
port 68 nsew default output
rlabel metal4 s 37462 66 37522 126 6 dout0[22]
port 67 nsew default output
rlabel metal4 s 38630 66 38690 126 6 dout0[23]
port 66 nsew default output
rlabel metal4 s 39798 66 39858 126 6 dout0[24]
port 65 nsew default output
rlabel metal4 s 40966 66 41026 126 6 dout0[25]
port 64 nsew default output
rlabel metal4 s 42134 66 42194 126 6 dout0[26]
port 63 nsew default output
rlabel metal4 s 43302 66 43362 126 6 dout0[27]
port 62 nsew default output
rlabel metal4 s 44470 66 44530 126 6 dout0[28]
port 61 nsew default output
rlabel metal4 s 45638 66 45698 126 6 dout0[29]
port 60 nsew default output
rlabel metal4 s 46806 66 46866 126 6 dout0[30]
port 59 nsew default output
rlabel metal4 s 47974 66 48034 126 6 dout0[31]
port 58 nsew default output
rlabel metal4 s 17805 89217 17865 89277 6 dout1[0]
port 121 nsew default output
rlabel metal4 s 19053 89217 19113 89277 6 dout1[1]
port 120 nsew default output
rlabel metal4 s 20301 89217 20361 89277 6 dout1[2]
port 119 nsew default output
rlabel metal4 s 21549 89217 21609 89277 6 dout1[3]
port 118 nsew default output
rlabel metal4 s 22797 89217 22857 89277 6 dout1[4]
port 117 nsew default output
rlabel metal4 s 24045 89217 24105 89277 6 dout1[5]
port 116 nsew default output
rlabel metal4 s 25293 89217 25353 89277 6 dout1[6]
port 115 nsew default output
rlabel metal4 s 26541 89217 26601 89277 6 dout1[7]
port 114 nsew default output
rlabel metal4 s 27789 89217 27849 89277 6 dout1[8]
port 113 nsew default output
rlabel metal4 s 29037 89217 29097 89277 6 dout1[9]
port 112 nsew default output
rlabel metal4 s 30285 89217 30345 89277 6 dout1[10]
port 111 nsew default output
rlabel metal4 s 31533 89217 31593 89277 6 dout1[11]
port 110 nsew default output
rlabel metal4 s 32781 89217 32841 89277 6 dout1[12]
port 109 nsew default output
rlabel metal4 s 34029 89217 34089 89277 6 dout1[13]
port 108 nsew default output
rlabel metal4 s 35277 89217 35337 89277 6 dout1[14]
port 107 nsew default output
rlabel metal4 s 36525 89217 36585 89277 6 dout1[15]
port 106 nsew default output
rlabel metal4 s 37773 89217 37833 89277 6 dout1[16]
port 105 nsew default output
rlabel metal4 s 39021 89217 39081 89277 6 dout1[17]
port 104 nsew default output
rlabel metal4 s 40269 89217 40329 89277 6 dout1[18]
port 103 nsew default output
rlabel metal4 s 41517 89217 41577 89277 6 dout1[19]
port 102 nsew default output
rlabel metal4 s 42765 89217 42825 89277 6 dout1[20]
port 101 nsew default output
rlabel metal4 s 44013 89217 44073 89277 6 dout1[21]
port 100 nsew default output
rlabel metal4 s 45261 89217 45321 89277 6 dout1[22]
port 99 nsew default output
rlabel metal4 s 46509 89217 46569 89277 6 dout1[23]
port 98 nsew default output
rlabel metal4 s 47757 89217 47817 89277 6 dout1[24]
port 97 nsew default output
rlabel metal4 s 49005 89217 49065 89277 6 dout1[25]
port 96 nsew default output
rlabel metal4 s 50253 89217 50313 89277 6 dout1[26]
port 95 nsew default output
rlabel metal4 s 51501 89217 51561 89277 6 dout1[27]
port 94 nsew default output
rlabel metal4 s 52749 89217 52809 89277 6 dout1[28]
port 93 nsew default output
rlabel metal4 s 53997 89217 54057 89277 6 dout1[29]
port 92 nsew default output
rlabel metal4 s 55245 89217 55305 89277 6 dout1[30]
port 91 nsew default output
rlabel metal4 s 56493 89217 56553 89277 6 dout1[31]
port 90 nsew default output
rlabel metal3 s 10863 51771 10961 51869 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 73868 63403 73966 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 63512 63316 63588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 31603 63403 31701 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 75208 75284 75284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 58888 52904 63316 52980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 38216 63316 38292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 55698 63403 55796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64328 82280 75284 82356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32828 28052 32926 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27350 28662 27410 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 30056 2992 30132 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 19720 816 19796 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 50456 63316 50532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 74681 64489 74779 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 53709 64057 53807 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 16709 1461 16807 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 18360 14552 18436 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 68338 12047 68436 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 5304 46180 5380 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 56511 64489 56609 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 68136 16396 68212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 52561 11393 52659 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 63598 12047 63696 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 31688 20808 31764 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 59160 16396 59236 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49914 80916 50012 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 44661 10961 44759 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 71879 11393 71977 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 38760 75284 38836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 51272 75284 51348 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 3861 83560 3959 83658 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51631 20592 51729 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 55352 16396 55428 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 68952 0 69028 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 79398 63403 79496 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 74681 11393 74779 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 54908 63403 55006 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 43848 63403 43946 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67681 34391 67779 34489 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38216 3128 75284 3204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 31688 16396 31764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8533 1461 8631 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 29651 11393 29749 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 61336 75284 61412 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 34136 0 34212 7964 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 65960 75284 66036 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 55721 64489 55819 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22982 80344 23042 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1360 28424 70388 28500 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 70299 64489 70397 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47077 1461 47175 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11424 23800 70116 23876 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 6936 25100 7012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 37119 64057 37217 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 64411 10961 64509 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38000 20149 38098 20247 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 36761 10961 36859 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 58463 12047 58561 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 48193 63403 48291 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 45832 58284 45908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 75053 12047 75151 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 78200 63316 78276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29557 1461 29655 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 14008 6664 14084 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 41859 64057 41957 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 46920 15776 46996 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 46648 63316 46724 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 62831 64057 62929 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 31144 75284 31220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 53351 64489 53449 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 51544 0 51620 4292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 28424 0 28500 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17347 28643 17445 28741 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 35553 12047 35651 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 50549 64057 50647 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 58072 16396 58148 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 39032 63316 39108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 43000 23094 43098 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 39032 16396 39108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17877 1461 17975 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36760 23094 36858 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21210 80916 21308 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 32393 12047 32491 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 33320 0 33396 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 64328 10140 64404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 67153 63403 67251 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 8840 34892 8916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49096 408 75284 484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25478 28662 25538 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 77409 11393 77507 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 49096 75284 49172 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 79288 63316 79364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 63784 0 63860 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 37944 63316 38020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 68719 64489 68817 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 61064 75284 61140 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41740 85036 41838 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42895 20592 42993 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26202 28052 26300 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49814 80344 49874 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 48280 0 48356 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 52561 64057 52659 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 53720 63316 53796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51816 12376 75284 12452 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 45428 12047 45526 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 39848 10140 39924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 64056 58284 64132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 70708 12047 70806 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36186 28052 36284 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 64411 64057 64509 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 69151 64489 69249 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 70040 10140 70116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 61608 10140 61684 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21210 28052 21308 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 45016 0 45092 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 46104 0 46180 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1904 30056 10140 30132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20524 85036 20622 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 69768 16396 69844 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51724 23932 51822 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 69941 64057 70039 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 55303 12047 55401 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38582 80344 38642 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 75208 10140 75284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 72760 10140 72836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29376 11560 75284 11636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 52904 10140 52980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 75843 12047 75941 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 42024 63316 42100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46070 28662 46130 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 76619 10961 76717 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 63784 75284 63860 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 29240 58284 29316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 41501 64057 41599 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 75471 64057 75569 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26053 1461 26151 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 47192 58284 47268 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 17272 11288 17348 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 56440 16396 56516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 28968 2856 29044 11364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22032 9656 75284 9732 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 70584 11364 70660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 78989 11393 79087 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 73891 64057 73989 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26928 17816 75284 17892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 33601 10961 33699 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 46104 75284 46180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 42291 11393 42389 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 67320 75284 67396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49814 28662 49874 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 13192 0 13268 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 67929 11393 68027 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 58068 12047 58166 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 44472 12784 44548 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 2312 0 2388 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 41752 75284 41828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42326 28662 42386 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 48280 75284 48356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 75752 10140 75828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 71089 64057 71187 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 45560 10140 45636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51548 80916 51646 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 10472 816 10548 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 62018 12047 62116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 46920 75284 46996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 68680 75284 68756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44123 21542 44221 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 39108 63403 39206 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 47821 64057 47919 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34076 80916 34174 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37958 28662 38018 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 34680 4080 34756 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 49759 64057 49857 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 49912 0 49988 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 53658 28052 53756 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 18088 0 18164 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 25704 18224 25780 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 58449 64489 58547 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 64769 11393 64867 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 35181 64057 35279 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 73576 16396 73652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 22440 0 22516 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45308 80916 45406 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 50191 64489 50289 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 33973 12047 34071 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 34136 16396 34212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 61609 64057 61707 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32342 80344 32402 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 75480 16396 75556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 54499 11393 54597 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 11832 15232 11908 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 79016 16396 79092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 21080 17620 21156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 41208 16396 41284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 2448 18904 17756 18980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44198 80344 44258 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52859 21542 52957 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 77656 75284 77732 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 53709 11393 53807 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44472 4760 75284 4836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 43112 63316 43188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 52538 12047 52636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8008 29635 8106 29733 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 52632 16396 52708 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27064 17544 75284 17620 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30415 20592 30513 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 34680 16396 34756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 5032 44956 5108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17915 21542 18013 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 38760 58284 38836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 41208 58284 41284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 7480 0 7556 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 40392 58284 40468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4361 24012 4459 24110 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40504 23094 40602 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 53723 63403 53821 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42812 80916 42910 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 72488 75284 72564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 272 19720 4156 19796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 17816 0 17892 14764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 37672 75284 37748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 56869 64489 56967 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 48824 58284 48900 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50488 23094 50586 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 74664 0 74740 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 3672 0 3748 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 73032 16396 73108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 31416 58284 31492 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 58449 64057 58547 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 31231 10961 31329 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 47736 10140 47812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 25976 11228 26052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36710 80344 36770 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 43384 75284 43460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 13464 10004 13540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24344 14552 75284 14628 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 64600 16396 64676 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 58616 10140 58692 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 59160 75284 59236 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 64411 11393 64509 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 79288 58284 79364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 36329 64057 36427 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 46599 11393 46697 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 36312 75284 36388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56603 21542 56701 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 22712 4156 22788 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 63993 12047 64091 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1191 34014 1289 34112 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 73032 63316 73108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 66504 63316 66580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71808 23256 75284 23332 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55292 80916 55390 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 65991 64057 66089 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 68136 0 68212 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 31589 64489 31687 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 60248 58284 60324 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37334 28662 37394 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 66504 16396 66580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 24888 0 24964 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 56712 16396 56788 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 44200 75284 44276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 58616 16396 58692 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 57800 16396 57876 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 32811 64489 32909 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 32811 64057 32909 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 56093 63403 56191 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 50728 75284 50804 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 53992 22984 54068 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 37944 20808 38020 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 51816 63316 51892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 31144 63316 31220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 58091 11393 58189 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 76840 3068 76916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 70856 16396 70932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31194 28052 31292 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1904 31144 10140 31220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 53328 63403 53426 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 33592 16396 33668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 34391 64057 34489 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4624 28152 75284 28228 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42426 80916 42524 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 45288 5304 45364 12860 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 53992 58284 54068 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 27608 4156 27684 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 71672 73788 71748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 75208 58284 75284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 52561 64489 52659 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 70312 0 70388 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27836 28052 27934 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46556 80916 46654 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 36761 64057 36859 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 59704 0 59780 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 49096 63316 49172 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48552 136 75284 212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 3861 77904 3959 78002 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22844 80916 22942 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 31589 11393 31687 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 19176 0 19252 1844 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 62424 0 62500 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 63784 16396 63860 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 43112 10140 43188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 88808 67668 88884 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21772 23932 21870 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 9701 1461 9799 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 73459 64057 73557 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 62696 0 62772 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 61609 11393 61707 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35387 21542 35485 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 49096 58284 49172 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 41208 63316 41284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 43081 10961 43179 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 37909 10961 38007 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34076 28052 34174 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 50549 10961 50647 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 63512 0 63588 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 22984 75284 23060 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 84184 17484 84260 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 48552 0 48628 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54182 28662 54242 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 56984 16396 57060 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 68719 64057 68817 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 76024 73788 76100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 46218 63403 46316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 58881 64057 58979 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 43573 1461 43671 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34214 80344 34274 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20213 1461 20311 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74063 74954 74161 75052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26764 23932 26862 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21659 21542 21757 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 50728 0 50804 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 35496 0 35572 2388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 48280 16396 48356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 65201 64057 65299 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 34952 58284 35028 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57120 22712 69980 22788 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55480 85874 55578 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 55624 75284 55700 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 55080 64540 55156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67246 32005 67344 32103 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 63598 63403 63696 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 52933 63403 53031 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 52088 0 52164 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26764 85036 26862 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 33601 11393 33699 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 63240 63316 63316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 45832 10140 45908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 55721 11393 55819 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 54808 10140 54884 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50438 80344 50498 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 44472 16396 44548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 680 0 756 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 49912 10140 49988 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 24072 0 24148 14084 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 16184 27608 75284 27684 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36748 23932 36846 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21596 28052 21694 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 39489 11393 39587 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 40120 58284 40196 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 50958 12047 51056 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 16728 0 16804 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 66595 35158 66693 35256 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 15640 46588 15716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34938 28052 35036 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 73304 89080 75012 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 88264 67260 88340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 52088 63316 52164 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 73576 63316 73652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 9928 0 10004 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 36312 63316 36388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 78631 11393 78729 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 31231 64057 31329 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 52088 58284 52164 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21734 80344 21794 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 42663 12047 42761 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 31589 64057 31687 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12240 25976 71204 26052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 1496 0 1572 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57907 80325 58005 80423 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47980 23932 48078 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 20264 22984 20340 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 78744 58284 78820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 43871 11393 43969 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 56079 64489 56177 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 79288 3612 79364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 56168 75284 56244 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1904 33320 10140 33396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 59160 58284 59236 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 12648 2040 12724 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 57301 11393 57399 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 35181 64489 35279 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57120 86088 75284 86164 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 54264 10140 54340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 50184 75284 50260 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 75829 10961 75927 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47418 28052 47516 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 55352 63316 55428 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52972 85036 53070 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 86632 75284 86708 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 71672 64540 71748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 66776 0 66852 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 78472 16396 78548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 41069 10961 41167 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 23800 0 23876 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 69224 29784 75284 29860 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 63979 64057 64077 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 53720 16396 53796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 43439 11393 43537 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 48611 10961 48709 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 48280 58284 48356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 73304 0 73380 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 35539 64489 35637 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 66232 75284 66308 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 57800 10140 57876 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40379 21542 40477 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26651 21542 26749 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 54536 61140 54612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 408 17544 2524 17620 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 15368 10064 15444 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 30009 64489 30107 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 40664 75284 40740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 73032 75284 73108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 35181 10961 35279 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8659 32788 8757 32886 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 43112 58284 43188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 45560 58284 45636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 78199 10961 78297 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 43081 64489 43179 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 74392 58284 74468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 70040 16396 70116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 65144 75284 65220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 33048 75284 33124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56728 85874 56826 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 40279 10961 40377 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51686 80344 51746 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 19992 71612 20068 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37434 28052 37532 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 72216 0 72292 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 66595 34368 66693 34466 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25528 85874 25626 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 50549 11393 50647 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 45016 16396 45092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 37551 64057 37649 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 56883 12047 56981 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 33048 16396 33124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 56511 10961 56609 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36572 80916 36670 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22844 28052 22942 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 45016 75284 45092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 50168 63403 50266 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28698 80916 28796 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 54808 75284 54884 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 59239 64057 59337 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 63203 12047 63301 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 50728 58284 50804 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 61228 63403 61326 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 35496 20808 35572 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 33048 58284 33124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 34368 63403 34466 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 27608 0 27684 8236 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21734 28662 21794 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39151 20592 39249 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 42568 16396 42644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 37128 58284 37204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 59432 64540 59508 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 30441 11393 30539 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 39032 58284 39108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74063 70474 74161 70572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 55289 64489 55387 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 2040 13540 2116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40454 28662 40514 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 66781 10961 66879 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46732 23932 46830 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 15368 23196 15444 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 70312 75284 70388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54906 80916 55004 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 39489 10961 39587 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23032 85874 23130 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 62152 63316 62228 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23120 11288 75284 11364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 33959 64489 34057 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 69496 75284 69572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 58616 58284 58692 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 56984 63316 57060 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 30799 64489 30897 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 55896 16396 55972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 37672 58284 37748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 55624 58284 55700 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 79398 12047 79496 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 59648 12047 59746 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51548 28052 51646 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57788 80916 57886 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30508 85036 30606 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 15541 1461 15639 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56540 28052 56638 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 48179 64489 48277 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30508 23932 30606 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 41478 12047 41576 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 42291 64057 42389 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 33592 75284 33668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 59239 11393 59337 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 83912 75284 83988 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 55896 58284 55972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 70856 63316 70932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 53328 12047 53426 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25516 85036 25614 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 50958 63403 51056 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 44229 11393 44327 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 55080 58284 55156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 63240 10140 63316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 59976 75284 60052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 54808 63316 54884 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 34749 11393 34847 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 37672 22984 37748 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 61251 11393 61349 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42988 23932 43086 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 30328 22984 30404 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 68408 36856 75284 36932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21679 20592 21777 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8659 36738 8757 36836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 29784 63316 29860 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23032 23094 23130 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 32811 10961 32909 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 54931 11393 55029 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 32232 16396 32308 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50363 21542 50461 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 18904 0 18980 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 44200 58284 44276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 23528 15504 23604 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 8568 0 8644 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 76024 10140 76100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47318 28662 47378 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 52360 58284 52436 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 43656 0 43732 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67249 36761 67347 36859 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 21080 10336 21156 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 46376 22984 46452 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55430 28662 55490 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 57659 64489 57757 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 57659 64057 57757 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 48179 11393 48277 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37996 23932 38094 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57392 82552 75284 82628 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 71128 10140 71204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 52632 0 52708 12316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 81464 3204 81540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 11560 21972 11636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 39576 10140 39652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33061 1461 33159 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37820 80916 37918 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 54499 64489 54597 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 52904 75284 52980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 71128 63316 71204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 50184 0 50260 11908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 69224 10140 69300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 23256 4156 23332 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 1224 75284 1300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 43674 28052 43772 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27899 21542 27997 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 61880 75284 61956 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29167 20592 29265 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 33864 63316 33940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35768 2584 75284 2660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 78744 73380 78820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 46241 10961 46339 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55292 28052 55390 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 6197 1461 6295 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 53992 75284 54068 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 47192 0 47268 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 272 17000 2252 17076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 49773 12047 49871 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 37400 16396 37476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42812 28052 42910 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 14008 24012 14084 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 53176 75284 53252 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34544 8296 75284 8372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 60248 75284 60324 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 65144 16396 65220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 43928 58284 44004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30600 15368 75284 15444 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 15096 816 15172 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 46104 58284 46180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 41480 10140 41556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 19992 17952 20068 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 57528 0 57604 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 46104 11364 46180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 40392 10140 40468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 54908 12047 55006 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 78200 73788 78276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24268 23932 24366 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17347 80325 17445 80423 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 51272 63316 51348 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32966 28662 33026 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 80648 70660 80724 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 77928 10140 78004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 66504 58284 66580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 66363 63403 66461 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44822 28662 44882 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 3128 0 3204 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 62041 64057 62139 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52410 80916 52508 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 69941 10961 70039 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 79288 16396 79364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 71400 10140 71476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 45451 10961 45549 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29272 23094 29370 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 50456 58284 50532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 58881 11393 58979 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 78989 64489 79087 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 76261 10961 76359 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 7573 35971 7671 36069 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 37133 63403 37231 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71264 84184 75284 84260 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 33320 63316 33396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 74664 58284 74740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 42840 22984 42916 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 47464 10140 47540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 69224 75284 69300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 51544 22984 51620 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 47389 64057 47487 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 51000 0 51076 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 67864 63316 67940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 53720 0 53796 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 39131 10961 39229 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 36584 0 36660 2660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 49401 11393 49499 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 76568 73380 76644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 67929 64489 68027 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47804 80916 47902 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 77841 64057 77939 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 50563 63403 50661 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 77112 75284 77188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 79016 75284 79092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 34952 75284 35028 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 31144 16396 31220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19238 28662 19298 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 68952 58284 69028 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28024 85874 28122 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 61608 0 61684 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45391 20592 45489 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 34952 816 35028 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 71521 64489 71619 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 59671 11393 59769 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57800 83640 70660 83716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 51339 64057 51437 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 61336 16396 61412 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 47031 64057 47129 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 31208 12047 31306 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 53448 16396 53524 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56984 21896 75284 21972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 24072 75284 24148 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 46241 64489 46339 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 76261 11393 76359 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 68569 31998 68667 32096 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 5440 85544 75284 85620 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 68361 10961 68459 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 70312 63316 70388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 75208 63316 75284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 62424 75284 62500 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 72760 16396 72836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 71672 16396 71748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 56869 11393 56967 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 72669 11393 72767 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 64388 63403 64486 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 73576 58284 73652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 36856 58284 36932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 34763 12047 34861 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 70312 58284 70388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30332 28052 30430 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 11016 22788 11092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 6120 48492 6196 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18040 85874 18138 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 33864 8160 33940 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25478 80344 25538 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 54931 10961 55029 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 30872 0 30948 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 29512 16396 29588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 32776 63316 32852 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 43574 28662 43634 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29222 80344 29282 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 9384 816 9460 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27974 28662 28034 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 66776 63316 66852 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 51816 0 51892 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 30600 58284 30676 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 62399 11393 62497 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 67864 10140 67940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 52919 10961 53017 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 40120 0 40196 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 53176 58284 53252 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 50168 12047 50266 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 49096 16396 49172 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 63979 64489 64077 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 70040 63316 70116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46744 85874 46842 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41078 28662 41138 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 69509 10961 69607 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 47008 63403 47106 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4361 18356 4459 18454 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 43871 64057 43969 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 73440 85816 75284 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 42840 10140 42916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 47736 16396 47812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67249 35181 67347 35279 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 40711 64489 40809 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67681 35971 67779 36069 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 44200 20808 44276 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 36584 16396 36660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 34391 10961 34489 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 37551 11393 37649 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 42291 10961 42389 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 74120 75284 74196 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 36584 58284 36660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 62424 58284 62500 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31756 85036 31854 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 38341 64489 38439 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 30872 75284 30948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 48552 10140 48628 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 65688 58284 65764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 71103 63403 71201 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4080 82280 63724 82356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 69496 58284 69572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38682 80916 38780 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 73459 11393 73557 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36086 28662 36146 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 35971 11393 36069 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23706 80916 23804 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56678 80344 56738 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 35496 63316 35572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 68272 88808 72564 88884 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40800 16728 75284 16804 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 57278 63403 57376 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 36856 16396 36932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45484 23932 45582 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54806 28662 54866 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56154 80916 56252 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 65559 64057 65657 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 40936 58284 41012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 38341 64057 38439 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 32504 58284 32580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 51816 58284 51892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20348 80916 20446 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 78199 64489 78297 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4361 26840 4459 26938 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 31416 16396 31492 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 69151 11393 69249 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40316 80916 40414 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 63979 11393 64077 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 27064 75284 27140 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 54808 16396 54884 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 70856 58284 70932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 49759 10961 49857 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 71498 12047 71596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27450 80916 27548 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 71521 10961 71619 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 42024 75284 42100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 79016 63316 79092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 35768 75284 35844 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 62424 63316 62500 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 22984 20808 23060 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 56168 63316 56244 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 43112 75284 43188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 33601 64489 33699 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40664 17000 75284 17076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 66595 30418 66693 30516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 40120 16396 40196 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20524 23932 20622 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 30799 10961 30897 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 35224 63316 35300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 39898 12047 39996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 50456 75284 50532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24175 20592 24273 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 59704 63316 59780 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 73101 11393 73199 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 69224 16396 69300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 66758 63403 66856 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 30056 58284 30132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 59704 10140 59780 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46639 20592 46737 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 30328 16396 30404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44822 80344 44882 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 14552 0 14628 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 46648 10140 46724 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 45832 75284 45908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 34749 64489 34847 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18360 19176 27412 19252 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 58888 0 58964 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 2856 17816 2932 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 69128 63403 69226 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 36040 58284 36116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48666 80916 48764 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 40664 63316 40740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 63621 11393 63719 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 49401 64489 49499 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 71400 75284 71476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 63240 16396 63316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48566 28662 48626 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 72669 64057 72767 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 56168 0 56244 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 41752 63316 41828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35462 80344 35522 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 37672 63316 37748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23020 85036 23118 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 62808 63403 62906 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 77112 58284 77188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 67592 16396 67668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 42296 58284 42372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 31688 75284 31764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 39108 12047 39206 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 9928 15036 10004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57936 19448 75284 19524 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 27336 1572 27412 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40492 23932 40590 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37733 1461 37831 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 62152 58284 62228 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 36856 0 36932 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 44472 58284 44548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 46376 75284 46452 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 66349 64489 66447 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 45560 16396 45636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49232 680 75284 756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 77928 58284 78004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 40664 16728 40740 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 54931 64057 55029 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 72683 63403 72781 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 62968 58284 63044 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52934 28662 52994 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 34749 10961 34847 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4080 85000 75284 85076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 75039 64057 75137 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 38760 16396 38836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 61336 10140 61412 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 71400 58284 71476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19276 85036 19374 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 61251 10961 61349 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 38216 13328 38292 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 61064 16396 61140 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 60043 63403 60141 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 58072 75284 58148 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31893 1461 31991 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 44200 10140 44276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 73576 10140 73652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32891 21542 32989 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4896 76840 16396 76916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 18088 25508 18164 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29846 28662 29906 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 28696 0 28772 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 77384 58284 77460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 39032 22984 39108 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33590 80344 33650 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 33973 63403 34071 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33016 85874 33114 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21596 80916 21694 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 60438 63403 60536 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 61609 10961 61707 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 42024 12376 42100 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 30009 64057 30107 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 40688 63403 40786 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 82280 3612 82356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 74658 12047 74756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 42024 16396 42100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 74664 10140 74740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 58888 16396 58964 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 65416 0 65492 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 46648 75284 46724 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 41859 64489 41957 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 33578 12047 33676 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34214 28662 34274 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 5032 78744 10140 78820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 48611 11393 48709 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67681 36761 67779 36859 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 39032 10140 39108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 65144 0 65220 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 65416 58284 65492 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52972 23932 53070 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 71944 63316 72020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 39898 63403 39996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 66232 0 66308 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 43656 75284 43732 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 18632 816 18708 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 32021 10961 32119 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33004 23932 33102 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 43453 12047 43551 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 56440 22984 56516 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 39503 12047 39601 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 50184 10140 50260 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 33592 63316 33668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40069 1461 40167 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 76296 10140 76372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 25160 0 25236 7284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 42840 64540 42916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 70040 0 70116 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27919 20592 28017 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 45832 0 45908 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 3808 18632 75284 18708 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 37400 13600 37476 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 44243 63403 44341 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 68569 29628 68667 29726 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 31960 0 32036 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 43928 0 44004 10140 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 36584 75284 36660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 59432 10140 59508 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 24072 22984 24148 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 13192 38020 13268 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 41752 16396 41828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24280 23094 24378 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 46376 58284 46452 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 44200 16396 44276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 47821 11393 47919 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 47403 63403 47501 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71477 27513 71575 27611 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 66595 32788 66693 32886 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 62696 10140 62772 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 89080 70660 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 57800 75284 57876 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 75480 63316 75556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 952 0 1028 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 75829 11393 75927 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 65688 75284 65764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 39131 64489 39229 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 58344 16396 58420 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 43656 16396 43732 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 43112 8840 75284 8916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45496 23094 45594 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 408 4292 484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 74664 75284 74740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 75448 12047 75546 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55355 21542 55453 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47887 20592 47985 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 72488 0 72564 88340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 75471 10961 75569 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 73473 12047 73571 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 73304 58284 73380 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 39848 75284 39924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 67592 0 67668 87932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20411 21542 20509 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19163 21542 19261 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49190 28662 49250 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 33959 11393 34057 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 29512 0 29588 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57402 28052 57500 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 41859 10961 41957 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 44472 75284 44548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22549 1461 22647 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 30056 63316 30132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 71672 58284 71748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 2584 28636 2660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 44229 64489 44327 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 1768 12316 1844 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 37923 63403 38021 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29946 80916 30044 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 62968 75284 63044 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 70584 0 70660 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 69509 64489 69607 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42405 1461 42503 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 10200 13736 10276 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4080 79288 10140 79364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 41873 12047 41971 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44248 85874 44346 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 5032 0 5108 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71808 28968 75284 29044 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 4488 43868 4564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 50184 63316 50260 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 57659 11393 57757 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 7573 34391 7671 34489 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 43674 80916 43772 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 65559 11393 65657 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 34391 64489 34489 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 67048 11364 67124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 55289 64057 55387 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38080 13736 75284 13812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 57673 63403 57771 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 65201 10961 65299 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 61064 58284 61140 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 54808 58284 54884 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 44200 63316 44276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 2992 17544 20476 17620 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 60520 58284 60596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 77841 11393 77939 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31094 80344 31154 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 31231 11393 31329 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 68733 63403 68831 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 74120 0 74196 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 52933 12047 53031 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 49368 0 49444 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 68680 16396 68756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 62696 75284 62772 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35500 23932 35598 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19238 80344 19298 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74063 79434 74161 79532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36565 1461 36663 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 41069 64489 41167 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 53709 10961 53807 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 60520 10140 60596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 46104 63316 46180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 46613 63403 46711 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 17272 26324 17348 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 55352 10140 55428 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46619 21542 46717 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 62696 16396 62772 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35397 1461 35495 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49228 23932 49326 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48245 1461 48343 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36992 2856 75284 2932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 79832 75284 79908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 36312 16396 36388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 73101 10961 73199 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 53448 75284 53524 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 43058 63403 43156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 75829 64489 75927 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 53720 75284 53796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 14552 17348 14628 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8659 35948 8757 36046 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 60461 64057 60559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 52919 64489 53017 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 46920 10140 46996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 85816 71748 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 47008 12047 47106 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 65968 63403 66066 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 51544 16396 51620 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12820 54468 12918 54566 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 88536 67124 88612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 36312 58284 36388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28012 85036 28110 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 31603 12047 31701 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 35539 10961 35637 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 52904 0 52980 4836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 43928 22984 44004 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 43848 12047 43946 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 78989 64057 79087 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 62968 10140 63044 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 63979 10961 64077 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 62424 10140 62500 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 43871 10961 43969 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 63189 10961 63287 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 47464 58284 47540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 22712 0 22788 11092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 64056 75284 64132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30470 80344 30530 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 82008 75284 82084 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 60029 64057 60127 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 39848 18360 39924 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 83368 17484 83444 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21772 85036 21870 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 54264 58284 54340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41702 28662 41762 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 57256 75284 57332 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 72288 12047 72386 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45909 1461 46007 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26776 23094 26874 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18714 28052 18812 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 38488 816 38564 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 42024 58284 42100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 12920 45364 12996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 55896 75284 55972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8659 34368 8757 34466 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 42840 16396 42916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 5848 11092 5924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 70584 75284 70660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54232 23094 54330 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 42663 63403 42761 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 6120 0 6196 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 42268 63403 42366 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 79003 12047 79101 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74799 74954 74897 75052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 79560 75284 79636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 67548 63403 67646 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 73101 64489 73199 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 77028 63403 77126 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24954 28052 25052 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42950 80344 43010 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29846 80344 29906 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 67571 11393 67669 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 80104 58284 80180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 50191 64057 50289 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 31960 63316 32036 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 65688 16396 65764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41888 8024 75284 8100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 66776 16396 66852 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48008 5848 75284 5924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 42649 64057 42747 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 84728 75284 84804 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 76633 12047 76731 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 78213 63403 78311 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 21896 4156 21972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51611 21542 51709 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51724 85036 51822 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 34680 58284 34756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 32504 16396 32580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 34952 10140 35028 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 40392 0 40468 16532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 56984 75284 57060 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67973 87364 68071 87462 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 29784 6196 29860 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 11288 16124 11364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31960 6936 75284 7012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29222 28662 29282 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47980 85036 48078 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 75039 10961 75137 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28598 28662 28658 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 46648 816 46724 15580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 60461 11393 60559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 78744 63316 78820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50476 23932 50574 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8659 31998 8757 32096 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 66776 10140 66852 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 59704 16396 59780 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 17000 0 17076 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 75480 58284 75556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 45019 64057 45117 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 25976 0 26052 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 61251 64489 61349 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 42649 11393 42747 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 59704 58284 59780 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 75039 11393 75137 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 75471 11393 75569 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 46920 63316 46996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 64769 10961 64867 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 76568 3612 76644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 71521 11393 71619 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 38318 63403 38416 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 40688 12047 40786 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59867 54484 59965 54582 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47056 15912 75284 15988 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 53992 11364 54068 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 37400 75284 37476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46170 28052 46268 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 16184 9928 16260 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 52360 16396 52436 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44922 80916 45020 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71264 81464 75284 81540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 43112 816 43188 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 73473 63403 73571 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 60029 10961 60127 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 62968 64540 63044 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 83096 63044 83172 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 52632 10140 52708 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 47798 63403 47896 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 52632 75284 52708 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 74664 16396 74740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 41480 58284 41556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 42296 63316 42372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28424 18904 37748 18980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 34952 16396 35028 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 46613 12047 46711 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 31416 75284 31492 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 60819 10961 60917 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 71103 12047 71201 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 77384 75284 77460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 72352 28696 75284 28772 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 14280 18164 14356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35512 23094 35610 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 71879 10961 71977 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1360 35224 6876 35300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 62041 11393 62139 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 43000 85874 43098 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 59253 12047 59351 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 55352 0 55428 5244 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 5304 0 5380 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 67864 16396 67940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 1224 0 1300 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 31144 58284 31220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 59432 16396 59508 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49504 3672 75284 3748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 46920 58284 46996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 68408 0 68484 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 64600 0 64676 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40454 80344 40514 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 60819 11393 60917 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57907 28643 58005 28741 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71264 19720 75284 19796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24092 80916 24190 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18032 20149 18130 20247 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18714 80916 18812 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 5440 84456 62908 84532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 31960 6196 32036 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 41083 12047 41181 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 57278 12047 57376 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 37944 58284 38020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 38341 10961 38439 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 77928 16396 78004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36655 20592 36753 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 34136 10140 34212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 68361 64057 68459 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 38488 10140 38564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 53448 0 53524 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 20536 1980 20612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 58858 12047 58956 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 35539 64057 35637 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 20264 75284 20340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 43384 63316 43460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 69224 29512 75284 29588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 50184 16396 50260 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 58888 63316 58964 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24268 85036 24366 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52796 28052 52894 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28598 80344 28658 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 75752 63316 75828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 5168 81464 17484 81540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 60520 16396 60596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 33320 58284 33396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 78631 64489 78729 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 64411 64489 64509 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 53720 10140 53796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 9112 27820 9188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37903 20592 38001 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 46104 16396 46180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 48008 75284 48084 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71808 26248 75284 26324 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37334 80344 37394 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 41752 20808 41828 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 33864 16396 33940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8005 36761 8103 36859 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 33048 0 33124 16940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 47464 63316 47540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 58091 64057 58189 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 32379 64057 32477 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 3672 79832 16396 79908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 42840 75284 42916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 44661 11393 44759 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 53351 10961 53449 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 68000 88264 72564 88340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 40392 75284 40468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 35948 63403 36046 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 60248 16396 60324 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 44638 63403 44736 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 22168 75284 22244 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 48193 12047 48291 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 47464 0 47540 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 48588 12047 48686 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 55698 12047 55796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 58072 10140 58148 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 3400 32172 3476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 43081 64057 43179 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 52904 20808 52980 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41237 1461 41335 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 73848 73788 73924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 7573 36761 7671 36859 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 69509 64057 69607 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25840 7208 75284 7284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 38699 64057 38797 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 86088 17484 86164 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 64056 63316 64132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20536 23094 20634 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 78472 11364 78548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 66504 0 66580 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23020 23932 23118 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 59671 64057 59769 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 51544 64540 51620 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 40711 11393 40809 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 29512 6196 29588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 68680 10140 68756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 36040 16396 36116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 77051 64057 77149 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 68408 10140 68484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 40120 75284 40196 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 74664 63316 74740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1904 28968 16396 29044 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25528 23094 25626 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24954 80916 25052 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64029 83736 64127 83834 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 51339 64489 51437 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 78989 10961 79087 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 7365 1461 7463 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 30023 63403 30121 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 30872 63316 30948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 62152 10140 62228 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 31589 10961 31687 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35512 85874 35610 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 72216 16396 72292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 60520 63316 60596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 53723 12047 53821 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 42296 10140 42372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 72669 10961 72767 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 56079 64057 56177 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31194 80916 31292 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 51272 58284 51348 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44236 85036 44334 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 2040 0 2116 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 30799 64057 30897 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 57800 58284 57876 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 52088 16396 52164 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 47736 75284 47812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 49640 75284 49716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28012 23932 28110 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 36584 22984 36660 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 9656 0 9732 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 74681 10961 74779 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 58888 58284 58964 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 46599 64489 46697 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 55289 10961 55387 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 29512 63316 29588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 40293 63403 40391 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 33169 10961 33267 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 34408 5516 34484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 13205 1461 13303 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32342 28662 32402 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38682 28052 38780 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 69128 12047 69226 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 33592 58284 33668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 40392 63316 40468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 62399 64057 62497 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 35224 16396 35300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 38488 64540 38564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 53448 58284 53524 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 55896 0 55972 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 79560 10140 79636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41564 28052 41662 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 42568 75284 42644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26726 80344 26786 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 70731 64489 70829 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 63512 58284 63588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 41859 11393 41957 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 71089 64489 71187 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 50563 12047 50661 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 45809 64057 45907 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 31144 3264 31220 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 60461 64489 60559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 77818 63403 77916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 71672 0 71748 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 77112 16396 77188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 44744 16396 44820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 54141 64489 54239 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 37923 12047 38021 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 39032 75284 39108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 43928 75284 44004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 1496 75284 1572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 34368 12047 34466 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32911 20592 33009 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29260 23932 29358 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23606 80344 23666 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 38699 64489 38797 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 70312 16396 70388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 67048 16396 67124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 53720 58284 53796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36760 85874 36858 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 68719 10961 68817 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 77112 63316 77188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 71128 0 71204 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 6664 31356 6740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24092 28052 24190 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 45809 10961 45907 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 56168 58284 56244 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 69768 34408 75284 34484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46694 80344 46754 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54044 80916 54142 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54806 80344 54866 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 56093 12047 56191 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64328 85272 75284 85348 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 51272 10140 51348 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39244 85036 39342 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42426 28052 42524 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 59671 64489 59769 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 70856 0 70932 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 64056 16396 64132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 74249 11393 74347 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 74249 64057 74347 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 21896 9656 21972 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48666 28052 48764 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25568 7480 75284 7556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32966 80344 33026 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 79016 10140 79092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 72216 58284 72292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54536 5304 75284 5380 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 40279 64489 40377 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 68136 58284 68212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 37672 16396 37748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 18632 1844 18708 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 45560 13056 45636 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55375 20592 55473 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 77384 16396 77460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 65991 11393 66089 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26202 80916 26300 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 74392 16396 74468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 70584 63316 70660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 62808 12047 62906 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 50184 22984 50260 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 71128 58284 71204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 42568 11364 42644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 30023 12047 30121 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24155 21542 24253 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 10744 24752 10820 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 58463 63403 58561 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 21624 75284 21700 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19100 28052 19198 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27350 80344 27410 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19183 20592 19281 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 64872 63316 64948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17852 80916 17950 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54182 80344 54242 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 76633 63403 76731 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 52919 64057 53017 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 72896 88536 74876 88612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4624 19720 69844 19796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 11832 40740 11908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 67571 10961 67669 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 35158 12047 35256 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37820 28052 37918 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 19176 20808 19252 22380 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56984 20536 71204 20612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 62831 11393 62929 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 22440 75284 22516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71477 21857 71575 21955 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30470 28662 30530 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67249 34391 67347 34489 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 44243 12047 44341 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 62968 16396 63044 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 36040 6876 36116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 33592 17000 33668 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 2856 29860 2932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24230 28662 24290 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47804 28052 47902 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 49640 58284 49716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56848 16184 75284 16260 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45560 13464 75284 13540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 29628 63403 29726 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 32232 75284 32308 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 33959 10961 34057 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 69165 34368 69263 34466 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 66781 11393 66879 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 3861 80732 3959 80830 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44060 80916 44158 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 61251 64057 61349 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 49378 12047 49476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 77384 63316 77460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 78631 64057 78729 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 72216 73380 72292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 46241 64057 46339 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 26792 816 26868 17212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36572 28052 36670 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 47403 12047 47501 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19100 80916 19198 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 25160 75284 25236 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34252 23932 34350 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 76840 58284 76916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 67048 75284 67124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 48552 63316 48628 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52984 23094 53082 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 5576 0 5652 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 37133 12047 37231 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 54513 12047 54611 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 49096 22984 49172 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39930 80916 40028 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 57301 64489 57399 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34838 28662 34898 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 3944 0 4020 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 78472 63316 78548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 72311 11393 72409 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45446 28662 45506 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 37128 63316 37204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 31960 58284 32036 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20672 6392 75284 6468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40399 20592 40497 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 64783 12047 64881 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 78608 63403 78706 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 41480 75284 41556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 455 34014 553 34112 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52796 80916 52894 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45696 13192 75284 13268 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 45288 22984 45364 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74799 72714 74897 72812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 51000 10140 51076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 79003 63403 79101 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1904 34680 10140 34756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 77656 58284 77732 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 65688 0 65764 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29084 80916 29182 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 30813 63403 30911 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 54141 11393 54239 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 73304 16396 73380 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 83640 17484 83716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 54536 10140 54612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29084 28052 29182 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 74249 10961 74347 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44248 23094 44346 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 24616 7888 24692 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17466 28052 17564 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41647 20592 41745 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 50184 58284 50260 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31756 23932 31854 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51952 4488 75284 4564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 58072 0 58148 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34838 80344 34898 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 30441 64489 30539 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 5576 47404 5652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 42568 0 42644 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 55080 16396 55156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37883 21542 37981 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44236 23932 44334 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 53709 64489 53807 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44922 28052 45020 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52310 80344 52370 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 74392 63316 74468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 75039 64489 75137 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 71128 73380 71204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 77841 10961 77939 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 73101 64057 73199 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 58881 10961 58979 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 26792 20808 26868 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 51544 58284 51620 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 52919 11393 53017 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 76296 16396 76372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36186 80916 36284 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 67864 0 67940 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 70977 84956 71075 85054 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 59239 64489 59337 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34264 85874 34362 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 72488 16396 72564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 73576 75284 73652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 53351 11393 53449 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 32788 63403 32886 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 67139 64489 67237 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 70856 75284 70932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 44744 10140 44820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 68680 63316 68756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 12104 41828 12180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 65144 58284 65220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 40936 12104 41012 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 48552 75284 48628 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 46648 58284 46724 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 10472 35980 10548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 67320 16396 67396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 30872 10140 30948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 36343 12047 36441 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 61880 0 61956 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 50456 20808 50532 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 67320 0 67396 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32828 80916 32926 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 56488 63403 56586 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 37528 63403 37626 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30520 85874 30618 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 78608 12047 78706 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 29240 20808 29316 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 44661 64057 44759 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46170 80916 46268 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 54264 63316 54340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 81192 75284 81268 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 59976 10140 60052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 47464 75284 47540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 53176 5032 75284 5108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 48824 75284 48900 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 41480 0 41556 7692 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 67864 58284 67940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 35496 75284 35572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 44638 12047 44736 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 76238 63403 76336 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 32788 12047 32886 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46694 28662 46754 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 56440 63316 56516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 41208 0 41284 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 68361 64489 68459 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36635 21542 36733 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 55080 75284 55156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37996 85036 38094 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 31688 58284 31764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 56869 64057 56967 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 64388 12047 64486 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 68408 35224 75284 35300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45371 21542 45469 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39576 3400 75284 3476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31580 80916 31678 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 50981 64057 51079 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 72288 63403 72386 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 67139 11393 67237 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 55624 63316 55700 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 68408 36040 75284 36116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56540 80916 56638 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 5304 82824 58828 82900 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 54141 10961 54239 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 59432 0 59508 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1360 30600 16396 30676 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 41873 63403 41971 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 76296 58284 76372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67246 32795 67344 32893 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 61623 63403 61721 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57936 24888 75284 24964 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 28968 58284 29044 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30332 80916 30430 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 78213 12047 78311 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 15912 0 15988 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 79560 64540 79636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20431 20592 20529 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 70299 10961 70397 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 63189 11393 63287 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71477 19029 71575 19127 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30395 21542 30493 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 39576 816 39652 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 43656 58284 43732 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39206 28662 39266 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 7 18356 105 18454 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26588 28052 26686 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 59671 10961 59769 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22358 80344 22418 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 53351 64057 53449 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 79560 58284 79636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 54264 20808 54340 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 60792 75284 60868 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 67153 12047 67251 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 59160 0 59236 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 50981 10961 51079 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 2312 14628 2388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 65559 10961 65657 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22458 28052 22556 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 61608 63316 61684 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 38760 10140 38836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52410 28052 52508 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54044 28052 54142 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19962 80916 20060 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57392 26520 75284 26596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22358 28662 22418 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67681 35181 67779 35279 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39830 80344 39890 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 27608 19584 27684 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 36738 63403 36836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21896 9928 75284 10004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45308 28052 45406 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 62696 58284 62772 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 26520 22984 26596 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 77928 63316 78004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 64872 16396 64948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40316 28052 40414 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41178 80916 41276 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 32504 63316 32580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 68952 75284 69028 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39131 21542 39229 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 60520 75284 60596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27450 28052 27548 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 27064 8840 27140 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 76024 58284 76100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28424 19176 37340 19252 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 35553 63403 35651 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 55624 0 55700 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 76568 16396 76644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 61608 58284 61684 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 21352 0 21428 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 41069 11393 41167 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 64872 10140 64948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 37528 12047 37626 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1904 37944 10140 38020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 14824 7692 14900 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 8024 33668 8100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 74936 75284 75012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20486 28662 20546 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 48588 63403 48686 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52934 80344 52994 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 68719 11393 68817 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 50191 10961 50289 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 25432 1708 25508 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 32504 3536 32580 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49115 21542 49213 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 69509 11393 69607 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 43384 58284 43460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 45451 64489 45549 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 60438 12047 60536 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57120 21352 75284 21428 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 75247 87784 75345 87882 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4361 21184 4459 21282 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 35539 11393 35637 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 51771 11393 51869 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 55352 58284 55428 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 40392 16396 40468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18028 85036 18126 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 61228 12047 61326 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 51816 75284 51892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 36329 10961 36427 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 66781 64057 66879 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 30799 11393 30897 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 78472 58284 78548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30520 23094 30618 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 20536 0 20612 2116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 34952 64540 35028 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 53558 28662 53618 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 83096 75284 83172 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 39131 64057 39229 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23717 1461 23815 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 45832 63316 45908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 51771 64489 51869 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 58616 63316 58692 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 60819 64489 60917 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 39576 58284 39652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 44229 10961 44327 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 77841 64489 77939 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 75829 64057 75927 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 74120 16396 74196 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 61880 58284 61956 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 70299 64057 70397 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8659 29628 8757 29726 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 52632 22984 52708 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 51000 63316 51076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 78200 58284 78276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31718 28662 31778 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 62018 63403 62116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 59976 63316 60052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 72760 63316 72836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 19176 86496 19252 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 29784 58284 29860 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19862 80344 19922 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 73168 86904 75284 86980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18614 80344 18674 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 66504 10140 66580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18028 23932 18126 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 51272 0 51348 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 37119 10961 37217 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 51748 63403 51846 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33320 17272 75284 17348 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 30441 10961 30539 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 70977 87784 71075 87882 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 77656 16396 77732 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57302 28662 57362 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 45033 63403 45131 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 55352 75284 55428 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 4760 36796 4836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 49773 63403 49871 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 59239 10961 59337 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31768 23094 31866 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42988 85036 43086 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19584 2040 75284 2116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 32021 11393 32119 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 12376 43052 12452 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 30328 7284 30404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 680 5516 756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 50549 64489 50647 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 77818 12047 77916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 26520 10820 26596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1191 31774 1289 31872 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 53040 12648 75284 12724 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 38216 75284 38292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 64600 75284 64676 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 87720 71476 87796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 79016 58284 79092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 19448 15716 19524 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 56079 10961 56177 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 47389 11393 47487 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27221 1461 27319 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 46599 10961 46697 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 31998 12047 32096 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29147 21542 29245 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54107 21542 54205 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 75471 64489 75569 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 75843 63403 75941 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 46376 63316 46452 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 39576 75284 39652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 54513 63403 54611 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31580 28052 31678 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 55289 11393 55387 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47867 21542 47965 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 68408 58284 68484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 73032 10140 73108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 136 0 212 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11101 25232 11199 25330 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 81736 57468 81812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 43112 16396 43188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 54499 64057 54597 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 49759 11393 49857 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 67571 64057 67669 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 47031 64489 47129 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 13464 0 13540 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 61880 16396 61956 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35407 20592 35505 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 50728 64540 50804 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 56883 63403 56981 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 38699 10961 38797 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 71400 16396 71476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 40279 11393 40377 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 48552 16396 48628 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 31688 10140 31764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 77423 63403 77521 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 34749 64057 34847 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 3128 30948 3204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57302 80344 57362 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54220 23932 54318 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 58072 63316 58148 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50488 85874 50586 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 68952 16396 69028 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 67943 63403 68041 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 14280 0 14356 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 53448 63316 53524 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 45560 75284 45636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12037 1461 12135 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40504 85874 40602 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 39921 10961 40019 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 36856 63316 36932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33048 18088 75284 18164 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 41752 58284 41828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 30600 75284 30676 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 48280 63316 48356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 56984 0 57060 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 37944 16396 38020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 66232 63316 66308 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 21624 0 21700 9460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 39489 64057 39587 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 77409 64489 77507 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 60792 0 60868 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 37672 0 37748 13268 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 56168 16396 56244 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51162 80916 51260 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 58449 10961 58547 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 49912 58284 49988 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8008 32795 8106 32893 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 65968 12047 66066 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 38216 58284 38292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 63621 10961 63719 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29512 11016 75284 11092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 39489 64489 39587 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 78744 16396 78820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 78200 10140 78276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 17544 19584 17620 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 72760 75284 72836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 66232 16396 66308 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26726 28662 26786 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 42649 64489 42747 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 51000 16396 51076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 6392 12724 6468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 36040 63316 36116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 68338 63403 68436 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 64783 63403 64881 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 32379 10961 32477 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 32811 11393 32909 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21784 85874 21882 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 56488 12047 56586 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 43928 10140 44004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 70731 10961 70829 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26102 28662 26162 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 67592 63316 67668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 40293 12047 40391 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 49640 0 49716 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44336 10472 75284 10548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 30056 16396 30132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25403 21542 25501 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34139 21542 34237 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46744 23094 46842 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 36738 12047 36836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19862 28662 19922 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 53176 0 53252 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 69768 75284 69844 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50300 80916 50398 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 44229 64057 44327 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32442 28052 32540 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 70312 10140 70388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34252 85036 34350 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 50728 10140 50804 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25423 20592 25521 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 33048 63316 33124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 43453 63403 43551 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 47736 22984 47812 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 65960 10140 66036 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 41501 10961 41599 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 74936 63316 75012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 53176 16396 53252 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19276 23932 19374 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 41478 63403 41576 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 74936 0 75012 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71808 25976 75284 26052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41564 80916 41662 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 79421 64057 79519 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 51816 16396 51892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 3536 20536 17620 20612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 64056 10140 64132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 33864 58284 33940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 34408 16396 34484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 48983 63403 49081 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 73078 63403 73176 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34938 80916 35036 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1191 36254 1289 36352 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 34408 63316 34484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 51339 11393 51437 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 27880 22984 27956 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 67864 75284 67940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41178 28052 41276 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 35496 16396 35572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 21624 22984 21700 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 4216 0 4292 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 32379 11393 32477 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 40711 64057 40809 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39256 23094 39354 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18360 1768 75284 1844 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 49640 16396 49716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 16184 47676 16260 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 39304 75284 39380 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 14280 54536 16396 54612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55468 85036 55566 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 70584 58284 70660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19962 28052 20060 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 48969 11393 49067 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48566 80344 48626 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 70708 63403 70806 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 62831 64489 62929 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1191 38494 1289 38592 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 43081 11393 43179 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 62413 12047 62511 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 41480 22984 41556 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 65991 10961 66089 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 29784 16396 29860 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 3861 86388 3959 86486 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 62041 10961 62139 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 66758 12047 66856 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 58091 64489 58189 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19288 23094 19386 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 60792 16396 60868 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 46376 16396 46452 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48280 19176 75284 19252 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 62399 10961 62497 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 29628 12047 29726 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 26248 71204 26324 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23706 28052 23804 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 63512 10140 63588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 34136 75284 34212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33004 85036 33102 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 43439 64489 43537 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 13736 2312 13812 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 2040 28696 70524 28772 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 30328 58284 30404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 20264 0 20340 6196 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 37551 10961 37649 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 49912 75284 49988 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47984 20149 48082 20247 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28016 20149 28114 20247 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 36329 11393 36427 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39068 80916 39166 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56623 20592 56721 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 45832 16396 45908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 10744 29044 10820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 57256 0 57332 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18088 15096 75284 15172 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67246 30425 67344 30523 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 4216 35708 4292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 63240 75284 63316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 62413 63403 62511 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39256 85874 39354 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 74658 63403 74756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8659 35158 8757 35256 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 15640 0 15716 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 67048 63316 67124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 36312 10608 36388 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 45823 63403 45921 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 73891 11393 73989 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 30600 0 30676 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 24888 15580 24964 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34229 1461 34327 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 71498 63403 71596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 56712 75284 56788 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 20536 20808 20612 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48280 18904 75284 18980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 31960 16396 32036 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 49368 63316 49444 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 62041 64489 62139 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 45288 58284 45364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55468 23932 55566 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38901 1461 38999 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 29784 0 29860 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 41208 75284 41284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 38318 12047 38416 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 39304 0 39380 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 37400 58284 37476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 57301 64057 57399 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 2720 17816 19660 17892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 42024 10140 42100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18040 23094 18138 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 73459 10961 73557 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1191 29534 1289 29632 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 24616 4156 24692 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 71128 16396 71204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 38488 75284 38564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55760 5576 75284 5652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 4760 0 4836 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 54536 75284 54612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 75208 0 75284 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 37551 64489 37649 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 33169 64057 33267 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11424 26792 70252 26868 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 38713 12047 38811 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56154 28052 56252 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 40492 85036 40590 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 70040 58284 70116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 63512 16396 63588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 52538 63403 52636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 76568 63316 76644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 18360 75284 18436 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30725 1461 30823 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 26792 10820 26868 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 23256 816 23332 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 69768 58284 69844 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49190 80344 49250 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 47736 63316 47812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 50728 16396 50804 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 87448 75284 87524 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 58344 75284 58420 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 77423 12047 77521 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63648 83368 75284 83444 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 80104 73380 80180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 67320 10140 67396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 42296 16396 42372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 35768 58284 35844 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 11560 816 11636 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 25160 22984 25236 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 26248 0 26324 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 72488 58284 72564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 12920 6528 12996 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 50981 64489 51079 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 74263 63403 74361 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 35224 22984 35300 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20486 80344 20546 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55430 80344 55490 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 7208 19388 7284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 63993 63403 64091 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 34391 11393 34489 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 31688 63316 31764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 65201 11393 65299 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 57528 16396 57604 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 60792 10140 60868 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 57528 58284 57604 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 74936 16396 75012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25340 80916 25438 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57936 25704 75284 25780 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 47192 75284 47268 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 68733 12047 68831 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 71944 10140 72020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 73459 64489 73557 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 32232 0 32308 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44060 28052 44158 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 29651 10961 29749 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17990 28662 18050 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 65573 63403 65671 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 65144 10140 65220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 32776 22984 32852 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71400 80648 73788 80724 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 58344 58284 58420 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 45288 16396 45364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55480 23094 55578 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 30736 14008 75284 14084 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 77928 73380 78004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31718 80344 31778 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 23800 10820 23876 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71264 82824 75284 82900 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 47389 10961 47487 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 34408 58284 34484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 52129 64489 52227 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 55352 22984 55428 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 35158 63403 35256 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 58858 63403 58956 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 41083 63403 41181 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 75053 63403 75151 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 36312 10140 36388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 30328 63316 30404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 36761 11393 36859 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 39921 11393 40019 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 71893 63403 71991 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 32393 63403 32491 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51162 28052 51260 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56716 85036 56814 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71400 83640 75284 83716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33016 23094 33114 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 49912 63316 49988 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1360 32776 7284 32852 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 29512 58284 29588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 76238 12047 76336 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56984 6120 75284 6196 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 54931 64489 55029 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 71089 10961 71187 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1904 36856 6876 36932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31094 28662 31154 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 47031 10961 47129 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 72216 10140 72292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 64872 58284 64948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 54141 64057 54239 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 67592 58284 67668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 33048 20808 33124 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71400 86360 75284 86436 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 64328 75284 64404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 45288 75284 45364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56728 23094 56826 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 47192 16396 47268 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 3944 34484 4020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 48008 20808 48084 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 55624 10140 55700 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 56712 20808 56788 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 25432 20808 25508 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 59704 75284 59780 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 54264 16396 54340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 65991 64489 66089 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26102 80344 26162 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 15387 54484 15485 54582 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38352 18904 47676 18980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 59253 63403 59351 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26588 80916 26686 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 57673 12047 57771 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 67139 10961 67237 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 64328 0 64404 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 48824 16396 48900 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 77384 10140 77460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47318 80344 47378 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 6089 34368 6187 34466 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 55721 10961 55819 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 52088 75284 52164 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 52360 0 52436 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49240 23094 49338 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 66363 12047 66461 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 43384 12512 43460 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 34763 63403 34861 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39930 28052 40028 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 75752 58284 75828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 60792 63316 60868 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 50191 11393 50289 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 66349 10961 66447 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 58344 63316 58420 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 61336 0 61412 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 69918 12047 70016 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 66776 58284 66852 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35324 28052 35422 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71477 24685 71575 24783 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 52904 16396 52980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 52632 58284 52708 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 71400 0 71476 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 66595 35948 66693 36046 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 76261 64489 76359 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56054 28662 56114 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 36343 63403 36441 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4624 17000 32580 17076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 41480 63316 41556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 45019 11393 45117 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67249 35971 67347 36069 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 53558 80344 53618 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 49368 10140 49444 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 64056 0 64132 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 455 38494 553 38592 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54127 20592 54225 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 38760 63316 38836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 79421 11393 79519 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 35768 0 35844 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 60043 12047 60141 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34159 20592 34257 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 59976 58284 60052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44741 1461 44839 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 35181 11393 35279 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 7752 24284 7828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 30872 58284 30948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 68136 64540 68212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 8568 8780 8644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8008 32005 8106 32103 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 72760 58284 72836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 70040 75284 70116 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 52129 11393 52227 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17952 14824 75284 14900 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 69496 0 69572 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 31416 22984 31492 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35324 80916 35422 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 39848 16396 39924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 67048 0 67124 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74063 77194 74161 77292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 38341 11393 38439 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 8296 0 8372 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 64872 75284 64948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 78631 10961 78729 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 71944 16396 72020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 74392 0 74468 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 51816 10140 51892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 65559 64489 65657 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 48552 58284 48628 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 64328 16396 64404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56678 28662 56738 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 66595 36738 66693 36836 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 41069 64057 41167 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33590 28662 33650 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 78199 11393 78297 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 73848 10140 73924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 7480 18436 7556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52879 20592 52977 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 37909 11393 38007 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 79832 58284 79908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 48983 12047 49081 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 63240 0 63316 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 6685 29628 6783 29726 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 65178 63403 65276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74799 79434 74897 79532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 63189 64057 63287 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 69941 64489 70039 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 25704 11500 25780 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 64328 58284 64404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 61336 63316 61412 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 29651 64489 29749 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 9384 21700 9460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 73032 0 73108 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 49640 11364 49716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 42291 64489 42389 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 47821 64489 47919 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 36329 64489 36427 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21784 23094 21882 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38008 85874 38106 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 61608 75284 61684 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 52561 10961 52659 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 29651 64057 29749 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 38488 16396 38564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 48611 64057 48709 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 39131 11393 39229 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22927 20592 23025 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 71879 64489 71977 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 71893 12047 71991 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24230 80344 24290 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 52129 64057 52227 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 7573 35181 7671 35279 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 79288 75284 79364 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 11016 0 11092 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 76619 64057 76717 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51736 23094 51834 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 73848 0 73924 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 66781 64489 66879 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33690 80916 33788 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 73440 87720 75284 87796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 51771 64057 51869 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39244 23932 39342 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 37944 75284 38020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 52632 63316 52708 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 30418 12047 30516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 74392 10140 74468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 67139 64057 67237 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 37119 64489 37217 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 36040 4488 36116 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25340 28052 25438 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 19176 22984 19252 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29946 28052 30044 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 48179 64057 48277 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74799 70474 74897 70572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 49401 10961 49499 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 33601 64057 33699 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 56440 0 56516 15988 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 45019 10961 45117 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 63189 64489 63287 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 68680 58284 68756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 59160 11364 59236 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 51000 58284 51076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27974 80344 28034 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 70313 12047 70411 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 54118 63403 54216 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 47821 10961 47919 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 76296 63316 76372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24854 80344 24914 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 60833 63403 60931 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 70731 64057 70829 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37434 80916 37532 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 28968 71204 29044 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 74936 11364 75012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19045 1461 19143 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 75448 63403 75546 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 43384 10140 43460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49368 11832 75284 11908 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 68136 75284 68212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 71521 64057 71619 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 37128 10140 37204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50383 20592 50481 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 49912 16396 49988 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 33169 11393 33267 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 44744 75284 44820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 69523 63403 69621 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 42649 10961 42747 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 87176 75284 87252 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 66349 64057 66447 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52984 85874 53082 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24480 14280 75284 14356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 66595 31998 66693 32096 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 55080 0 55156 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 49096 0 49172 3340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 33578 63403 33676 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 62831 10961 62929 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 38760 0 38836 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 69496 16396 69572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28288 9384 75284 9460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 27336 0 27412 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 57528 75284 57604 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 40392 20808 40468 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 33320 16396 33396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1360 37400 11364 37476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 7752 0 7828 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 64600 58284 64676 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 30056 75284 30132 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 58449 11393 58547 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 74936 58284 75012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 60248 0 60324 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8008 30425 8106 30523 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 45428 63403 45526 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57120 21080 69980 21156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 62968 0 63044 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74799 77194 74897 77292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 34408 0 34484 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36856 10744 75284 10820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 42840 58284 42916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 27836 80916 27934 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 40711 10961 40809 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 63621 64489 63719 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 73032 58284 73108 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 30872 16396 30948 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 28968 22984 29044 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 408 0 484 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 60029 64489 60127 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 76296 75284 76372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56716 23932 56814 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 52904 58420 52980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 56869 10961 56967 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 50456 16396 50532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 45033 12047 45131 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46556 28052 46654 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 45451 64057 45549 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 35971 64489 36069 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49052 28052 49150 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 55624 16396 55700 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 72760 0 72836 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 57800 0 57876 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 70731 11393 70829 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51736 85874 51834 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 33169 64489 33267 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42326 80344 42386 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22907 21542 23005 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 49759 64489 49857 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 56984 10140 57060 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47942 80344 48002 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 75480 10140 75556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 37128 75284 37204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28389 1461 28487 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 65416 75284 65492 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 43574 80344 43634 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 48280 16456 75284 16532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41078 80344 41138 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 52143 12047 52241 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 9112 8704 9188 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 85000 3612 85076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 53992 16396 54068 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 46920 16396 46996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 45823 12047 45921 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 12648 44140 12724 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 64769 64489 64867 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 9656 15852 9732 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 30009 11393 30107 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 76619 64489 76717 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 69224 31960 75284 32036 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 56511 11393 56609 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 65144 63316 65220 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 56511 64057 56609 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 60792 58284 60868 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57402 80916 57500 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50476 85036 50574 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 56440 58284 56516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 67592 10140 67668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 29240 16396 29316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 57256 10140 57332 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41752 85874 41850 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 77409 10961 77507 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21381 1461 21479 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24885 1461 24983 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10869 1461 10967 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47992 85874 48090 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 37909 64489 38007 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 51544 10140 51620 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35462 28662 35522 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 65960 0 66036 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 53992 63316 54068 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35500 85036 35598 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 31208 63403 31306 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1904 35768 16396 35844 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4624 22712 17484 22788 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51686 28662 51746 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 33183 12047 33281 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 51353 12047 51451 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 49368 75284 49444 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 43439 64057 43537 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 59432 58284 59508 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 54264 75284 54340 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 46218 12047 46316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 42268 12047 42366 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 77051 10961 77149 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 60819 64057 60917 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 51000 75284 51076 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 58888 75284 58964 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8005 35971 8103 36069 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 20808 75284 20884 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 7208 0 7284 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 10200 20884 10276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 37128 16396 37204 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 45016 63316 45092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31643 21542 31741 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 16320 23256 71204 23332 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 455 31774 553 31872 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 75208 16396 75284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 23606 28662 23666 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 71944 58284 72020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39304 6664 75284 6740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51062 28662 51122 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 54536 58284 54612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 46648 20808 46724 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 34136 22984 34212 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 1768 0 1844 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 40664 10140 40740 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39830 28662 39890 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 76024 16396 76100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41740 23932 41838 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50438 28662 50498 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 23528 75284 23604 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 47389 64489 47487 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 59160 63316 59236 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36748 85036 36846 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 8024 14960 8100 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 69224 63316 69300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36710 28662 36770 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 61609 64489 61707 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 16456 11560 16532 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 68680 0 68756 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 11288 5984 11364 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29272 85874 29370 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 35971 64057 36069 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 66349 11393 66447 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 39304 16396 39380 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 15912 38292 15988 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 68408 63316 68484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 57659 10961 57757 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1904 32504 10140 32580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 68408 75284 68484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 51272 16396 51348 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 45809 11393 45907 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 45451 11393 45549 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 56440 10140 56516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 43928 16396 44004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 46376 5440 46452 15716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 68136 10140 68212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 65178 12047 65276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 34136 64540 34212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 30441 64057 30539 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 5848 816 5924 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 41501 64489 41599 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 60520 0 60596 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 37400 63316 37476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 52143 63403 52241 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 3536 19176 17348 19252 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 60029 11393 60127 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 75752 16396 75828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 14373 1461 14471 1559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 85272 63724 85348 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 58091 10961 58189 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 73891 64489 73989 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 25516 23932 25614 24030 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 67048 58284 67124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20348 28052 20446 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 52129 10961 52227 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 32379 64489 32477 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 56712 0 56788 5788 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 54264 0 54340 4972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 37672 10140 37748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 12376 0 12452 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 74681 64057 74779 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57936 27336 75284 27412 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 62152 75284 62228 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 32021 64057 32119 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 40936 16396 41012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 70856 10140 70932 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 39921 64489 40019 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 59648 63403 59746 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 69768 0 69844 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 74120 58284 74196 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 21352 17756 21428 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54220 85036 54318 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22982 28662 23042 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 59976 0 60052 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 58616 0 58692 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50728 3944 75284 4020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 69523 12047 69621 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 43871 64489 43969 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 31416 816 31492 7420 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 65688 10140 65764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 44744 0 44820 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 49096 10140 49172 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 13736 30132 13812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26776 85874 26874 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 76024 64540 76100 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 32504 75284 32580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 51062 80344 51122 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 69224 0 69300 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 51544 75284 51620 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46732 85036 46830 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 41480 16396 41556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 70299 11393 70397 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 62696 63316 62772 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 48179 10961 48277 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 46376 10140 46452 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 73891 10961 73989 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 71400 63316 71476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 41208 10140 41284 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 86360 70660 86436 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 17816 22984 17892 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 48008 58284 48084 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 19448 0 19524 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 57256 63316 57332 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17935 20592 18033 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 6936 816 7012 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 33320 75284 33396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 72311 10961 72409 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 63621 64057 63719 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 19288 85874 19386 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 43928 63316 44004 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 68000 32776 75284 32852 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 82552 18028 82628 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18614 28662 18674 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38352 19176 47268 19252 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 39848 58284 39924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50592 12104 75284 12180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 46599 64057 46697 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 73576 0 73652 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 80104 16396 80180 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 20808 17680 20884 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 39576 63316 39652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20536 85874 20634 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 65201 64489 65299 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 44744 58284 44820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 56712 58284 56788 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 67548 12047 67646 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 47464 16396 47540 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 62152 0 62228 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 62152 16396 62228 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 55303 63403 55401 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 72669 64489 72767 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45496 85874 45594 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42950 28662 43010 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 45019 64489 45117 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 56984 58284 57060 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49240 85874 49338 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 24344 75284 24420 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 60833 12047 60931 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 76261 64057 76359 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 44661 64489 44759 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 50456 11364 50532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 3672 41556 3748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 63512 75284 63588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 39921 64057 40019 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 42568 63316 42644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 67943 12047 68041 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 46070 80344 46130 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 26671 20592 26769 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 68000 30328 75284 30404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 62434 54468 62532 54566 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 61623 12047 61721 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 71944 0 72020 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 49640 63316 49716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 77051 64489 77149 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 67320 64540 67396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10744 79560 16396 79636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 33864 75284 33940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 39848 63316 39924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24854 28662 24914 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 73712 88808 75284 88884 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 49378 63403 49476 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 22458 80916 22556 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 18360 18904 27684 18980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 48280 10140 48356 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 56079 11393 56177 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45484 85036 45582 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 42296 75284 42372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 73848 63316 73924 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44143 20592 44241 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 51339 10961 51437 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 72311 64057 72409 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 86904 71748 86980 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 71089 11393 71187 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 8296 27548 8372 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 60461 10961 60559 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 12104 0 12180 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 52310 28662 52370 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 35224 58284 35300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47942 28662 48002 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 70977 82128 71075 82226 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 55080 10140 55156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 41752 11364 41828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 52360 75284 52436 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 38488 58284 38564 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8704 29512 11364 29588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 76619 11393 76717 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 39032 0 39108 6468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 36761 64489 36859 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 63240 58284 63316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 45560 63316 45636 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57800 25432 70252 25508 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 40936 75284 41012 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 455 29534 553 29632 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 78199 64057 78297 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49914 28052 50012 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 59976 16396 60052 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 65960 63316 66036 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 65416 16396 65492 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 28152 4156 28228 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 69496 63316 69572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 69918 63403 70016 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 55624 15640 75284 15716 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 37958 80344 38018 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 48969 64057 49067 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 78200 16396 78276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 43248 4216 75284 4292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 71808 20536 75284 20612 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 38216 16396 38292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 77028 12047 77126 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 61336 58284 61412 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8659 30418 8757 30516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 45016 58284 45092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 42568 58284 42644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 78472 73788 78548 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 3400 0 3476 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 29240 75284 29316 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 69151 10961 69249 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 47798 12047 47896 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 69151 64057 69249 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 80376 73244 80452 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 56054 80344 56114 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 58888 10140 58964 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 32442 80916 32540 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 31998 63403 32096 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 69224 58284 69300 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 66595 29628 66693 29726 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 53448 10140 53524 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 61608 16396 61684 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 46648 16396 46724 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 47736 58284 47812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 16456 40332 16532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 67929 64057 68027 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 16728 33396 16804 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 73078 12047 73176 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 37909 64057 38007 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 52088 10140 52164 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 6664 1768 6740 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 67320 58284 67396 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 62424 16396 62500 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 38713 63403 38811 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 55721 64057 55819 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 14824 2584 14900 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 15096 11500 15172 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 30418 63403 30516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 22168 11832 22244 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28016 8568 75284 8644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17852 28052 17950 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 44744 63316 44820 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 50981 11393 51079 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 75480 73380 75556 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 65573 12047 65671 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31768 85874 31866 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 76840 75284 76916 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 455 36254 553 36352 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 30009 10961 30107 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 24280 85874 24378 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 50300 28052 50398 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 22712 22984 22788 85892 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 33690 28052 33788 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 46241 11393 46339 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 43058 12047 43156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 84456 75284 84532 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 54118 12047 54216 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 34136 58284 34212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 33959 64057 34057 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 67592 75284 67668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 71672 10140 71748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 66232 58284 66308 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 20808 2312 75284 2388 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11424 26520 18028 26596 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 37119 11393 37217 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 42875 21542 42973 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 136 5924 212 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47992 23094 48090 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 72311 64489 72409 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 37128 5032 37204 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 35971 10961 36069 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 77409 64057 77507 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 62399 64489 62497 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 37944 0 38020 2796 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 5032 77112 10140 77188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 45809 64489 45907 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 36086 80344 36146 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4080 76568 10140 76644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41627 21542 41725 21640 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38582 28662 38642 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 79421 64489 79519 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 4488 0 4564 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 74249 64489 74347 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 35948 12047 36046 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 66504 75284 66580 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 74263 12047 74361 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 45016 10140 45092 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 54499 10961 54597 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 48969 10961 49067 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31824 7752 75284 7828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 28152 9384 28228 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 69496 10140 69572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 39304 58284 39380 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 70584 16396 70660 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41752 23094 41850 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 33183 63403 33281 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 71944 75284 72020 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8005 34391 8103 34489 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17990 80344 18050 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 48824 6256 48900 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 56440 75284 56516 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 63203 63403 63301 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 6685 31998 6783 32096 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 58344 0 58420 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 87992 75284 88068 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 31663 20592 31761 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 51748 12047 51846 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 29260 85036 29358 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 35496 58284 35572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 54536 0 54612 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 32232 58284 32308 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 44198 28662 44258 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 48969 64489 49067 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 34680 63316 34756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 70313 63403 70411 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 68408 16396 68484 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 58344 11364 58420 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21110 28662 21170 28722 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 47418 80916 47516 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 59432 75284 59508 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 1360 33048 11364 33124 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 58616 75284 58692 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 53992 0 54068 12588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 76568 58284 76644 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 63784 58284 63860 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39206 80344 39266 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 4624 25432 17484 25508 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 21110 80344 21170 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49228 85036 49326 85134 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 8005 35181 8103 35279 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 67571 64489 67669 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63920 29512 66580 29588 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 6392 0 6468 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 33592 10140 33668 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54264 12920 75284 12996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 66776 75284 66852 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 57800 63316 57876 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 74063 72714 74161 72812 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 58881 64489 58979 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 67246 29635 67344 29733 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 54808 0 54884 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 48008 16396 48084 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 38216 10140 38292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 73304 73380 73380 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28152 10200 75284 10276 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54906 28052 55004 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 67929 10961 68027 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 39068 28052 39166 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 64328 63316 64404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 24344 14280 24420 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 72216 63316 72292 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 69941 11393 70039 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 30813 12047 30911 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 27880 75284 27956 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 41702 80344 41762 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 71879 64057 71977 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 39503 63403 39601 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49135 20592 49233 20690 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 17000 58072 58284 58148 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 53658 80916 53756 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 66232 11364 66308 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 41501 11393 41599 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 38699 11393 38797 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 40279 64057 40377 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 50456 0 50532 3748 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 54232 85874 54330 85972 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28698 28052 28796 28150 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 58068 63403 58166 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 42296 0 42372 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 43439 10961 43537 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 75752 75284 75828 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 49052 80916 49150 81014 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 34680 75284 34756 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 952 75284 1028 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 48611 64489 48709 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 47031 11393 47129 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 61064 0 61140 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 64872 0 64948 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 39576 16396 39652 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 64769 64057 64867 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 77051 11393 77149 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 2584 0 2660 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 31231 64489 31329 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 56168 10140 56244 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63305 51353 63403 51451 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 8840 0 8916 89156 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 80920 75284 80996 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 12104 43384 16396 43460 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 34264 23094 34362 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 45446 80344 45506 80404 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 79421 10961 79519 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 35496 10140 35572 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 59024 65688 63316 65764 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 0 33864 11364 33940 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 35632 9112 75284 9188 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 65144 74392 73380 74468 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 72683 12047 72781 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 28024 23094 28122 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 63959 49401 64057 49499 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 64391 32021 64489 32119 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11949 73868 12047 73966 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 10863 57301 10961 57399 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 38008 23094 38106 23192 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 57120 24616 75284 24692 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal3 s 11295 68361 11393 68459 6 vdd
port 122 nsew power bidirectional abutment
rlabel metal4 s 55488 20808 55564 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 32011 82489 32109 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 71808 10548 71884 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 27472 4156 27548 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 32393 63675 32491 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 68816 75284 68892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41748 21210 41846 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 70977 80714 71075 80812 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 47872 22984 47948 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 58453 16730 58513 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 60928 0 61004 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 54931 64914 55029 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 37913 58682 37973 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50731 26479 50829 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 53351 64914 53449 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 66640 0 66716 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 83776 18028 83852 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 64464 10548 64540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 69918 63675 70016 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 39108 63675 39206 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4624 23936 17756 24012 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 73463 58682 73523 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8387 35948 8485 36046 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28094 84262 28192 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 272 18496 1844 18572 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 48588 11775 48686 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 32383 58682 32443 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49236 21210 49334 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 76677 10536 76775 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 43070 84262 43168 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 36448 75284 36524 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 27910 21979 28008 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 75344 63044 75420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31960 7072 75284 7148 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 86224 17484 86300 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68841 31998 68939 32096 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 62457 10536 62555 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 37264 10548 37340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 52984 22772 53082 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 69904 75284 69980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20213 47 20311 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 37264 75284 37340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 34753 16730 34813 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31838 84262 31936 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 59568 75284 59644 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 60112 0 60188 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 45968 11636 46044 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 32788 63675 32886 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 70731 10536 70829 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 46784 20808 46860 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 62403 16730 62463 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 53312 75284 53388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 50958 11775 51056 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 68733 63675 68831 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 56576 63044 56652 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 67153 11775 67251 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 32640 816 32716 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 37676 16730 37736 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 40256 22984 40332 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 11152 0 11228 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 38624 16184 38700 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 29920 0 29996 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 24208 75284 24284 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 76704 73380 76780 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 79783 16730 79843 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 64037 64914 64135 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8976 34272 10548 34348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 58690 16730 58750 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 67184 10548 67260 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 48588 63675 48686 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74799 73834 74897 73932 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 61613 58682 61673 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 41873 11775 41971 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 60270 16730 60330 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 81872 75284 81948 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 52224 10548 52300 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39576 3264 75284 3340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 24752 4156 24828 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51736 22772 51834 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 39131 64914 39229 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 37536 63044 37612 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 50553 58682 50613 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55723 26479 55821 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 13872 2312 13948 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 68960 58682 69020 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 39921 64914 40019 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 42100 58682 42160 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45560 13328 75284 13404 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 32437 64914 32535 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 31231 10536 31329 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39499 82489 39597 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 40528 20808 40604 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 31552 63044 31628 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 43000 22772 43098 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 2992 30948 3068 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49240 86196 49338 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 33184 63044 33260 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 32096 66308 32172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38352 20128 47676 20204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 50320 75284 50396 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 73440 0 73516 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 53040 75284 53116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 2992 17680 19660 17756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 38352 13328 38428 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 16320 47676 16396 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 19584 7480 19660 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 21670 21979 21768 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55760 5440 75284 5516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 49401 64914 49499 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 43520 63044 43596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 79546 16730 79606 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 272 4292 348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 58091 10536 58189 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 52133 58682 52193 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 86496 3612 86572 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 30566 16730 30626 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 60033 58682 60093 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 32368 3536 32444 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 66116 16730 66176 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35397 47 35495 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 57900 58682 57960 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 32897 21008 32995 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40500 21210 40598 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 51680 20808 51756 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 40293 11775 40391 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40747 82489 40845 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 48193 63675 48291 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 70357 64914 70455 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 69750 16730 69810 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23032 86196 23130 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 68000 0 68076 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 43081 10536 43179 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 60656 75284 60732 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 65563 58682 65623 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 72683 63675 72781 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 67933 16730 67993 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 73517 64914 73615 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 47156 16730 47216 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51806 24706 51904 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 36738 11775 36836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 78631 64914 78729 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 63648 63044 63724 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 80020 16730 80080 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 57664 63044 57740 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 55698 11775 55796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 71646 16730 71706 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 54931 10536 55029 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 54128 10548 54204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4488 17136 26324 17212 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 80512 75284 80588 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 56488 11775 56586 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 27200 0 27276 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 63746 58682 63806 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56848 16320 75284 16396 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 75471 64914 75569 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 61850 16730 61910 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 14416 0 14492 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 54672 75284 54748 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 46218 63675 46316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74799 71594 74897 71692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 22549 47 22647 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 36387 10536 36485 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35512 22772 35610 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 48183 58682 48243 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 63993 63675 64091 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20532 21210 20630 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 45968 0 46044 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24161 21008 24259 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8976 35088 10548 35164 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 31008 0 31084 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 44233 16730 44293 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 56488 63675 56586 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 42663 11775 42761 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 39493 58682 39553 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 73226 58682 73286 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 2720 17816 2796 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 34368 11775 34466 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 50048 0 50124 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74063 78314 74161 78412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 67728 75284 67804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 77520 10548 77596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 62016 10548 62092 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 37536 19584 37612 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 61228 63675 61326 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 47008 63675 47106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54232 86196 54330 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20606 24706 20704 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 13205 47 13303 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 3808 34484 3884 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 41616 22984 41692 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 13056 0 13132 6060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39142 21979 39240 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 43243 26479 43341 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 63920 0 63996 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 30464 63044 30540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1191 37374 1289 37472 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 68816 63044 68892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28024 86196 28122 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 57301 10536 57399 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28020 21210 28118 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 64773 16730 64833 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 36333 58682 36393 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 34990 58682 35050 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 79696 75284 79772 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 42976 75284 43052 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 60823 16730 60883 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 11696 21972 11772 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50488 22772 50586 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 67143 58682 67203 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 70540 58682 70600 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19174 21979 19272 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 70856 16730 70916 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55624 15504 75284 15580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 56304 75284 56380 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 60384 75284 60460 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 61744 63044 61820 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 52187 10536 52285 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28094 24706 28192 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33259 82489 33357 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 35553 11775 35651 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 36570 16730 36630 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 55760 0 55836 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 30192 2992 30268 15036 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 45696 10548 45772 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 70313 63675 70411 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25528 86196 25626 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 69151 10536 69249 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 49027 64914 49125 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 48960 75284 49036 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 64783 63675 64881 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 51397 64914 51495 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 55530 58682 55590 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 38080 75284 38156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 88672 72564 88748 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 49763 58682 49823 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 38896 22984 38972 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19448 6256 75284 6332 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 33578 11775 33676 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 54944 75284 55020 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55361 21008 55459 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 74800 0 74876 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 26112 75284 26188 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 40256 75284 40332 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 76160 75284 76236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 52224 75284 52300 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 14416 18164 14492 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 63648 0 63724 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 29776 58682 29836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 42890 58682 42950 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56728 86196 56826 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 37177 10536 37275 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 66758 11775 66856 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 6528 0 6604 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 46512 10548 46588 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 26662 21979 26760 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 49776 75284 49852 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 58208 10548 58284 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 84592 75284 84668 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35512 86196 35610 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 816 0 892 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 35553 63675 35651 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 47393 16730 47453 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 77028 11775 77126 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1191 35134 1289 35232 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 61060 58682 61120 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 79424 63044 79500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 41626 16730 41686 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 63920 10548 63996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68841 29628 68939 29726 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 43792 75284 43868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71400 84864 75284 84940 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 70708 63675 70806 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 29648 0 29724 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 62560 63044 62636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 72288 11775 72386 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74799 78314 74897 78412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 5304 82688 75284 82764 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 38713 11775 38811 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33320 17136 75284 17212 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 0 0 76 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 53160 58682 53220 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19358 24706 19456 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 79152 11636 79228 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 54908 11775 55006 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 51580 58682 51640 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 72352 28560 75284 28636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 38318 11775 38416 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30763 26479 30861 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 32368 75284 32444 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 59006 16730 59066 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 66096 63044 66172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 73984 0 74060 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 51771 64914 51869 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 71093 16730 71153 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 67571 64914 67669 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 43792 63044 43868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33086 84262 33184 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 35904 63044 35980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 4352 0 4428 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 59297 10536 59395 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 35360 22984 35436 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46814 84262 46912 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 67696 16730 67756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50558 84262 50656 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 50048 75284 50124 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 73868 63675 73966 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30763 82489 30861 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 64736 75284 64812 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8387 29628 8485 29726 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 30857 10536 30955 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 56320 16730 56380 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 62859 54469 62957 54567 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 66096 75284 66172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28267 82489 28365 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 47946 16730 48006 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30516 21210 30614 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 67943 63675 68041 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 77423 63675 77521 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 60823 58682 60883 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 47056 0 47132 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54475 82489 54573 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 78756 16730 78816 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 33728 10548 33804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 63430 58682 63490 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 57664 75284 57740 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 34017 10536 34115 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 66368 10548 66444 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 77966 16730 78026 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54475 26479 54573 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 34200 16730 34260 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35508 21210 35606 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 17952 20808 18028 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 32146 16730 32206 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 64536 58682 64596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 49504 63044 49580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 34272 20808 34348 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 47328 75284 47404 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 47872 63044 47948 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4624 26928 75284 27004 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 75887 64914 75985 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 31280 3264 31356 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 79230 16730 79290 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 73891 64914 73989 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 1632 6468 1708 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 48416 75284 48492 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19531 82489 19629 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 62413 63675 62511 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 6413 29628 6511 29726 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 16592 40332 16668 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11101 23818 11199 23916 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 57278 11775 57376 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 28288 0 28364 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 46241 10536 46339 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 46240 0 46316 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 50864 75284 50940 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 35971 64914 36069 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35582 24706 35680 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 42432 63724 42508 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 29376 75284 29452 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 56137 10536 56235 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71808 24752 75284 24828 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34507 26479 34605 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 45152 22984 45228 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46744 22772 46842 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 29104 816 29180 10684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 47992 86196 48090 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 53767 10536 53865 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44336 10336 75284 10412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 47878 21979 47976 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 42416 58682 42476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35582 84262 35680 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30590 84262 30688 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 52143 11775 52241 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 68777 64914 68875 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 76261 64914 76359 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 64192 75284 64268 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 72311 64914 72409 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 32640 75284 32716 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48235 26479 48333 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 36720 20808 36796 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 75344 75284 75420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 66781 10536 66879 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 29648 66308 29724 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 63203 63675 63301 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 27744 75284 27820 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 63920 75284 63996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 45077 10536 45175 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 49232 0 49308 3340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 69904 10548 69980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 3861 84974 3959 85072 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 45023 16730 45083 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 70977 86370 71075 86468 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 31824 0 31900 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 52496 75284 52572 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1191 32894 1289 32992 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 54141 10536 54239 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 54128 0 54204 4972 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 58480 63044 58556 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 40337 10536 40435 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 82416 75284 82492 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 47328 10548 47404 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 64411 64914 64509 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 13328 37204 13404 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 13192 54400 15172 54476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 72624 0 72700 88340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33016 22772 33114 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 33173 58682 33233 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 37676 58682 37736 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 36830 24706 36928 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 23392 4156 23468 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 29920 75284 29996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48235 82489 48333 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 74016 58682 74076 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 53227 82489 53325 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 62831 64914 62929 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40504 86196 40602 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 57120 75284 57196 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 44233 58682 44293 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 35632 75284 35708 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8976 29648 10548 29724 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 27064 17408 75284 17484 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 63376 75284 63452 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 44786 58682 44846 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 60877 10536 60975 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 18496 14552 18572 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 69941 64914 70039 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41822 84262 41920 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 78756 58682 78816 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 28986 16730 29046 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 31552 22984 31628 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 4352 35708 4428 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 31356 58682 31416 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28152 10064 75284 10140 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 5032 77248 73788 77324 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 60461 64914 60559 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 41310 16730 41370 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 40337 64914 40435 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 59480 16730 59540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 41072 75284 41148 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50558 24706 50656 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 53584 0 53660 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57936 24752 71204 24828 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 45152 75284 45228 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 38703 16730 38763 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74063 76074 74161 76172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 44880 0 44956 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 75072 63044 75148 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 53950 58682 54010 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 61251 64914 61349 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34229 47 34327 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 56873 16730 56933 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45377 21008 45475 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 60438 63675 60536 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 71498 11775 71596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 9520 0 9596 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 77423 11775 77521 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 32811 10536 32909 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 23120 11152 23196 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63512 83504 75284 83580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 45152 63044 45228 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 53723 11775 53821 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 79424 10548 79500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 66758 63675 66856 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 16048 9928 16124 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 70992 63044 71068 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 72352 75284 72428 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 68272 63044 68348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39304 6800 75284 6876 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 65280 75284 65356 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 49232 75284 49308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 34544 63724 34620 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 26384 75284 26460 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 61200 10548 61276 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30406 21979 30504 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 63104 63044 63180 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 31830 58682 31890 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 54944 10548 55020 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 63247 10536 63345 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 28832 2856 28908 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 41873 63675 41971 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 35181 64914 35279 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24480 14416 75284 14492 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 47984 19029 48082 19127 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 61200 75284 61276 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4361 25426 4459 25524 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74063 71594 74161 71692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 31552 75284 31628 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 52224 0 52300 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29272 86196 29370 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 45260 58682 45320 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 61744 75284 61820 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 13863 54484 13961 54582 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 43058 11775 43156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 47946 58682 48006 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35768 2720 75284 2796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 61228 11775 61326 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 3264 32172 3340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23275 82489 23373 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 75072 0 75148 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 26656 22984 26732 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 21488 17620 21564 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 71521 64914 71619 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 65178 11775 65276 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 46240 10548 46316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 53040 0 53116 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39499 26479 39597 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 52984 86196 53082 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 68361 10536 68459 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 41478 11775 41576 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 36343 63675 36441 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 74253 58682 74313 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 57664 10548 57740 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 18768 7752 18844 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 76238 63675 76336 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 55216 22984 55292 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 3536 19312 17348 19388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 9248 816 9324 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 53476 16730 53536 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 19040 71204 19116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 41616 63044 41692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28424 20128 37748 20204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 32383 16730 32443 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 34391 64914 34489 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 11696 15232 11772 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 43243 82489 43341 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34260 21210 34358 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 21784 86196 21882 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38078 84262 38176 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 56320 58682 56380 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 10064 0 10140 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 53227 26479 53325 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 54503 16730 54563 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 1360 0 1436 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 62560 0 62636 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 78336 10548 78412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 63104 10548 63180 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 48237 10536 48335 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 76704 3068 76780 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 3536 41556 3612 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 21854 24706 21952 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25771 26479 25869 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 47447 10536 47545 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45496 86196 45594 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 56304 0 56380 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 37536 75284 37612 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 67197 64914 67295 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 45696 63044 45772 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19358 84262 19456 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 16048 38292 16124 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56984 21488 75284 21564 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 52370 16730 52430 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 27019 26479 27117 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 55216 10548 55292 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 46784 75284 46860 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28016 19312 37340 19388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 43848 63675 43946 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 36760 22772 36858 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 47056 10548 47132 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 45823 11775 45921 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 58752 63044 58828 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 75843 63675 75941 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 56576 0 56652 5788 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 13056 6528 13132 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4624 18496 75284 18572 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 41863 58682 41923 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 60112 75284 60188 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 54128 20808 54204 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 54400 0 54476 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 62016 0 62092 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 57120 0 57196 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34150 21979 34248 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 16864 0 16940 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 71498 63675 71596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40574 24706 40672 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 51106 16730 51166 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 23936 22984 24012 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 64827 10536 64925 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 66407 10536 66505 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 35597 64914 35695 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 62288 75284 62364 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 42100 16730 42160 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 41127 10536 41225 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45492 21210 45590 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 50864 63044 50940 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 51408 0 51484 12044 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 42024 3808 75284 3884 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 75448 11775 75546 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 58881 64914 58979 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49096 272 75284 348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40574 84262 40672 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 53160 16730 53220 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 21760 71204 21836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46987 26479 47085 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 44243 63675 44341 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 35632 0 35708 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 31552 10548 31628 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20808 2448 75284 2524 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 55721 10536 55819 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 29104 22984 29180 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71808 27472 75284 27548 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 6528 13812 6604 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 72080 0 72156 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44491 82489 44589 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 43871 10536 43969 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 48183 16730 48243 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 66407 64914 66505 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 48611 10536 48709 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 58752 75284 58828 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 78440 16730 78500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 63104 75284 63180 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 36176 10608 36252 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 62560 11636 62636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 23936 0 24012 14356 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 52933 63675 53031 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 68723 58682 68783 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 42160 10548 42236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 58068 11775 58166 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 52768 22984 52844 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 54118 63675 54216 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 42707 10536 42805 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1904 33456 11636 33532 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 49773 63675 49871 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8387 32788 8485 32886 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 65552 75284 65628 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 20944 71612 21020 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34264 22772 34362 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 15776 54400 59644 54476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 42432 75284 42508 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 36992 63724 37068 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 16320 11560 16396 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 34000 22984 34076 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 28288 70388 28364 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 45813 58682 45873 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 39503 63675 39601 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 43497 10536 43595 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 47077 47 47175 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 19312 20808 19388 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 39503 11775 39601 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 85136 17756 85212 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56984 20400 75284 20476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 66116 58682 66176 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 25296 10820 25372 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 78993 16730 79053 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4080 80784 17620 80860 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 72120 16730 72180 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 68338 11775 68436 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 60461 10536 60559 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29376 11696 75284 11772 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 32912 7692 32988 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 74658 11775 74756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 70708 11775 70806 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55480 22772 55578 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 72624 63044 72700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 40256 63044 40332 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 39730 58682 39790 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 22576 0 22652 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34544 8160 75284 8236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 49027 10536 49125 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 67671 32005 67769 32103 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 57663 16730 57723 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 58480 75284 58556 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 72288 63675 72386 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 26776 22772 26874 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 68000 63044 68076 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41822 24706 41920 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 9520 21700 9596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28288 9520 75284 9596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 61376 16730 61436 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 55846 16730 55906 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 40688 11775 40786 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16709 47 16807 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20536 86196 20634 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 62041 64914 62139 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 31830 16730 31890 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49504 3536 75284 3612 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 41888 10548 41964 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 22848 22984 22924 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68952 29648 75284 29724 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55480 86196 55578 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 58091 64914 58189 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10869 47 10967 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20417 21008 20515 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35755 26479 35853 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49310 84262 49408 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 48420 58682 48480 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 43453 11775 43551 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 272 18224 4156 18300 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 36096 58682 36156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 39712 75284 39788 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49232 816 75284 892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 60087 64914 60185 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 8976 34892 9052 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30520 86196 30618 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 38624 63044 38700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50488 86196 50586 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 2448 14628 2524 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 78440 58682 78500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 31647 10536 31745 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 72080 73380 72156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 63247 64914 63345 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 39168 75284 39244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 51580 16730 51640 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 5168 0 5244 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 30013 16730 30073 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 76432 75284 76508 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 65991 64914 66089 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 30250 16730 30310 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 75888 10548 75964 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 47403 11775 47501 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31764 21210 31862 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 44661 10536 44759 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 48420 16730 48480 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 67184 63044 67260 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 41072 63044 41148 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 66590 58682 66650 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 47798 63675 47896 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 47992 22772 48090 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 75596 16730 75656 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 60438 11775 60536 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 36886 16730 36946 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33016 86196 33114 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 4624 0 4700 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 33963 16730 34023 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 42976 10548 43052 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 36641 21008 36739 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 59796 58682 59856 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18088 14960 75284 15036 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 52561 64914 52659 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71400 82144 75284 82220 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 59796 16730 59856 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56798 84262 56896 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 78257 64914 78355 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 4080 42644 4156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 78608 75284 78684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38901 47 38999 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 42996 21210 43094 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 44608 63044 44684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71477 20443 71575 20541 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 69567 64914 69665 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 15776 0 15852 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31838 24706 31936 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 42416 16730 42476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 43792 10548 43868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 36992 5032 37068 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 25568 1708 25644 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 74800 63044 74876 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44472 4896 75284 4972 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 31603 11775 31701 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 69513 58682 69573 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68952 32096 75284 32172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68000 36720 75284 36796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 61623 63675 61721 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 43248 4352 75284 4428 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71264 21216 75284 21292 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 59253 63675 59351 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 75616 10548 75692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 65573 11775 65671 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 31603 63675 31701 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 40046 16730 40106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 41073 16730 41133 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 41083 11775 41181 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 48960 0 49036 11636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 16592 0 16668 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 34000 63044 34076 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71808 19040 75284 19116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28389 47 28487 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25528 22772 25626 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57392 83776 63724 83852 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 9248 27820 9324 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 67671 30425 67769 30523 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 272 0 348 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 66353 58682 66413 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 44661 64914 44759 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 70176 63724 70252 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 3536 0 3612 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 23936 4156 24012 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 65617 10536 65715 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57120 85952 75284 86028 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1904 36992 10548 37068 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 74263 63675 74361 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18360 20128 27684 20204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 79783 58682 79843 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 62640 58682 62700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20672 6528 75284 6604 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 67548 11775 67646 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 22027 26479 22125 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 58216 58682 58276 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 32096 6468 32172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 73101 10536 73199 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 68544 0 68620 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 47872 75284 47948 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 87584 71476 87660 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 73168 75284 73244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31824 7616 75284 7692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 59006 58682 59066 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 63983 58682 64043 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39326 84262 39424 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 60043 63675 60141 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 62016 63044 62092 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 17926 21979 18024 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 47630 16730 47690 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38000 19029 38098 19127 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29515 26479 29613 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 58507 64914 58605 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 62018 63675 62116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 56848 63044 56924 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 78064 63724 78140 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45566 24706 45664 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 49504 75284 49580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 56927 10536 57025 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 51106 58682 51166 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 31998 63675 32096 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 69088 10548 69164 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1904 32368 10548 32444 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 63598 11775 63696 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29512 10880 75284 10956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 41501 64914 41599 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 49210 58682 49270 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 69128 63675 69226 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 69904 63044 69980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 37536 10548 37612 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 3536 20400 17620 20476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51816 12240 75284 12316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 64388 11775 64486 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 32096 63044 32172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 50320 22984 50396 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 63993 11775 64091 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20536 22772 20634 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56971 82489 57069 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34334 84262 34432 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 41072 10548 41148 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44248 22772 44346 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 50168 11775 50266 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 64220 16730 64280 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18040 86196 18138 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 46050 58682 46110 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 33410 58682 33470 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 22848 71612 22924 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 37264 63044 37340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 33183 11775 33281 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 30566 58682 30626 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48280 20128 75284 20204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35393 21008 35491 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 73712 0 73788 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 56093 63675 56191 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18040 22772 18138 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 34990 16730 35050 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39256 86196 39354 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 34816 4080 34892 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 69632 75284 69708 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 69360 75284 69436 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 34763 11775 34861 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57120 23936 70116 24012 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 44336 75284 44412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 10880 0 10956 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 50000 16730 50060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19284 21210 19382 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 68960 16730 69020 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 73984 10548 74060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19045 47 19143 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38008 86196 38106 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 65991 10536 66089 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 74658 63675 74756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 77467 10536 77565 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 35904 4488 35980 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 68170 16730 68230 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 73473 63675 73571 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 55056 16730 55116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 79398 11775 79496 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 52870 21979 52968 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 55347 64914 55445 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 66912 75284 66988 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 455 30654 553 30752 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50731 82489 50829 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 58858 11775 58956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 35306 16730 35366 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 76238 11775 76336 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 57717 10536 57815 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 1360 5924 1436 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 80784 3612 80860 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 72120 58682 72180 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 20400 0 20476 2116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 47600 75284 47676 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 74528 11636 74604 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25598 84262 25696 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 73700 16730 73760 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 28016 20808 28092 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7365 47 7463 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 74490 58682 74550 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 79421 10536 79519 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 62832 75284 62908 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 21780 21210 21878 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 68816 10548 68892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 30441 64914 30539 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8387 35158 8485 35256 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 65552 63044 65628 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54302 84262 54400 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 22032 9792 75284 9868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 41344 0 41420 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 60248 54400 62228 54476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 59648 63675 59746 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31768 86196 31866 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 47798 11775 47896 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 33601 64914 33699 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 50048 63044 50124 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 40836 16730 40896 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 50981 64914 51079 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 38352 63044 38428 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 79546 58682 79606 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33086 24706 33184 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 29460 58682 29520 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 53856 0 53932 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19531 26479 19629 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 70992 0 71068 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20422 21979 20520 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 42268 11775 42366 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 44638 11775 44736 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 23392 15504 23468 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25414 21979 25512 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71477 28927 71575 29025 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 37177 64914 37275 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 38940 16730 39000 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 44243 11775 44341 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 30067 10536 30165 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 42160 63044 42236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 32011 26479 32109 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 53584 10548 53660 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23275 26479 23373 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 70540 16730 70600 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54113 21008 54211 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 42432 0 42508 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 43443 16730 43503 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 79230 58682 79290 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 43070 24706 43168 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51622 21979 51720 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 55293 16730 55353 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 73984 63044 74060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 6256 12724 6332 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 56636 16730 56696 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 66912 0 66988 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 5984 0 6060 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 8160 816 8236 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 42160 12376 42236 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 72727 10536 72825 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 42291 64914 42389 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19169 21008 19267 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45739 26479 45837 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 67728 0 67804 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 70720 0 70796 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 13328 0 13404 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 29651 64914 29749 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31649 21008 31747 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41237 47 41335 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 76160 10548 76236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 34544 66988 34620 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 50048 11636 50124 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 38150 16730 38210 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 50592 0 50668 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 75833 16730 75893 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 19584 15716 19660 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 41344 63044 41420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 34807 10536 34905 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 65326 58682 65386 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71264 81328 75284 81404 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 56873 58682 56933 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 65008 75284 65084 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71264 84320 75284 84396 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34264 86196 34362 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 35088 63044 35164 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 58480 0 58556 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 34391 10536 34489 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 67696 58682 67756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 43520 10548 43596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 46218 11775 46316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 36720 0 36796 2660 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7583 29635 7681 29733 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 74528 75284 74604 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7 16940 105 17038 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 75888 63044 75964 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 7072 816 7148 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 46512 75284 46588 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 43497 64914 43595 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 72673 16730 72733 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 76386 16730 76446 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 34763 63675 34861 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 46657 64914 46755 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55723 82489 55821 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 49378 63675 49476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 60833 63675 60931 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 36646 21979 36744 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 48688 10548 48764 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 65552 10548 65628 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 77413 16730 77473 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 72910 58682 72970 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 72673 58682 72733 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 50168 63675 50266 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 65617 64914 65715 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28024 22772 28122 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 5984 48492 6060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 37123 58682 37183 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 73440 10548 73516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 39131 10536 39229 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 13600 0 13676 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 13872 30132 13948 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 39168 10548 39244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 48237 64914 48335 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25409 21008 25507 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44318 84262 44416 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 43443 58682 43503 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 55488 0 55564 5244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 67143 16730 67203 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 2720 28636 2796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 75280 16730 75340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 66368 0 66444 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 53856 63044 53932 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 22918 21979 23016 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20606 84262 20704 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 48960 10548 49036 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 35948 63675 36046 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 455 35134 553 35232 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25598 24706 25696 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 81056 17620 81132 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 75097 10536 75195 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54264 12784 75284 12860 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 77051 64914 77149 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 12240 41828 12316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 73440 85680 75284 85756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 41616 10548 41692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 44608 10548 44684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 55530 16730 55590 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 57426 16730 57486 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 57426 58682 57486 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 14960 11500 15036 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 72896 0 72972 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 65008 0 65084 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 43000 86196 43098 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 55216 63044 55292 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12240 78608 63044 78684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 37894 21979 37992 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 83232 17484 83308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 68272 10548 68348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 49776 0 49852 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 45424 816 45500 12860 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 73440 63044 73516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 56083 58682 56143 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 60112 10548 60188 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 43248 12512 43324 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 29104 75284 29180 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 11424 16124 11500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39326 24706 39424 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 47873 21008 47971 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 3264 0 3340 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33061 47 33159 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 62457 64914 62555 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 58752 10548 58828 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54302 24706 54400 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 54266 16730 54326 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58208 80784 75284 80860 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51806 84262 51904 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34145 21008 34243 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4080 77792 10548 77868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38080 13872 75284 13948 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46814 24706 46912 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40747 26479 40845 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 21381 47 21479 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39256 22772 39354 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 58507 10536 58605 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 51353 63675 51451 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 36570 58682 36630 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 45968 63044 46044 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 67728 10548 67804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 53054 84262 53152 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 50320 0 50396 3748 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 45867 64914 45965 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 70720 75284 70796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 6800 31356 6876 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 47447 64914 47545 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 35904 7284 35980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 81328 58964 81404 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 50316 16730 50376 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 30067 64914 30165 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 69632 63044 69708 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8432 34544 10548 34620 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 49526 16730 49586 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 56848 75284 56924 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4624 21216 69980 21292 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 53767 64914 53865 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 66096 0 66172 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 3861 79318 3959 79416 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 75344 10548 75420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 33728 63044 33804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24166 21979 24264 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 76860 16730 76920 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 21760 20808 21836 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 33456 63044 33532 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 36387 64914 36485 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 72727 64914 72825 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 52561 10536 52659 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54536 5168 75284 5244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 45033 63675 45131 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 52768 0 52844 12316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 48960 22984 49036 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64328 83776 75284 83852 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30520 22772 30618 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 51680 63044 51756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 36096 16730 36156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 53040 10548 53116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 76633 11775 76731 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 55846 58682 55906 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 70856 58682 70916 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 66640 75284 66716 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68000 35904 75284 35980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 75596 58682 75656 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 47031 10536 47129 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 57900 16730 57960 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 43206 58682 43266 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 14373 47 14471 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 67456 0 67532 87932 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 63104 0 63180 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 44064 75284 44140 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 75043 58682 75103 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 54266 58682 54326 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 73440 87584 75284 87660 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 52686 58682 52746 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 50607 10536 50705 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 42704 0 42780 8644 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 41888 3808 41964 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 50191 64914 50289 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8387 34368 8485 34466 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 69918 11775 70016 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 33227 10536 33325 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 57936 11636 58012 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 46240 75284 46316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 84048 17484 84124 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 71646 58682 71706 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 55760 63044 55836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 73078 63675 73176 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 42653 16730 42713 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 71808 75284 71884 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 39168 20808 39244 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 55216 0 55292 15308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 20128 0 20204 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 50864 0 50940 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 78213 11775 78311 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 61251 10536 61349 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 65800 58682 65860 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 68361 64914 68459 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 31356 16730 31416 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 79424 73788 79500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 42704 63044 42780 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 50958 63675 51056 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 4896 0 4972 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 72352 10548 72428 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 75843 11775 75941 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 39108 11775 39206 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 74307 10536 74405 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41633 21008 41731 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35632 9248 75284 9324 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 26776 86196 26874 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 49378 11775 49476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 36448 22984 36524 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1360 38624 10548 38700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 30803 16730 30863 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18283 26479 18381 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 43680 16730 43740 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 48736 58682 48796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 37733 47 37831 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 25024 0 25100 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 40688 63675 40786 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48008 19312 75284 19388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 67987 64914 68085 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 60384 10548 60460 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 70977 89198 71075 89296 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 69128 11775 69226 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 74528 0 74604 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 35948 11775 36046 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 61060 16730 61120 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11424 25296 18028 25372 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 61744 0 61820 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 44786 16730 44846 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 84864 70660 84940 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57800 28016 75284 28092 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4624 18224 39516 18300 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 71521 10536 71619 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 15232 10064 15308 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 64220 58682 64280 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18088 19312 27412 19388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 45424 75284 45500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 43112 8976 75284 9052 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 67380 16730 67440 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 43871 64914 43969 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 43520 0 43596 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 61667 64914 61765 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30401 21008 30499 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 5440 84320 58692 84396 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 59568 10548 59644 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24280 86196 24378 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48062 24706 48160 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 24208 20808 24284 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 66912 63044 66988 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 66640 11636 66716 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 7616 0 7692 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56971 26479 57069 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34507 82489 34605 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 66590 16730 66650 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 48736 16730 48796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 47056 15776 75284 15852 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 29376 10880 29452 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 67548 63675 67646 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12037 47 12135 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 75097 64914 75195 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71264 22576 75284 22652 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 16864 33396 16940 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 36830 84262 36928 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 53328 63675 53426 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 34272 63044 34348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29153 21008 29251 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1360 36176 75284 36252 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 19856 69844 19932 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 45576 16730 45636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 67671 32795 67769 32893 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28016 19029 28114 19127 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 71883 16730 71943 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 71264 75284 71340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 66867 36738 66965 36836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49368 11968 75284 12044 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 35632 63044 35708 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56798 24706 56896 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23028 21210 23126 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 31208 11775 31306 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 74800 10548 74876 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 52187 64914 52285 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18283 82489 18381 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 30803 58682 30863 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 64388 63675 64486 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 30736 75284 30812 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 544 5516 620 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 79421 64914 79519 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 62041 10536 62139 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 12240 0 12316 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 10336 35980 10412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 71147 64914 71245 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 71808 0 71884 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 67592 32912 75284 32988 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 48983 11775 49081 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 56576 75284 56652 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34408 8704 75284 8780 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 31593 58682 31653 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7583 32795 7681 32893 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 17921 21008 18019 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 73440 73380 73516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 65201 64914 65299 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 52977 10536 53075 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 63920 63044 63996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 62640 16730 62700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 47328 63044 47404 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 62288 0 62364 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 58463 11775 58561 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 61472 0 61548 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 54400 10548 54476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35398 21979 35496 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 66867 35158 66965 35256 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 79047 64914 79145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 78203 58682 78263 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 66363 63675 66461 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 76623 16730 76683 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 35360 75284 35436 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 88128 67260 88204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 31280 75284 31356 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 69513 16730 69573 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 62560 75284 62636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 42653 58682 42713 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 61472 75284 61548 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 39984 63044 40060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 76633 63675 76731 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54118 21979 54216 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68106 34391 68204 34489 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 41083 63675 41181 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 72352 63044 72428 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 25024 75284 25100 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 61376 58682 61436 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40385 21008 40483 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 45424 63044 45500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 77176 58682 77236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41638 21979 41736 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 34753 58682 34813 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 59296 63044 59372 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48280 544 75284 620 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 31008 75284 31084 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 31998 11775 32096 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 66640 63044 66716 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 59568 63044 59644 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 77841 10536 77939 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55366 21979 55464 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 33728 17000 33804 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 53950 16730 54010 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45739 82489 45837 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 9792 15852 9868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 28016 17212 28092 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 15504 0 15580 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 85952 17756 86028 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 36720 63044 36796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 46840 58682 46900 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 66906 16730 66966 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44248 86196 44346 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 77650 16730 77710 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44741 47 44839 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 43680 58682 43740 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 67380 58682 67440 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 70720 63044 70796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 70176 0 70252 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 36738 63675 36836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57936 19584 75284 19660 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 45867 10536 45965 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 61200 0 61276 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 36720 66308 36796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 59296 0 59372 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 45077 64914 45175 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 58216 16730 58276 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 21488 22984 21564 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30736 14144 75284 14220 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 455 37374 553 37472 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 48611 64914 48709 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71808 21760 75284 21836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 60384 63044 60460 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 83232 75284 83308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56984 5984 75284 6060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 66368 63044 66444 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 60112 63044 60188 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 33173 16730 33233 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45696 13056 75284 13132 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 68544 75284 68620 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 32936 58682 32996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 36343 11775 36441 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 55488 75284 55564 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 36565 47 36663 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 51353 11775 51451 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 51408 10548 51484 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 39984 10548 40060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 61200 63044 61276 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51617 21008 51715 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 65573 63675 65671 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 49232 20808 49308 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 55216 75284 55292 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 13600 10004 13676 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33259 26479 33357 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 34000 75284 34076 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 52923 58682 52983 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 27905 21008 28003 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 43206 16730 43266 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 59480 58682 59540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 11152 16940 11228 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 54503 58682 54563 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 31647 64914 31745 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 65280 10548 65356 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 70176 75284 70252 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 46603 16730 46663 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7583 30425 7681 30523 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 44608 75284 44684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 78213 63675 78311 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 22304 11832 22380 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 33963 58682 34023 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 31593 16730 31653 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 44336 12784 44412 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 14144 24012 14220 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 42881 21008 42979 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 21760 0 21836 9460 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 30813 11775 30911 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4361 16942 4459 17040 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28016 8432 75284 8508 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12395 54469 12493 54567 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 77792 3612 77868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 53584 75284 53660 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 66867 29628 66965 29726 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 35158 63675 35256 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 59024 63724 59100 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 70066 58682 70126 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 52933 11775 53031 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 36333 16730 36393 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 1904 12316 1980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 25840 11228 25916 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 56093 11775 56191 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 33726 58682 33786 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1904 28832 75284 28908 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4361 19770 4459 19868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24350 84262 24448 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 20944 816 21020 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 71893 11775 71991 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 65968 63675 66066 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 35158 11775 35256 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8976 36720 10548 36796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 37967 64914 38065 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19288 86196 19386 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 73226 16730 73286 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 86768 75284 86844 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 44470 16730 44530 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 45023 58682 45083 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 37360 16730 37420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 59840 0 59916 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 43848 11775 43946 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 12784 45364 12860 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 37808 22984 37884 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 53856 75284 53932 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 77818 11775 77916 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 34017 64914 34115 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 42704 10548 42780 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 73473 11775 73571 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 15541 47 15639 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 73517 10536 73615 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 53723 63675 53821 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 56083 16730 56143 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 35904 66308 35980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 74307 64914 74405 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 79047 10536 79145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 57673 11775 57771 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 48193 11775 48291 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 61613 16730 61673 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 65563 16730 65623 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57936 25568 70252 25644 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 61667 10536 61765 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 42886 21979 42984 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 27744 22984 27820 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25771 82489 25869 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1904 31280 10548 31356 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 50607 64914 50705 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 9792 0 9868 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 74016 16730 74076 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 68777 10536 68875 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 65178 63675 65276 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 38896 0 38972 6468 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 51408 63044 51484 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 52538 11775 52636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 37133 63675 37231 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 52133 16730 52193 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 13056 38020 13132 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 56848 10548 56924 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 69276 16730 69336 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 37123 16730 37183 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68000 88128 75284 88204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64029 85150 64127 85248 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 72624 10548 72700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 62288 63044 62364 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 67571 10536 67669 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 70448 10548 70524 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 26112 0 26188 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 54513 11775 54611 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 38466 58682 38526 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 59243 58682 59303 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 51343 16730 51403 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 71937 64914 72035 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 34807 64914 34905 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 53312 63044 53388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8976 32912 10548 32988 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23102 84262 23200 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 67456 63044 67532 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 27472 0 27548 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 25296 22984 25372 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54228 21210 54326 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 31208 63675 31306 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 40800 75284 40876 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 57301 64914 57399 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 50000 58682 50060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 44336 63044 44412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 62403 58682 62463 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74063 73834 74161 73932 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 73868 11775 73966 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 40256 0 40332 16804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 37923 11775 38021 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 39256 58682 39316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 53040 63044 53116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 64783 11775 64881 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 51343 58682 51403 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 45451 64914 45549 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 10880 22788 10956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 38341 10536 38439 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 8432 8780 8508 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1904 30192 75284 30268 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29268 21210 29366 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 26846 24706 26944 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 72436 58682 72496 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 48144 10548 48220 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 40800 10548 40876 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 59568 0 59644 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 48144 63044 48220 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 3128 25568 11500 25644 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 39168 0 39244 3068 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 52977 64914 53075 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 8976 8704 9052 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 22304 75284 22380 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 20400 22984 20476 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 70176 10548 70252 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57120 23120 75284 23196 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 65201 10536 65299 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 39547 10536 39645 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 39440 75284 39516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 34272 5788 34348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 77248 4156 77324 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 79003 63675 79101 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 49776 63044 49852 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 37923 63675 38021 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 38150 58682 38210 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 22913 21008 23011 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16456 22032 75284 22108 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46740 21210 46838 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 40283 16730 40343 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 51680 10548 51756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 52496 63044 52572 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 30250 58682 30310 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 42890 16730 42950 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 69151 64914 69249 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 75280 58682 75340 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41752 86196 41850 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 60033 16730 60093 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 19040 22984 19116 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 70303 16730 70363 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 75888 75284 75964 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 43248 75284 43324 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1360 34000 10548 34076 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 29776 16730 29836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 62166 58682 62226 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 62808 11775 62906 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 21665 21008 21763 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 63376 0 63452 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 39898 11775 39996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 7072 25100 7148 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64029 82322 64127 82420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 64736 63044 64812 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 15232 23196 15308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 65280 0 65356 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4624 22032 15988 22108 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 33601 10536 33699 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 30192 22984 30268 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 85408 75284 85484 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 23664 0 23740 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 37360 58682 37420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 73168 10548 73244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 57673 63675 57771 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 29628 63675 29726 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 33183 63675 33281 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 45428 63675 45526 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 39256 16730 39316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 65010 16730 65070 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 49504 0 49580 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 6800 1768 6876 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24350 24706 24448 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 40800 63044 40876 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31893 47 31991 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57936 27472 71204 27548 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 21216 4156 21292 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68106 35971 68204 36069 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38216 2992 75284 3068 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 74256 73380 74332 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 65552 0 65628 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 48688 75284 48764 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 71264 0 71340 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 59296 75284 59372 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 32620 58682 32680 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 75887 10536 75985 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 41072 12104 41148 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 60928 75284 61004 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 78880 73380 78956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24523 26479 24621 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 49401 10536 49499 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 46613 11775 46711 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 41478 63675 41576 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 30813 63675 30911 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1191 30654 1289 30752 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 64464 75284 64540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48245 47 48343 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 29628 11775 29726 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 38896 75284 38972 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 43520 75284 43596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 46050 16730 46110 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 56636 58682 56696 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8387 31998 8485 32096 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 47031 64914 47129 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7148 36761 7246 36859 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 5168 79968 73380 80044 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 45813 16730 45873 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 65326 16730 65386 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 74256 63044 74332 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 39730 16730 39790 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 35088 7284 35164 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 27221 47 27319 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 87040 75284 87116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 66353 16730 66413 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45382 21979 45480 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 64192 0 64268 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 88400 67124 88476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 5440 85680 71748 85756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 75053 63675 75151 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 71937 10536 72035 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 77467 64914 77565 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 58463 63675 58561 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 49763 16730 49823 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19288 22772 19386 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 17408 816 17484 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 68338 63675 68436 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 37133 11775 37231 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 70720 10548 70796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 37264 816 37340 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 61623 11775 61721 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 75043 16730 75103 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 55698 63675 55796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 32021 64914 32119 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45566 84262 45664 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 7888 33668 7964 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 26846 84262 26944 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 31280 63044 31356 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 75247 89200 75345 89298 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 25840 18224 25916 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 74256 10548 74332 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 58208 63044 58284 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 50592 75284 50668 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 35597 10536 35695 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 57392 75284 57468 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25524 21210 25622 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 39440 16048 39516 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 39712 18360 39788 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55550 24706 55648 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 54740 58682 54800 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 66867 31998 66965 32096 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 6197 47 6295 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 29648 63044 29724 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 58858 63675 58956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58208 28560 70524 28636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 79152 63044 79228 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 51408 22984 51484 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 50553 16730 50613 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 56848 0 56924 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 44880 75284 44956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 61391 54484 61489 54582 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 69632 0 69708 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 6413 31998 6511 32096 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 32902 21979 33000 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 43081 64914 43179 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 59671 10536 59769 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 71893 63675 71991 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 73304 88944 75284 89020 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 72683 11775 72781 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 43996 58682 44056 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 50592 10548 50668 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 5712 11092 5788 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 30464 20808 30540 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 77413 58682 77473 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 38703 58682 38763 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23717 47 23815 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 51397 10536 51495 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 85680 3204 85756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 11968 0 12044 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49310 24706 49408 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56609 21008 56707 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 51136 0 51212 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 7616 18436 7692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68000 35088 75284 35164 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 41888 63044 41964 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40800 16864 75284 16940 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 37003 26479 37101 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 32788 11775 32886 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 75053 11775 75151 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 35543 16730 35603 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 20400 1980 20476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 47056 63044 47132 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 75616 73380 75692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 62808 63675 62906 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 30464 66308 30540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 56032 10548 56108 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 45152 10548 45228 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 32912 66308 32988 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 67592 30464 75284 30540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 59243 16730 59303 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 66867 32788 66965 32886 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 51680 75284 51756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 5440 47404 5516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 71536 75284 71612 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 61850 58682 61910 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 26657 21008 26755 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 66912 10548 66988 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 79152 75284 79228 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 76070 58682 76130 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18110 24706 18208 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 49773 11775 49871 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 77818 63675 77916 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68106 36761 68204 36859 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 69360 0 69436 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 57392 63044 57468 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 55347 10536 55445 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 47630 58682 47690 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 58068 63675 58166 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 38080 63044 38156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 1088 75284 1164 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 46241 64914 46339 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 28267 26479 28365 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 56576 10548 56652 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 40256 10548 40332 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 67933 58682 67993 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 68000 10548 68076 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 70066 16730 70126 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 26772 21210 26870 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 70448 63044 70524 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 41626 58682 41686 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 57392 0 57468 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 66363 11775 66461 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 65800 16730 65860 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 32811 64914 32909 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 62288 10548 62364 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18360 1904 75284 1980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46784 16048 75284 16124 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 36856 10608 75284 10684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 41344 75284 41420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 5817 34368 5915 34466 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 62166 16730 62226 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 10608 24752 10684 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 72436 16730 72496 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 79003 11775 79101 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24280 22772 24378 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 37808 0 37884 2796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 73168 63044 73244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 65824 0 65900 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 38352 10548 38428 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 1904 0 1980 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 55056 58682 55116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 73168 0 73244 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4080 83504 17484 83580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 73463 16730 73523 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 38940 58682 39000 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 71536 63044 71612 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 62413 11775 62511 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 50864 10548 50940 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 55293 58682 55353 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 41888 75284 41964 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74063 80554 74161 80652 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 72311 10536 72409 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 34816 63044 34892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 60586 16730 60646 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 77028 63675 77126 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 47328 0 47404 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 60928 63044 61004 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 44287 64914 44385 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 40800 816 40876 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 57392 10548 57468 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 70992 73380 71068 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 66096 10548 66172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 70977 83542 71075 83640 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30725 47 30823 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48144 18224 75284 18300 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 45696 13056 45772 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 38352 75284 38428 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 43573 47 43671 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 57664 0 57740 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 61744 10548 61820 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 5712 816 5788 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 77176 16730 77236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 15776 39244 15852 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 74800 75284 74876 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 54557 64914 54655 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 59568 84048 75284 84124 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 36760 86196 36858 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 56032 75284 56108 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 408 17408 20476 17484 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 68486 16730 68546 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 69437 34368 69535 34466 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 21784 22772 21882 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 39493 16730 39553 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 68816 0 68892 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 32912 20808 32988 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 60384 0 60460 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30590 24706 30688 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 29651 10536 29749 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 70731 64914 70829 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 78608 4156 78684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 12512 44140 12588 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 53713 58682 53773 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 21488 0 21564 9732 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 53312 10548 53388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 82144 70660 82220 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 33227 64914 33325 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 54908 63675 55006 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44134 21979 44232 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 0 75284 76 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 42268 63675 42366 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 54944 63044 55020 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 71147 10536 71245 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 60087 10536 60185 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 64736 0 64812 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 43453 63675 43551 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8976 32096 10548 32172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 51952 0 52028 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 67943 11775 68041 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 67197 10536 67295 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 76976 63044 77052 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 38080 11636 38156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 2992 0 3068 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 63983 16730 64043 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 50563 11775 50661 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 2176 13540 2252 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38078 24706 38176 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 52224 63044 52300 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 50191 10536 50289 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1360 29648 6468 29724 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24276 21210 24374 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 48416 0 48492 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 3861 76490 3959 76588 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 18224 0 18300 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 51136 63724 51212 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 63746 16730 63806 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 52538 63675 52636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 72896 75284 72972 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 8704 0 8780 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 63598 63675 63696 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 72216 22848 75284 22924 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 80020 58682 80080 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 66867 35948 66965 36046 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 3861 82146 3959 82244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 46366 58682 46426 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 57663 58682 57723 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 36992 75284 37068 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29557 47 29655 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51736 86196 51834 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 73891 10536 73989 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 25568 816 25644 7012 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58208 80240 73244 80316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 30023 63675 30121 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18110 84262 18208 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 53328 11775 53426 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 29460 16730 29520 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 78336 75284 78412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 76070 16730 76130 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 73101 64914 73199 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 66906 58682 66966 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 63648 10548 63724 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 66368 75284 66444 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 8432 0 8508 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48280 16592 75284 16668 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 17136 2252 17212 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 52865 21008 52963 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 70448 0 70524 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 5168 44956 5244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 57110 58682 57170 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 77966 58682 78026 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51979 82489 52077 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49240 22772 49338 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74799 76074 74897 76172 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 21854 84262 21952 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 24480 7888 24556 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 70992 10548 71068 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 30736 10548 30812 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 53312 0 53388 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 44336 10548 44412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 60877 64914 60975 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 32912 0 32988 16804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29272 22772 29370 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 12784 816 12860 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 45696 75284 45772 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50369 21008 50467 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 52370 58682 52430 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71477 23271 71575 23369 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 71883 58682 71943 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 44638 63675 44736 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 66867 30418 66965 30516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 60270 58682 60330 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 51136 75284 51212 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 30023 11775 30121 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 62832 10548 62908 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 36761 64914 36859 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 45968 75284 46044 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 34334 24706 34432 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 62832 63044 62908 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8976 35904 10548 35980 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 52686 16730 52746 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 19856 17952 19932 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 544 0 620 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 65968 11775 66066 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 41917 64914 42015 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 64037 10536 64135 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 78608 11775 78706 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 40711 64914 40809 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 52923 16730 52983 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 28560 0 28636 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48008 5712 75284 5788 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 25296 0 25372 7284 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 75833 58682 75893 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44318 24706 44416 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18032 19029 18130 19127 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 42976 63044 43052 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 78993 58682 79053 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 73078 11775 73176 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 69276 58682 69336 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4361 28254 4459 28352 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 47872 10548 47948 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 42704 75284 42780 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 77650 58682 77710 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 26656 70252 26732 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24523 82489 24621 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 17680 22984 17756 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 44608 0 44684 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19584 2176 75284 2252 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11016 1632 75284 1708 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49126 21979 49224 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 68272 0 68348 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 62831 10536 62929 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 54944 0 55020 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 9701 47 9799 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 20128 17756 20204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 58690 58682 58750 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 77051 10536 77149 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 52496 0 52572 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 33456 75284 33532 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 49817 10536 49915 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 77792 63044 77868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 33184 0 33260 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 47393 58682 47453 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7 19772 105 19870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57392 25296 75284 25372 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 55760 75284 55836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 53351 10536 53449 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 62018 11775 62116 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 57278 63675 57376 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 64827 64914 64925 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 51896 58682 51956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 3808 0 3884 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 29920 10548 29996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 55303 63675 55401 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 74806 16730 74866 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 455 28414 553 28512 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 51680 0 51756 4292 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 39440 10548 39516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4361 22598 4459 22696 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23102 24706 23200 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 68486 58682 68546 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 38624 75284 38700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23032 22772 23130 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 35543 58682 35603 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 67184 75284 67260 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 62956 58682 63016 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 59253 11775 59351 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38008 22772 38106 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38004 21210 38102 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 65280 63044 65356 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 6256 0 6332 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44491 26479 44589 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 38757 10536 38855 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 41127 64914 41225 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 64536 16730 64596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 44470 58682 44530 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 7344 0 7420 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 35360 0 35436 2388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 37003 82489 37101 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1360 31824 75284 31900 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 52980 21210 53078 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 82960 58828 83036 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 49504 10548 49580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 33728 75284 33804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 69496 34272 75284 34348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29342 84262 29440 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 36448 0 36524 10412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 46840 16730 46900 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 455 32894 553 32992 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12104 24480 75284 24556 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 64736 10548 64812 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 59024 75284 59100 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 4624 43868 4700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 43058 63675 43156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 65824 75284 65900 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71264 82960 75284 83036 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51979 26479 52077 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63648 57936 75284 58012 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 14688 7692 14764 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 59024 10548 59100 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 34816 10548 34892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 46512 63044 46588 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56848 22576 69980 22652 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8387 30418 8485 30516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 47821 64914 47919 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 27200 1572 27276 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 34272 66308 34348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24344 14688 75284 14764 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1904 37808 10548 37884 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 66781 64914 66879 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 56511 10536 56609 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 59648 11775 59746 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 56032 0 56108 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 53040 12512 75284 12588 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 34816 75284 34892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49483 82489 49581 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 53856 10548 53932 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 2448 18768 75284 18844 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 59296 10548 59372 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 70303 58682 70363 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 54128 75284 54204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8976 30464 10548 30540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1191 28414 1289 28512 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 78064 75284 78140 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 41616 75284 41692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48062 84262 48160 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 37967 10536 38065 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 45260 16730 45320 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49121 21008 49219 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 2720 17952 25508 18028 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 40283 58682 40343 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 56576 22984 56652 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 41616 0 41692 3612 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31768 22772 31866 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 47008 11775 47106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 10064 20884 10140 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45496 22772 45594 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8533 47 8631 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23120 11424 75284 11500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 57936 0 58012 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 33973 11775 34071 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 78608 63675 78706 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 2040 28560 17076 28636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 48973 16730 49033 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 69904 0 69980 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 44287 10536 44385 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 46613 63675 46711 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 42160 75284 42236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 70313 11775 70411 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 43792 0 43868 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 48983 63675 49081 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 55303 11775 55401 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 47156 58682 47216 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 63203 11775 63301 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 26928 4156 27004 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 37889 21008 37987 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 2448 0 2524 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 20672 17620 20748 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 50563 63675 50661 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 38713 63675 38811 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 43996 16730 44056 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 30418 63675 30516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 41863 16730 41923 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 78336 63044 78412 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 57110 16730 57170 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46630 21979 46728 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 51748 63675 51846 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 41501 10536 41599 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 36756 21210 36854 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50484 21210 50582 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 55760 10548 55836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 36720 7284 36796 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33048 17952 75284 18028 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 11968 40740 12044 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56724 21210 56822 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40069 47 40167 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55476 21210 55574 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 44064 22984 44140 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 60656 0 60732 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 74490 16730 74550 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 77520 75284 77596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 32912 63044 32988 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 38757 64914 38855 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 78880 63044 78956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 51408 75284 51484 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 76623 58682 76683 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 64464 0 64540 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 73712 75284 73788 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 47988 21210 48086 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 48688 63044 48764 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 77841 64914 77939 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4080 86496 75284 86572 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 74263 11775 74361 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 45033 11775 45131 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 55550 84262 55648 84360 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 46657 10536 46755 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 72624 73788 72700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 35780 58682 35840 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 27019 82489 27117 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 33726 16730 33786 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 60043 11775 60141 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 54232 22772 54330 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 72910 16730 72970 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7148 34391 7246 34489 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 42704 22984 42780 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 76976 75284 77052 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 52768 75284 52844 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 34272 0 34348 7964 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 54513 63675 54611 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 11424 5984 11500 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 58752 0 58828 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 59840 75284 59916 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 24480 10276 24556 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 29223 16730 29283 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 59024 0 59100 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 60833 11775 60931 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 40528 75284 40604 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 75471 10536 75569 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 34544 0 34620 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 30441 10536 30539 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 51896 16730 51956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7148 35181 7246 35279 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 40046 58682 40106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 32437 10536 32535 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 30418 11775 30516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71477 26099 71575 26197 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 23664 75284 23740 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 76704 63044 76780 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 45424 10548 45500 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 68272 75284 68348 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 4896 76704 10548 76780 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 37551 10536 37649 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 17952 0 18028 1572 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 19312 0 19388 1844 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 31231 64914 31329 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 21216 10336 21292 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 22848 0 22924 10956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 36886 58682 36946 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 63621 64914 63719 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 74806 58682 74866 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 71093 58682 71153 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 64773 58682 64833 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 78064 10548 78140 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 50981 10536 51079 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 69523 11775 69621 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 30600 15232 75284 15308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 49776 10548 49852 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 56511 64914 56609 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12240 25840 18300 25916 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 76677 64914 76775 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51952 4624 75284 4700 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 67456 75284 67532 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 47056 75284 47132 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44244 21210 44342 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 87312 67668 87388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 38318 63675 38416 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 35088 66308 35164 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57664 25840 75284 25916 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 17136 11288 17212 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 58453 58682 58513 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 74799 80554 74897 80652 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 69088 0 69164 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39252 21210 39350 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 33973 63675 34071 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 49526 58682 49586 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 37808 75284 37884 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1904 34544 7284 34620 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 23256 11152 75284 11228 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 45909 47 46007 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 26053 47 26151 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 34200 58682 34260 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 38080 0 38156 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 56927 64914 57025 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 47403 63675 47501 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 1904 35632 10548 35708 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 39921 10536 40019 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 30736 63044 30812 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11101 26646 11199 26744 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 31040 16730 31100 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 74681 10536 74779 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 37551 64914 37649 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 73700 58682 73760 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 76386 58682 76446 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 55721 64914 55819 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 69088 75284 69164 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 75616 63724 75692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68000 34544 75284 34620 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 83504 3612 83580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 71330 16730 71390 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 53054 24706 53152 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 22027 82489 22125 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 51771 10536 51869 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29342 24706 29440 24804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 41344 11636 41420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 67456 10548 67532 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 8704 26732 8780 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56614 21979 56712 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56848 86224 75284 86300 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 75072 10548 75148 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 34516 58682 34576 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 35088 9112 35164 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 63430 16730 63490 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 30464 7692 30540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 42405 47 42503 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 58480 10548 58556 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 53476 58682 53536 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 25568 20808 25644 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58208 81056 75284 81132 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 65010 58682 65070 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 63648 75284 63724 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 34368 63675 34466 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 50316 58682 50376 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68272 87312 75284 87388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 67728 63724 67804 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 29223 58682 29283 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 36448 63044 36524 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 69523 63675 69621 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 44129 21008 44227 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 33456 0 33532 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 7888 14960 7964 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 48973 58682 49033 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 67671 29635 67769 29733 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 41917 10536 42015 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 17877 47 17975 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 49483 26479 49581 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 4080 0 4156 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16320 23392 75284 23468 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38251 82489 38349 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 51748 11775 51846 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 39547 64914 39645 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20779 82489 20877 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56728 22772 56826 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 45152 0 45228 13132 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 19040 0 19116 6060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 54128 63044 54204 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 46512 22984 46588 85892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 56032 63044 56108 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 80240 17076 80316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38080 19312 47268 19388 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 32096 0 32172 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 77792 73380 77868 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 54400 75284 54476 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 38251 26479 38349 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 22032 9656 22108 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 31654 21979 31752 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 76160 63044 76236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 52496 10548 52572 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 23120 17756 23196 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 64464 63044 64540 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41995 82489 42093 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 60928 10548 61004 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 51136 10548 51212 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 76860 58682 76920 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7583 32005 7681 32103 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 68106 35181 68204 35279 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 50320 63044 50396 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 48552 1360 75284 1436 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12240 46240 63044 46316 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 54740 16730 54800 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 46512 5440 46588 15716 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 78257 10536 78355 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 39898 63675 39996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 59671 64914 59769 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 69750 58682 69810 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 30736 0 30812 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 71400 87856 75012 87932 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 42707 64914 42805 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41752 22772 41850 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 71536 10548 71612 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 25840 7344 75284 7420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 37528 63675 37626 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 32393 11775 32491 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 50790 58682 50850 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 69567 10536 69665 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 75448 63675 75546 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 87856 70660 87932 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 63193 58682 63253 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 22576 17484 22652 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 28986 58682 29046 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 48960 63044 49036 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 32368 63044 32444 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 37528 11775 37626 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 42663 63675 42761 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 24752 0 24828 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 54672 0 54748 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40504 22772 40602 22870 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 74681 64914 74779 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 45428 11775 45526 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41888 7888 75284 7964 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 71808 63044 71884 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 42976 20808 43052 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 46366 16730 46426 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 37944 13600 75284 13676 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 59297 64914 59395 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 24885 47 24983 145 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29515 82489 29613 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 67973 88778 68071 88876 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 69088 63044 69164 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 8160 27548 8236 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 32146 58682 32206 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 67184 0 67260 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 5168 81600 17484 81676 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 72352 0 72428 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 33184 10548 33260 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 40711 10536 40809 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 48144 75284 48220 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 67987 10536 68085 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 5032 78608 10548 78684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 34516 16730 34576 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46987 82489 47085 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 41995 26479 42093 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 50790 16730 50850 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 38466 16730 38526 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 48688 6256 48764 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 26384 0 26460 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46744 86196 46842 86294 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 48144 0 48220 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 15504 46588 15580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 40293 63675 40391 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 57120 85136 75284 85212 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 20779 26479 20877 26577 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 35780 16730 35840 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 50592 63044 50668 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 1632 0 1708 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 20672 17680 20748 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 68733 11775 68831 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 50320 10548 50396 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 7148 35971 7246 36069 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 54118 11775 54216 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 51732 21210 51830 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 14688 0 14764 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 14144 6664 14220 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 37913 16730 37973 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11696 53584 63724 53660 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 40836 58682 40896 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 35755 82489 35853 82587 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 26928 17680 75284 17756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 36761 10536 36859 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 67153 63675 67251 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 56883 63675 56981 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 32620 16730 32680 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 69941 10536 70039 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 56883 11775 56981 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 51952 75284 52028 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 26928 8840 27004 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 77520 63044 77596 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 63193 16730 63253 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 29158 21979 29256 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 49210 16730 49270 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 31040 58682 31100 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 70448 73788 70524 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 5440 0 5516 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 73984 75284 74060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 68170 58682 68230 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 47600 19584 47676 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 39440 63044 39516 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 35971 10536 36069 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 19040 7616 24284 7692 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 41310 58682 41370 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 37808 63044 37884 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 62956 16730 63016 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 76261 10536 76359 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 40390 21979 40488 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 32936 16730 32996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 45823 63675 45921 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 39137 21008 39235 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 816 6468 892 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 8387 36738 8485 36836 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 40520 16730 40580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 12512 2040 12588 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 29920 63044 29996 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 52143 63675 52241 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 49817 64914 49915 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 33012 21210 33110 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 62016 75284 62092 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 45424 20808 45500 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 33184 75284 33260 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 3672 76976 10548 77052 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 11677 71103 11775 71201 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 79398 63675 79496 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 35306 58682 35366 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 74253 16730 74313 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 57936 63044 58012 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 53713 16730 53773 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 71536 0 71612 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 38341 64914 38439 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 36448 10548 36524 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 68000 75284 68076 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 54141 64914 54239 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 30013 58682 30073 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 58208 0 58284 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 17680 2524 17756 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 10608 29044 10684 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 46603 58682 46663 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 45576 58682 45636 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 42291 10536 42389 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 39168 63044 39244 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 39984 0 40060 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 54557 10536 54655 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 4896 36796 4972 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 10336 13736 10412 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 17952 27200 75284 27276 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 69632 10548 69708 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 45451 10536 45549 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 40520 58682 40580 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 70357 10536 70455 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 46625 21008 46723 21106 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 57717 64914 57815 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 71103 63675 71201 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 7344 19388 7420 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 14960 2584 15036 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 47821 10536 47919 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 74256 0 74332 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 60586 58682 60646 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 42432 10548 42508 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50728 4080 75284 4156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 3672 78880 10548 78956 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 68723 16730 68783 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 58881 10536 58979 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 66867 34368 66965 34466 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 18036 21210 18134 21308 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 75072 73788 75148 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 41073 58682 41133 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 56984 20672 75284 20748 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 32021 10536 32119 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 62832 0 62908 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 58208 75284 58284 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64736 39984 75284 40060 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 30857 64914 30955 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 78631 10536 78729 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 12376 74528 63044 74604 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 78203 16730 78263 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 50374 21979 50472 22077 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 58622 71330 58682 71390 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 64816 56137 64914 56235 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 35181 10536 35279 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 22032 4156 22108 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 64411 10536 64509 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 0 88944 70796 89020 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 10438 63621 10536 63719 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 2176 0 2252 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 16670 33410 16730 33470 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal4 s 1088 0 1164 89156 6 gnd
port 123 nsew ground bidirectional abutment
rlabel metal3 s 63577 33578 63675 33676 6 gnd
port 123 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 75296 89247
string LEFclass BLOCK
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 12810894
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sram_1rw1r_32_256_8_sky130.gds
string GDS_START 6490168
<< end >>
