magic
tech sky130B
timestamp 1644511149
<< properties >>
string GDS_END 3514710
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3514258
<< end >>
