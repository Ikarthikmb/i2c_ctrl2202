magic
tech sky130A
magscale 1 2
timestamp 1647938899
<< checkpaint >>
rect -12658 -11586 596582 715522
<< metal1 >>
rect 331214 702992 331220 703044
rect 331272 703032 331278 703044
rect 332502 703032 332508 703044
rect 331272 703004 332508 703032
rect 331272 702992 331278 703004
rect 332502 702992 332508 703004
rect 332560 702992 332566 703044
rect 318794 700952 318800 701004
rect 318852 700992 318858 701004
rect 413646 700992 413652 701004
rect 318852 700964 413652 700992
rect 318852 700952 318858 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 218974 700884 218980 700936
rect 219032 700924 219038 700936
rect 327902 700924 327908 700936
rect 219032 700896 327908 700924
rect 219032 700884 219038 700896
rect 327902 700884 327908 700896
rect 327960 700884 327966 700936
rect 314654 700816 314660 700868
rect 314712 700856 314718 700868
rect 478506 700856 478512 700868
rect 314712 700828 478512 700856
rect 314712 700816 314718 700828
rect 478506 700816 478512 700828
rect 478564 700816 478570 700868
rect 154114 700748 154120 700800
rect 154172 700788 154178 700800
rect 333238 700788 333244 700800
rect 154172 700760 333244 700788
rect 154172 700748 154178 700760
rect 333238 700748 333244 700760
rect 333296 700748 333302 700800
rect 137830 700680 137836 700732
rect 137888 700720 137894 700732
rect 329098 700720 329104 700732
rect 137888 700692 329104 700720
rect 137888 700680 137894 700692
rect 329098 700680 329104 700692
rect 329156 700680 329162 700732
rect 202782 700612 202788 700664
rect 202840 700652 202846 700664
rect 327718 700652 327724 700664
rect 202840 700624 327724 700652
rect 202840 700612 202846 700624
rect 327718 700612 327724 700624
rect 327776 700612 327782 700664
rect 327810 700612 327816 700664
rect 327868 700652 327874 700664
rect 527174 700652 527180 700664
rect 327868 700624 527180 700652
rect 327868 700612 327874 700624
rect 527174 700612 527180 700624
rect 527232 700612 527238 700664
rect 309134 700544 309140 700596
rect 309192 700584 309198 700596
rect 543458 700584 543464 700596
rect 309192 700556 543464 700584
rect 309192 700544 309198 700556
rect 543458 700544 543464 700556
rect 543516 700544 543522 700596
rect 89162 700476 89168 700528
rect 89220 700516 89226 700528
rect 338758 700516 338764 700528
rect 89220 700488 338764 700516
rect 89220 700476 89226 700488
rect 338758 700476 338764 700488
rect 338816 700476 338822 700528
rect 72970 700408 72976 700460
rect 73028 700448 73034 700460
rect 331858 700448 331864 700460
rect 73028 700420 331864 700448
rect 73028 700408 73034 700420
rect 331858 700408 331864 700420
rect 331916 700408 331922 700460
rect 24302 700340 24308 700392
rect 24360 700380 24366 700392
rect 342898 700380 342904 700392
rect 24360 700352 342904 700380
rect 24360 700340 24366 700352
rect 342898 700340 342904 700352
rect 342956 700340 342962 700392
rect 8110 700272 8116 700324
rect 8168 700312 8174 700324
rect 331950 700312 331956 700324
rect 8168 700284 331956 700312
rect 8168 700272 8174 700284
rect 331950 700272 331956 700284
rect 332008 700272 332014 700324
rect 317414 700204 317420 700256
rect 317472 700244 317478 700256
rect 397454 700244 397460 700256
rect 317472 700216 397460 700244
rect 317472 700204 317478 700216
rect 397454 700204 397460 700216
rect 397512 700204 397518 700256
rect 267642 700136 267648 700188
rect 267700 700176 267706 700188
rect 324958 700176 324964 700188
rect 267700 700148 324964 700176
rect 267700 700136 267706 700148
rect 324958 700136 324964 700148
rect 325016 700136 325022 700188
rect 322934 700068 322940 700120
rect 322992 700108 322998 700120
rect 348786 700108 348792 700120
rect 322992 700080 348792 700108
rect 322992 700068 322998 700080
rect 348786 700068 348792 700080
rect 348844 700068 348850 700120
rect 303614 696940 303620 696992
rect 303672 696980 303678 696992
rect 580166 696980 580172 696992
rect 303672 696952 580172 696980
rect 303672 696940 303678 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 304994 683204 305000 683256
rect 305052 683244 305058 683256
rect 580166 683244 580172 683256
rect 305052 683216 580172 683244
rect 305052 683204 305058 683216
rect 580166 683204 580172 683216
rect 580224 683204 580230 683256
rect 3418 683136 3424 683188
rect 3476 683176 3482 683188
rect 349154 683176 349160 683188
rect 3476 683148 349160 683176
rect 3476 683136 3482 683148
rect 349154 683136 349160 683148
rect 349212 683136 349218 683188
rect 300854 670760 300860 670812
rect 300912 670800 300918 670812
rect 580166 670800 580172 670812
rect 300912 670772 580172 670800
rect 300912 670760 300918 670772
rect 580166 670760 580172 670772
rect 580224 670760 580230 670812
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 351914 670732 351920 670744
rect 3568 670704 351920 670732
rect 3568 670692 3574 670704
rect 351914 670692 351920 670704
rect 351972 670692 351978 670744
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 350534 656928 350540 656940
rect 3476 656900 350540 656928
rect 3476 656888 3482 656900
rect 350534 656888 350540 656900
rect 350592 656888 350598 656940
rect 298094 643084 298100 643136
rect 298152 643124 298158 643136
rect 580166 643124 580172 643136
rect 298152 643096 580172 643124
rect 298152 643084 298158 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 353294 632108 353300 632120
rect 3476 632080 353300 632108
rect 3476 632068 3482 632080
rect 353294 632068 353300 632080
rect 353352 632068 353358 632120
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 580166 630680 580172 630692
rect 299624 630652 580172 630680
rect 299624 630640 299630 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 356054 618304 356060 618316
rect 3200 618276 356060 618304
rect 3200 618264 3206 618276
rect 356054 618264 356060 618276
rect 356112 618264 356118 618316
rect 296714 616836 296720 616888
rect 296772 616876 296778 616888
rect 580166 616876 580172 616888
rect 296772 616848 580172 616876
rect 296772 616836 296778 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 354674 605860 354680 605872
rect 3292 605832 354680 605860
rect 3292 605820 3298 605832
rect 354674 605820 354680 605832
rect 354732 605820 354738 605872
rect 293954 590656 293960 590708
rect 294012 590696 294018 590708
rect 579798 590696 579804 590708
rect 294012 590668 579804 590696
rect 294012 590656 294018 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 358814 579680 358820 579692
rect 3384 579652 358820 579680
rect 3384 579640 3390 579652
rect 358814 579640 358820 579652
rect 358872 579640 358878 579692
rect 295334 576852 295340 576904
rect 295392 576892 295398 576904
rect 580166 576892 580172 576904
rect 295392 576864 580172 576892
rect 295392 576852 295398 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 361574 565876 361580 565888
rect 3476 565848 361580 565876
rect 3476 565836 3482 565848
rect 361574 565836 361580 565848
rect 361632 565836 361638 565888
rect 292574 563048 292580 563100
rect 292632 563088 292638 563100
rect 579798 563088 579804 563100
rect 292632 563060 579804 563088
rect 292632 563048 292638 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 337378 553432 337384 553444
rect 3476 553404 337384 553432
rect 3476 553392 3482 553404
rect 337378 553392 337384 553404
rect 337436 553392 337442 553444
rect 288434 536800 288440 536852
rect 288492 536840 288498 536852
rect 580166 536840 580172 536852
rect 288492 536812 580172 536840
rect 288492 536800 288498 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 362954 527184 362960 527196
rect 3476 527156 362960 527184
rect 3476 527144 3482 527156
rect 362954 527144 362960 527156
rect 363012 527144 363018 527196
rect 289814 524424 289820 524476
rect 289872 524464 289878 524476
rect 580166 524464 580172 524476
rect 289872 524436 580172 524464
rect 289872 524424 289878 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 345658 514808 345664 514820
rect 3476 514780 345664 514808
rect 3476 514768 3482 514780
rect 345658 514768 345664 514780
rect 345716 514768 345722 514820
rect 287054 510620 287060 510672
rect 287112 510660 287118 510672
rect 580166 510660 580172 510672
rect 287112 510632 580172 510660
rect 287112 510620 287118 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 341518 501004 341524 501016
rect 3108 500976 341524 501004
rect 3108 500964 3114 500976
rect 341518 500964 341524 500976
rect 341576 500964 341582 501016
rect 284294 484372 284300 484424
rect 284352 484412 284358 484424
rect 580166 484412 580172 484424
rect 284352 484384 580172 484412
rect 284352 484372 284358 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 252646 478864 252652 478916
rect 252704 478904 252710 478916
rect 577590 478904 577596 478916
rect 252704 478876 577596 478904
rect 252704 478864 252710 478876
rect 577590 478864 577596 478876
rect 577648 478864 577654 478916
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 368014 474756 368020 474768
rect 3476 474728 368020 474756
rect 3476 474716 3482 474728
rect 368014 474716 368020 474728
rect 368072 474716 368078 474768
rect 285858 470568 285864 470620
rect 285916 470608 285922 470620
rect 579982 470608 579988 470620
rect 285916 470580 579988 470608
rect 285916 470568 285922 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 349062 462380 349068 462392
rect 3292 462352 349068 462380
rect 3292 462340 3298 462352
rect 349062 462340 349068 462352
rect 349120 462340 349126 462392
rect 299474 462204 299480 462256
rect 299532 462244 299538 462256
rect 325694 462244 325700 462256
rect 299532 462216 325700 462244
rect 299532 462204 299538 462216
rect 325694 462204 325700 462216
rect 325752 462204 325758 462256
rect 321370 462136 321376 462188
rect 321428 462176 321434 462188
rect 364334 462176 364340 462188
rect 321428 462148 364340 462176
rect 321428 462136 321434 462148
rect 364334 462136 364340 462148
rect 364392 462136 364398 462188
rect 234614 462068 234620 462120
rect 234672 462108 234678 462120
rect 330202 462108 330208 462120
rect 234672 462080 330208 462108
rect 234672 462068 234678 462080
rect 330202 462068 330208 462080
rect 330260 462068 330266 462120
rect 316586 462000 316592 462052
rect 316644 462040 316650 462052
rect 429194 462040 429200 462052
rect 316644 462012 429200 462040
rect 316644 462000 316650 462012
rect 429194 462000 429200 462012
rect 429252 462000 429258 462052
rect 313182 461932 313188 461984
rect 313240 461972 313246 461984
rect 462314 461972 462320 461984
rect 313240 461944 462320 461972
rect 313240 461932 313246 461944
rect 462314 461932 462320 461944
rect 462372 461932 462378 461984
rect 169754 461864 169760 461916
rect 169812 461904 169818 461916
rect 334894 461904 334900 461916
rect 169812 461876 334900 461904
rect 169812 461864 169818 461876
rect 334894 461864 334900 461876
rect 334952 461864 334958 461916
rect 311802 461796 311808 461848
rect 311860 461836 311866 461848
rect 494054 461836 494060 461848
rect 311860 461808 494060 461836
rect 311860 461796 311866 461808
rect 494054 461796 494060 461808
rect 494112 461796 494118 461848
rect 104894 461728 104900 461780
rect 104952 461768 104958 461780
rect 339678 461768 339684 461780
rect 104952 461740 339684 461768
rect 104952 461728 104958 461740
rect 339678 461728 339684 461740
rect 339736 461728 339742 461780
rect 307110 461660 307116 461712
rect 307168 461700 307174 461712
rect 558914 461700 558920 461712
rect 307168 461672 558920 461700
rect 307168 461660 307174 461672
rect 558914 461660 558920 461672
rect 558972 461660 558978 461712
rect 40034 461592 40040 461644
rect 40092 461632 40098 461644
rect 344370 461632 344376 461644
rect 40092 461604 344376 461632
rect 40092 461592 40098 461604
rect 344370 461592 344376 461604
rect 344428 461592 344434 461644
rect 272334 460912 272340 460964
rect 272392 460952 272398 460964
rect 578878 460952 578884 460964
rect 272392 460924 578884 460952
rect 272392 460912 272398 460924
rect 578878 460912 578884 460924
rect 578936 460912 578942 460964
rect 3878 460640 3884 460692
rect 3936 460680 3942 460692
rect 380894 460680 380900 460692
rect 3936 460652 380900 460680
rect 3936 460640 3942 460652
rect 380894 460640 380900 460652
rect 380952 460640 380958 460692
rect 3602 460572 3608 460624
rect 3660 460612 3666 460624
rect 383930 460612 383936 460624
rect 3660 460584 383936 460612
rect 3660 460572 3666 460584
rect 383930 460572 383936 460584
rect 383988 460572 383994 460624
rect 324958 460504 324964 460556
rect 325016 460544 325022 460556
rect 327074 460544 327080 460556
rect 325016 460516 327080 460544
rect 325016 460504 325022 460516
rect 327074 460504 327080 460516
rect 327132 460504 327138 460556
rect 329098 460504 329104 460556
rect 329156 460544 329162 460556
rect 336734 460544 336740 460556
rect 329156 460516 336740 460544
rect 329156 460504 329162 460516
rect 336734 460504 336740 460516
rect 336792 460504 336798 460556
rect 342898 460504 342904 460556
rect 342956 460544 342962 460556
rect 347774 460544 347780 460556
rect 342956 460516 347780 460544
rect 342956 460504 342962 460516
rect 347774 460504 347780 460516
rect 347832 460504 347838 460556
rect 308674 460436 308680 460488
rect 308732 460476 308738 460488
rect 327810 460476 327816 460488
rect 308732 460448 327816 460476
rect 308732 460436 308738 460448
rect 327810 460436 327816 460448
rect 327868 460436 327874 460488
rect 333238 460436 333244 460488
rect 333296 460476 333302 460488
rect 338114 460476 338120 460488
rect 333296 460448 338120 460476
rect 333296 460436 333302 460448
rect 338114 460436 338120 460448
rect 338172 460436 338178 460488
rect 345658 460436 345664 460488
rect 345716 460476 345722 460488
rect 366450 460476 366456 460488
rect 345716 460448 366456 460476
rect 345716 460436 345722 460448
rect 366450 460436 366456 460448
rect 366508 460436 366514 460488
rect 282914 460368 282920 460420
rect 282972 460408 282978 460420
rect 328546 460408 328552 460420
rect 282972 460380 328552 460408
rect 282972 460368 282978 460380
rect 328546 460368 328552 460380
rect 328604 460368 328610 460420
rect 331858 460368 331864 460420
rect 331916 460408 331922 460420
rect 341242 460408 341248 460420
rect 331916 460380 341248 460408
rect 331916 460368 331922 460380
rect 341242 460368 341248 460380
rect 341300 460368 341306 460420
rect 341518 460368 341524 460420
rect 341576 460408 341582 460420
rect 364886 460408 364892 460420
rect 341576 460380 364892 460408
rect 341576 460368 341582 460380
rect 364886 460368 364892 460380
rect 364944 460368 364950 460420
rect 255038 460300 255044 460352
rect 255096 460340 255102 460352
rect 308950 460340 308956 460352
rect 255096 460312 308956 460340
rect 255096 460300 255102 460312
rect 308950 460300 308956 460312
rect 309008 460300 309014 460352
rect 322842 460300 322848 460352
rect 322900 460340 322906 460352
rect 331214 460340 331220 460352
rect 322900 460312 331220 460340
rect 322900 460300 322906 460312
rect 331214 460300 331220 460312
rect 331272 460300 331278 460352
rect 331950 460300 331956 460352
rect 332008 460340 332014 460352
rect 345934 460340 345940 460352
rect 332008 460312 345940 460340
rect 332008 460300 332014 460312
rect 345934 460300 345940 460312
rect 345992 460300 345998 460352
rect 349062 460300 349068 460352
rect 349120 460340 349126 460352
rect 371234 460340 371240 460352
rect 349120 460312 371240 460340
rect 349120 460300 349126 460312
rect 371234 460300 371240 460312
rect 371292 460300 371298 460352
rect 250254 460232 250260 460284
rect 250312 460272 250318 460284
rect 321554 460272 321560 460284
rect 250312 460244 321560 460272
rect 250312 460232 250318 460244
rect 321554 460232 321560 460244
rect 321612 460232 321618 460284
rect 337378 460232 337384 460284
rect 337436 460272 337442 460284
rect 360194 460272 360200 460284
rect 337436 460244 360200 460272
rect 337436 460232 337442 460244
rect 360194 460232 360200 460244
rect 360252 460232 360258 460284
rect 277118 460164 277124 460216
rect 277176 460204 277182 460216
rect 378042 460204 378048 460216
rect 277176 460176 378048 460204
rect 277176 460164 277182 460176
rect 378042 460164 378048 460176
rect 378100 460164 378106 460216
rect 281442 460096 281448 460148
rect 281500 460136 281506 460148
rect 415026 460136 415032 460148
rect 281500 460108 415032 460136
rect 281500 460096 281506 460108
rect 415026 460096 415032 460108
rect 415084 460096 415090 460148
rect 280062 460028 280068 460080
rect 280120 460068 280126 460080
rect 580074 460068 580080 460080
rect 280120 460040 580080 460068
rect 280120 460028 280126 460040
rect 580074 460028 580080 460040
rect 580132 460028 580138 460080
rect 269022 459960 269028 460012
rect 269080 460000 269086 460012
rect 577406 460000 577412 460012
rect 269080 459972 577412 460000
rect 269080 459960 269086 459972
rect 577406 459960 577412 459972
rect 577464 459960 577470 460012
rect 234338 459892 234344 459944
rect 234396 459932 234402 459944
rect 248046 459932 248052 459944
rect 234396 459904 248052 459932
rect 234396 459892 234402 459904
rect 248046 459892 248052 459904
rect 248104 459892 248110 459944
rect 264514 459892 264520 459944
rect 264572 459932 264578 459944
rect 580626 459932 580632 459944
rect 264572 459904 580632 459932
rect 264572 459892 264578 459904
rect 580626 459892 580632 459904
rect 580684 459892 580690 459944
rect 4982 459824 4988 459876
rect 5040 459864 5046 459876
rect 369854 459864 369860 459876
rect 5040 459836 369860 459864
rect 5040 459824 5046 459836
rect 369854 459824 369860 459836
rect 369912 459824 369918 459876
rect 3326 459756 3332 459808
rect 3384 459796 3390 459808
rect 375926 459796 375932 459808
rect 3384 459768 375932 459796
rect 3384 459756 3390 459768
rect 375926 459756 375932 459768
rect 375984 459756 375990 459808
rect 3786 459688 3792 459740
rect 3844 459728 3850 459740
rect 379146 459728 379152 459740
rect 3844 459700 379152 459728
rect 3844 459688 3850 459700
rect 379146 459688 379152 459700
rect 379204 459688 379210 459740
rect 234430 459620 234436 459672
rect 234488 459660 234494 459672
rect 243262 459660 243268 459672
rect 234488 459632 243268 459660
rect 234488 459620 234494 459632
rect 243262 459620 243268 459632
rect 243320 459620 243326 459672
rect 327902 459620 327908 459672
rect 327960 459660 327966 459672
rect 333330 459660 333336 459672
rect 327960 459632 333336 459660
rect 327960 459620 327966 459632
rect 333330 459620 333336 459632
rect 333388 459620 333394 459672
rect 234522 459552 234528 459604
rect 234580 459592 234586 459604
rect 238846 459592 238852 459604
rect 234580 459564 238852 459592
rect 234580 459552 234586 459564
rect 238846 459552 238852 459564
rect 238904 459552 238910 459604
rect 327718 459552 327724 459604
rect 327776 459592 327782 459604
rect 331766 459592 331772 459604
rect 327776 459564 331772 459592
rect 327776 459552 327782 459564
rect 331766 459552 331772 459564
rect 331824 459552 331830 459604
rect 338758 459552 338764 459604
rect 338816 459592 338822 459604
rect 342806 459592 342812 459604
rect 338816 459564 342812 459592
rect 338816 459552 338822 459564
rect 342806 459552 342812 459564
rect 342864 459552 342870 459604
rect 360654 459552 360660 459604
rect 360712 459592 360718 459604
rect 374362 459592 374368 459604
rect 360712 459564 374368 459592
rect 360712 459552 360718 459564
rect 374362 459552 374368 459564
rect 374420 459552 374426 459604
rect 231210 459144 231216 459196
rect 231268 459184 231274 459196
rect 399662 459184 399668 459196
rect 231268 459156 399668 459184
rect 231268 459144 231274 459156
rect 399662 459144 399668 459156
rect 399720 459144 399726 459196
rect 231118 459076 231124 459128
rect 231176 459116 231182 459128
rect 404354 459116 404360 459128
rect 231176 459088 404360 459116
rect 231176 459076 231182 459088
rect 404354 459076 404360 459088
rect 404412 459076 404418 459128
rect 378042 459008 378048 459060
rect 378100 459048 378106 459060
rect 580810 459048 580816 459060
rect 378100 459020 580816 459048
rect 378100 459008 378106 459020
rect 580810 459008 580816 459020
rect 580868 459008 580874 459060
rect 321554 458940 321560 458992
rect 321612 458980 321618 458992
rect 580258 458980 580264 458992
rect 321612 458952 580264 458980
rect 321612 458940 321618 458952
rect 580258 458940 580264 458952
rect 580316 458940 580322 458992
rect 283466 458872 283472 458924
rect 283524 458912 283530 458924
rect 580166 458912 580172 458924
rect 283524 458884 580172 458912
rect 283524 458872 283530 458884
rect 580166 458872 580172 458884
rect 580224 458872 580230 458924
rect 270402 458804 270408 458856
rect 270460 458844 270466 458856
rect 577314 458844 577320 458856
rect 270460 458816 577320 458844
rect 270460 458804 270466 458816
rect 577314 458804 577320 458816
rect 577372 458804 577378 458856
rect 267642 458736 267648 458788
rect 267700 458776 267706 458788
rect 574830 458776 574836 458788
rect 267700 458748 574836 458776
rect 267700 458736 267706 458748
rect 574830 458736 574836 458748
rect 574888 458736 574894 458788
rect 262858 458668 262864 458720
rect 262916 458708 262922 458720
rect 574738 458708 574744 458720
rect 262916 458680 574744 458708
rect 262916 458668 262922 458680
rect 574738 458668 574744 458680
rect 574796 458668 574802 458720
rect 257982 458600 257988 458652
rect 258040 458640 258046 458652
rect 577774 458640 577780 458652
rect 258040 458612 577780 458640
rect 258040 458600 258046 458612
rect 577774 458600 577780 458612
rect 577832 458600 577838 458652
rect 3234 458532 3240 458584
rect 3292 458572 3298 458584
rect 372798 458572 372804 458584
rect 3292 458544 372804 458572
rect 3292 458532 3298 458544
rect 372798 458532 372804 458544
rect 372856 458532 372862 458584
rect 3970 458464 3976 458516
rect 4028 458504 4034 458516
rect 377582 458504 377588 458516
rect 4028 458476 377588 458504
rect 4028 458464 4034 458476
rect 377582 458464 377588 458476
rect 377640 458464 377646 458516
rect 3694 458396 3700 458448
rect 3752 458436 3758 458448
rect 382274 458436 382280 458448
rect 3752 458408 382280 458436
rect 3752 458396 3758 458408
rect 382274 458396 382280 458408
rect 382332 458396 382338 458448
rect 3510 458328 3516 458380
rect 3568 458368 3574 458380
rect 387058 458368 387064 458380
rect 3568 458340 387064 458368
rect 3568 458328 3574 458340
rect 387058 458328 387064 458340
rect 387116 458328 387122 458380
rect 3418 458260 3424 458312
rect 3476 458300 3482 458312
rect 391934 458300 391940 458312
rect 3476 458272 391940 458300
rect 3476 458260 3482 458272
rect 391934 458260 391940 458272
rect 391992 458260 391998 458312
rect 4890 458192 4896 458244
rect 4948 458232 4954 458244
rect 396856 458232 396862 458244
rect 4948 458204 396862 458232
rect 4948 458192 4954 458204
rect 396856 458192 396862 458204
rect 396914 458192 396920 458244
rect 258046 457592 287054 457620
rect 4062 457444 4068 457496
rect 4120 457484 4126 457496
rect 258046 457484 258074 457592
rect 4120 457456 258074 457484
rect 260806 457524 270494 457552
rect 4120 457444 4126 457456
rect 260806 457212 260834 457524
rect 261294 457444 261300 457496
rect 261352 457444 261358 457496
rect 266078 457444 266084 457496
rect 266136 457444 266142 457496
rect 258046 457184 260834 457212
rect 234154 457104 234160 457156
rect 234212 457144 234218 457156
rect 258046 457144 258074 457184
rect 234212 457116 258074 457144
rect 234212 457104 234218 457116
rect 261312 456804 261340 457444
rect 266096 456872 266124 457444
rect 270466 457212 270494 457524
rect 273226 457524 282914 457552
rect 273226 457212 273254 457524
rect 273990 457444 273996 457496
rect 274048 457444 274054 457496
rect 275554 457444 275560 457496
rect 275612 457444 275618 457496
rect 278590 457444 278596 457496
rect 278648 457444 278654 457496
rect 270466 457184 273254 457212
rect 274008 456940 274036 457444
rect 275572 457008 275600 457444
rect 278608 457076 278636 457444
rect 282886 457212 282914 457524
rect 287026 457484 287054 457592
rect 360654 457484 360660 457496
rect 287026 457456 360660 457484
rect 360654 457444 360660 457456
rect 360712 457444 360718 457496
rect 388622 457484 388628 457496
rect 373966 457456 388628 457484
rect 282886 457184 287054 457212
rect 287026 457144 287054 457184
rect 373966 457144 373994 457456
rect 388622 457444 388628 457456
rect 388680 457444 388686 457496
rect 287026 457116 373994 457144
rect 580166 457076 580172 457088
rect 278608 457048 580172 457076
rect 580166 457036 580172 457048
rect 580224 457036 580230 457088
rect 580902 457008 580908 457020
rect 275572 456980 580908 457008
rect 580902 456968 580908 456980
rect 580960 456968 580966 457020
rect 580718 456940 580724 456952
rect 274008 456912 580724 456940
rect 580718 456900 580724 456912
rect 580776 456900 580782 456952
rect 578142 456872 578148 456884
rect 266096 456844 578148 456872
rect 578142 456832 578148 456844
rect 578200 456832 578206 456884
rect 577958 456804 577964 456816
rect 261312 456776 577964 456804
rect 577958 456764 577964 456776
rect 578016 456764 578022 456816
rect 2774 449828 2780 449880
rect 2832 449868 2838 449880
rect 4982 449868 4988 449880
rect 2832 449840 4988 449868
rect 2832 449828 2838 449840
rect 4982 449828 4988 449840
rect 5040 449828 5046 449880
rect 415026 419432 415032 419484
rect 415084 419472 415090 419484
rect 579982 419472 579988 419484
rect 415084 419444 579988 419472
rect 415084 419432 415090 419444
rect 579982 419432 579988 419444
rect 580040 419432 580046 419484
rect 341012 337764 341018 337816
rect 341070 337804 341076 337816
rect 341242 337804 341248 337816
rect 341070 337776 341248 337804
rect 341070 337764 341076 337776
rect 341242 337764 341248 337776
rect 341300 337764 341306 337816
rect 252554 336744 252560 336796
rect 252612 336784 252618 336796
rect 252830 336784 252836 336796
rect 252612 336756 252836 336784
rect 252612 336744 252618 336756
rect 252830 336744 252836 336756
rect 252888 336744 252894 336796
rect 265158 336744 265164 336796
rect 265216 336784 265222 336796
rect 265342 336784 265348 336796
rect 265216 336756 265348 336784
rect 265216 336744 265222 336756
rect 265342 336744 265348 336756
rect 265400 336744 265406 336796
rect 306558 336744 306564 336796
rect 306616 336784 306622 336796
rect 307202 336784 307208 336796
rect 306616 336756 307208 336784
rect 306616 336744 306622 336756
rect 307202 336744 307208 336756
rect 307260 336744 307266 336796
rect 309226 336744 309232 336796
rect 309284 336784 309290 336796
rect 309502 336784 309508 336796
rect 309284 336756 309508 336784
rect 309284 336744 309290 336756
rect 309502 336744 309508 336756
rect 309560 336744 309566 336796
rect 361758 336744 361764 336796
rect 361816 336784 361822 336796
rect 362310 336784 362316 336796
rect 361816 336756 362316 336784
rect 361816 336744 361822 336756
rect 362310 336744 362316 336756
rect 362368 336744 362374 336796
rect 390646 336744 390652 336796
rect 390704 336784 390710 336796
rect 391198 336784 391204 336796
rect 390704 336756 391204 336784
rect 390704 336744 390710 336756
rect 391198 336744 391204 336756
rect 391256 336744 391262 336796
rect 177298 336676 177304 336728
rect 177356 336716 177362 336728
rect 268838 336716 268844 336728
rect 177356 336688 268844 336716
rect 177356 336676 177362 336688
rect 268838 336676 268844 336688
rect 268896 336676 268902 336728
rect 305638 336676 305644 336728
rect 305696 336716 305702 336728
rect 325418 336716 325424 336728
rect 305696 336688 325424 336716
rect 305696 336676 305702 336688
rect 325418 336676 325424 336688
rect 325476 336676 325482 336728
rect 340782 336676 340788 336728
rect 340840 336716 340846 336728
rect 341334 336716 341340 336728
rect 340840 336688 341340 336716
rect 340840 336676 340846 336688
rect 341334 336676 341340 336688
rect 341392 336676 341398 336728
rect 361574 336676 361580 336728
rect 361632 336716 361638 336728
rect 361942 336716 361948 336728
rect 361632 336688 361948 336716
rect 361632 336676 361638 336688
rect 361942 336676 361948 336688
rect 362000 336676 362006 336728
rect 365622 336676 365628 336728
rect 365680 336716 365686 336728
rect 388530 336716 388536 336728
rect 365680 336688 388536 336716
rect 365680 336676 365686 336688
rect 388530 336676 388536 336688
rect 388588 336676 388594 336728
rect 390554 336676 390560 336728
rect 390612 336716 390618 336728
rect 390830 336716 390836 336728
rect 390612 336688 390836 336716
rect 390612 336676 390618 336688
rect 390830 336676 390836 336688
rect 390888 336676 390894 336728
rect 396074 336676 396080 336728
rect 396132 336716 396138 336728
rect 396350 336716 396356 336728
rect 396132 336688 396356 336716
rect 396132 336676 396138 336688
rect 396350 336676 396356 336688
rect 396408 336676 396414 336728
rect 401594 336676 401600 336728
rect 401652 336716 401658 336728
rect 401870 336716 401876 336728
rect 401652 336688 401876 336716
rect 401652 336676 401658 336688
rect 401870 336676 401876 336688
rect 401928 336676 401934 336728
rect 414014 336676 414020 336728
rect 414072 336716 414078 336728
rect 450538 336716 450544 336728
rect 414072 336688 450544 336716
rect 414072 336676 414078 336688
rect 450538 336676 450544 336688
rect 450596 336676 450602 336728
rect 173158 336608 173164 336660
rect 173216 336648 173222 336660
rect 266630 336648 266636 336660
rect 173216 336620 266636 336648
rect 173216 336608 173222 336620
rect 266630 336608 266636 336620
rect 266688 336608 266694 336660
rect 290274 336608 290280 336660
rect 290332 336648 290338 336660
rect 324314 336648 324320 336660
rect 290332 336620 324320 336648
rect 290332 336608 290338 336620
rect 324314 336608 324320 336620
rect 324372 336608 324378 336660
rect 346394 336608 346400 336660
rect 346452 336648 346458 336660
rect 358078 336648 358084 336660
rect 346452 336620 358084 336648
rect 346452 336608 346458 336620
rect 358078 336608 358084 336620
rect 358136 336608 358142 336660
rect 360102 336608 360108 336660
rect 360160 336648 360166 336660
rect 373074 336648 373080 336660
rect 360160 336620 373080 336648
rect 360160 336608 360166 336620
rect 373074 336608 373080 336620
rect 373132 336608 373138 336660
rect 376754 336608 376760 336660
rect 376812 336648 376818 336660
rect 377030 336648 377036 336660
rect 376812 336620 377036 336648
rect 376812 336608 376818 336620
rect 377030 336608 377036 336620
rect 377088 336608 377094 336660
rect 378962 336608 378968 336660
rect 379020 336648 379026 336660
rect 428458 336648 428464 336660
rect 379020 336620 428464 336648
rect 379020 336608 379026 336620
rect 428458 336608 428464 336620
rect 428516 336608 428522 336660
rect 163498 336540 163504 336592
rect 163556 336580 163562 336592
rect 264422 336580 264428 336592
rect 163556 336552 264428 336580
rect 163556 336540 163562 336552
rect 264422 336540 264428 336552
rect 264480 336540 264486 336592
rect 284294 336540 284300 336592
rect 284352 336580 284358 336592
rect 322474 336580 322480 336592
rect 284352 336552 322480 336580
rect 284352 336540 284358 336552
rect 322474 336540 322480 336552
rect 322532 336540 322538 336592
rect 355870 336540 355876 336592
rect 355928 336580 355934 336592
rect 366450 336580 366456 336592
rect 355928 336552 366456 336580
rect 355928 336540 355934 336552
rect 366450 336540 366456 336552
rect 366508 336540 366514 336592
rect 367554 336540 367560 336592
rect 367612 336580 367618 336592
rect 422938 336580 422944 336592
rect 367612 336552 422944 336580
rect 367612 336540 367618 336552
rect 422938 336540 422944 336552
rect 422996 336540 423002 336592
rect 153838 336472 153844 336524
rect 153896 336512 153902 336524
rect 262214 336512 262220 336524
rect 153896 336484 262220 336512
rect 153896 336472 153902 336484
rect 262214 336472 262220 336484
rect 262272 336472 262278 336524
rect 268378 336472 268384 336524
rect 268436 336512 268442 336524
rect 314102 336512 314108 336524
rect 268436 336484 314108 336512
rect 268436 336472 268442 336484
rect 314102 336472 314108 336484
rect 314160 336472 314166 336524
rect 315022 336472 315028 336524
rect 315080 336512 315086 336524
rect 331950 336512 331956 336524
rect 315080 336484 331956 336512
rect 315080 336472 315086 336484
rect 331950 336472 331956 336484
rect 332008 336472 332014 336524
rect 353754 336472 353760 336524
rect 353812 336512 353818 336524
rect 362126 336512 362132 336524
rect 353812 336484 362132 336512
rect 353812 336472 353818 336484
rect 362126 336472 362132 336484
rect 362184 336472 362190 336524
rect 371142 336472 371148 336524
rect 371200 336512 371206 336524
rect 425790 336512 425796 336524
rect 371200 336484 425796 336512
rect 371200 336472 371206 336484
rect 425790 336472 425796 336484
rect 425848 336472 425854 336524
rect 149698 336404 149704 336456
rect 149756 336444 149762 336456
rect 261110 336444 261116 336456
rect 149756 336416 261116 336444
rect 149756 336404 149762 336416
rect 261110 336404 261116 336416
rect 261168 336404 261174 336456
rect 273622 336404 273628 336456
rect 273680 336444 273686 336456
rect 319254 336444 319260 336456
rect 273680 336416 319260 336444
rect 273680 336404 273686 336416
rect 319254 336404 319260 336416
rect 319312 336404 319318 336456
rect 331214 336404 331220 336456
rect 331272 336444 331278 336456
rect 337102 336444 337108 336456
rect 331272 336416 337108 336444
rect 331272 336404 331278 336416
rect 337102 336404 337108 336416
rect 337160 336404 337166 336456
rect 355778 336404 355784 336456
rect 355836 336444 355842 336456
rect 367646 336444 367652 336456
rect 355836 336416 367652 336444
rect 355836 336404 355842 336416
rect 367646 336404 367652 336416
rect 367704 336404 367710 336456
rect 368658 336404 368664 336456
rect 368716 336444 368722 336456
rect 425698 336444 425704 336456
rect 368716 336416 425704 336444
rect 368716 336404 368722 336416
rect 425698 336404 425704 336416
rect 425756 336404 425762 336456
rect 145558 336336 145564 336388
rect 145616 336376 145622 336388
rect 258994 336376 259000 336388
rect 145616 336348 259000 336376
rect 145616 336336 145622 336348
rect 258994 336336 259000 336348
rect 259052 336336 259058 336388
rect 265618 336336 265624 336388
rect 265676 336376 265682 336388
rect 265676 336348 309824 336376
rect 265676 336336 265682 336348
rect 45554 336268 45560 336320
rect 45612 336308 45618 336320
rect 249058 336308 249064 336320
rect 45612 336280 249064 336308
rect 45612 336268 45618 336280
rect 249058 336268 249064 336280
rect 249116 336268 249122 336320
rect 268562 336268 268568 336320
rect 268620 336308 268626 336320
rect 309594 336308 309600 336320
rect 268620 336280 309600 336308
rect 268620 336268 268626 336280
rect 309594 336268 309600 336280
rect 309652 336268 309658 336320
rect 309796 336308 309824 336348
rect 312538 336336 312544 336388
rect 312596 336376 312602 336388
rect 324682 336376 324688 336388
rect 312596 336348 324688 336376
rect 312596 336336 312602 336348
rect 324682 336336 324688 336348
rect 324740 336336 324746 336388
rect 347682 336336 347688 336388
rect 347740 336376 347746 336388
rect 362310 336376 362316 336388
rect 347740 336348 362316 336376
rect 347740 336336 347746 336348
rect 362310 336336 362316 336348
rect 362368 336336 362374 336388
rect 374178 336336 374184 336388
rect 374236 336376 374242 336388
rect 378962 336376 378968 336388
rect 374236 336348 378968 336376
rect 374236 336336 374242 336348
rect 378962 336336 378968 336348
rect 379020 336336 379026 336388
rect 379606 336336 379612 336388
rect 379664 336376 379670 336388
rect 442258 336376 442264 336388
rect 379664 336348 442264 336376
rect 379664 336336 379670 336348
rect 442258 336336 442264 336348
rect 442316 336336 442322 336388
rect 312998 336308 313004 336320
rect 309796 336280 313004 336308
rect 312998 336268 313004 336280
rect 313056 336268 313062 336320
rect 316402 336268 316408 336320
rect 316460 336308 316466 336320
rect 332686 336308 332692 336320
rect 316460 336280 332692 336308
rect 316460 336268 316466 336280
rect 332686 336268 332692 336280
rect 332744 336268 332750 336320
rect 348602 336268 348608 336320
rect 348660 336308 348666 336320
rect 364978 336308 364984 336320
rect 348660 336280 364984 336308
rect 348660 336268 348666 336280
rect 364978 336268 364984 336280
rect 365036 336268 365042 336320
rect 373166 336268 373172 336320
rect 373224 336308 373230 336320
rect 436738 336308 436744 336320
rect 373224 336280 436744 336308
rect 373224 336268 373230 336280
rect 436738 336268 436744 336280
rect 436796 336268 436802 336320
rect 31754 336200 31760 336252
rect 31812 336240 31818 336252
rect 244734 336240 244740 336252
rect 31812 336212 244740 336240
rect 31812 336200 31818 336212
rect 244734 336200 244740 336212
rect 244792 336200 244798 336252
rect 264238 336200 264244 336252
rect 264296 336240 264302 336252
rect 311894 336240 311900 336252
rect 264296 336212 311900 336240
rect 264296 336200 264302 336212
rect 311894 336200 311900 336212
rect 311952 336200 311958 336252
rect 312722 336200 312728 336252
rect 312780 336240 312786 336252
rect 330570 336240 330576 336252
rect 312780 336212 330576 336240
rect 312780 336200 312786 336212
rect 330570 336200 330576 336212
rect 330628 336200 330634 336252
rect 345290 336200 345296 336252
rect 345348 336240 345354 336252
rect 355410 336240 355416 336252
rect 345348 336212 355416 336240
rect 345348 336200 345354 336212
rect 355410 336200 355416 336212
rect 355468 336200 355474 336252
rect 356882 336200 356888 336252
rect 356940 336240 356946 336252
rect 373350 336240 373356 336252
rect 356940 336212 373356 336240
rect 356940 336200 356946 336212
rect 373350 336200 373356 336212
rect 373408 336200 373414 336252
rect 376662 336200 376668 336252
rect 376720 336240 376726 336252
rect 439498 336240 439504 336252
rect 376720 336212 439504 336240
rect 376720 336200 376726 336212
rect 439498 336200 439504 336212
rect 439556 336200 439562 336252
rect 24854 336132 24860 336184
rect 24912 336172 24918 336184
rect 242526 336172 242532 336184
rect 24912 336144 242532 336172
rect 24912 336132 24918 336144
rect 242526 336132 242532 336144
rect 242584 336132 242590 336184
rect 262858 336132 262864 336184
rect 262916 336172 262922 336184
rect 310790 336172 310796 336184
rect 262916 336144 310796 336172
rect 262916 336132 262922 336144
rect 310790 336132 310796 336144
rect 310848 336132 310854 336184
rect 313274 336132 313280 336184
rect 313332 336172 313338 336184
rect 331582 336172 331588 336184
rect 313332 336144 331588 336172
rect 313332 336132 313338 336144
rect 331582 336132 331588 336144
rect 331640 336132 331646 336184
rect 350350 336132 350356 336184
rect 350408 336172 350414 336184
rect 367830 336172 367836 336184
rect 350408 336144 367836 336172
rect 350408 336132 350414 336144
rect 367830 336132 367836 336144
rect 367888 336132 367894 336184
rect 381814 336132 381820 336184
rect 381872 336172 381878 336184
rect 447778 336172 447784 336184
rect 381872 336144 447784 336172
rect 381872 336132 381878 336144
rect 447778 336132 447784 336144
rect 447836 336132 447842 336184
rect 15194 336064 15200 336116
rect 15252 336104 15258 336116
rect 239582 336104 239588 336116
rect 15252 336076 239588 336104
rect 15252 336064 15258 336076
rect 239582 336064 239588 336076
rect 239640 336064 239646 336116
rect 265526 336104 265532 336116
rect 248386 336076 265532 336104
rect 5534 335996 5540 336048
rect 5592 336036 5598 336048
rect 236638 336036 236644 336048
rect 5592 336008 236644 336036
rect 5592 335996 5598 336008
rect 236638 335996 236644 336008
rect 236696 335996 236702 336048
rect 239398 335996 239404 336048
rect 239456 336036 239462 336048
rect 248386 336036 248414 336076
rect 265526 336064 265532 336076
rect 265584 336064 265590 336116
rect 269390 336064 269396 336116
rect 269448 336104 269454 336116
rect 318150 336104 318156 336116
rect 269448 336076 318156 336104
rect 269448 336064 269454 336076
rect 318150 336064 318156 336076
rect 318208 336064 318214 336116
rect 352558 336064 352564 336116
rect 352616 336104 352622 336116
rect 371878 336104 371884 336116
rect 352616 336076 371884 336104
rect 352616 336064 352622 336076
rect 371878 336064 371884 336076
rect 371936 336064 371942 336116
rect 377490 336064 377496 336116
rect 377548 336104 377554 336116
rect 443638 336104 443644 336116
rect 377548 336076 443644 336104
rect 377548 336064 377554 336076
rect 443638 336064 443644 336076
rect 443696 336064 443702 336116
rect 239456 336008 248414 336036
rect 239456 335996 239462 336008
rect 262214 335996 262220 336048
rect 262272 336036 262278 336048
rect 316034 336036 316040 336048
rect 262272 336008 316040 336036
rect 262272 335996 262278 336008
rect 316034 335996 316040 336008
rect 316092 335996 316098 336048
rect 319438 335996 319444 336048
rect 319496 336036 319502 336048
rect 330202 336036 330208 336048
rect 319496 336008 330208 336036
rect 319496 335996 319502 336008
rect 330202 335996 330208 336008
rect 330260 335996 330266 336048
rect 349982 335996 349988 336048
rect 350040 336036 350046 336048
rect 370498 336036 370504 336048
rect 350040 336008 370504 336036
rect 350040 335996 350046 336008
rect 370498 335996 370504 336008
rect 370556 335996 370562 336048
rect 375282 335996 375288 336048
rect 375340 336036 375346 336048
rect 440878 336036 440884 336048
rect 375340 336008 440884 336036
rect 375340 335996 375346 336008
rect 440878 335996 440884 336008
rect 440936 335996 440942 336048
rect 185578 335928 185584 335980
rect 185636 335968 185642 335980
rect 271046 335968 271052 335980
rect 185636 335940 271052 335968
rect 185636 335928 185642 335940
rect 271046 335928 271052 335940
rect 271104 335928 271110 335980
rect 307018 335928 307024 335980
rect 307076 335968 307082 335980
rect 326522 335968 326528 335980
rect 307076 335940 326528 335968
rect 307076 335928 307082 335940
rect 326522 335928 326528 335940
rect 326580 335928 326586 335980
rect 363230 335928 363236 335980
rect 363288 335968 363294 335980
rect 388438 335968 388444 335980
rect 363288 335940 388444 335968
rect 363288 335928 363294 335940
rect 388438 335928 388444 335940
rect 388496 335928 388502 335980
rect 388530 335928 388536 335980
rect 388588 335968 388594 335980
rect 391198 335968 391204 335980
rect 388588 335940 391204 335968
rect 388588 335928 388594 335940
rect 391198 335928 391204 335940
rect 391256 335928 391262 335980
rect 412542 335928 412548 335980
rect 412600 335968 412606 335980
rect 431218 335968 431224 335980
rect 412600 335940 431224 335968
rect 412600 335928 412606 335940
rect 431218 335928 431224 335940
rect 431276 335928 431282 335980
rect 188338 335860 188344 335912
rect 188396 335900 188402 335912
rect 272150 335900 272156 335912
rect 188396 335872 272156 335900
rect 188396 335860 188402 335872
rect 272150 335860 272156 335872
rect 272208 335860 272214 335912
rect 311250 335860 311256 335912
rect 311308 335900 311314 335912
rect 329466 335900 329472 335912
rect 311308 335872 329472 335900
rect 311308 335860 311314 335872
rect 329466 335860 329472 335872
rect 329524 335860 329530 335912
rect 358814 335860 358820 335912
rect 358872 335900 358878 335912
rect 374638 335900 374644 335912
rect 358872 335872 374644 335900
rect 358872 335860 358878 335872
rect 374638 335860 374644 335872
rect 374696 335860 374702 335912
rect 408402 335860 408408 335912
rect 408460 335900 408466 335912
rect 418890 335900 418896 335912
rect 408460 335872 418896 335900
rect 408460 335860 408466 335872
rect 418890 335860 418896 335872
rect 418948 335860 418954 335912
rect 261570 335792 261576 335844
rect 261628 335832 261634 335844
rect 261628 335804 296714 335832
rect 261628 335792 261634 335804
rect 258810 335724 258816 335776
rect 258868 335764 258874 335776
rect 290182 335764 290188 335776
rect 258868 335736 290188 335764
rect 258868 335724 258874 335736
rect 290182 335724 290188 335736
rect 290240 335724 290246 335776
rect 258718 335656 258724 335708
rect 258776 335696 258782 335708
rect 288894 335696 288900 335708
rect 258776 335668 288900 335696
rect 258776 335656 258782 335668
rect 288894 335656 288900 335668
rect 288952 335656 288958 335708
rect 296686 335696 296714 335804
rect 309594 335792 309600 335844
rect 309652 335832 309658 335844
rect 314838 335832 314844 335844
rect 309652 335804 314844 335832
rect 309652 335792 309658 335804
rect 314838 335792 314844 335804
rect 314896 335792 314902 335844
rect 317414 335792 317420 335844
rect 317472 335832 317478 335844
rect 333054 335832 333060 335844
rect 317472 335804 333060 335832
rect 317472 335792 317478 335804
rect 333054 335792 333060 335804
rect 333112 335792 333118 335844
rect 357158 335792 357164 335844
rect 357216 335832 357222 335844
rect 369118 335832 369124 335844
rect 357216 335804 369124 335832
rect 357216 335792 357222 335804
rect 369118 335792 369124 335804
rect 369176 335792 369182 335844
rect 410334 335792 410340 335844
rect 410392 335832 410398 335844
rect 418798 335832 418804 335844
rect 410392 335804 418804 335832
rect 410392 335792 410398 335804
rect 418798 335792 418804 335804
rect 418856 335792 418862 335844
rect 307110 335724 307116 335776
rect 307168 335764 307174 335776
rect 322106 335764 322112 335776
rect 307168 335736 322112 335764
rect 307168 335724 307174 335736
rect 322106 335724 322112 335736
rect 322164 335724 322170 335776
rect 350810 335724 350816 335776
rect 350868 335764 350874 335776
rect 363598 335764 363604 335776
rect 350868 335736 363604 335764
rect 350868 335724 350874 335736
rect 363598 335724 363604 335736
rect 363656 335724 363662 335776
rect 366266 335764 366272 335776
rect 364306 335736 366272 335764
rect 307478 335696 307484 335708
rect 296686 335668 307484 335696
rect 307478 335656 307484 335668
rect 307536 335656 307542 335708
rect 315298 335656 315304 335708
rect 315356 335696 315362 335708
rect 327074 335696 327080 335708
rect 315356 335668 327080 335696
rect 315356 335656 315362 335668
rect 327074 335656 327080 335668
rect 327132 335656 327138 335708
rect 244918 335588 244924 335640
rect 244976 335628 244982 335640
rect 273254 335628 273260 335640
rect 244976 335600 273260 335628
rect 244976 335588 244982 335600
rect 273254 335588 273260 335600
rect 273312 335588 273318 335640
rect 307202 335588 307208 335640
rect 307260 335628 307266 335640
rect 315206 335628 315212 335640
rect 307260 335600 315212 335628
rect 307260 335588 307266 335600
rect 315206 335588 315212 335600
rect 315264 335588 315270 335640
rect 354858 335588 354864 335640
rect 354916 335628 354922 335640
rect 364306 335628 364334 335736
rect 366266 335724 366272 335736
rect 366324 335724 366330 335776
rect 354916 335600 364334 335628
rect 354916 335588 354922 335600
rect 242158 335520 242164 335572
rect 242216 335560 242222 335572
rect 269942 335560 269948 335572
rect 242216 335532 269948 335560
rect 242216 335520 242222 335532
rect 269942 335520 269948 335532
rect 270000 335520 270006 335572
rect 236638 335452 236644 335504
rect 236696 335492 236702 335504
rect 263318 335492 263324 335504
rect 236696 335464 263324 335492
rect 236696 335452 236702 335464
rect 263318 335452 263324 335464
rect 263376 335452 263382 335504
rect 352650 335452 352656 335504
rect 352708 335492 352714 335504
rect 358170 335492 358176 335504
rect 352708 335464 358176 335492
rect 352708 335452 352714 335464
rect 358170 335452 358176 335464
rect 358228 335452 358234 335504
rect 242250 335384 242256 335436
rect 242308 335424 242314 335436
rect 267826 335424 267832 335436
rect 242308 335396 267832 335424
rect 242308 335384 242314 335396
rect 267826 335384 267832 335396
rect 267884 335384 267890 335436
rect 351822 335384 351828 335436
rect 351880 335424 351886 335436
rect 356698 335424 356704 335436
rect 351880 335396 356704 335424
rect 351880 335384 351886 335396
rect 356698 335384 356704 335396
rect 356756 335384 356762 335436
rect 330202 335316 330208 335368
rect 330260 335356 330266 335368
rect 336734 335356 336740 335368
rect 330260 335328 336740 335356
rect 330260 335316 330266 335328
rect 336734 335316 336740 335328
rect 336792 335316 336798 335368
rect 350442 335316 350448 335368
rect 350500 335356 350506 335368
rect 355318 335356 355324 335368
rect 350500 335328 355324 335356
rect 350500 335316 350506 335328
rect 355318 335316 355324 335328
rect 355376 335316 355382 335368
rect 371970 335316 371976 335368
rect 372028 335356 372034 335368
rect 376018 335356 376024 335368
rect 372028 335328 376024 335356
rect 372028 335316 372034 335328
rect 376018 335316 376024 335328
rect 376076 335316 376082 335368
rect 278958 330760 278964 330812
rect 279016 330760 279022 330812
rect 280246 330760 280252 330812
rect 280304 330760 280310 330812
rect 339678 330760 339684 330812
rect 339736 330760 339742 330812
rect 342438 330760 342444 330812
rect 342496 330760 342502 330812
rect 386598 330760 386604 330812
rect 386656 330760 386662 330812
rect 404446 330760 404452 330812
rect 404504 330760 404510 330812
rect 234614 330624 234620 330676
rect 234672 330664 234678 330676
rect 234798 330664 234804 330676
rect 234672 330636 234804 330664
rect 234672 330624 234678 330636
rect 234798 330624 234804 330636
rect 234856 330624 234862 330676
rect 278976 330608 279004 330760
rect 280264 330608 280292 330760
rect 339696 330608 339724 330760
rect 342456 330608 342484 330760
rect 386616 330608 386644 330760
rect 404464 330608 404492 330760
rect 278958 330556 278964 330608
rect 279016 330556 279022 330608
rect 280246 330556 280252 330608
rect 280304 330556 280310 330608
rect 285674 330556 285680 330608
rect 285732 330596 285738 330608
rect 286042 330596 286048 330608
rect 285732 330568 286048 330596
rect 285732 330556 285738 330568
rect 286042 330556 286048 330568
rect 286100 330556 286106 330608
rect 302234 330556 302240 330608
rect 302292 330596 302298 330608
rect 302602 330596 302608 330608
rect 302292 330568 302608 330596
rect 302292 330556 302298 330568
rect 302602 330556 302608 330568
rect 302660 330556 302666 330608
rect 304994 330556 305000 330608
rect 305052 330596 305058 330608
rect 305362 330596 305368 330608
rect 305052 330568 305368 330596
rect 305052 330556 305058 330568
rect 305362 330556 305368 330568
rect 305420 330556 305426 330608
rect 339678 330556 339684 330608
rect 339736 330556 339742 330608
rect 342438 330556 342444 330608
rect 342496 330556 342502 330608
rect 386598 330556 386604 330608
rect 386656 330556 386662 330608
rect 404446 330556 404452 330608
rect 404504 330556 404510 330608
rect 405734 330556 405740 330608
rect 405792 330596 405798 330608
rect 406838 330596 406844 330608
rect 405792 330568 406844 330596
rect 405792 330556 405798 330568
rect 406838 330556 406844 330568
rect 406896 330556 406902 330608
rect 236086 330488 236092 330540
rect 236144 330528 236150 330540
rect 237006 330528 237012 330540
rect 236144 330500 237012 330528
rect 236144 330488 236150 330500
rect 237006 330488 237012 330500
rect 237064 330488 237070 330540
rect 237466 330488 237472 330540
rect 237524 330528 237530 330540
rect 238478 330528 238484 330540
rect 237524 330500 238484 330528
rect 237524 330488 237530 330500
rect 238478 330488 238484 330500
rect 238536 330488 238542 330540
rect 240134 330488 240140 330540
rect 240192 330528 240198 330540
rect 240686 330528 240692 330540
rect 240192 330500 240692 330528
rect 240192 330488 240198 330500
rect 240686 330488 240692 330500
rect 240744 330488 240750 330540
rect 254026 330488 254032 330540
rect 254084 330528 254090 330540
rect 254946 330528 254952 330540
rect 254084 330500 254952 330528
rect 254084 330488 254090 330500
rect 254946 330488 254952 330500
rect 255004 330488 255010 330540
rect 255498 330488 255504 330540
rect 255556 330528 255562 330540
rect 256418 330528 256424 330540
rect 255556 330500 256424 330528
rect 255556 330488 255562 330500
rect 256418 330488 256424 330500
rect 256476 330488 256482 330540
rect 256694 330488 256700 330540
rect 256752 330528 256758 330540
rect 257154 330528 257160 330540
rect 256752 330500 257160 330528
rect 256752 330488 256758 330500
rect 257154 330488 257160 330500
rect 257212 330488 257218 330540
rect 258166 330488 258172 330540
rect 258224 330528 258230 330540
rect 258626 330528 258632 330540
rect 258224 330500 258632 330528
rect 258224 330488 258230 330500
rect 258626 330488 258632 330500
rect 258684 330488 258690 330540
rect 259638 330488 259644 330540
rect 259696 330528 259702 330540
rect 260374 330528 260380 330540
rect 259696 330500 260380 330528
rect 259696 330488 259702 330500
rect 260374 330488 260380 330500
rect 260432 330488 260438 330540
rect 261018 330488 261024 330540
rect 261076 330528 261082 330540
rect 261846 330528 261852 330540
rect 261076 330500 261852 330528
rect 261076 330488 261082 330500
rect 261846 330488 261852 330500
rect 261904 330488 261910 330540
rect 262398 330488 262404 330540
rect 262456 330528 262462 330540
rect 262950 330528 262956 330540
rect 262456 330500 262956 330528
rect 262456 330488 262462 330500
rect 262950 330488 262956 330500
rect 263008 330488 263014 330540
rect 266538 330488 266544 330540
rect 266596 330528 266602 330540
rect 267366 330528 267372 330540
rect 266596 330500 267372 330528
rect 266596 330488 266602 330500
rect 267366 330488 267372 330500
rect 267424 330488 267430 330540
rect 271966 330488 271972 330540
rect 272024 330528 272030 330540
rect 272794 330528 272800 330540
rect 272024 330500 272800 330528
rect 272024 330488 272030 330500
rect 272794 330488 272800 330500
rect 272852 330488 272858 330540
rect 273346 330488 273352 330540
rect 273404 330528 273410 330540
rect 273898 330528 273904 330540
rect 273404 330500 273904 330528
rect 273404 330488 273410 330500
rect 273898 330488 273904 330500
rect 273956 330488 273962 330540
rect 274634 330488 274640 330540
rect 274692 330528 274698 330540
rect 275738 330528 275744 330540
rect 274692 330500 275744 330528
rect 274692 330488 274698 330500
rect 275738 330488 275744 330500
rect 275796 330488 275802 330540
rect 276106 330488 276112 330540
rect 276164 330528 276170 330540
rect 276842 330528 276848 330540
rect 276164 330500 276848 330528
rect 276164 330488 276170 330500
rect 276842 330488 276848 330500
rect 276900 330488 276906 330540
rect 277578 330488 277584 330540
rect 277636 330528 277642 330540
rect 278314 330528 278320 330540
rect 277636 330500 278320 330528
rect 277636 330488 277642 330500
rect 278314 330488 278320 330500
rect 278372 330488 278378 330540
rect 278866 330488 278872 330540
rect 278924 330528 278930 330540
rect 279418 330528 279424 330540
rect 278924 330500 279424 330528
rect 278924 330488 278930 330500
rect 279418 330488 279424 330500
rect 279476 330488 279482 330540
rect 280338 330488 280344 330540
rect 280396 330528 280402 330540
rect 281258 330528 281264 330540
rect 280396 330500 281264 330528
rect 280396 330488 280402 330500
rect 281258 330488 281264 330500
rect 281316 330488 281322 330540
rect 283098 330488 283104 330540
rect 283156 330528 283162 330540
rect 283742 330528 283748 330540
rect 283156 330500 283748 330528
rect 283156 330488 283162 330500
rect 283742 330488 283748 330500
rect 283800 330488 283806 330540
rect 284386 330488 284392 330540
rect 284444 330528 284450 330540
rect 284846 330528 284852 330540
rect 284444 330500 284852 330528
rect 284444 330488 284450 330500
rect 284846 330488 284852 330500
rect 284904 330488 284910 330540
rect 285766 330488 285772 330540
rect 285824 330528 285830 330540
rect 286318 330528 286324 330540
rect 285824 330500 286324 330528
rect 285824 330488 285830 330500
rect 286318 330488 286324 330500
rect 286376 330488 286382 330540
rect 287054 330488 287060 330540
rect 287112 330528 287118 330540
rect 288158 330528 288164 330540
rect 287112 330500 288164 330528
rect 287112 330488 287118 330500
rect 288158 330488 288164 330500
rect 288216 330488 288222 330540
rect 289906 330488 289912 330540
rect 289964 330528 289970 330540
rect 290366 330528 290372 330540
rect 289964 330500 290372 330528
rect 289964 330488 289970 330500
rect 290366 330488 290372 330500
rect 290424 330488 290430 330540
rect 291286 330488 291292 330540
rect 291344 330528 291350 330540
rect 292206 330528 292212 330540
rect 291344 330500 292212 330528
rect 291344 330488 291350 330500
rect 292206 330488 292212 330500
rect 292264 330488 292270 330540
rect 302326 330488 302332 330540
rect 302384 330528 302390 330540
rect 302786 330528 302792 330540
rect 302384 330500 302792 330528
rect 302384 330488 302390 330500
rect 302786 330488 302792 330500
rect 302844 330488 302850 330540
rect 303706 330488 303712 330540
rect 303764 330528 303770 330540
rect 304626 330528 304632 330540
rect 303764 330500 304632 330528
rect 303764 330488 303770 330500
rect 304626 330488 304632 330500
rect 304684 330488 304690 330540
rect 305086 330488 305092 330540
rect 305144 330528 305150 330540
rect 305730 330528 305736 330540
rect 305144 330500 305736 330528
rect 305144 330488 305150 330500
rect 305730 330488 305736 330500
rect 305788 330488 305794 330540
rect 306466 330488 306472 330540
rect 306524 330528 306530 330540
rect 306834 330528 306840 330540
rect 306524 330500 306840 330528
rect 306524 330488 306530 330500
rect 306834 330488 306840 330500
rect 306892 330488 306898 330540
rect 307846 330488 307852 330540
rect 307904 330528 307910 330540
rect 308582 330528 308588 330540
rect 307904 330500 308588 330528
rect 307904 330488 307910 330500
rect 308582 330488 308588 330500
rect 308640 330488 308646 330540
rect 309318 330488 309324 330540
rect 309376 330528 309382 330540
rect 310054 330528 310060 330540
rect 309376 330500 310060 330528
rect 309376 330488 309382 330500
rect 310054 330488 310060 330500
rect 310112 330488 310118 330540
rect 314838 330488 314844 330540
rect 314896 330528 314902 330540
rect 315574 330528 315580 330540
rect 314896 330500 315580 330528
rect 314896 330488 314902 330500
rect 315574 330488 315580 330500
rect 315632 330488 315638 330540
rect 318886 330488 318892 330540
rect 318944 330528 318950 330540
rect 319898 330528 319904 330540
rect 318944 330500 319904 330528
rect 318944 330488 318950 330500
rect 319898 330488 319904 330500
rect 319956 330488 319962 330540
rect 333974 330488 333980 330540
rect 334032 330528 334038 330540
rect 334526 330528 334532 330540
rect 334032 330500 334532 330528
rect 334032 330488 334038 330500
rect 334526 330488 334532 330500
rect 334584 330488 334590 330540
rect 336826 330488 336832 330540
rect 336884 330528 336890 330540
rect 337838 330528 337844 330540
rect 336884 330500 337844 330528
rect 336884 330488 336890 330500
rect 337838 330488 337844 330500
rect 337896 330488 337902 330540
rect 339586 330488 339592 330540
rect 339644 330528 339650 330540
rect 340046 330528 340052 330540
rect 339644 330500 340052 330528
rect 339644 330488 339650 330500
rect 340046 330488 340052 330500
rect 340104 330488 340110 330540
rect 341058 330488 341064 330540
rect 341116 330528 341122 330540
rect 341518 330528 341524 330540
rect 341116 330500 341524 330528
rect 341116 330488 341122 330500
rect 341518 330488 341524 330500
rect 341576 330488 341582 330540
rect 342346 330488 342352 330540
rect 342404 330528 342410 330540
rect 342990 330528 342996 330540
rect 342404 330500 342996 330528
rect 342404 330488 342410 330500
rect 342990 330488 342996 330500
rect 343048 330488 343054 330540
rect 343634 330488 343640 330540
rect 343692 330528 343698 330540
rect 344738 330528 344744 330540
rect 343692 330500 344744 330528
rect 343692 330488 343698 330500
rect 344738 330488 344744 330500
rect 344796 330488 344802 330540
rect 345014 330488 345020 330540
rect 345072 330528 345078 330540
rect 345842 330528 345848 330540
rect 345072 330500 345848 330528
rect 345072 330488 345078 330500
rect 345842 330488 345848 330500
rect 345900 330488 345906 330540
rect 351914 330488 351920 330540
rect 351972 330528 351978 330540
rect 352834 330528 352840 330540
rect 351972 330500 352840 330528
rect 351972 330488 351978 330500
rect 352834 330488 352840 330500
rect 352892 330488 352898 330540
rect 356054 330488 356060 330540
rect 356112 330528 356118 330540
rect 357250 330528 357256 330540
rect 356112 330500 357256 330528
rect 356112 330488 356118 330500
rect 357250 330488 357256 330500
rect 357308 330488 357314 330540
rect 357526 330488 357532 330540
rect 357584 330528 357590 330540
rect 358262 330528 358268 330540
rect 357584 330500 358268 330528
rect 357584 330488 357590 330500
rect 358262 330488 358268 330500
rect 358320 330488 358326 330540
rect 363046 330488 363052 330540
rect 363104 330528 363110 330540
rect 363782 330528 363788 330540
rect 363104 330500 363788 330528
rect 363104 330488 363110 330500
rect 363782 330488 363788 330500
rect 363840 330488 363846 330540
rect 365806 330488 365812 330540
rect 365864 330528 365870 330540
rect 366358 330528 366364 330540
rect 365864 330500 366364 330528
rect 365864 330488 365870 330500
rect 366358 330488 366364 330500
rect 366416 330488 366422 330540
rect 367094 330488 367100 330540
rect 367152 330528 367158 330540
rect 367738 330528 367744 330540
rect 367152 330500 367744 330528
rect 367152 330488 367158 330500
rect 367738 330488 367744 330500
rect 367796 330488 367802 330540
rect 368566 330488 368572 330540
rect 368624 330528 368630 330540
rect 369210 330528 369216 330540
rect 368624 330500 369216 330528
rect 368624 330488 368630 330500
rect 369210 330488 369216 330500
rect 369268 330488 369274 330540
rect 371234 330488 371240 330540
rect 371292 330528 371298 330540
rect 372154 330528 372160 330540
rect 371292 330500 372160 330528
rect 371292 330488 371298 330500
rect 372154 330488 372160 330500
rect 372212 330488 372218 330540
rect 372798 330488 372804 330540
rect 372856 330528 372862 330540
rect 373258 330528 373264 330540
rect 372856 330500 373264 330528
rect 372856 330488 372862 330500
rect 373258 330488 373264 330500
rect 373316 330488 373322 330540
rect 373994 330488 374000 330540
rect 374052 330528 374058 330540
rect 374730 330528 374736 330540
rect 374052 330500 374736 330528
rect 374052 330488 374058 330500
rect 374730 330488 374736 330500
rect 374788 330488 374794 330540
rect 376846 330488 376852 330540
rect 376904 330528 376910 330540
rect 377674 330528 377680 330540
rect 376904 330500 377680 330528
rect 376904 330488 376910 330500
rect 377674 330488 377680 330500
rect 377732 330488 377738 330540
rect 378318 330488 378324 330540
rect 378376 330528 378382 330540
rect 379146 330528 379152 330540
rect 378376 330500 379152 330528
rect 378376 330488 378382 330500
rect 379146 330488 379152 330500
rect 379204 330488 379210 330540
rect 379514 330488 379520 330540
rect 379572 330528 379578 330540
rect 380526 330528 380532 330540
rect 379572 330500 380532 330528
rect 379572 330488 379578 330500
rect 380526 330488 380532 330500
rect 380584 330488 380590 330540
rect 382274 330488 382280 330540
rect 382332 330528 382338 330540
rect 382734 330528 382740 330540
rect 382332 330500 382740 330528
rect 382332 330488 382338 330500
rect 382734 330488 382740 330500
rect 382792 330488 382798 330540
rect 383746 330488 383752 330540
rect 383804 330528 383810 330540
rect 384574 330528 384580 330540
rect 383804 330500 384580 330528
rect 383804 330488 383810 330500
rect 384574 330488 384580 330500
rect 384632 330488 384638 330540
rect 385034 330488 385040 330540
rect 385092 330528 385098 330540
rect 385678 330528 385684 330540
rect 385092 330500 385684 330528
rect 385092 330488 385098 330500
rect 385678 330488 385684 330500
rect 385736 330488 385742 330540
rect 386506 330488 386512 330540
rect 386564 330528 386570 330540
rect 387518 330528 387524 330540
rect 386564 330500 387524 330528
rect 386564 330488 386570 330500
rect 387518 330488 387524 330500
rect 387576 330488 387582 330540
rect 387794 330488 387800 330540
rect 387852 330528 387858 330540
rect 388622 330528 388628 330540
rect 387852 330500 388628 330528
rect 387852 330488 387858 330500
rect 388622 330488 388628 330500
rect 388680 330488 388686 330540
rect 389174 330488 389180 330540
rect 389232 330528 389238 330540
rect 389726 330528 389732 330540
rect 389232 330500 389732 330528
rect 389232 330488 389238 330500
rect 389726 330488 389732 330500
rect 389784 330488 389790 330540
rect 390830 330488 390836 330540
rect 390888 330528 390894 330540
rect 391474 330528 391480 330540
rect 390888 330500 391480 330528
rect 390888 330488 390894 330500
rect 391474 330488 391480 330500
rect 391532 330488 391538 330540
rect 391934 330488 391940 330540
rect 391992 330528 391998 330540
rect 392946 330528 392952 330540
rect 391992 330500 392952 330528
rect 391992 330488 391998 330500
rect 392946 330488 392952 330500
rect 393004 330488 393010 330540
rect 393498 330488 393504 330540
rect 393556 330528 393562 330540
rect 394418 330528 394424 330540
rect 393556 330500 394424 330528
rect 393556 330488 393562 330500
rect 394418 330488 394424 330500
rect 394476 330488 394482 330540
rect 394694 330488 394700 330540
rect 394752 330528 394758 330540
rect 395154 330528 395160 330540
rect 394752 330500 395160 330528
rect 394752 330488 394758 330500
rect 395154 330488 395160 330500
rect 395212 330488 395218 330540
rect 396166 330488 396172 330540
rect 396224 330528 396230 330540
rect 396626 330528 396632 330540
rect 396224 330500 396632 330528
rect 396224 330488 396230 330500
rect 396626 330488 396632 330500
rect 396684 330488 396690 330540
rect 397454 330488 397460 330540
rect 397512 330528 397518 330540
rect 398466 330528 398472 330540
rect 397512 330500 398472 330528
rect 397512 330488 397518 330500
rect 398466 330488 398472 330500
rect 398524 330488 398530 330540
rect 399018 330488 399024 330540
rect 399076 330528 399082 330540
rect 399938 330528 399944 330540
rect 399076 330500 399944 330528
rect 399076 330488 399082 330500
rect 399938 330488 399944 330500
rect 399996 330488 400002 330540
rect 400214 330488 400220 330540
rect 400272 330528 400278 330540
rect 400674 330528 400680 330540
rect 400272 330500 400680 330528
rect 400272 330488 400278 330500
rect 400674 330488 400680 330500
rect 400732 330488 400738 330540
rect 401686 330488 401692 330540
rect 401744 330528 401750 330540
rect 402146 330528 402152 330540
rect 401744 330500 402152 330528
rect 401744 330488 401750 330500
rect 402146 330488 402152 330500
rect 402204 330488 402210 330540
rect 403158 330488 403164 330540
rect 403216 330528 403222 330540
rect 403894 330528 403900 330540
rect 403216 330500 403900 330528
rect 403216 330488 403222 330500
rect 403894 330488 403900 330500
rect 403952 330488 403958 330540
rect 404538 330488 404544 330540
rect 404596 330528 404602 330540
rect 405366 330528 405372 330540
rect 404596 330500 405372 330528
rect 404596 330488 404602 330500
rect 405366 330488 405372 330500
rect 405424 330488 405430 330540
rect 405918 330488 405924 330540
rect 405976 330528 405982 330540
rect 406102 330528 406108 330540
rect 405976 330500 406108 330528
rect 405976 330488 405982 330500
rect 406102 330488 406108 330500
rect 406160 330488 406166 330540
rect 408494 330488 408500 330540
rect 408552 330528 408558 330540
rect 409414 330528 409420 330540
rect 408552 330500 409420 330528
rect 408552 330488 408558 330500
rect 409414 330488 409420 330500
rect 409472 330488 409478 330540
rect 409874 330488 409880 330540
rect 409932 330528 409938 330540
rect 410518 330528 410524 330540
rect 409932 330500 410524 330528
rect 409932 330488 409938 330500
rect 410518 330488 410524 330500
rect 410576 330488 410582 330540
rect 240226 330420 240232 330472
rect 240284 330460 240290 330472
rect 241054 330460 241060 330472
rect 240284 330432 241060 330460
rect 240284 330420 240290 330432
rect 241054 330420 241060 330432
rect 241112 330420 241118 330472
rect 255314 330420 255320 330472
rect 255372 330460 255378 330472
rect 256050 330460 256056 330472
rect 255372 330432 256056 330460
rect 255372 330420 255378 330432
rect 256050 330420 256056 330432
rect 256108 330420 256114 330472
rect 256786 330420 256792 330472
rect 256844 330460 256850 330472
rect 257522 330460 257528 330472
rect 256844 330432 257528 330460
rect 256844 330420 256850 330432
rect 257522 330420 257528 330432
rect 257580 330420 257586 330472
rect 259454 330420 259460 330472
rect 259512 330460 259518 330472
rect 260006 330460 260012 330472
rect 259512 330432 260012 330460
rect 259512 330420 259518 330432
rect 260006 330420 260012 330432
rect 260064 330420 260070 330472
rect 273438 330420 273444 330472
rect 273496 330460 273502 330472
rect 274266 330460 274272 330472
rect 273496 330432 274272 330460
rect 273496 330420 273502 330432
rect 274266 330420 274272 330432
rect 274324 330420 274330 330472
rect 277394 330420 277400 330472
rect 277452 330460 277458 330472
rect 277946 330460 277952 330472
rect 277452 330432 277952 330460
rect 277452 330420 277458 330432
rect 277946 330420 277952 330432
rect 278004 330420 278010 330472
rect 282914 330420 282920 330472
rect 282972 330460 282978 330472
rect 283374 330460 283380 330472
rect 282972 330432 283380 330460
rect 282972 330420 282978 330432
rect 283374 330420 283380 330432
rect 283432 330420 283438 330472
rect 284478 330420 284484 330472
rect 284536 330460 284542 330472
rect 285214 330460 285220 330472
rect 284536 330432 285220 330460
rect 284536 330420 284542 330432
rect 285214 330420 285220 330432
rect 285272 330420 285278 330472
rect 285858 330420 285864 330472
rect 285916 330460 285922 330472
rect 286686 330460 286692 330472
rect 285916 330432 286692 330460
rect 285916 330420 285922 330432
rect 286686 330420 286692 330432
rect 286744 330420 286750 330472
rect 289998 330420 290004 330472
rect 290056 330460 290062 330472
rect 290734 330460 290740 330472
rect 290056 330432 290740 330460
rect 290056 330420 290062 330432
rect 290734 330420 290740 330432
rect 290792 330420 290798 330472
rect 302418 330420 302424 330472
rect 302476 330460 302482 330472
rect 303154 330460 303160 330472
rect 302476 330432 303160 330460
rect 302476 330420 302482 330432
rect 303154 330420 303160 330432
rect 303212 330420 303218 330472
rect 305178 330420 305184 330472
rect 305236 330460 305242 330472
rect 306098 330460 306104 330472
rect 305236 330432 306104 330460
rect 305236 330420 305242 330432
rect 306098 330420 306104 330432
rect 306156 330420 306162 330472
rect 309134 330420 309140 330472
rect 309192 330460 309198 330472
rect 309686 330460 309692 330472
rect 309192 330432 309692 330460
rect 309192 330420 309198 330432
rect 309686 330420 309692 330432
rect 309744 330420 309750 330472
rect 340966 330420 340972 330472
rect 341024 330460 341030 330472
rect 341886 330460 341892 330472
rect 341024 330432 341892 330460
rect 341024 330420 341030 330432
rect 341886 330420 341892 330432
rect 341944 330420 341950 330472
rect 365714 330420 365720 330472
rect 365772 330460 365778 330472
rect 366726 330460 366732 330472
rect 365772 330432 366732 330460
rect 365772 330420 365778 330432
rect 366726 330420 366732 330432
rect 366784 330420 366790 330472
rect 368658 330420 368664 330472
rect 368716 330460 368722 330472
rect 369578 330460 369584 330472
rect 368716 330432 369584 330460
rect 368716 330420 368722 330432
rect 369578 330420 369584 330432
rect 369636 330420 369642 330472
rect 372614 330420 372620 330472
rect 372672 330460 372678 330472
rect 373626 330460 373632 330472
rect 372672 330432 373632 330460
rect 372672 330420 372678 330432
rect 373626 330420 373632 330432
rect 373684 330420 373690 330472
rect 378134 330420 378140 330472
rect 378192 330460 378198 330472
rect 378778 330460 378784 330472
rect 378192 330432 378784 330460
rect 378192 330420 378198 330432
rect 378778 330420 378784 330432
rect 378836 330420 378842 330472
rect 385126 330420 385132 330472
rect 385184 330460 385190 330472
rect 386046 330460 386052 330472
rect 385184 330432 386052 330460
rect 385184 330420 385190 330432
rect 386046 330420 386052 330432
rect 386104 330420 386110 330472
rect 389266 330420 389272 330472
rect 389324 330460 389330 330472
rect 390094 330460 390100 330472
rect 389324 330432 390100 330460
rect 389324 330420 389330 330432
rect 390094 330420 390100 330432
rect 390152 330420 390158 330472
rect 405826 330420 405832 330472
rect 405884 330460 405890 330472
rect 406470 330460 406476 330472
rect 405884 330432 406476 330460
rect 405884 330420 405890 330432
rect 406470 330420 406476 330432
rect 406528 330420 406534 330472
rect 409966 330420 409972 330472
rect 410024 330460 410030 330472
rect 410886 330460 410892 330472
rect 410024 330432 410892 330460
rect 410024 330420 410030 330432
rect 410886 330420 410892 330432
rect 410944 330420 410950 330472
rect 310698 329944 310704 329996
rect 310756 329984 310762 329996
rect 311526 329984 311532 329996
rect 310756 329956 311532 329984
rect 310756 329944 310762 329956
rect 311526 329944 311532 329956
rect 311584 329944 311590 329996
rect 281534 329808 281540 329860
rect 281592 329848 281598 329860
rect 282362 329848 282368 329860
rect 281592 329820 282368 329848
rect 281592 329808 281598 329820
rect 282362 329808 282368 329820
rect 282420 329808 282426 329860
rect 234798 329400 234804 329452
rect 234856 329440 234862 329452
rect 235534 329440 235540 329452
rect 234856 329412 235540 329440
rect 234856 329400 234862 329412
rect 235534 329400 235540 329412
rect 235592 329400 235598 329452
rect 367278 329400 367284 329452
rect 367336 329440 367342 329452
rect 368106 329440 368112 329452
rect 367336 329412 368112 329440
rect 367336 329400 367342 329412
rect 368106 329400 368112 329412
rect 368164 329400 368170 329452
rect 237374 329264 237380 329316
rect 237432 329304 237438 329316
rect 238110 329304 238116 329316
rect 237432 329276 238116 329304
rect 237432 329264 237438 329276
rect 238110 329264 238116 329276
rect 238168 329264 238174 329316
rect 243078 329128 243084 329180
rect 243136 329168 243142 329180
rect 243998 329168 244004 329180
rect 243136 329140 244004 329168
rect 243136 329128 243142 329140
rect 243998 329128 244004 329140
rect 244056 329128 244062 329180
rect 317598 328924 317604 328976
rect 317656 328964 317662 328976
rect 318518 328964 318524 328976
rect 317656 328936 318524 328964
rect 317656 328924 317662 328936
rect 318518 328924 318524 328936
rect 318576 328924 318582 328976
rect 265066 328788 265072 328840
rect 265124 328828 265130 328840
rect 265894 328828 265900 328840
rect 265124 328800 265900 328828
rect 265124 328788 265130 328800
rect 265894 328788 265900 328800
rect 265952 328788 265958 328840
rect 375374 328720 375380 328772
rect 375432 328760 375438 328772
rect 375834 328760 375840 328772
rect 375432 328732 375840 328760
rect 375432 328720 375438 328732
rect 375834 328720 375840 328732
rect 375892 328720 375898 328772
rect 316310 328584 316316 328636
rect 316368 328624 316374 328636
rect 317046 328624 317052 328636
rect 316368 328596 317052 328624
rect 316368 328584 316374 328596
rect 317046 328584 317052 328596
rect 317104 328584 317110 328636
rect 393314 328448 393320 328500
rect 393372 328488 393378 328500
rect 394050 328488 394056 328500
rect 393372 328460 394056 328488
rect 393372 328448 393378 328460
rect 394050 328448 394056 328460
rect 394108 328448 394114 328500
rect 398834 328448 398840 328500
rect 398892 328488 398898 328500
rect 399570 328488 399576 328500
rect 398892 328460 399576 328488
rect 398892 328448 398898 328460
rect 399570 328448 399576 328460
rect 399628 328448 399634 328500
rect 263686 327496 263692 327548
rect 263744 327536 263750 327548
rect 264054 327536 264060 327548
rect 263744 327508 264060 327536
rect 263744 327496 263750 327508
rect 264054 327496 264060 327508
rect 264112 327496 264118 327548
rect 380986 327428 380992 327480
rect 381044 327468 381050 327480
rect 381998 327468 382004 327480
rect 381044 327440 382004 327468
rect 381044 327428 381050 327440
rect 381998 327428 382004 327440
rect 382056 327428 382062 327480
rect 245838 326816 245844 326868
rect 245896 326816 245902 326868
rect 267826 326816 267832 326868
rect 267884 326856 267890 326868
rect 268470 326856 268476 326868
rect 267884 326828 268476 326856
rect 267884 326816 267890 326828
rect 268470 326816 268476 326828
rect 268528 326816 268534 326868
rect 311986 326816 311992 326868
rect 312044 326856 312050 326868
rect 312630 326856 312636 326868
rect 312044 326828 312636 326856
rect 312044 326816 312050 326828
rect 312630 326816 312636 326828
rect 312688 326816 312694 326868
rect 245856 326664 245884 326816
rect 245838 326612 245844 326664
rect 245896 326612 245902 326664
rect 292666 326408 292672 326460
rect 292724 326448 292730 326460
rect 293678 326448 293684 326460
rect 292724 326420 293684 326448
rect 292724 326408 292730 326420
rect 293678 326408 293684 326420
rect 293736 326408 293742 326460
rect 294046 326408 294052 326460
rect 294104 326448 294110 326460
rect 294782 326448 294788 326460
rect 294104 326420 294788 326448
rect 294104 326408 294110 326420
rect 294782 326408 294788 326420
rect 294840 326408 294846 326460
rect 298278 326408 298284 326460
rect 298336 326448 298342 326460
rect 298462 326448 298468 326460
rect 298336 326420 298468 326448
rect 298336 326408 298342 326420
rect 298462 326408 298468 326420
rect 298520 326408 298526 326460
rect 299566 326408 299572 326460
rect 299624 326448 299630 326460
rect 300578 326448 300584 326460
rect 299624 326420 300584 326448
rect 299624 326408 299630 326420
rect 300578 326408 300584 326420
rect 300636 326408 300642 326460
rect 245746 326340 245752 326392
rect 245804 326380 245810 326392
rect 246206 326380 246212 326392
rect 245804 326352 246212 326380
rect 245804 326340 245810 326352
rect 246206 326340 246212 326352
rect 246264 326340 246270 326392
rect 247034 326340 247040 326392
rect 247092 326380 247098 326392
rect 247954 326380 247960 326392
rect 247092 326352 247960 326380
rect 247092 326340 247098 326352
rect 247954 326340 247960 326352
rect 248012 326340 248018 326392
rect 249886 326340 249892 326392
rect 249944 326380 249950 326392
rect 250898 326380 250904 326392
rect 249944 326352 250904 326380
rect 249944 326340 249950 326352
rect 250898 326340 250904 326352
rect 250956 326340 250962 326392
rect 251174 326340 251180 326392
rect 251232 326380 251238 326392
rect 251634 326380 251640 326392
rect 251232 326352 251640 326380
rect 251232 326340 251238 326352
rect 251634 326340 251640 326352
rect 251692 326340 251698 326392
rect 292574 326340 292580 326392
rect 292632 326380 292638 326392
rect 293310 326380 293316 326392
rect 292632 326352 293316 326380
rect 292632 326340 292638 326352
rect 293310 326340 293316 326352
rect 293368 326340 293374 326392
rect 293954 326340 293960 326392
rect 294012 326380 294018 326392
rect 294414 326380 294420 326392
rect 294012 326352 294420 326380
rect 294012 326340 294018 326352
rect 294414 326340 294420 326352
rect 294472 326340 294478 326392
rect 298094 326340 298100 326392
rect 298152 326380 298158 326392
rect 298738 326380 298744 326392
rect 298152 326352 298744 326380
rect 298152 326340 298158 326352
rect 298738 326340 298744 326352
rect 298796 326340 298802 326392
rect 299474 326340 299480 326392
rect 299532 326380 299538 326392
rect 299842 326380 299848 326392
rect 299532 326352 299848 326380
rect 299532 326340 299538 326352
rect 299842 326340 299848 326352
rect 299900 326340 299906 326392
rect 300946 326340 300952 326392
rect 301004 326380 301010 326392
rect 301682 326380 301688 326392
rect 301004 326352 301688 326380
rect 301004 326340 301010 326352
rect 301682 326340 301688 326352
rect 301740 326340 301746 326392
rect 321646 326340 321652 326392
rect 321704 326380 321710 326392
rect 321830 326380 321836 326392
rect 321704 326352 321836 326380
rect 321704 326340 321710 326352
rect 321830 326340 321836 326352
rect 321888 326340 321894 326392
rect 322934 326340 322940 326392
rect 322992 326380 322998 326392
rect 323578 326380 323584 326392
rect 322992 326352 323584 326380
rect 322992 326340 322998 326352
rect 323578 326340 323584 326352
rect 323636 326340 323642 326392
rect 327166 326340 327172 326392
rect 327224 326380 327230 326392
rect 327626 326380 327632 326392
rect 327224 326352 327632 326380
rect 327224 326340 327230 326352
rect 327626 326340 327632 326352
rect 327684 326340 327690 326392
rect 329926 326340 329932 326392
rect 329984 326380 329990 326392
rect 330938 326380 330944 326392
rect 329984 326352 330944 326380
rect 329984 326340 329990 326352
rect 330938 326340 330944 326352
rect 330996 326340 331002 326392
rect 294138 326272 294144 326324
rect 294196 326312 294202 326324
rect 295150 326312 295156 326324
rect 294196 326284 295156 326312
rect 294196 326272 294202 326284
rect 295150 326272 295156 326284
rect 295208 326272 295214 326324
rect 296714 326136 296720 326188
rect 296772 326176 296778 326188
rect 297634 326176 297640 326188
rect 296772 326148 297640 326176
rect 296772 326136 296778 326148
rect 297634 326136 297640 326148
rect 297692 326136 297698 326188
rect 394786 326068 394792 326120
rect 394844 326108 394850 326120
rect 395522 326108 395528 326120
rect 394844 326080 395528 326108
rect 394844 326068 394850 326080
rect 395522 326068 395528 326080
rect 395580 326068 395586 326120
rect 400306 326068 400312 326120
rect 400364 326108 400370 326120
rect 401042 326108 401048 326120
rect 400364 326080 401048 326108
rect 400364 326068 400370 326080
rect 401042 326068 401048 326080
rect 401100 326068 401106 326120
rect 252646 326000 252652 326052
rect 252704 326040 252710 326052
rect 253106 326040 253112 326052
rect 252704 326012 253112 326040
rect 252704 326000 252710 326012
rect 253106 326000 253112 326012
rect 253164 326000 253170 326052
rect 242894 325728 242900 325780
rect 242952 325768 242958 325780
rect 243630 325768 243636 325780
rect 242952 325740 243636 325768
rect 242952 325728 242958 325740
rect 243630 325728 243636 325740
rect 243688 325728 243694 325780
rect 577314 325456 577320 325508
rect 577372 325496 577378 325508
rect 580718 325496 580724 325508
rect 577372 325468 580724 325496
rect 577372 325456 577378 325468
rect 580718 325456 580724 325468
rect 580776 325456 580782 325508
rect 249794 323824 249800 323876
rect 249852 323864 249858 323876
rect 250530 323864 250536 323876
rect 249852 323836 250536 323864
rect 249852 323824 249858 323836
rect 250530 323824 250536 323836
rect 250588 323824 250594 323876
rect 325786 323552 325792 323604
rect 325844 323592 325850 323604
rect 325970 323592 325976 323604
rect 325844 323564 325976 323592
rect 325844 323552 325850 323564
rect 325970 323552 325976 323564
rect 326028 323552 326034 323604
rect 323118 323212 323124 323264
rect 323176 323252 323182 323264
rect 323946 323252 323952 323264
rect 323176 323224 323952 323252
rect 323176 323212 323182 323224
rect 323946 323212 323952 323224
rect 324004 323212 324010 323264
rect 251266 322192 251272 322244
rect 251324 322232 251330 322244
rect 252002 322232 252008 322244
rect 251324 322204 252008 322232
rect 251324 322192 251330 322204
rect 252002 322192 252008 322204
rect 252060 322192 252066 322244
rect 328454 320832 328460 320884
rect 328512 320872 328518 320884
rect 328638 320872 328644 320884
rect 328512 320844 328644 320872
rect 328512 320832 328518 320844
rect 328638 320832 328644 320844
rect 328696 320832 328702 320884
rect 245654 319200 245660 319252
rect 245712 319240 245718 319252
rect 245930 319240 245936 319252
rect 245712 319212 245936 319240
rect 245712 319200 245718 319212
rect 245930 319200 245936 319212
rect 245988 319200 245994 319252
rect 3326 306280 3332 306332
rect 3384 306320 3390 306332
rect 233602 306320 233608 306332
rect 3384 306292 233608 306320
rect 3384 306280 3390 306292
rect 233602 306280 233608 306292
rect 233660 306280 233666 306332
rect 577406 299412 577412 299464
rect 577464 299452 577470 299464
rect 579614 299452 579620 299464
rect 577464 299424 579620 299452
rect 577464 299412 577470 299424
rect 579614 299412 579620 299424
rect 579672 299412 579678 299464
rect 578142 273164 578148 273216
rect 578200 273204 578206 273216
rect 579614 273204 579620 273216
rect 578200 273176 579620 273204
rect 578200 273164 578206 273176
rect 579614 273164 579620 273176
rect 579672 273164 579678 273216
rect 574830 259360 574836 259412
rect 574888 259400 574894 259412
rect 579798 259400 579804 259412
rect 574888 259372 579804 259400
rect 574888 259360 574894 259372
rect 579798 259360 579804 259372
rect 579856 259360 579862 259412
rect 3142 255212 3148 255264
rect 3200 255252 3206 255264
rect 233786 255252 233792 255264
rect 3200 255224 233792 255252
rect 3200 255212 3206 255224
rect 233786 255212 233792 255224
rect 233844 255212 233850 255264
rect 3510 241408 3516 241460
rect 3568 241448 3574 241460
rect 234154 241448 234160 241460
rect 3568 241420 234160 241448
rect 3568 241408 3574 241420
rect 234154 241408 234160 241420
rect 234212 241408 234218 241460
rect 577958 233180 577964 233232
rect 578016 233220 578022 233232
rect 579614 233220 579620 233232
rect 578016 233192 579620 233220
rect 578016 233180 578022 233192
rect 579614 233180 579620 233192
rect 579672 233180 579678 233232
rect 574738 219376 574744 219428
rect 574796 219416 574802 219428
rect 580166 219416 580172 219428
rect 574796 219388 580172 219416
rect 574796 219376 574802 219388
rect 580166 219376 580172 219388
rect 580224 219376 580230 219428
rect 3418 202784 3424 202836
rect 3476 202824 3482 202836
rect 233970 202824 233976 202836
rect 3476 202796 233976 202824
rect 3476 202784 3482 202796
rect 233970 202784 233976 202796
rect 234028 202784 234034 202836
rect 578050 193128 578056 193180
rect 578108 193168 578114 193180
rect 579614 193168 579620 193180
rect 578108 193140 579620 193168
rect 578108 193128 578114 193140
rect 579614 193128 579620 193140
rect 579672 193128 579678 193180
rect 3418 188980 3424 189032
rect 3476 189020 3482 189032
rect 234246 189020 234252 189032
rect 3476 188992 234252 189020
rect 3476 188980 3482 188992
rect 234246 188980 234252 188992
rect 234304 188980 234310 189032
rect 577774 179324 577780 179376
rect 577832 179364 577838 179376
rect 580074 179364 580080 179376
rect 577832 179336 580080 179364
rect 577832 179324 577838 179336
rect 580074 179324 580080 179336
rect 580132 179324 580138 179376
rect 2774 163752 2780 163804
rect 2832 163792 2838 163804
rect 4890 163792 4896 163804
rect 2832 163764 4896 163792
rect 2832 163752 2838 163764
rect 4890 163752 4896 163764
rect 4948 163752 4954 163804
rect 3418 150356 3424 150408
rect 3476 150396 3482 150408
rect 231210 150396 231216 150408
rect 3476 150368 231216 150396
rect 3476 150356 3482 150368
rect 231210 150356 231216 150368
rect 231268 150356 231274 150408
rect 577590 139340 577596 139392
rect 577648 139380 577654 139392
rect 579614 139380 579620 139392
rect 577648 139352 579620 139380
rect 577648 139340 577654 139352
rect 579614 139340 579620 139352
rect 579672 139340 579678 139392
rect 3234 137912 3240 137964
rect 3292 137952 3298 137964
rect 234062 137952 234068 137964
rect 3292 137924 234068 137952
rect 3292 137912 3298 137924
rect 234062 137912 234068 137924
rect 234120 137912 234126 137964
rect 577866 112956 577872 113008
rect 577924 112996 577930 113008
rect 580534 112996 580540 113008
rect 577924 112968 580540 112996
rect 577924 112956 577930 112968
rect 580534 112956 580540 112968
rect 580592 112956 580598 113008
rect 234338 100648 234344 100700
rect 234396 100688 234402 100700
rect 580166 100688 580172 100700
rect 234396 100660 580172 100688
rect 234396 100648 234402 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3418 97928 3424 97980
rect 3476 97968 3482 97980
rect 231118 97968 231124 97980
rect 3476 97940 231124 97968
rect 3476 97928 3482 97940
rect 231118 97928 231124 97940
rect 231176 97928 231182 97980
rect 3142 85484 3148 85536
rect 3200 85524 3206 85536
rect 233878 85524 233884 85536
rect 3200 85496 233884 85524
rect 3200 85484 3206 85496
rect 233878 85484 233884 85496
rect 233936 85484 233942 85536
rect 577682 73108 577688 73160
rect 577740 73148 577746 73160
rect 579706 73148 579712 73160
rect 577740 73120 579712 73148
rect 577740 73108 577746 73120
rect 579706 73108 579712 73120
rect 579764 73108 579770 73160
rect 2774 71612 2780 71664
rect 2832 71652 2838 71664
rect 4798 71652 4804 71664
rect 2832 71624 4804 71652
rect 2832 71612 2838 71624
rect 4798 71612 4804 71624
rect 4856 71612 4862 71664
rect 234430 60664 234436 60716
rect 234488 60704 234494 60716
rect 580166 60704 580172 60716
rect 234488 60676 580172 60704
rect 234488 60664 234494 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 577498 33056 577504 33108
rect 577556 33096 577562 33108
rect 579614 33096 579620 33108
rect 577556 33068 579620 33096
rect 577556 33056 577562 33068
rect 579614 33056 579620 33068
rect 579672 33056 579678 33108
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 414934 20652 414940 20664
rect 3476 20624 414940 20652
rect 3476 20612 3482 20624
rect 414934 20612 414940 20624
rect 414992 20612 414998 20664
rect 234522 20544 234528 20596
rect 234580 20584 234586 20596
rect 580166 20584 580172 20596
rect 234580 20556 580172 20584
rect 234580 20544 234586 20556
rect 580166 20544 580172 20556
rect 580224 20544 580230 20596
rect 74534 20272 74540 20324
rect 74592 20312 74598 20324
rect 258258 20312 258264 20324
rect 74592 20284 258264 20312
rect 74592 20272 74598 20284
rect 258258 20272 258264 20284
rect 258316 20272 258322 20324
rect 70394 20204 70400 20256
rect 70452 20244 70458 20256
rect 256878 20244 256884 20256
rect 70452 20216 256884 20244
rect 70452 20204 70458 20216
rect 256878 20204 256884 20216
rect 256936 20204 256942 20256
rect 67634 20136 67640 20188
rect 67692 20176 67698 20188
rect 255590 20176 255596 20188
rect 67692 20148 255596 20176
rect 67692 20136 67698 20148
rect 255590 20136 255596 20148
rect 255648 20136 255654 20188
rect 63494 20068 63500 20120
rect 63552 20108 63558 20120
rect 254210 20108 254216 20120
rect 63552 20080 254216 20108
rect 63552 20068 63558 20080
rect 254210 20068 254216 20080
rect 254268 20068 254274 20120
rect 60734 20000 60740 20052
rect 60792 20040 60798 20052
rect 252830 20040 252836 20052
rect 60792 20012 252836 20040
rect 60792 20000 60798 20012
rect 252830 20000 252836 20012
rect 252888 20000 252894 20052
rect 234706 19932 234712 19984
rect 234764 19972 234770 19984
rect 580258 19972 580264 19984
rect 234764 19944 580264 19972
rect 234764 19932 234770 19944
rect 580258 19932 580264 19944
rect 580316 19932 580322 19984
rect 149054 19252 149060 19304
rect 149112 19292 149118 19304
rect 280430 19292 280436 19304
rect 149112 19264 280436 19292
rect 149112 19252 149118 19264
rect 280430 19252 280436 19264
rect 280488 19252 280494 19304
rect 144914 19184 144920 19236
rect 144972 19224 144978 19236
rect 279050 19224 279056 19236
rect 144972 19196 279056 19224
rect 144972 19184 144978 19196
rect 279050 19184 279056 19196
rect 279108 19184 279114 19236
rect 62114 19116 62120 19168
rect 62172 19156 62178 19168
rect 254118 19156 254124 19168
rect 62172 19128 254124 19156
rect 62172 19116 62178 19128
rect 254118 19116 254124 19128
rect 254176 19116 254182 19168
rect 59354 19048 59360 19100
rect 59412 19088 59418 19100
rect 252646 19088 252652 19100
rect 59412 19060 252652 19088
rect 59412 19048 59418 19060
rect 252646 19048 252652 19060
rect 252704 19048 252710 19100
rect 55214 18980 55220 19032
rect 55272 19020 55278 19032
rect 251266 19020 251272 19032
rect 55272 18992 251272 19020
rect 55272 18980 55278 18992
rect 251266 18980 251272 18992
rect 251324 18980 251330 19032
rect 56594 18912 56600 18964
rect 56652 18952 56658 18964
rect 252738 18952 252744 18964
rect 56652 18924 252744 18952
rect 56652 18912 56658 18924
rect 252738 18912 252744 18924
rect 252796 18912 252802 18964
rect 52454 18844 52460 18896
rect 52512 18884 52518 18896
rect 251358 18884 251364 18896
rect 52512 18856 251364 18884
rect 52512 18844 52518 18856
rect 251358 18844 251364 18856
rect 251416 18844 251422 18896
rect 49694 18776 49700 18828
rect 49752 18816 49758 18828
rect 250070 18816 250076 18828
rect 49752 18788 250076 18816
rect 49752 18776 49758 18788
rect 250070 18776 250076 18788
rect 250128 18776 250134 18828
rect 44174 18708 44180 18760
rect 44232 18748 44238 18760
rect 248598 18748 248604 18760
rect 44232 18720 248604 18748
rect 44232 18708 44238 18720
rect 248598 18708 248604 18720
rect 248656 18708 248662 18760
rect 41414 18640 41420 18692
rect 41472 18680 41478 18692
rect 247218 18680 247224 18692
rect 41472 18652 247224 18680
rect 41472 18640 41478 18652
rect 247218 18640 247224 18652
rect 247276 18640 247282 18692
rect 37274 18572 37280 18624
rect 37332 18612 37338 18624
rect 245930 18612 245936 18624
rect 37332 18584 245936 18612
rect 37332 18572 37338 18584
rect 245930 18572 245936 18584
rect 245988 18572 245994 18624
rect 151814 18504 151820 18556
rect 151872 18544 151878 18556
rect 281718 18544 281724 18556
rect 151872 18516 281724 18544
rect 151872 18504 151878 18516
rect 281718 18504 281724 18516
rect 281776 18504 281782 18556
rect 198734 18436 198740 18488
rect 198792 18476 198798 18488
rect 295518 18476 295524 18488
rect 198792 18448 295524 18476
rect 198792 18436 198798 18448
rect 295518 18436 295524 18448
rect 295576 18436 295582 18488
rect 201494 18368 201500 18420
rect 201552 18408 201558 18420
rect 296990 18408 296996 18420
rect 201552 18380 296996 18408
rect 201552 18368 201558 18380
rect 296990 18368 296996 18380
rect 297048 18368 297054 18420
rect 204254 17892 204260 17944
rect 204312 17932 204318 17944
rect 298278 17932 298284 17944
rect 204312 17904 298284 17932
rect 204312 17892 204318 17904
rect 298278 17892 298284 17904
rect 298336 17892 298342 17944
rect 201586 17824 201592 17876
rect 201644 17864 201650 17876
rect 296898 17864 296904 17876
rect 201644 17836 296904 17864
rect 201644 17824 201650 17836
rect 296898 17824 296904 17836
rect 296956 17824 296962 17876
rect 194594 17756 194600 17808
rect 194652 17796 194658 17808
rect 294138 17796 294144 17808
rect 194652 17768 294144 17796
rect 194652 17756 194658 17768
rect 294138 17756 294144 17768
rect 294196 17756 294202 17808
rect 191834 17688 191840 17740
rect 191892 17728 191898 17740
rect 294230 17728 294236 17740
rect 191892 17700 294236 17728
rect 191892 17688 191898 17700
rect 294230 17688 294236 17700
rect 294288 17688 294294 17740
rect 153194 17620 153200 17672
rect 153252 17660 153258 17672
rect 281534 17660 281540 17672
rect 153252 17632 281540 17660
rect 153252 17620 153258 17632
rect 281534 17620 281540 17632
rect 281592 17620 281598 17672
rect 151906 17552 151912 17604
rect 151964 17592 151970 17604
rect 281626 17592 281632 17604
rect 151964 17564 281632 17592
rect 151964 17552 151970 17564
rect 281626 17552 281632 17564
rect 281684 17552 281690 17604
rect 150434 17484 150440 17536
rect 150492 17524 150498 17536
rect 280338 17524 280344 17536
rect 150492 17496 280344 17524
rect 150492 17484 150498 17496
rect 280338 17484 280344 17496
rect 280396 17484 280402 17536
rect 147674 17416 147680 17468
rect 147732 17456 147738 17468
rect 280154 17456 280160 17468
rect 147732 17428 280160 17456
rect 147732 17416 147738 17428
rect 280154 17416 280160 17428
rect 280212 17416 280218 17468
rect 146294 17348 146300 17400
rect 146352 17388 146358 17400
rect 280246 17388 280252 17400
rect 146352 17360 280252 17388
rect 146352 17348 146358 17360
rect 280246 17348 280252 17360
rect 280304 17348 280310 17400
rect 143534 17280 143540 17332
rect 143592 17320 143598 17332
rect 278866 17320 278872 17332
rect 143592 17292 278872 17320
rect 143592 17280 143598 17292
rect 278866 17280 278872 17292
rect 278924 17280 278930 17332
rect 142154 17212 142160 17264
rect 142212 17252 142218 17264
rect 278958 17252 278964 17264
rect 142212 17224 278964 17252
rect 142212 17212 142218 17224
rect 278958 17212 278964 17224
rect 279016 17212 279022 17264
rect 208394 17144 208400 17196
rect 208452 17184 208458 17196
rect 298370 17184 298376 17196
rect 208452 17156 298376 17184
rect 208452 17144 208458 17156
rect 298370 17144 298376 17156
rect 298428 17144 298434 17196
rect 211154 17076 211160 17128
rect 211212 17116 211218 17128
rect 299750 17116 299756 17128
rect 211212 17088 299756 17116
rect 211212 17076 211218 17088
rect 299750 17076 299756 17088
rect 299808 17076 299814 17128
rect 215294 17008 215300 17060
rect 215352 17048 215358 17060
rect 301038 17048 301044 17060
rect 215352 17020 301044 17048
rect 215352 17008 215358 17020
rect 301038 17008 301044 17020
rect 301096 17008 301102 17060
rect 171962 16532 171968 16584
rect 172020 16572 172026 16584
rect 287330 16572 287336 16584
rect 172020 16544 287336 16572
rect 172020 16532 172026 16544
rect 287330 16532 287336 16544
rect 287388 16532 287394 16584
rect 168374 16464 168380 16516
rect 168432 16504 168438 16516
rect 285858 16504 285864 16516
rect 168432 16476 285864 16504
rect 168432 16464 168438 16476
rect 285858 16464 285864 16476
rect 285916 16464 285922 16516
rect 164418 16396 164424 16448
rect 164476 16436 164482 16448
rect 285950 16436 285956 16448
rect 164476 16408 285956 16436
rect 164476 16396 164482 16408
rect 285950 16396 285956 16408
rect 286008 16396 286014 16448
rect 161290 16328 161296 16380
rect 161348 16368 161354 16380
rect 284662 16368 284668 16380
rect 161348 16340 284668 16368
rect 161348 16328 161354 16340
rect 284662 16328 284668 16340
rect 284720 16328 284726 16380
rect 125594 16260 125600 16312
rect 125652 16300 125658 16312
rect 273530 16300 273536 16312
rect 125652 16272 273536 16300
rect 125652 16260 125658 16272
rect 273530 16260 273536 16272
rect 273588 16260 273594 16312
rect 123018 16192 123024 16244
rect 123076 16232 123082 16244
rect 271966 16232 271972 16244
rect 123076 16204 271972 16232
rect 123076 16192 123082 16204
rect 271966 16192 271972 16204
rect 272024 16192 272030 16244
rect 118694 16124 118700 16176
rect 118752 16164 118758 16176
rect 272058 16164 272064 16176
rect 118752 16136 272064 16164
rect 118752 16124 118758 16136
rect 272058 16124 272064 16136
rect 272116 16124 272122 16176
rect 116394 16056 116400 16108
rect 116452 16096 116458 16108
rect 270678 16096 270684 16108
rect 116452 16068 270684 16096
rect 116452 16056 116458 16068
rect 270678 16056 270684 16068
rect 270736 16056 270742 16108
rect 34514 15988 34520 16040
rect 34572 16028 34578 16040
rect 245838 16028 245844 16040
rect 34572 16000 245844 16028
rect 34572 15988 34578 16000
rect 245838 15988 245844 16000
rect 245896 15988 245902 16040
rect 368658 15988 368664 16040
rect 368716 16028 368722 16040
rect 436738 16028 436744 16040
rect 368716 16000 436744 16028
rect 368716 15988 368722 16000
rect 436738 15988 436744 16000
rect 436796 15988 436802 16040
rect 30834 15920 30840 15972
rect 30892 15960 30898 15972
rect 244366 15960 244372 15972
rect 30892 15932 244372 15960
rect 30892 15920 30898 15932
rect 244366 15920 244372 15932
rect 244424 15920 244430 15972
rect 378410 15920 378416 15972
rect 378468 15960 378474 15972
rect 465166 15960 465172 15972
rect 378468 15932 465172 15960
rect 378468 15920 378474 15932
rect 465166 15920 465172 15932
rect 465224 15920 465230 15972
rect 27706 15852 27712 15904
rect 27764 15892 27770 15904
rect 243170 15892 243176 15904
rect 27764 15864 243176 15892
rect 27764 15852 27770 15864
rect 243170 15852 243176 15864
rect 243228 15852 243234 15904
rect 412818 15852 412824 15904
rect 412876 15892 412882 15904
rect 578602 15892 578608 15904
rect 412876 15864 578608 15892
rect 412876 15852 412882 15864
rect 578602 15852 578608 15864
rect 578660 15852 578666 15904
rect 218054 15784 218060 15836
rect 218112 15824 218118 15836
rect 302510 15824 302516 15836
rect 218112 15796 302516 15824
rect 218112 15784 218118 15796
rect 302510 15784 302516 15796
rect 302568 15784 302574 15836
rect 221090 15716 221096 15768
rect 221148 15756 221154 15768
rect 302418 15756 302424 15768
rect 221148 15728 302424 15756
rect 221148 15716 221154 15728
rect 302418 15716 302424 15728
rect 302476 15716 302482 15768
rect 225138 15648 225144 15700
rect 225196 15688 225202 15700
rect 303890 15688 303896 15700
rect 225196 15660 303896 15688
rect 225196 15648 225202 15660
rect 303890 15648 303896 15660
rect 303948 15648 303954 15700
rect 102226 15104 102232 15156
rect 102284 15144 102290 15156
rect 266446 15144 266452 15156
rect 102284 15116 266452 15144
rect 102284 15104 102290 15116
rect 266446 15104 266452 15116
rect 266504 15104 266510 15156
rect 394878 15104 394884 15156
rect 394936 15144 394942 15156
rect 517882 15144 517888 15156
rect 394936 15116 517888 15144
rect 394936 15104 394942 15116
rect 517882 15104 517888 15116
rect 517940 15104 517946 15156
rect 98178 15036 98184 15088
rect 98236 15076 98242 15088
rect 265158 15076 265164 15088
rect 98236 15048 265164 15076
rect 98236 15036 98242 15048
rect 265158 15036 265164 15048
rect 265216 15036 265222 15088
rect 396258 15036 396264 15088
rect 396316 15076 396322 15088
rect 521654 15076 521660 15088
rect 396316 15048 521660 15076
rect 396316 15036 396322 15048
rect 521654 15036 521660 15048
rect 521712 15036 521718 15088
rect 93854 14968 93860 15020
rect 93912 15008 93918 15020
rect 263686 15008 263692 15020
rect 93912 14980 263692 15008
rect 93912 14968 93918 14980
rect 263686 14968 263692 14980
rect 263744 14968 263750 15020
rect 396350 14968 396356 15020
rect 396408 15008 396414 15020
rect 525426 15008 525432 15020
rect 396408 14980 525432 15008
rect 396408 14968 396414 14980
rect 525426 14968 525432 14980
rect 525484 14968 525490 15020
rect 91554 14900 91560 14952
rect 91612 14940 91618 14952
rect 262398 14940 262404 14952
rect 91612 14912 262404 14940
rect 91612 14900 91618 14912
rect 262398 14900 262404 14912
rect 262456 14900 262462 14952
rect 397730 14900 397736 14952
rect 397788 14940 397794 14952
rect 528554 14940 528560 14952
rect 397788 14912 528560 14940
rect 397788 14900 397794 14912
rect 528554 14900 528560 14912
rect 528612 14900 528618 14952
rect 87506 14832 87512 14884
rect 87564 14872 87570 14884
rect 261018 14872 261024 14884
rect 87564 14844 261024 14872
rect 87564 14832 87570 14844
rect 261018 14832 261024 14844
rect 261076 14832 261082 14884
rect 399110 14832 399116 14884
rect 399168 14872 399174 14884
rect 532050 14872 532056 14884
rect 399168 14844 532056 14872
rect 399168 14832 399174 14844
rect 532050 14832 532056 14844
rect 532108 14832 532114 14884
rect 84194 14764 84200 14816
rect 84252 14804 84258 14816
rect 260926 14804 260932 14816
rect 84252 14776 260932 14804
rect 84252 14764 84258 14776
rect 260926 14764 260932 14776
rect 260984 14764 260990 14816
rect 400398 14764 400404 14816
rect 400456 14804 400462 14816
rect 536098 14804 536104 14816
rect 400456 14776 536104 14804
rect 400456 14764 400462 14776
rect 536098 14764 536104 14776
rect 536156 14764 536162 14816
rect 80882 14696 80888 14748
rect 80940 14736 80946 14748
rect 259730 14736 259736 14748
rect 80940 14708 259736 14736
rect 80940 14696 80946 14708
rect 259730 14696 259736 14708
rect 259788 14696 259794 14748
rect 401778 14696 401784 14748
rect 401836 14736 401842 14748
rect 539594 14736 539600 14748
rect 401836 14708 539600 14736
rect 401836 14696 401842 14708
rect 539594 14696 539600 14708
rect 539652 14696 539658 14748
rect 77386 14628 77392 14680
rect 77444 14668 77450 14680
rect 258166 14668 258172 14680
rect 77444 14640 258172 14668
rect 77444 14628 77450 14640
rect 258166 14628 258172 14640
rect 258224 14628 258230 14680
rect 401870 14628 401876 14680
rect 401928 14668 401934 14680
rect 542722 14668 542728 14680
rect 401928 14640 542728 14668
rect 401928 14628 401934 14640
rect 542722 14628 542728 14640
rect 542780 14628 542786 14680
rect 73338 14560 73344 14612
rect 73396 14600 73402 14612
rect 256786 14600 256792 14612
rect 73396 14572 256792 14600
rect 73396 14560 73402 14572
rect 256786 14560 256792 14572
rect 256844 14560 256850 14612
rect 403250 14560 403256 14612
rect 403308 14600 403314 14612
rect 546494 14600 546500 14612
rect 403308 14572 546500 14600
rect 403308 14560 403314 14572
rect 546494 14560 546500 14572
rect 546552 14560 546558 14612
rect 69842 14492 69848 14544
rect 69900 14532 69906 14544
rect 255498 14532 255504 14544
rect 69900 14504 255504 14532
rect 69900 14492 69906 14504
rect 255498 14492 255504 14504
rect 255556 14492 255562 14544
rect 406010 14492 406016 14544
rect 406068 14532 406074 14544
rect 553762 14532 553768 14544
rect 406068 14504 553768 14532
rect 406068 14492 406074 14504
rect 553762 14492 553768 14504
rect 553820 14492 553826 14544
rect 66714 14424 66720 14476
rect 66772 14464 66778 14476
rect 255406 14464 255412 14476
rect 66772 14436 255412 14464
rect 66772 14424 66778 14436
rect 255406 14424 255412 14436
rect 255464 14424 255470 14476
rect 408770 14424 408776 14476
rect 408828 14464 408834 14476
rect 564434 14464 564440 14476
rect 408828 14436 564440 14464
rect 408828 14424 408834 14436
rect 564434 14424 564440 14436
rect 564492 14424 564498 14476
rect 105722 14356 105728 14408
rect 105780 14396 105786 14408
rect 266538 14396 266544 14408
rect 105780 14368 266544 14396
rect 105780 14356 105786 14368
rect 266538 14356 266544 14368
rect 266596 14356 266602 14408
rect 393590 14356 393596 14408
rect 393648 14396 393654 14408
rect 514754 14396 514760 14408
rect 393648 14368 514760 14396
rect 393648 14356 393654 14368
rect 514754 14356 514760 14368
rect 514812 14356 514818 14408
rect 109034 14288 109040 14340
rect 109092 14328 109098 14340
rect 267826 14328 267832 14340
rect 109092 14300 267832 14328
rect 109092 14288 109098 14300
rect 267826 14288 267832 14300
rect 267884 14288 267890 14340
rect 390830 14288 390836 14340
rect 390888 14328 390894 14340
rect 507210 14328 507216 14340
rect 390888 14300 507216 14328
rect 390888 14288 390894 14300
rect 507210 14288 507216 14300
rect 507268 14288 507274 14340
rect 112346 14220 112352 14272
rect 112404 14260 112410 14272
rect 269298 14260 269304 14272
rect 112404 14232 269304 14260
rect 112404 14220 112410 14232
rect 269298 14220 269304 14232
rect 269356 14220 269362 14272
rect 367278 14220 367284 14272
rect 367336 14260 367342 14272
rect 432046 14260 432052 14272
rect 367336 14232 432052 14260
rect 367336 14220 367342 14232
rect 432046 14220 432052 14232
rect 432104 14220 432110 14272
rect 118786 13744 118792 13796
rect 118844 13784 118850 13796
rect 270770 13784 270776 13796
rect 118844 13756 270776 13784
rect 118844 13744 118850 13756
rect 270770 13744 270776 13756
rect 270828 13744 270834 13796
rect 367186 13744 367192 13796
rect 367244 13784 367250 13796
rect 428458 13784 428464 13796
rect 367244 13756 428464 13784
rect 367244 13744 367250 13756
rect 428458 13744 428464 13756
rect 428516 13744 428522 13796
rect 114738 13676 114744 13728
rect 114796 13716 114802 13728
rect 270586 13716 270592 13728
rect 114796 13688 270592 13716
rect 114796 13676 114802 13688
rect 270586 13676 270592 13688
rect 270644 13676 270650 13728
rect 372798 13676 372804 13728
rect 372856 13716 372862 13728
rect 448514 13716 448520 13728
rect 372856 13688 448520 13716
rect 372856 13676 372862 13688
rect 448514 13676 448520 13688
rect 448572 13676 448578 13728
rect 110414 13608 110420 13660
rect 110472 13648 110478 13660
rect 269206 13648 269212 13660
rect 110472 13620 269212 13648
rect 110472 13608 110478 13620
rect 269206 13608 269212 13620
rect 269264 13608 269270 13660
rect 374086 13608 374092 13660
rect 374144 13648 374150 13660
rect 451642 13648 451648 13660
rect 374144 13620 451648 13648
rect 374144 13608 374150 13620
rect 451642 13608 451648 13620
rect 451700 13608 451706 13660
rect 108114 13540 108120 13592
rect 108172 13580 108178 13592
rect 267918 13580 267924 13592
rect 108172 13552 267924 13580
rect 108172 13540 108178 13552
rect 267918 13540 267924 13552
rect 267976 13540 267982 13592
rect 375466 13540 375472 13592
rect 375524 13580 375530 13592
rect 455690 13580 455696 13592
rect 375524 13552 455696 13580
rect 375524 13540 375530 13552
rect 455690 13540 455696 13552
rect 455748 13540 455754 13592
rect 104066 13472 104072 13524
rect 104124 13512 104130 13524
rect 266630 13512 266636 13524
rect 104124 13484 266636 13512
rect 104124 13472 104130 13484
rect 266630 13472 266636 13484
rect 266688 13472 266694 13524
rect 376938 13472 376944 13524
rect 376996 13512 377002 13524
rect 459186 13512 459192 13524
rect 376996 13484 459192 13512
rect 376996 13472 377002 13484
rect 459186 13472 459192 13484
rect 459244 13472 459250 13524
rect 100754 13404 100760 13456
rect 100812 13444 100818 13456
rect 265066 13444 265072 13456
rect 100812 13416 265072 13444
rect 100812 13404 100818 13416
rect 265066 13404 265072 13416
rect 265124 13404 265130 13456
rect 376846 13404 376852 13456
rect 376904 13444 376910 13456
rect 462314 13444 462320 13456
rect 376904 13416 462320 13444
rect 376904 13404 376910 13416
rect 462314 13404 462320 13416
rect 462372 13404 462378 13456
rect 97442 13336 97448 13388
rect 97500 13376 97506 13388
rect 265250 13376 265256 13388
rect 97500 13348 265256 13376
rect 97500 13336 97506 13348
rect 265250 13336 265256 13348
rect 265308 13336 265314 13388
rect 393498 13336 393504 13388
rect 393556 13376 393562 13388
rect 517146 13376 517152 13388
rect 393556 13348 517152 13376
rect 393556 13336 393562 13348
rect 517146 13336 517152 13348
rect 517204 13336 517210 13388
rect 93946 13268 93952 13320
rect 94004 13308 94010 13320
rect 263778 13308 263784 13320
rect 94004 13280 263784 13308
rect 94004 13268 94010 13280
rect 263778 13268 263784 13280
rect 263836 13268 263842 13320
rect 394786 13268 394792 13320
rect 394844 13308 394850 13320
rect 520274 13308 520280 13320
rect 394844 13280 520280 13308
rect 394844 13268 394850 13280
rect 520274 13268 520280 13280
rect 520332 13268 520338 13320
rect 52546 13200 52552 13252
rect 52604 13240 52610 13252
rect 249886 13240 249892 13252
rect 52604 13212 249892 13240
rect 52604 13200 52610 13212
rect 249886 13200 249892 13212
rect 249944 13200 249950 13252
rect 396166 13200 396172 13252
rect 396224 13240 396230 13252
rect 523770 13240 523776 13252
rect 396224 13212 523776 13240
rect 396224 13200 396230 13212
rect 523770 13200 523776 13212
rect 523828 13200 523834 13252
rect 48498 13132 48504 13184
rect 48556 13172 48562 13184
rect 249978 13172 249984 13184
rect 48556 13144 249984 13172
rect 48556 13132 48562 13144
rect 249978 13132 249984 13144
rect 250036 13132 250042 13184
rect 397638 13132 397644 13184
rect 397696 13172 397702 13184
rect 527818 13172 527824 13184
rect 397696 13144 527824 13172
rect 397696 13132 397702 13144
rect 527818 13132 527824 13144
rect 527876 13132 527882 13184
rect 44266 13064 44272 13116
rect 44324 13104 44330 13116
rect 248506 13104 248512 13116
rect 44324 13076 248512 13104
rect 44324 13064 44330 13076
rect 248506 13064 248512 13076
rect 248564 13064 248570 13116
rect 405918 13064 405924 13116
rect 405976 13104 405982 13116
rect 554774 13104 554780 13116
rect 405976 13076 554780 13104
rect 405976 13064 405982 13076
rect 554774 13064 554780 13076
rect 554832 13064 554838 13116
rect 122282 12996 122288 13048
rect 122340 13036 122346 13048
rect 272150 13036 272156 13048
rect 122340 13008 272156 13036
rect 122340 12996 122346 13008
rect 272150 12996 272156 13008
rect 272208 12996 272214 13048
rect 365990 12996 365996 13048
rect 366048 13036 366054 13048
rect 423674 13036 423680 13048
rect 366048 13008 423680 13036
rect 366048 12996 366054 13008
rect 423674 12996 423680 13008
rect 423732 12996 423738 13048
rect 156138 12928 156144 12980
rect 156196 12968 156202 12980
rect 283190 12968 283196 12980
rect 156196 12940 283196 12968
rect 156196 12928 156202 12940
rect 283190 12928 283196 12940
rect 283248 12928 283254 12980
rect 364518 12928 364524 12980
rect 364576 12968 364582 12980
rect 420914 12968 420920 12980
rect 364576 12940 420920 12968
rect 364576 12928 364582 12940
rect 420914 12928 420920 12940
rect 420972 12928 420978 12980
rect 160094 12860 160100 12912
rect 160152 12900 160158 12912
rect 284570 12900 284576 12912
rect 160152 12872 284576 12900
rect 160152 12860 160158 12872
rect 284570 12860 284576 12872
rect 284628 12860 284634 12912
rect 363046 12860 363052 12912
rect 363104 12900 363110 12912
rect 417418 12900 417424 12912
rect 363104 12872 417424 12900
rect 363104 12860 363110 12872
rect 417418 12860 417424 12872
rect 417476 12860 417482 12912
rect 223574 12384 223580 12436
rect 223632 12424 223638 12436
rect 303798 12424 303804 12436
rect 223632 12396 303804 12424
rect 223632 12384 223638 12396
rect 303798 12384 303804 12396
rect 303856 12384 303862 12436
rect 385310 12384 385316 12436
rect 385368 12424 385374 12436
rect 487154 12424 487160 12436
rect 385368 12396 487160 12424
rect 385368 12384 385374 12396
rect 487154 12384 487160 12396
rect 487212 12384 487218 12436
rect 219986 12316 219992 12368
rect 220044 12356 220050 12368
rect 302326 12356 302332 12368
rect 220044 12328 302332 12356
rect 220044 12316 220050 12328
rect 302326 12316 302332 12328
rect 302384 12316 302390 12368
rect 386598 12316 386604 12368
rect 386656 12356 386662 12368
rect 489914 12356 489920 12368
rect 386656 12328 489920 12356
rect 386656 12316 386662 12328
rect 489914 12316 489920 12328
rect 489972 12316 489978 12368
rect 216858 12248 216864 12300
rect 216916 12288 216922 12300
rect 300946 12288 300952 12300
rect 216916 12260 300952 12288
rect 216916 12248 216922 12260
rect 300946 12248 300952 12260
rect 301004 12248 301010 12300
rect 385126 12248 385132 12300
rect 385184 12288 385190 12300
rect 490006 12288 490012 12300
rect 385184 12260 490012 12288
rect 385184 12248 385190 12260
rect 490006 12248 490012 12260
rect 490064 12248 490070 12300
rect 213362 12180 213368 12232
rect 213420 12220 213426 12232
rect 299566 12220 299572 12232
rect 213420 12192 299572 12220
rect 213420 12180 213426 12192
rect 299566 12180 299572 12192
rect 299624 12180 299630 12232
rect 386690 12180 386696 12232
rect 386748 12220 386754 12232
rect 493042 12220 493048 12232
rect 386748 12192 493048 12220
rect 386748 12180 386754 12192
rect 493042 12180 493048 12192
rect 493100 12180 493106 12232
rect 209774 12112 209780 12164
rect 209832 12152 209838 12164
rect 299658 12152 299664 12164
rect 209832 12124 299664 12152
rect 209832 12112 209838 12124
rect 299658 12112 299664 12124
rect 299716 12112 299722 12164
rect 386506 12112 386512 12164
rect 386564 12152 386570 12164
rect 494698 12152 494704 12164
rect 386564 12124 494704 12152
rect 386564 12112 386570 12124
rect 494698 12112 494704 12124
rect 494756 12112 494762 12164
rect 206186 12044 206192 12096
rect 206244 12084 206250 12096
rect 298186 12084 298192 12096
rect 206244 12056 298192 12084
rect 206244 12044 206250 12056
rect 298186 12044 298192 12056
rect 298244 12044 298250 12096
rect 387978 12044 387984 12096
rect 388036 12084 388042 12096
rect 497090 12084 497096 12096
rect 388036 12056 497096 12084
rect 388036 12044 388042 12056
rect 497090 12044 497096 12056
rect 497148 12044 497154 12096
rect 138842 11976 138848 12028
rect 138900 12016 138906 12028
rect 277670 12016 277676 12028
rect 138900 11988 277676 12016
rect 138900 11976 138906 11988
rect 277670 11976 277676 11988
rect 277728 11976 277734 12028
rect 389450 11976 389456 12028
rect 389508 12016 389514 12028
rect 500586 12016 500592 12028
rect 389508 11988 500592 12016
rect 389508 11976 389514 11988
rect 500586 11976 500592 11988
rect 500644 11976 500650 12028
rect 135254 11908 135260 11960
rect 135312 11948 135318 11960
rect 276290 11948 276296 11960
rect 135312 11920 276296 11948
rect 135312 11908 135318 11920
rect 276290 11908 276296 11920
rect 276348 11908 276354 11960
rect 390738 11908 390744 11960
rect 390796 11948 390802 11960
rect 503714 11948 503720 11960
rect 390796 11920 503720 11948
rect 390796 11908 390802 11920
rect 503714 11908 503720 11920
rect 503772 11908 503778 11960
rect 36722 11840 36728 11892
rect 36780 11880 36786 11892
rect 245746 11880 245752 11892
rect 36780 11852 245752 11880
rect 36780 11840 36786 11852
rect 245746 11840 245752 11852
rect 245804 11840 245810 11892
rect 392210 11840 392216 11892
rect 392268 11880 392274 11892
rect 511258 11880 511264 11892
rect 392268 11852 511264 11880
rect 392268 11840 392274 11852
rect 511258 11840 511264 11852
rect 511316 11840 511322 11892
rect 17954 11772 17960 11824
rect 18012 11812 18018 11824
rect 240410 11812 240416 11824
rect 18012 11784 240416 11812
rect 18012 11772 18018 11784
rect 240410 11772 240416 11784
rect 240468 11772 240474 11824
rect 403158 11772 403164 11824
rect 403216 11812 403222 11824
rect 547874 11812 547880 11824
rect 403216 11784 547880 11812
rect 403216 11772 403222 11784
rect 547874 11772 547880 11784
rect 547932 11772 547938 11824
rect 13538 11704 13544 11756
rect 13596 11744 13602 11756
rect 238846 11744 238852 11756
rect 13596 11716 238852 11744
rect 13596 11704 13602 11716
rect 238846 11704 238852 11716
rect 238904 11704 238910 11756
rect 276014 11704 276020 11756
rect 276072 11744 276078 11756
rect 276750 11744 276756 11756
rect 276072 11716 276756 11744
rect 276072 11704 276078 11716
rect 276750 11704 276756 11716
rect 276808 11704 276814 11756
rect 404630 11704 404636 11756
rect 404688 11744 404694 11756
rect 551002 11744 551008 11756
rect 404688 11716 551008 11744
rect 404688 11704 404694 11716
rect 551002 11704 551008 11716
rect 551060 11704 551066 11756
rect 201494 11636 201500 11688
rect 201552 11676 201558 11688
rect 202690 11676 202696 11688
rect 201552 11648 202696 11676
rect 201552 11636 201558 11648
rect 202690 11636 202696 11648
rect 202748 11636 202754 11688
rect 226334 11636 226340 11688
rect 226392 11676 226398 11688
rect 305270 11676 305276 11688
rect 226392 11648 305276 11676
rect 226392 11636 226398 11648
rect 305270 11636 305276 11648
rect 305328 11636 305334 11688
rect 385218 11636 385224 11688
rect 385276 11676 385282 11688
rect 486418 11676 486424 11688
rect 385276 11648 486424 11676
rect 385276 11636 385282 11648
rect 486418 11636 486424 11648
rect 486476 11636 486482 11688
rect 231026 11568 231032 11620
rect 231084 11608 231090 11620
rect 305178 11608 305184 11620
rect 231084 11580 305184 11608
rect 231084 11568 231090 11580
rect 305178 11568 305184 11580
rect 305236 11568 305242 11620
rect 383930 11568 383936 11620
rect 383988 11608 383994 11620
rect 484026 11608 484032 11620
rect 383988 11580 484032 11608
rect 383988 11568 383994 11580
rect 484026 11568 484032 11580
rect 484084 11568 484090 11620
rect 234614 11500 234620 11552
rect 234672 11540 234678 11552
rect 306558 11540 306564 11552
rect 234672 11512 306564 11540
rect 234672 11500 234678 11512
rect 306558 11500 306564 11512
rect 306616 11500 306622 11552
rect 382458 11500 382464 11552
rect 382516 11540 382522 11552
rect 480530 11540 480536 11552
rect 382516 11512 480536 11540
rect 382516 11500 382522 11512
rect 480530 11500 480536 11512
rect 480588 11500 480594 11552
rect 176654 10956 176660 11008
rect 176712 10996 176718 11008
rect 290090 10996 290096 11008
rect 176712 10968 290096 10996
rect 176712 10956 176718 10968
rect 290090 10956 290096 10968
rect 290148 10956 290154 11008
rect 372706 10956 372712 11008
rect 372764 10996 372770 11008
rect 445754 10996 445760 11008
rect 372764 10968 445760 10996
rect 372764 10956 372770 10968
rect 445754 10956 445760 10968
rect 445812 10956 445818 11008
rect 173894 10888 173900 10940
rect 173952 10928 173958 10940
rect 288526 10928 288532 10940
rect 173952 10900 288532 10928
rect 173952 10888 173958 10900
rect 288526 10888 288532 10900
rect 288584 10888 288590 10940
rect 372614 10888 372620 10940
rect 372672 10928 372678 10940
rect 448606 10928 448612 10940
rect 372672 10900 448612 10928
rect 372672 10888 372678 10900
rect 448606 10888 448612 10900
rect 448664 10888 448670 10940
rect 170306 10820 170312 10872
rect 170364 10860 170370 10872
rect 287238 10860 287244 10872
rect 170364 10832 287244 10860
rect 170364 10820 170370 10832
rect 287238 10820 287244 10832
rect 287296 10820 287302 10872
rect 373994 10820 374000 10872
rect 374052 10860 374058 10872
rect 453298 10860 453304 10872
rect 374052 10832 453304 10860
rect 374052 10820 374058 10832
rect 453298 10820 453304 10832
rect 453356 10820 453362 10872
rect 167178 10752 167184 10804
rect 167236 10792 167242 10804
rect 285766 10792 285772 10804
rect 167236 10764 285772 10792
rect 167236 10752 167242 10764
rect 285766 10752 285772 10764
rect 285824 10752 285830 10804
rect 375374 10752 375380 10804
rect 375432 10792 375438 10804
rect 456886 10792 456892 10804
rect 375432 10764 456892 10792
rect 375432 10752 375438 10764
rect 456886 10752 456892 10764
rect 456944 10752 456950 10804
rect 163406 10684 163412 10736
rect 163464 10724 163470 10736
rect 284478 10724 284484 10736
rect 163464 10696 284484 10724
rect 163464 10684 163470 10696
rect 284478 10684 284484 10696
rect 284536 10684 284542 10736
rect 376754 10684 376760 10736
rect 376812 10724 376818 10736
rect 459922 10724 459928 10736
rect 376812 10696 459928 10724
rect 376812 10684 376818 10696
rect 459922 10684 459928 10696
rect 459980 10684 459986 10736
rect 158898 10616 158904 10668
rect 158956 10656 158962 10668
rect 283098 10656 283104 10668
rect 158956 10628 283104 10656
rect 158956 10616 158962 10628
rect 283098 10616 283104 10628
rect 283156 10616 283162 10668
rect 378226 10616 378232 10668
rect 378284 10656 378290 10668
rect 463970 10656 463976 10668
rect 378284 10628 463976 10656
rect 378284 10616 378290 10628
rect 463970 10616 463976 10628
rect 464028 10616 464034 10668
rect 155402 10548 155408 10600
rect 155460 10588 155466 10600
rect 283006 10588 283012 10600
rect 155460 10560 283012 10588
rect 155460 10548 155466 10560
rect 283006 10548 283012 10560
rect 283064 10548 283070 10600
rect 378318 10548 378324 10600
rect 378376 10588 378382 10600
rect 467466 10588 467472 10600
rect 378376 10560 467472 10588
rect 378376 10548 378382 10560
rect 467466 10548 467472 10560
rect 467524 10548 467530 10600
rect 126974 10480 126980 10532
rect 127032 10520 127038 10532
rect 273438 10520 273444 10532
rect 127032 10492 273444 10520
rect 127032 10480 127038 10492
rect 273438 10480 273444 10492
rect 273496 10480 273502 10532
rect 379698 10480 379704 10532
rect 379756 10520 379762 10532
rect 470594 10520 470600 10532
rect 379756 10492 470600 10520
rect 379756 10480 379762 10492
rect 470594 10480 470600 10492
rect 470652 10480 470658 10532
rect 89898 10412 89904 10464
rect 89956 10452 89962 10464
rect 262306 10452 262312 10464
rect 89956 10424 262312 10452
rect 89956 10412 89962 10424
rect 262306 10412 262312 10424
rect 262364 10412 262370 10464
rect 381078 10412 381084 10464
rect 381136 10452 381142 10464
rect 474090 10452 474096 10464
rect 381136 10424 474096 10452
rect 381136 10412 381142 10424
rect 474090 10412 474096 10424
rect 474148 10412 474154 10464
rect 86402 10344 86408 10396
rect 86460 10384 86466 10396
rect 261110 10384 261116 10396
rect 86460 10356 261116 10384
rect 86460 10344 86466 10356
rect 261110 10344 261116 10356
rect 261168 10344 261174 10396
rect 382366 10344 382372 10396
rect 382424 10384 382430 10396
rect 478138 10384 478144 10396
rect 382424 10356 478144 10384
rect 382424 10344 382430 10356
rect 478138 10344 478144 10356
rect 478196 10344 478202 10396
rect 83274 10276 83280 10328
rect 83332 10316 83338 10328
rect 259638 10316 259644 10328
rect 83332 10288 259644 10316
rect 83332 10276 83338 10288
rect 259638 10276 259644 10288
rect 259696 10276 259702 10328
rect 383838 10276 383844 10328
rect 383896 10316 383902 10328
rect 482370 10316 482376 10328
rect 383896 10288 482376 10316
rect 383896 10276 383902 10288
rect 482370 10276 482376 10288
rect 482428 10276 482434 10328
rect 180978 10208 180984 10260
rect 181036 10248 181042 10260
rect 289998 10248 290004 10260
rect 181036 10220 290004 10248
rect 181036 10208 181042 10220
rect 289998 10208 290004 10220
rect 290056 10208 290062 10260
rect 371418 10208 371424 10260
rect 371476 10248 371482 10260
rect 442166 10248 442172 10260
rect 371476 10220 442172 10248
rect 371476 10208 371482 10220
rect 442166 10208 442172 10220
rect 442224 10208 442230 10260
rect 184934 10140 184940 10192
rect 184992 10180 184998 10192
rect 291470 10180 291476 10192
rect 184992 10152 291476 10180
rect 184992 10140 184998 10152
rect 291470 10140 291476 10152
rect 291528 10140 291534 10192
rect 369946 10140 369952 10192
rect 370004 10180 370010 10192
rect 439130 10180 439136 10192
rect 370004 10152 439136 10180
rect 370004 10140 370010 10152
rect 439130 10140 439136 10152
rect 439188 10140 439194 10192
rect 188246 10072 188252 10124
rect 188304 10112 188310 10124
rect 292850 10112 292856 10124
rect 188304 10084 292856 10112
rect 188304 10072 188310 10084
rect 292850 10072 292856 10084
rect 292908 10072 292914 10124
rect 368566 10072 368572 10124
rect 368624 10112 368630 10124
rect 435082 10112 435088 10124
rect 368624 10084 435088 10112
rect 368624 10072 368630 10084
rect 435082 10072 435088 10084
rect 435140 10072 435146 10124
rect 151722 9596 151728 9648
rect 151780 9636 151786 9648
rect 153010 9636 153016 9648
rect 151780 9608 153016 9636
rect 151780 9596 151786 9608
rect 153010 9596 153016 9608
rect 153068 9596 153074 9648
rect 222746 9596 222752 9648
rect 222804 9636 222810 9648
rect 303614 9636 303620 9648
rect 222804 9608 303620 9636
rect 222804 9596 222810 9608
rect 303614 9596 303620 9608
rect 303672 9596 303678 9648
rect 400306 9596 400312 9648
rect 400364 9636 400370 9648
rect 538398 9636 538404 9648
rect 400364 9608 538404 9636
rect 400364 9596 400370 9608
rect 538398 9596 538404 9608
rect 538456 9596 538462 9648
rect 219250 9528 219256 9580
rect 219308 9568 219314 9580
rect 302234 9568 302240 9580
rect 219308 9540 302240 9568
rect 219308 9528 219314 9540
rect 302234 9528 302240 9540
rect 302292 9528 302298 9580
rect 401686 9528 401692 9580
rect 401744 9568 401750 9580
rect 541986 9568 541992 9580
rect 401744 9540 541992 9568
rect 401744 9528 401750 9540
rect 541986 9528 541992 9540
rect 542044 9528 542050 9580
rect 141234 9460 141240 9512
rect 141292 9500 141298 9512
rect 277578 9500 277584 9512
rect 141292 9472 277584 9500
rect 141292 9460 141298 9472
rect 277578 9460 277584 9472
rect 277636 9460 277642 9512
rect 403066 9460 403072 9512
rect 403124 9500 403130 9512
rect 545482 9500 545488 9512
rect 403124 9472 545488 9500
rect 403124 9460 403130 9472
rect 545482 9460 545488 9472
rect 545540 9460 545546 9512
rect 137646 9392 137652 9444
rect 137704 9432 137710 9444
rect 277486 9432 277492 9444
rect 137704 9404 277492 9432
rect 137704 9392 137710 9404
rect 277486 9392 277492 9404
rect 277544 9392 277550 9444
rect 404446 9392 404452 9444
rect 404504 9432 404510 9444
rect 549070 9432 549076 9444
rect 404504 9404 549076 9432
rect 404504 9392 404510 9404
rect 549070 9392 549076 9404
rect 549128 9392 549134 9444
rect 76190 9324 76196 9376
rect 76248 9364 76254 9376
rect 258350 9364 258356 9376
rect 76248 9336 258356 9364
rect 76248 9324 76254 9336
rect 258350 9324 258356 9336
rect 258408 9324 258414 9376
rect 404538 9324 404544 9376
rect 404596 9364 404602 9376
rect 552658 9364 552664 9376
rect 404596 9336 552664 9364
rect 404596 9324 404602 9336
rect 552658 9324 552664 9336
rect 552716 9324 552722 9376
rect 72602 9256 72608 9308
rect 72660 9296 72666 9308
rect 256694 9296 256700 9308
rect 72660 9268 256700 9296
rect 72660 9256 72666 9268
rect 256694 9256 256700 9268
rect 256752 9256 256758 9308
rect 405826 9256 405832 9308
rect 405884 9296 405890 9308
rect 556154 9296 556160 9308
rect 405884 9268 556160 9296
rect 405884 9256 405890 9268
rect 556154 9256 556160 9268
rect 556212 9256 556218 9308
rect 33594 9188 33600 9240
rect 33652 9228 33658 9240
rect 244458 9228 244464 9240
rect 33652 9200 244464 9228
rect 33652 9188 33658 9200
rect 244458 9188 244464 9200
rect 244516 9188 244522 9240
rect 407206 9188 407212 9240
rect 407264 9228 407270 9240
rect 559742 9228 559748 9240
rect 407264 9200 559748 9228
rect 407264 9188 407270 9200
rect 559742 9188 559748 9200
rect 559800 9188 559806 9240
rect 30098 9120 30104 9172
rect 30156 9160 30162 9172
rect 243078 9160 243084 9172
rect 30156 9132 243084 9160
rect 30156 9120 30162 9132
rect 243078 9120 243084 9132
rect 243136 9120 243142 9172
rect 408678 9120 408684 9172
rect 408736 9160 408742 9172
rect 563238 9160 563244 9172
rect 408736 9132 563244 9160
rect 408736 9120 408742 9132
rect 563238 9120 563244 9132
rect 563296 9120 563302 9172
rect 26510 9052 26516 9104
rect 26568 9092 26574 9104
rect 242986 9092 242992 9104
rect 26568 9064 242992 9092
rect 26568 9052 26574 9064
rect 242986 9052 242992 9064
rect 243044 9052 243050 9104
rect 410058 9052 410064 9104
rect 410116 9092 410122 9104
rect 566826 9092 566832 9104
rect 410116 9064 566832 9092
rect 410116 9052 410122 9064
rect 566826 9052 566832 9064
rect 566884 9052 566890 9104
rect 21818 8984 21824 9036
rect 21876 9024 21882 9036
rect 241606 9024 241612 9036
rect 21876 8996 241612 9024
rect 21876 8984 21882 8996
rect 241606 8984 241612 8996
rect 241664 8984 241670 9036
rect 409966 8984 409972 9036
rect 410024 9024 410030 9036
rect 570322 9024 570328 9036
rect 410024 8996 570328 9024
rect 410024 8984 410030 8996
rect 570322 8984 570328 8996
rect 570380 8984 570386 9036
rect 4062 8916 4068 8968
rect 4120 8956 4126 8968
rect 236178 8956 236184 8968
rect 4120 8928 236184 8956
rect 4120 8916 4126 8928
rect 236178 8916 236184 8928
rect 236236 8916 236242 8968
rect 238110 8916 238116 8968
rect 238168 8956 238174 8968
rect 307938 8956 307944 8968
rect 238168 8928 307944 8956
rect 238168 8916 238174 8928
rect 307938 8916 307944 8928
rect 307996 8916 308002 8968
rect 411438 8916 411444 8968
rect 411496 8956 411502 8968
rect 573910 8956 573916 8968
rect 411496 8928 573916 8956
rect 411496 8916 411502 8928
rect 573910 8916 573916 8928
rect 573968 8916 573974 8968
rect 226426 8848 226432 8900
rect 226484 8888 226490 8900
rect 303706 8888 303712 8900
rect 226484 8860 303712 8888
rect 226484 8848 226490 8860
rect 303706 8848 303712 8860
rect 303764 8848 303770 8900
rect 399018 8848 399024 8900
rect 399076 8888 399082 8900
rect 534902 8888 534908 8900
rect 399076 8860 534908 8888
rect 399076 8848 399082 8860
rect 534902 8848 534908 8860
rect 534960 8848 534966 8900
rect 229830 8780 229836 8832
rect 229888 8820 229894 8832
rect 305086 8820 305092 8832
rect 229888 8792 305092 8820
rect 229888 8780 229894 8792
rect 305086 8780 305092 8792
rect 305144 8780 305150 8832
rect 398926 8780 398932 8832
rect 398984 8820 398990 8832
rect 531314 8820 531320 8832
rect 398984 8792 531320 8820
rect 398984 8780 398990 8792
rect 531314 8780 531320 8792
rect 531372 8780 531378 8832
rect 233418 8712 233424 8764
rect 233476 8752 233482 8764
rect 306466 8752 306472 8764
rect 233476 8724 306472 8752
rect 233476 8712 233482 8724
rect 306466 8712 306472 8724
rect 306524 8712 306530 8764
rect 361850 8712 361856 8764
rect 361908 8752 361914 8764
rect 414290 8752 414296 8764
rect 361908 8724 414296 8752
rect 361908 8712 361914 8724
rect 414290 8712 414296 8724
rect 414348 8712 414354 8764
rect 187326 8236 187332 8288
rect 187384 8276 187390 8288
rect 292758 8276 292764 8288
rect 187384 8248 292764 8276
rect 187384 8236 187390 8248
rect 292758 8236 292764 8248
rect 292816 8236 292822 8288
rect 380986 8236 380992 8288
rect 381044 8276 381050 8288
rect 476942 8276 476948 8288
rect 381044 8248 476948 8276
rect 381044 8236 381050 8248
rect 476942 8236 476948 8248
rect 477000 8236 477006 8288
rect 183738 8168 183744 8220
rect 183796 8208 183802 8220
rect 291378 8208 291384 8220
rect 183796 8180 291384 8208
rect 183796 8168 183802 8180
rect 291378 8168 291384 8180
rect 291436 8168 291442 8220
rect 383654 8168 383660 8220
rect 383712 8208 383718 8220
rect 481726 8208 481732 8220
rect 383712 8180 481732 8208
rect 383712 8168 383718 8180
rect 481726 8168 481732 8180
rect 481784 8168 481790 8220
rect 180242 8100 180248 8152
rect 180300 8140 180306 8152
rect 289906 8140 289912 8152
rect 180300 8112 289912 8140
rect 180300 8100 180306 8112
rect 289906 8100 289912 8112
rect 289964 8100 289970 8152
rect 383746 8100 383752 8152
rect 383804 8140 383810 8152
rect 485222 8140 485228 8152
rect 383804 8112 485228 8140
rect 383804 8100 383810 8112
rect 485222 8100 485228 8112
rect 485280 8100 485286 8152
rect 176746 8032 176752 8084
rect 176804 8072 176810 8084
rect 288618 8072 288624 8084
rect 176804 8044 288624 8072
rect 176804 8032 176810 8044
rect 288618 8032 288624 8044
rect 288676 8032 288682 8084
rect 385034 8032 385040 8084
rect 385092 8072 385098 8084
rect 488810 8072 488816 8084
rect 385092 8044 488816 8072
rect 385092 8032 385098 8044
rect 488810 8032 488816 8044
rect 488868 8032 488874 8084
rect 173066 7964 173072 8016
rect 173124 8004 173130 8016
rect 287054 8004 287060 8016
rect 173124 7976 287060 8004
rect 173124 7964 173130 7976
rect 287054 7964 287060 7976
rect 287112 7964 287118 8016
rect 386414 7964 386420 8016
rect 386472 8004 386478 8016
rect 492306 8004 492312 8016
rect 386472 7976 492312 8004
rect 386472 7964 386478 7976
rect 492306 7964 492312 7976
rect 492364 7964 492370 8016
rect 169570 7896 169576 7948
rect 169628 7936 169634 7948
rect 287146 7936 287152 7948
rect 169628 7908 287152 7936
rect 169628 7896 169634 7908
rect 287146 7896 287152 7908
rect 287204 7896 287210 7948
rect 387886 7896 387892 7948
rect 387944 7936 387950 7948
rect 495894 7936 495900 7948
rect 387944 7908 495900 7936
rect 387944 7896 387950 7908
rect 495894 7896 495900 7908
rect 495952 7896 495958 7948
rect 166074 7828 166080 7880
rect 166132 7868 166138 7880
rect 285674 7868 285680 7880
rect 166132 7840 285680 7868
rect 166132 7828 166138 7840
rect 285674 7828 285680 7840
rect 285732 7828 285738 7880
rect 389358 7828 389364 7880
rect 389416 7868 389422 7880
rect 499390 7868 499396 7880
rect 389416 7840 499396 7868
rect 389416 7828 389422 7840
rect 499390 7828 499396 7840
rect 499448 7828 499454 7880
rect 157794 7760 157800 7812
rect 157852 7800 157858 7812
rect 282914 7800 282920 7812
rect 157852 7772 282920 7800
rect 157852 7760 157858 7772
rect 282914 7760 282920 7772
rect 282972 7760 282978 7812
rect 283650 7760 283656 7812
rect 283708 7800 283714 7812
rect 316310 7800 316316 7812
rect 283708 7772 316316 7800
rect 283708 7760 283714 7772
rect 316310 7760 316316 7772
rect 316368 7760 316374 7812
rect 389266 7760 389272 7812
rect 389324 7800 389330 7812
rect 502978 7800 502984 7812
rect 389324 7772 502984 7800
rect 389324 7760 389330 7772
rect 502978 7760 502984 7772
rect 503036 7760 503042 7812
rect 134150 7692 134156 7744
rect 134208 7732 134214 7744
rect 276198 7732 276204 7744
rect 134208 7704 276204 7732
rect 134208 7692 134214 7704
rect 276198 7692 276204 7704
rect 276256 7692 276262 7744
rect 277486 7692 277492 7744
rect 277544 7732 277550 7744
rect 313458 7732 313464 7744
rect 277544 7704 313464 7732
rect 277544 7692 277550 7704
rect 313458 7692 313464 7704
rect 313516 7692 313522 7744
rect 390646 7692 390652 7744
rect 390704 7732 390710 7744
rect 506474 7732 506480 7744
rect 390704 7704 506480 7732
rect 390704 7692 390710 7704
rect 506474 7692 506480 7704
rect 506532 7692 506538 7744
rect 130562 7624 130568 7676
rect 130620 7664 130626 7676
rect 274818 7664 274824 7676
rect 130620 7636 274824 7664
rect 130620 7624 130626 7636
rect 274818 7624 274824 7636
rect 274876 7624 274882 7676
rect 275186 7624 275192 7676
rect 275244 7664 275250 7676
rect 311986 7664 311992 7676
rect 275244 7636 311992 7664
rect 275244 7624 275250 7636
rect 311986 7624 311992 7636
rect 312044 7624 312050 7676
rect 392118 7624 392124 7676
rect 392176 7664 392182 7676
rect 510062 7664 510068 7676
rect 392176 7636 510068 7664
rect 392176 7624 392182 7636
rect 510062 7624 510068 7636
rect 510120 7624 510126 7676
rect 127066 7556 127072 7608
rect 127124 7596 127130 7608
rect 273346 7596 273352 7608
rect 127124 7568 273352 7596
rect 127124 7556 127130 7568
rect 273346 7556 273352 7568
rect 273404 7556 273410 7608
rect 274542 7556 274548 7608
rect 274600 7596 274606 7608
rect 310698 7596 310704 7608
rect 274600 7568 310704 7596
rect 274600 7556 274606 7568
rect 310698 7556 310704 7568
rect 310756 7556 310762 7608
rect 393406 7556 393412 7608
rect 393464 7596 393470 7608
rect 513558 7596 513564 7608
rect 393464 7568 513564 7596
rect 393464 7556 393470 7568
rect 513558 7556 513564 7568
rect 513616 7556 513622 7608
rect 190822 7488 190828 7540
rect 190880 7528 190886 7540
rect 292666 7528 292672 7540
rect 190880 7500 292672 7528
rect 190880 7488 190886 7500
rect 292666 7488 292672 7500
rect 292724 7488 292730 7540
rect 380894 7488 380900 7540
rect 380952 7528 380958 7540
rect 473446 7528 473452 7540
rect 380952 7500 473452 7528
rect 380952 7488 380958 7500
rect 473446 7488 473452 7500
rect 473504 7488 473510 7540
rect 194410 7420 194416 7472
rect 194468 7460 194474 7472
rect 294046 7460 294052 7472
rect 194468 7432 294052 7460
rect 194468 7420 194474 7432
rect 294046 7420 294052 7432
rect 294104 7420 294110 7472
rect 379606 7420 379612 7472
rect 379664 7460 379670 7472
rect 469858 7460 469864 7472
rect 379664 7432 469864 7460
rect 379664 7420 379670 7432
rect 469858 7420 469864 7432
rect 469916 7420 469922 7472
rect 197906 7352 197912 7404
rect 197964 7392 197970 7404
rect 295426 7392 295432 7404
rect 197964 7364 295432 7392
rect 197964 7352 197970 7364
rect 295426 7352 295432 7364
rect 295484 7352 295490 7404
rect 378134 7352 378140 7404
rect 378192 7392 378198 7404
rect 466270 7392 466276 7404
rect 378192 7364 466276 7392
rect 378192 7352 378198 7364
rect 466270 7352 466276 7364
rect 466328 7352 466334 7404
rect 69106 6808 69112 6860
rect 69164 6848 69170 6860
rect 255314 6848 255320 6860
rect 69164 6820 255320 6848
rect 69164 6808 69170 6820
rect 255314 6808 255320 6820
rect 255372 6808 255378 6860
rect 279510 6808 279516 6860
rect 279568 6848 279574 6860
rect 320266 6848 320272 6860
rect 279568 6820 320272 6848
rect 279568 6808 279574 6820
rect 320266 6808 320272 6820
rect 320324 6808 320330 6860
rect 365714 6808 365720 6860
rect 365772 6848 365778 6860
rect 427262 6848 427268 6860
rect 365772 6820 427268 6848
rect 365772 6808 365778 6820
rect 427262 6808 427268 6820
rect 427320 6808 427326 6860
rect 65518 6740 65524 6792
rect 65576 6780 65582 6792
rect 254026 6780 254032 6792
rect 65576 6752 254032 6780
rect 65576 6740 65582 6752
rect 254026 6740 254032 6752
rect 254084 6740 254090 6792
rect 276014 6740 276020 6792
rect 276072 6780 276078 6792
rect 318886 6780 318892 6792
rect 276072 6752 318892 6780
rect 276072 6740 276078 6752
rect 318886 6740 318892 6752
rect 318944 6740 318950 6792
rect 367094 6740 367100 6792
rect 367152 6780 367158 6792
rect 430850 6780 430856 6792
rect 367152 6752 430856 6780
rect 367152 6740 367158 6752
rect 430850 6740 430856 6752
rect 430908 6740 430914 6792
rect 62022 6672 62028 6724
rect 62080 6712 62086 6724
rect 253934 6712 253940 6724
rect 62080 6684 253940 6712
rect 62080 6672 62086 6684
rect 253934 6672 253940 6684
rect 253992 6672 253998 6724
rect 272426 6672 272432 6724
rect 272484 6712 272490 6724
rect 318978 6712 318984 6724
rect 272484 6684 318984 6712
rect 272484 6672 272490 6684
rect 318978 6672 318984 6684
rect 319036 6672 319042 6724
rect 368474 6672 368480 6724
rect 368532 6712 368538 6724
rect 434438 6712 434444 6724
rect 368532 6684 434444 6712
rect 368532 6672 368538 6684
rect 434438 6672 434444 6684
rect 434496 6672 434502 6724
rect 58434 6604 58440 6656
rect 58492 6644 58498 6656
rect 252554 6644 252560 6656
rect 58492 6616 252560 6644
rect 58492 6604 58498 6616
rect 252554 6604 252560 6616
rect 252612 6604 252618 6656
rect 268838 6604 268844 6656
rect 268896 6644 268902 6656
rect 317690 6644 317696 6656
rect 268896 6616 317696 6644
rect 268896 6604 268902 6616
rect 317690 6604 317696 6616
rect 317748 6604 317754 6656
rect 369854 6604 369860 6656
rect 369912 6644 369918 6656
rect 437934 6644 437940 6656
rect 369912 6616 437940 6644
rect 369912 6604 369918 6616
rect 437934 6604 437940 6616
rect 437992 6604 437998 6656
rect 54938 6536 54944 6588
rect 54996 6576 55002 6588
rect 251174 6576 251180 6588
rect 54996 6548 251180 6576
rect 54996 6536 55002 6548
rect 251174 6536 251180 6548
rect 251232 6536 251238 6588
rect 265342 6536 265348 6588
rect 265400 6576 265406 6588
rect 316218 6576 316224 6588
rect 265400 6548 316224 6576
rect 265400 6536 265406 6548
rect 316218 6536 316224 6548
rect 316276 6536 316282 6588
rect 371326 6536 371332 6588
rect 371384 6576 371390 6588
rect 441522 6576 441528 6588
rect 371384 6548 441528 6576
rect 371384 6536 371390 6548
rect 441522 6536 441528 6548
rect 441580 6536 441586 6588
rect 51350 6468 51356 6520
rect 51408 6508 51414 6520
rect 249794 6508 249800 6520
rect 51408 6480 249800 6508
rect 51408 6468 51414 6480
rect 249794 6468 249800 6480
rect 249852 6468 249858 6520
rect 261754 6468 261760 6520
rect 261812 6508 261818 6520
rect 314838 6508 314844 6520
rect 261812 6480 314844 6508
rect 261812 6468 261818 6480
rect 314838 6468 314844 6480
rect 314896 6468 314902 6520
rect 371234 6468 371240 6520
rect 371292 6508 371298 6520
rect 445018 6508 445024 6520
rect 371292 6480 445024 6508
rect 371292 6468 371298 6480
rect 445018 6468 445024 6480
rect 445076 6468 445082 6520
rect 47854 6400 47860 6452
rect 47912 6440 47918 6452
rect 248690 6440 248696 6452
rect 47912 6412 248696 6440
rect 47912 6400 47918 6412
rect 248690 6400 248696 6412
rect 248748 6400 248754 6452
rect 258258 6400 258264 6452
rect 258316 6440 258322 6452
rect 314746 6440 314752 6452
rect 258316 6412 314752 6440
rect 258316 6400 258322 6412
rect 314746 6400 314752 6412
rect 314804 6400 314810 6452
rect 407114 6400 407120 6452
rect 407172 6440 407178 6452
rect 558546 6440 558552 6452
rect 407172 6412 558552 6440
rect 407172 6400 407178 6412
rect 558546 6400 558552 6412
rect 558604 6400 558610 6452
rect 12342 6332 12348 6384
rect 12400 6372 12406 6384
rect 237466 6372 237472 6384
rect 12400 6344 237472 6372
rect 12400 6332 12406 6344
rect 237466 6332 237472 6344
rect 237524 6332 237530 6384
rect 254670 6332 254676 6384
rect 254728 6372 254734 6384
rect 313366 6372 313372 6384
rect 254728 6344 313372 6372
rect 254728 6332 254734 6344
rect 313366 6332 313372 6344
rect 313424 6332 313430 6384
rect 408586 6332 408592 6384
rect 408644 6372 408650 6384
rect 562042 6372 562048 6384
rect 408644 6344 562048 6372
rect 408644 6332 408650 6344
rect 562042 6332 562048 6344
rect 562100 6332 562106 6384
rect 7650 6264 7656 6316
rect 7708 6304 7714 6316
rect 236086 6304 236092 6316
rect 7708 6276 236092 6304
rect 7708 6264 7714 6276
rect 236086 6264 236092 6276
rect 236144 6264 236150 6316
rect 239306 6264 239312 6316
rect 239364 6304 239370 6316
rect 307846 6304 307852 6316
rect 239364 6276 307852 6304
rect 239364 6264 239370 6276
rect 307846 6264 307852 6276
rect 307904 6264 307910 6316
rect 365806 6264 365812 6316
rect 365864 6304 365870 6316
rect 391842 6304 391848 6316
rect 365864 6276 391848 6304
rect 365864 6264 365870 6276
rect 391842 6264 391848 6276
rect 391900 6264 391906 6316
rect 408494 6264 408500 6316
rect 408552 6304 408558 6316
rect 565630 6304 565636 6316
rect 408552 6276 565636 6304
rect 408552 6264 408558 6276
rect 565630 6264 565636 6276
rect 565688 6264 565694 6316
rect 2866 6196 2872 6248
rect 2924 6236 2930 6248
rect 234798 6236 234804 6248
rect 2924 6208 234804 6236
rect 2924 6196 2930 6208
rect 234798 6196 234804 6208
rect 234856 6196 234862 6248
rect 240502 6196 240508 6248
rect 240560 6236 240566 6248
rect 309410 6236 309416 6248
rect 240560 6208 309416 6236
rect 240560 6196 240566 6208
rect 309410 6196 309416 6208
rect 309468 6196 309474 6248
rect 360286 6196 360292 6248
rect 360344 6236 360350 6248
rect 407206 6236 407212 6248
rect 360344 6208 407212 6236
rect 360344 6196 360350 6208
rect 407206 6196 407212 6208
rect 407264 6196 407270 6248
rect 409874 6196 409880 6248
rect 409932 6236 409938 6248
rect 569126 6236 569132 6248
rect 409932 6208 569132 6236
rect 409932 6196 409938 6208
rect 569126 6196 569132 6208
rect 569184 6196 569190 6248
rect 1670 6128 1676 6180
rect 1728 6168 1734 6180
rect 234890 6168 234896 6180
rect 1728 6140 234896 6168
rect 1728 6128 1734 6140
rect 234890 6128 234896 6140
rect 234948 6128 234954 6180
rect 237006 6128 237012 6180
rect 237064 6168 237070 6180
rect 307754 6168 307760 6180
rect 237064 6140 307760 6168
rect 237064 6128 237070 6140
rect 307754 6128 307760 6140
rect 307812 6128 307818 6180
rect 360378 6128 360384 6180
rect 360436 6168 360442 6180
rect 409598 6168 409604 6180
rect 360436 6140 409604 6168
rect 360436 6128 360442 6140
rect 409598 6128 409604 6140
rect 409656 6128 409662 6180
rect 412634 6128 412640 6180
rect 412692 6168 412698 6180
rect 576302 6168 576308 6180
rect 412692 6140 576308 6168
rect 412692 6128 412698 6140
rect 576302 6128 576308 6140
rect 576360 6128 576366 6180
rect 140038 6060 140044 6112
rect 140096 6100 140102 6112
rect 277394 6100 277400 6112
rect 140096 6072 277400 6100
rect 140096 6060 140102 6072
rect 277394 6060 277400 6072
rect 277452 6060 277458 6112
rect 286594 6060 286600 6112
rect 286652 6100 286658 6112
rect 323210 6100 323216 6112
rect 286652 6072 323216 6100
rect 286652 6060 286658 6072
rect 323210 6060 323216 6072
rect 323268 6060 323274 6112
rect 365898 6060 365904 6112
rect 365956 6100 365962 6112
rect 423766 6100 423772 6112
rect 365956 6072 423772 6100
rect 365956 6060 365962 6072
rect 423766 6060 423772 6072
rect 423824 6060 423830 6112
rect 143626 5992 143632 6044
rect 143684 6032 143690 6044
rect 278774 6032 278780 6044
rect 143684 6004 278780 6032
rect 143684 5992 143690 6004
rect 278774 5992 278780 6004
rect 278832 5992 278838 6044
rect 299290 5992 299296 6044
rect 299348 6032 299354 6044
rect 310606 6032 310612 6044
rect 299348 6004 310612 6032
rect 299348 5992 299354 6004
rect 310606 5992 310612 6004
rect 310664 5992 310670 6044
rect 364426 5992 364432 6044
rect 364484 6032 364490 6044
rect 420178 6032 420184 6044
rect 364484 6004 420184 6032
rect 364484 5992 364490 6004
rect 420178 5992 420184 6004
rect 420236 5992 420242 6044
rect 232222 5924 232228 5976
rect 232280 5964 232286 5976
rect 306650 5964 306656 5976
rect 232280 5936 306656 5964
rect 232280 5924 232286 5936
rect 306650 5924 306656 5936
rect 306708 5924 306714 5976
rect 362954 5924 362960 5976
rect 363012 5964 363018 5976
rect 416682 5964 416688 5976
rect 363012 5936 416688 5964
rect 363012 5924 363018 5936
rect 416682 5924 416688 5936
rect 416740 5924 416746 5976
rect 235810 5856 235816 5908
rect 235868 5896 235874 5908
rect 261478 5896 261484 5908
rect 235868 5868 261484 5896
rect 235868 5856 235874 5868
rect 261478 5856 261484 5868
rect 261536 5856 261542 5908
rect 361758 5856 361764 5908
rect 361816 5896 361822 5908
rect 413094 5896 413100 5908
rect 361816 5868 413100 5896
rect 361816 5856 361822 5868
rect 413094 5856 413100 5868
rect 413152 5856 413158 5908
rect 361666 5788 361672 5840
rect 361724 5828 361730 5840
rect 410794 5828 410800 5840
rect 361724 5800 410800 5828
rect 361724 5788 361730 5800
rect 410794 5788 410800 5800
rect 410852 5788 410858 5840
rect 85666 5448 85672 5500
rect 85724 5488 85730 5500
rect 149698 5488 149704 5500
rect 85724 5460 149704 5488
rect 85724 5448 85730 5460
rect 149698 5448 149704 5460
rect 149756 5448 149762 5500
rect 210970 5448 210976 5500
rect 211028 5488 211034 5500
rect 299474 5488 299480 5500
rect 211028 5460 299480 5488
rect 211028 5448 211034 5460
rect 299474 5448 299480 5460
rect 299532 5448 299538 5500
rect 364334 5448 364340 5500
rect 364392 5488 364398 5500
rect 384942 5488 384948 5500
rect 364392 5460 384948 5488
rect 364392 5448 364398 5460
rect 384942 5448 384948 5460
rect 385000 5448 385006 5500
rect 390554 5448 390560 5500
rect 390612 5488 390618 5500
rect 505370 5488 505376 5500
rect 390612 5460 505376 5488
rect 390612 5448 390618 5460
rect 505370 5448 505376 5460
rect 505428 5448 505434 5500
rect 89162 5380 89168 5432
rect 89220 5420 89226 5432
rect 153838 5420 153844 5432
rect 89220 5392 153844 5420
rect 89220 5380 89226 5392
rect 153838 5380 153844 5392
rect 153896 5380 153902 5432
rect 207382 5380 207388 5432
rect 207440 5420 207446 5432
rect 298094 5420 298100 5432
rect 207440 5392 298100 5420
rect 207440 5380 207446 5392
rect 298094 5380 298100 5392
rect 298152 5380 298158 5432
rect 301498 5380 301504 5432
rect 301556 5420 301562 5432
rect 312078 5420 312084 5432
rect 301556 5392 312084 5420
rect 301556 5380 301562 5392
rect 312078 5380 312084 5392
rect 312136 5380 312142 5432
rect 361574 5380 361580 5432
rect 361632 5420 361638 5432
rect 382274 5420 382280 5432
rect 361632 5392 382280 5420
rect 361632 5380 361638 5392
rect 382274 5380 382280 5392
rect 382332 5380 382338 5432
rect 392026 5380 392032 5432
rect 392084 5420 392090 5432
rect 508866 5420 508872 5432
rect 392084 5392 508872 5420
rect 392084 5380 392090 5392
rect 508866 5380 508872 5392
rect 508924 5380 508930 5432
rect 110506 5312 110512 5364
rect 110564 5352 110570 5364
rect 177298 5352 177304 5364
rect 110564 5324 177304 5352
rect 110564 5312 110570 5324
rect 177298 5312 177304 5324
rect 177356 5312 177362 5364
rect 203886 5312 203892 5364
rect 203944 5352 203950 5364
rect 296714 5352 296720 5364
rect 203944 5324 296720 5352
rect 203944 5312 203950 5324
rect 296714 5312 296720 5324
rect 296772 5312 296778 5364
rect 297174 5312 297180 5364
rect 297232 5352 297238 5364
rect 310790 5352 310796 5364
rect 297232 5324 310796 5352
rect 297232 5312 297238 5324
rect 310790 5312 310796 5324
rect 310848 5312 310854 5364
rect 352006 5312 352012 5364
rect 352064 5352 352070 5364
rect 378870 5352 378876 5364
rect 352064 5324 378876 5352
rect 352064 5312 352070 5324
rect 378870 5312 378876 5324
rect 378928 5312 378934 5364
rect 391934 5312 391940 5364
rect 391992 5352 391998 5364
rect 512454 5352 512460 5364
rect 391992 5324 512460 5352
rect 391992 5312 391998 5324
rect 512454 5312 512460 5324
rect 512512 5312 512518 5364
rect 78582 5244 78588 5296
rect 78640 5284 78646 5296
rect 145558 5284 145564 5296
rect 78640 5256 145564 5284
rect 78640 5244 78646 5256
rect 145558 5244 145564 5256
rect 145616 5244 145622 5296
rect 196802 5244 196808 5296
rect 196860 5284 196866 5296
rect 295334 5284 295340 5296
rect 196860 5256 295340 5284
rect 196860 5244 196866 5256
rect 295334 5244 295340 5256
rect 295392 5244 295398 5296
rect 303154 5244 303160 5296
rect 303212 5284 303218 5296
rect 328638 5284 328644 5296
rect 303212 5256 328644 5284
rect 303212 5244 303218 5256
rect 328638 5244 328644 5256
rect 328696 5244 328702 5296
rect 351914 5244 351920 5296
rect 351972 5284 351978 5296
rect 382366 5284 382372 5296
rect 351972 5256 382372 5284
rect 351972 5244 351978 5256
rect 382366 5244 382372 5256
rect 382424 5244 382430 5296
rect 393314 5244 393320 5296
rect 393372 5284 393378 5296
rect 515950 5284 515956 5296
rect 393372 5256 515956 5284
rect 393372 5244 393378 5256
rect 515950 5244 515956 5256
rect 516008 5244 516014 5296
rect 117590 5176 117596 5228
rect 117648 5216 117654 5228
rect 185578 5216 185584 5228
rect 117648 5188 185584 5216
rect 117648 5176 117654 5188
rect 185578 5176 185584 5188
rect 185636 5176 185642 5228
rect 193214 5176 193220 5228
rect 193272 5216 193278 5228
rect 293954 5216 293960 5228
rect 193272 5188 293960 5216
rect 193272 5176 193278 5188
rect 293954 5176 293960 5188
rect 294012 5176 294018 5228
rect 294046 5176 294052 5228
rect 294104 5216 294110 5228
rect 321646 5216 321652 5228
rect 294104 5188 321652 5216
rect 294104 5176 294110 5188
rect 321646 5176 321652 5188
rect 321704 5176 321710 5228
rect 353386 5176 353392 5228
rect 353444 5216 353450 5228
rect 385954 5216 385960 5228
rect 353444 5188 385960 5216
rect 353444 5176 353450 5188
rect 385954 5176 385960 5188
rect 386012 5176 386018 5228
rect 394694 5176 394700 5228
rect 394752 5216 394758 5228
rect 519538 5216 519544 5228
rect 394752 5188 519544 5216
rect 394752 5176 394758 5188
rect 519538 5176 519544 5188
rect 519596 5176 519602 5228
rect 121086 5108 121092 5160
rect 121144 5148 121150 5160
rect 188338 5148 188344 5160
rect 121144 5120 188344 5148
rect 121144 5108 121150 5120
rect 188338 5108 188344 5120
rect 188396 5108 188402 5160
rect 189718 5108 189724 5160
rect 189776 5148 189782 5160
rect 292574 5148 292580 5160
rect 189776 5120 292580 5148
rect 189776 5108 189782 5120
rect 292574 5108 292580 5120
rect 292632 5108 292638 5160
rect 299658 5108 299664 5160
rect 299716 5148 299722 5160
rect 327258 5148 327264 5160
rect 299716 5120 327264 5148
rect 299716 5108 299722 5120
rect 327258 5108 327264 5120
rect 327316 5108 327322 5160
rect 353478 5108 353484 5160
rect 353536 5148 353542 5160
rect 387150 5148 387156 5160
rect 353536 5120 387156 5148
rect 353536 5108 353542 5120
rect 387150 5108 387156 5120
rect 387208 5108 387214 5160
rect 396074 5108 396080 5160
rect 396132 5148 396138 5160
rect 523034 5148 523040 5160
rect 396132 5120 523040 5148
rect 396132 5108 396138 5120
rect 523034 5108 523040 5120
rect 523092 5108 523098 5160
rect 96246 5040 96252 5092
rect 96304 5080 96310 5092
rect 163498 5080 163504 5092
rect 96304 5052 163504 5080
rect 96304 5040 96310 5052
rect 163498 5040 163504 5052
rect 163556 5040 163562 5092
rect 186130 5040 186136 5092
rect 186188 5080 186194 5092
rect 291286 5080 291292 5092
rect 186188 5052 291292 5080
rect 186188 5040 186194 5052
rect 291286 5040 291292 5052
rect 291344 5040 291350 5092
rect 296070 5040 296076 5092
rect 296128 5080 296134 5092
rect 325786 5080 325792 5092
rect 296128 5052 325792 5080
rect 296128 5040 296134 5052
rect 325786 5040 325792 5052
rect 325844 5040 325850 5092
rect 354674 5040 354680 5092
rect 354732 5080 354738 5092
rect 389450 5080 389456 5092
rect 354732 5052 389456 5080
rect 354732 5040 354738 5052
rect 389450 5040 389456 5052
rect 389508 5040 389514 5092
rect 397546 5040 397552 5092
rect 397604 5080 397610 5092
rect 526622 5080 526628 5092
rect 397604 5052 526628 5080
rect 397604 5040 397610 5052
rect 526622 5040 526628 5052
rect 526680 5040 526686 5092
rect 103330 4972 103336 5024
rect 103388 5012 103394 5024
rect 173158 5012 173164 5024
rect 103388 4984 173164 5012
rect 103388 4972 103394 4984
rect 173158 4972 173164 4984
rect 173216 4972 173222 5024
rect 182542 4972 182548 5024
rect 182600 5012 182606 5024
rect 291194 5012 291200 5024
rect 182600 4984 291200 5012
rect 182600 4972 182606 4984
rect 291194 4972 291200 4984
rect 291252 4972 291258 5024
rect 292574 4972 292580 5024
rect 292632 5012 292638 5024
rect 324498 5012 324504 5024
rect 292632 4984 324504 5012
rect 292632 4972 292638 4984
rect 324498 4972 324504 4984
rect 324556 4972 324562 5024
rect 356146 4972 356152 5024
rect 356204 5012 356210 5024
rect 393038 5012 393044 5024
rect 356204 4984 393044 5012
rect 356204 4972 356210 4984
rect 393038 4972 393044 4984
rect 393096 4972 393102 5024
rect 398834 4972 398840 5024
rect 398892 5012 398898 5024
rect 533706 5012 533712 5024
rect 398892 4984 533712 5012
rect 398892 4972 398898 4984
rect 533706 4972 533712 4984
rect 533764 4972 533770 5024
rect 146938 4904 146944 4956
rect 146996 4944 147002 4956
rect 276106 4944 276112 4956
rect 146996 4916 276112 4944
rect 146996 4904 147002 4916
rect 276106 4904 276112 4916
rect 276164 4904 276170 4956
rect 285398 4904 285404 4956
rect 285456 4944 285462 4956
rect 323026 4944 323032 4956
rect 285456 4916 323032 4944
rect 285456 4904 285462 4916
rect 323026 4904 323032 4916
rect 323084 4904 323090 4956
rect 356054 4904 356060 4956
rect 356112 4944 356118 4956
rect 396534 4944 396540 4956
rect 356112 4916 396540 4944
rect 356112 4904 356118 4916
rect 396534 4904 396540 4916
rect 396592 4904 396598 4956
rect 400214 4904 400220 4956
rect 400272 4944 400278 4956
rect 537202 4944 537208 4956
rect 400272 4916 537208 4944
rect 400272 4904 400278 4916
rect 537202 4904 537208 4916
rect 537260 4904 537266 4956
rect 132954 4836 132960 4888
rect 133012 4876 133018 4888
rect 274634 4876 274640 4888
rect 133012 4848 274640 4876
rect 133012 4836 133018 4848
rect 274634 4836 274640 4848
rect 274692 4836 274698 4888
rect 278314 4836 278320 4888
rect 278372 4876 278378 4888
rect 320174 4876 320180 4888
rect 278372 4848 320180 4876
rect 278372 4836 278378 4848
rect 320174 4836 320180 4848
rect 320232 4836 320238 4888
rect 357618 4836 357624 4888
rect 357676 4876 357682 4888
rect 398926 4876 398932 4888
rect 357676 4848 398932 4876
rect 357676 4836 357682 4848
rect 398926 4836 398932 4848
rect 398984 4836 398990 4888
rect 401594 4836 401600 4888
rect 401652 4876 401658 4888
rect 540790 4876 540796 4888
rect 401652 4848 540796 4876
rect 401652 4836 401658 4848
rect 540790 4836 540796 4848
rect 540848 4836 540854 4888
rect 129366 4768 129372 4820
rect 129424 4808 129430 4820
rect 274726 4808 274732 4820
rect 129424 4780 274732 4808
rect 129424 4768 129430 4780
rect 274726 4768 274732 4780
rect 274784 4768 274790 4820
rect 274818 4768 274824 4820
rect 274876 4808 274882 4820
rect 319070 4808 319076 4820
rect 274876 4780 319076 4808
rect 274876 4768 274882 4780
rect 319070 4768 319076 4780
rect 319128 4768 319134 4820
rect 357526 4768 357532 4820
rect 357584 4808 357590 4820
rect 400122 4808 400128 4820
rect 357584 4780 400128 4808
rect 357584 4768 357590 4780
rect 400122 4768 400128 4780
rect 400180 4768 400186 4820
rect 402974 4768 402980 4820
rect 403032 4808 403038 4820
rect 544378 4808 544384 4820
rect 403032 4780 544384 4808
rect 403032 4768 403038 4780
rect 544378 4768 544384 4780
rect 544436 4768 544442 4820
rect 136450 4700 136456 4752
rect 136508 4740 136514 4752
rect 146938 4740 146944 4752
rect 136508 4712 146944 4740
rect 136508 4700 136514 4712
rect 146938 4700 146944 4712
rect 146996 4700 147002 4752
rect 214466 4700 214472 4752
rect 214524 4740 214530 4752
rect 300854 4740 300860 4752
rect 214524 4712 300860 4740
rect 214524 4700 214530 4712
rect 300854 4700 300860 4712
rect 300912 4700 300918 4752
rect 389174 4700 389180 4752
rect 389232 4740 389238 4752
rect 501782 4740 501788 4752
rect 389232 4712 501788 4740
rect 389232 4700 389238 4712
rect 501782 4700 501788 4712
rect 501840 4700 501846 4752
rect 175458 4632 175464 4684
rect 175516 4672 175522 4684
rect 258718 4672 258724 4684
rect 175516 4644 258724 4672
rect 175516 4632 175522 4644
rect 258718 4632 258724 4644
rect 258776 4632 258782 4684
rect 264146 4632 264152 4684
rect 264204 4672 264210 4684
rect 316126 4672 316132 4684
rect 264204 4644 316132 4672
rect 264204 4632 264210 4644
rect 316126 4632 316132 4644
rect 316184 4632 316190 4684
rect 387794 4632 387800 4684
rect 387852 4672 387858 4684
rect 498194 4672 498200 4684
rect 387852 4644 498200 4672
rect 387852 4632 387858 4644
rect 498194 4632 498200 4644
rect 498252 4632 498258 4684
rect 179046 4564 179052 4616
rect 179104 4604 179110 4616
rect 258810 4604 258816 4616
rect 179104 4576 258816 4604
rect 179104 4564 179110 4576
rect 258810 4564 258816 4576
rect 258868 4564 258874 4616
rect 288986 4564 288992 4616
rect 289044 4604 289050 4616
rect 323118 4604 323124 4616
rect 289044 4576 323124 4604
rect 289044 4564 289050 4576
rect 323118 4564 323124 4576
rect 323176 4564 323182 4616
rect 360194 4564 360200 4616
rect 360252 4604 360258 4616
rect 406010 4604 406016 4616
rect 360252 4576 406016 4604
rect 360252 4564 360258 4576
rect 406010 4564 406016 4576
rect 406068 4564 406074 4616
rect 291838 4496 291844 4548
rect 291896 4536 291902 4548
rect 317598 4536 317604 4548
rect 291896 4508 317604 4536
rect 291896 4496 291902 4508
rect 317598 4496 317604 4508
rect 317656 4496 317662 4548
rect 358906 4496 358912 4548
rect 358964 4536 358970 4548
rect 403618 4536 403624 4548
rect 358964 4508 403624 4536
rect 358964 4496 358970 4508
rect 403618 4496 403624 4508
rect 403676 4496 403682 4548
rect 291746 4428 291752 4480
rect 291804 4468 291810 4480
rect 317506 4468 317512 4480
rect 291804 4440 317512 4468
rect 291804 4428 291810 4440
rect 317506 4428 317512 4440
rect 317564 4428 317570 4480
rect 358814 4428 358820 4480
rect 358872 4468 358878 4480
rect 402514 4468 402520 4480
rect 358872 4440 402520 4468
rect 358872 4428 358878 4440
rect 402514 4428 402520 4440
rect 402572 4428 402578 4480
rect 126974 4156 126980 4208
rect 127032 4196 127038 4208
rect 128170 4196 128176 4208
rect 127032 4168 128176 4196
rect 127032 4156 127038 4168
rect 128170 4156 128176 4168
rect 128228 4156 128234 4208
rect 176654 4156 176660 4208
rect 176712 4196 176718 4208
rect 177850 4196 177856 4208
rect 176712 4168 177856 4196
rect 176712 4156 176718 4168
rect 177850 4156 177856 4168
rect 177908 4156 177914 4208
rect 226334 4156 226340 4208
rect 226392 4196 226398 4208
rect 227530 4196 227536 4208
rect 226392 4168 227536 4196
rect 226392 4156 226398 4168
rect 227530 4156 227536 4168
rect 227588 4156 227594 4208
rect 361758 4156 361764 4208
rect 361816 4196 361822 4208
rect 361816 4168 361988 4196
rect 361816 4156 361822 4168
rect 99834 4088 99840 4140
rect 99892 4128 99898 4140
rect 239398 4128 239404 4140
rect 99892 4100 239404 4128
rect 99892 4088 99898 4100
rect 239398 4088 239404 4100
rect 239456 4088 239462 4140
rect 246390 4088 246396 4140
rect 246448 4128 246454 4140
rect 262858 4128 262864 4140
rect 246448 4100 262864 4128
rect 246448 4088 246454 4100
rect 262858 4088 262864 4100
rect 262916 4088 262922 4140
rect 271230 4088 271236 4140
rect 271288 4128 271294 4140
rect 291838 4128 291844 4140
rect 271288 4100 291844 4128
rect 271288 4088 271294 4100
rect 291838 4088 291844 4100
rect 291896 4088 291902 4140
rect 298462 4088 298468 4140
rect 298520 4128 298526 4140
rect 315298 4128 315304 4140
rect 298520 4100 315304 4128
rect 298520 4088 298526 4100
rect 315298 4088 315304 4100
rect 315356 4088 315362 4140
rect 320910 4088 320916 4140
rect 320968 4128 320974 4140
rect 320968 4100 331536 4128
rect 320968 4088 320974 4100
rect 92750 4020 92756 4072
rect 92808 4060 92814 4072
rect 236638 4060 236644 4072
rect 92808 4032 236644 4060
rect 92808 4020 92814 4032
rect 236638 4020 236644 4032
rect 236696 4020 236702 4072
rect 255866 4020 255872 4072
rect 255924 4060 255930 4072
rect 277486 4060 277492 4072
rect 255924 4032 277492 4060
rect 255924 4020 255930 4032
rect 277486 4020 277492 4032
rect 277544 4020 277550 4072
rect 283098 4020 283104 4072
rect 283156 4060 283162 4072
rect 307110 4060 307116 4072
rect 283156 4032 307116 4060
rect 283156 4020 283162 4032
rect 307110 4020 307116 4032
rect 307168 4020 307174 4072
rect 316218 4020 316224 4072
rect 316276 4060 316282 4072
rect 331398 4060 331404 4072
rect 316276 4032 331404 4060
rect 316276 4020 316282 4032
rect 331398 4020 331404 4032
rect 331456 4020 331462 4072
rect 331508 4060 331536 4100
rect 333882 4088 333888 4140
rect 333940 4128 333946 4140
rect 336826 4128 336832 4140
rect 333940 4100 336832 4128
rect 333940 4088 333946 4100
rect 336826 4088 336832 4100
rect 336884 4088 336890 4140
rect 346486 4088 346492 4140
rect 346544 4128 346550 4140
rect 361850 4128 361856 4140
rect 346544 4100 361856 4128
rect 346544 4088 346550 4100
rect 361850 4088 361856 4100
rect 361908 4088 361914 4140
rect 334066 4060 334072 4072
rect 331508 4032 334072 4060
rect 334066 4020 334072 4032
rect 334124 4020 334130 4072
rect 343818 4020 343824 4072
rect 343876 4060 343882 4072
rect 354030 4060 354036 4072
rect 343876 4032 354036 4060
rect 343876 4020 343882 4032
rect 354030 4020 354036 4032
rect 354088 4020 354094 4072
rect 358170 4020 358176 4072
rect 358228 4060 358234 4072
rect 361960 4060 361988 4168
rect 362310 4088 362316 4140
rect 362368 4128 362374 4140
rect 364334 4128 364340 4140
rect 362368 4100 364340 4128
rect 362368 4088 362374 4100
rect 364334 4088 364340 4100
rect 364392 4088 364398 4140
rect 364978 4088 364984 4140
rect 365036 4128 365042 4140
rect 368198 4128 368204 4140
rect 365036 4100 368204 4128
rect 365036 4088 365042 4100
rect 368198 4088 368204 4100
rect 368256 4088 368262 4140
rect 382274 4088 382280 4140
rect 382332 4128 382338 4140
rect 411898 4128 411904 4140
rect 382332 4100 411904 4128
rect 382332 4088 382338 4100
rect 411898 4088 411904 4100
rect 411956 4088 411962 4140
rect 418798 4088 418804 4140
rect 418856 4128 418862 4140
rect 419074 4128 419080 4140
rect 418856 4100 419080 4128
rect 418856 4088 418862 4100
rect 419074 4088 419080 4100
rect 419132 4088 419138 4140
rect 425790 4088 425796 4140
rect 425848 4128 425854 4140
rect 440326 4128 440332 4140
rect 425848 4100 440332 4128
rect 425848 4088 425854 4100
rect 440326 4088 440332 4100
rect 440384 4088 440390 4140
rect 442258 4088 442264 4140
rect 442316 4128 442322 4140
rect 442718 4128 442724 4140
rect 442316 4100 442724 4128
rect 442316 4088 442322 4100
rect 442718 4088 442724 4100
rect 442776 4088 442782 4140
rect 447778 4088 447784 4140
rect 447836 4128 447842 4140
rect 475746 4128 475752 4140
rect 447836 4100 475752 4128
rect 447836 4088 447842 4100
rect 475746 4088 475752 4100
rect 475804 4088 475810 4140
rect 377674 4060 377680 4072
rect 358228 4032 358860 4060
rect 358228 4020 358234 4032
rect 82078 3952 82084 4004
rect 82136 3992 82142 4004
rect 259454 3992 259460 4004
rect 82136 3964 259460 3992
rect 82136 3952 82142 3964
rect 259454 3952 259460 3964
rect 259512 3952 259518 4004
rect 267734 3952 267740 4004
rect 267792 3992 267798 4004
rect 291746 3992 291752 4004
rect 267792 3964 291752 3992
rect 267792 3952 267798 3964
rect 291746 3952 291752 3964
rect 291804 3952 291810 4004
rect 294874 3952 294880 4004
rect 294932 3992 294938 4004
rect 325878 3992 325884 4004
rect 294932 3964 325884 3992
rect 294932 3952 294938 3964
rect 325878 3952 325884 3964
rect 325936 3952 325942 4004
rect 345106 3952 345112 4004
rect 345164 3992 345170 4004
rect 358722 3992 358728 4004
rect 345164 3964 358728 3992
rect 345164 3952 345170 3964
rect 358722 3952 358728 3964
rect 358780 3952 358786 4004
rect 358832 3992 358860 4032
rect 360166 4032 361896 4060
rect 361960 4032 377680 4060
rect 360166 3992 360194 4032
rect 358832 3964 360194 3992
rect 361868 3992 361896 4032
rect 377674 4020 377680 4032
rect 377732 4020 377738 4072
rect 379514 4020 379520 4072
rect 379572 4060 379578 4072
rect 472250 4060 472256 4072
rect 379572 4032 472256 4060
rect 379572 4020 379578 4032
rect 472250 4020 472256 4032
rect 472308 4020 472314 4072
rect 381170 3992 381176 4004
rect 361868 3964 381176 3992
rect 381170 3952 381176 3964
rect 381228 3952 381234 4004
rect 382458 3952 382464 4004
rect 382516 3992 382522 4004
rect 479334 3992 479340 4004
rect 382516 3964 479340 3992
rect 382516 3952 382522 3964
rect 479334 3952 479340 3964
rect 479392 3952 479398 4004
rect 43070 3884 43076 3936
rect 43128 3924 43134 3936
rect 247034 3924 247040 3936
rect 43128 3896 247040 3924
rect 43128 3884 43134 3896
rect 247034 3884 247040 3896
rect 247092 3884 247098 3936
rect 252370 3884 252376 3936
rect 252428 3924 252434 3936
rect 275186 3924 275192 3936
rect 252428 3896 275192 3924
rect 252428 3884 252434 3896
rect 275186 3884 275192 3896
rect 275244 3884 275250 3936
rect 287790 3884 287796 3936
rect 287848 3924 287854 3936
rect 322934 3924 322940 3936
rect 287848 3896 322940 3924
rect 287848 3884 287854 3896
rect 322934 3884 322940 3896
rect 322992 3884 322998 3936
rect 325602 3884 325608 3936
rect 325660 3924 325666 3936
rect 335354 3924 335360 3936
rect 325660 3896 335360 3924
rect 325660 3884 325666 3896
rect 335354 3884 335360 3896
rect 335412 3884 335418 3936
rect 340966 3884 340972 3936
rect 341024 3924 341030 3936
rect 346946 3924 346952 3936
rect 341024 3896 346952 3924
rect 341024 3884 341030 3896
rect 346946 3884 346952 3896
rect 347004 3884 347010 3936
rect 347866 3884 347872 3936
rect 347924 3924 347930 3936
rect 359458 3924 359464 3936
rect 347924 3896 359464 3924
rect 347924 3884 347930 3896
rect 359458 3884 359464 3896
rect 359516 3884 359522 3936
rect 361758 3924 361764 3936
rect 359568 3896 361764 3924
rect 35986 3816 35992 3868
rect 36044 3856 36050 3868
rect 245654 3856 245660 3868
rect 36044 3828 245660 3856
rect 36044 3816 36050 3828
rect 245654 3816 245660 3828
rect 245712 3816 245718 3868
rect 248782 3816 248788 3868
rect 248840 3856 248846 3868
rect 274542 3856 274548 3868
rect 248840 3828 274548 3856
rect 248840 3816 248846 3828
rect 274542 3816 274548 3828
rect 274600 3816 274606 3868
rect 280706 3816 280712 3868
rect 280764 3856 280770 3868
rect 321738 3856 321744 3868
rect 280764 3828 321744 3856
rect 280764 3816 280770 3828
rect 321738 3816 321744 3828
rect 321796 3816 321802 3868
rect 326798 3816 326804 3868
rect 326856 3856 326862 3868
rect 335446 3856 335452 3868
rect 326856 3828 335452 3856
rect 326856 3816 326862 3828
rect 335446 3816 335452 3828
rect 335504 3816 335510 3868
rect 343910 3816 343916 3868
rect 343968 3856 343974 3868
rect 355226 3856 355232 3868
rect 343968 3828 355232 3856
rect 343968 3816 343974 3828
rect 355226 3816 355232 3828
rect 355284 3816 355290 3868
rect 356698 3816 356704 3868
rect 356756 3856 356762 3868
rect 359568 3856 359596 3896
rect 361758 3884 361764 3896
rect 361816 3884 361822 3936
rect 361850 3884 361856 3936
rect 361908 3924 361914 3936
rect 363506 3924 363512 3936
rect 361908 3896 363512 3924
rect 361908 3884 361914 3896
rect 363506 3884 363512 3896
rect 363564 3884 363570 3936
rect 367738 3884 367744 3936
rect 367796 3924 367802 3936
rect 390646 3924 390652 3936
rect 367796 3896 390652 3924
rect 367796 3884 367802 3896
rect 390646 3884 390652 3896
rect 390704 3884 390710 3936
rect 391198 3884 391204 3936
rect 391256 3924 391262 3936
rect 422570 3924 422576 3936
rect 391256 3896 422576 3924
rect 391256 3884 391262 3896
rect 422570 3884 422576 3896
rect 422628 3884 422634 3936
rect 428550 3884 428556 3936
rect 428608 3924 428614 3936
rect 450906 3924 450912 3936
rect 428608 3896 450912 3924
rect 428608 3884 428614 3896
rect 450906 3884 450912 3896
rect 450964 3884 450970 3936
rect 454678 3884 454684 3936
rect 454736 3924 454742 3936
rect 583386 3924 583392 3936
rect 454736 3896 583392 3924
rect 454736 3884 454742 3896
rect 583386 3884 583392 3896
rect 583444 3884 583450 3936
rect 356756 3828 359596 3856
rect 356756 3816 356762 3828
rect 361482 3816 361488 3868
rect 361540 3856 361546 3868
rect 374086 3856 374092 3868
rect 361540 3828 374092 3856
rect 361540 3816 361546 3828
rect 374086 3816 374092 3828
rect 374144 3816 374150 3868
rect 376018 3816 376024 3868
rect 376076 3856 376082 3868
rect 443822 3856 443828 3868
rect 376076 3828 443828 3856
rect 376076 3816 376082 3828
rect 443822 3816 443828 3828
rect 443880 3816 443886 3868
rect 450538 3816 450544 3868
rect 450596 3856 450602 3868
rect 580994 3856 581000 3868
rect 450596 3828 581000 3856
rect 450596 3816 450602 3828
rect 580994 3816 581000 3828
rect 581052 3816 581058 3868
rect 28902 3748 28908 3800
rect 28960 3788 28966 3800
rect 242894 3788 242900 3800
rect 28960 3760 242900 3788
rect 28960 3748 28966 3760
rect 242894 3748 242900 3760
rect 242952 3748 242958 3800
rect 260650 3748 260656 3800
rect 260708 3788 260714 3800
rect 307202 3788 307208 3800
rect 260708 3760 307208 3788
rect 260708 3748 260714 3760
rect 307202 3748 307208 3760
rect 307260 3748 307266 3800
rect 311434 3748 311440 3800
rect 311492 3788 311498 3800
rect 329926 3788 329932 3800
rect 311492 3760 329932 3788
rect 311492 3748 311498 3760
rect 329926 3748 329932 3760
rect 329984 3748 329990 3800
rect 347958 3748 347964 3800
rect 348016 3788 348022 3800
rect 369394 3788 369400 3800
rect 348016 3760 369400 3788
rect 348016 3748 348022 3760
rect 369394 3748 369400 3760
rect 369452 3748 369458 3800
rect 369486 3748 369492 3800
rect 369544 3788 369550 3800
rect 375282 3788 375288 3800
rect 369544 3760 375288 3788
rect 369544 3748 369550 3760
rect 375282 3748 375288 3760
rect 375340 3748 375346 3800
rect 377398 3748 377404 3800
rect 377456 3788 377462 3800
rect 408402 3788 408408 3800
rect 377456 3760 408408 3788
rect 377456 3748 377462 3760
rect 408402 3748 408408 3760
rect 408460 3748 408466 3800
rect 418890 3748 418896 3800
rect 418948 3788 418954 3800
rect 560846 3788 560852 3800
rect 418948 3760 560852 3788
rect 418948 3748 418954 3760
rect 560846 3748 560852 3760
rect 560904 3748 560910 3800
rect 24210 3680 24216 3732
rect 24268 3720 24274 3732
rect 241790 3720 241796 3732
rect 24268 3692 241796 3720
rect 24268 3680 24274 3692
rect 241790 3680 241796 3692
rect 241848 3680 241854 3732
rect 247586 3680 247592 3732
rect 247644 3720 247650 3732
rect 297174 3720 297180 3732
rect 247644 3692 297180 3720
rect 247644 3680 247650 3692
rect 297174 3680 297180 3692
rect 297232 3680 297238 3732
rect 310238 3680 310244 3732
rect 310296 3720 310302 3732
rect 312630 3720 312636 3732
rect 310296 3692 312636 3720
rect 310296 3680 310302 3692
rect 312630 3680 312636 3692
rect 312688 3680 312694 3732
rect 312722 3680 312728 3732
rect 312780 3720 312786 3732
rect 330018 3720 330024 3732
rect 312780 3692 330024 3720
rect 312780 3680 312786 3692
rect 330018 3680 330024 3692
rect 330076 3680 330082 3732
rect 335078 3680 335084 3732
rect 335136 3720 335142 3732
rect 338114 3720 338120 3732
rect 335136 3692 338120 3720
rect 335136 3680 335142 3692
rect 338114 3680 338120 3692
rect 338172 3680 338178 3732
rect 341058 3680 341064 3732
rect 341116 3720 341122 3732
rect 345750 3720 345756 3732
rect 341116 3692 345756 3720
rect 341116 3680 341122 3692
rect 345750 3680 345756 3692
rect 345808 3680 345814 3732
rect 347774 3680 347780 3732
rect 347832 3720 347838 3732
rect 365806 3720 365812 3732
rect 347832 3692 365812 3720
rect 347832 3680 347838 3692
rect 365806 3680 365812 3692
rect 365864 3680 365870 3732
rect 366450 3680 366456 3732
rect 366508 3720 366514 3732
rect 391842 3720 391848 3732
rect 366508 3692 391848 3720
rect 366508 3680 366514 3692
rect 391842 3680 391848 3692
rect 391900 3680 391906 3732
rect 391934 3680 391940 3732
rect 391992 3720 391998 3732
rect 426158 3720 426164 3732
rect 391992 3692 426164 3720
rect 391992 3680 391998 3692
rect 426158 3680 426164 3692
rect 426216 3680 426222 3732
rect 431218 3680 431224 3732
rect 431276 3720 431282 3732
rect 575106 3720 575112 3732
rect 431276 3692 575112 3720
rect 431276 3680 431282 3692
rect 575106 3680 575112 3692
rect 575164 3680 575170 3732
rect 19426 3612 19432 3664
rect 19484 3652 19490 3664
rect 240134 3652 240140 3664
rect 19484 3624 240140 3652
rect 19484 3612 19490 3624
rect 240134 3612 240140 3624
rect 240192 3612 240198 3664
rect 251174 3612 251180 3664
rect 251232 3652 251238 3664
rect 301498 3652 301504 3664
rect 251232 3624 301504 3652
rect 251232 3612 251238 3624
rect 301498 3612 301504 3624
rect 301556 3612 301562 3664
rect 305546 3612 305552 3664
rect 305604 3652 305610 3664
rect 328730 3652 328736 3664
rect 305604 3624 328736 3652
rect 305604 3612 305610 3624
rect 328730 3612 328736 3624
rect 328788 3612 328794 3664
rect 349154 3612 349160 3664
rect 349212 3652 349218 3664
rect 370590 3652 370596 3664
rect 349212 3624 370596 3652
rect 349212 3612 349218 3624
rect 370590 3612 370596 3624
rect 370648 3612 370654 3664
rect 374638 3612 374644 3664
rect 374696 3652 374702 3664
rect 401318 3652 401324 3664
rect 374696 3624 401324 3652
rect 374696 3612 374702 3624
rect 401318 3612 401324 3624
rect 401376 3612 401382 3664
rect 404354 3612 404360 3664
rect 404412 3652 404418 3664
rect 550266 3652 550272 3664
rect 404412 3624 550272 3652
rect 404412 3612 404418 3624
rect 550266 3612 550272 3624
rect 550324 3612 550330 3664
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 240226 3584 240232 3596
rect 20680 3556 240232 3584
rect 20680 3544 20686 3556
rect 240226 3544 240232 3556
rect 240284 3544 240290 3596
rect 244090 3544 244096 3596
rect 244148 3584 244154 3596
rect 297726 3584 297732 3596
rect 244148 3556 297732 3584
rect 244148 3544 244154 3556
rect 297726 3544 297732 3556
rect 297784 3544 297790 3596
rect 304350 3544 304356 3596
rect 304408 3584 304414 3596
rect 328546 3584 328552 3596
rect 304408 3556 328552 3584
rect 304408 3544 304414 3556
rect 328546 3544 328552 3556
rect 328604 3544 328610 3596
rect 332686 3544 332692 3596
rect 332744 3584 332750 3596
rect 336918 3584 336924 3596
rect 332744 3556 336924 3584
rect 332744 3544 332750 3556
rect 336918 3544 336924 3556
rect 336976 3544 336982 3596
rect 350534 3544 350540 3596
rect 350592 3584 350598 3596
rect 376478 3584 376484 3596
rect 350592 3556 376484 3584
rect 350592 3544 350598 3556
rect 376478 3544 376484 3556
rect 376536 3544 376542 3596
rect 384942 3544 384948 3596
rect 385000 3584 385006 3596
rect 418982 3584 418988 3596
rect 385000 3556 418988 3584
rect 385000 3544 385006 3556
rect 418982 3544 418988 3556
rect 419040 3544 419046 3596
rect 419074 3544 419080 3596
rect 419132 3584 419138 3596
rect 568022 3584 568028 3596
rect 419132 3556 568028 3584
rect 419132 3544 419138 3556
rect 568022 3544 568028 3556
rect 568080 3544 568086 3596
rect 14734 3476 14740 3528
rect 14792 3516 14798 3528
rect 238938 3516 238944 3528
rect 14792 3488 238944 3516
rect 14792 3476 14798 3488
rect 238938 3476 238944 3488
rect 238996 3476 239002 3528
rect 245194 3476 245200 3528
rect 245252 3516 245258 3528
rect 299290 3516 299296 3528
rect 245252 3488 299296 3516
rect 245252 3476 245258 3488
rect 299290 3476 299296 3488
rect 299348 3476 299354 3528
rect 301958 3476 301964 3528
rect 302016 3516 302022 3528
rect 327350 3516 327356 3528
rect 302016 3488 327356 3516
rect 302016 3476 302022 3488
rect 327350 3476 327356 3488
rect 327408 3476 327414 3528
rect 343726 3476 343732 3528
rect 343784 3516 343790 3528
rect 352834 3516 352840 3528
rect 343784 3488 352840 3516
rect 343784 3476 343790 3488
rect 352834 3476 352840 3488
rect 352892 3476 352898 3528
rect 353294 3476 353300 3528
rect 353352 3516 353358 3528
rect 383562 3516 383568 3528
rect 353352 3488 383568 3516
rect 353352 3476 353358 3488
rect 383562 3476 383568 3488
rect 383620 3476 383626 3528
rect 405734 3476 405740 3528
rect 405792 3516 405798 3528
rect 557350 3516 557356 3528
rect 405792 3488 557356 3516
rect 405792 3476 405798 3488
rect 557350 3476 557356 3488
rect 557408 3476 557414 3528
rect 11146 3408 11152 3460
rect 11204 3448 11210 3460
rect 237374 3448 237380 3460
rect 11204 3420 237380 3448
rect 11204 3408 11210 3420
rect 237374 3408 237380 3420
rect 237432 3408 237438 3460
rect 242894 3408 242900 3460
rect 242952 3448 242958 3460
rect 242952 3420 306696 3448
rect 242952 3408 242958 3420
rect 44174 3340 44180 3392
rect 44232 3380 44238 3392
rect 45094 3380 45100 3392
rect 44232 3352 45100 3380
rect 44232 3340 44238 3352
rect 45094 3340 45100 3352
rect 45152 3340 45158 3392
rect 52454 3340 52460 3392
rect 52512 3380 52518 3392
rect 53374 3380 53380 3392
rect 52512 3352 53380 3380
rect 52512 3340 52518 3352
rect 53374 3340 53380 3352
rect 53432 3340 53438 3392
rect 93854 3340 93860 3392
rect 93912 3380 93918 3392
rect 94774 3380 94780 3392
rect 93912 3352 94780 3380
rect 93912 3340 93918 3352
rect 94774 3340 94780 3352
rect 94832 3340 94838 3392
rect 110414 3340 110420 3392
rect 110472 3380 110478 3392
rect 111610 3380 111616 3392
rect 110472 3352 111616 3380
rect 110472 3340 110478 3352
rect 111610 3340 111616 3352
rect 111668 3340 111674 3392
rect 242250 3380 242256 3392
rect 113146 3352 242256 3380
rect 106918 3272 106924 3324
rect 106976 3312 106982 3324
rect 113146 3312 113174 3352
rect 242250 3340 242256 3352
rect 242308 3340 242314 3392
rect 249978 3340 249984 3392
rect 250036 3380 250042 3392
rect 264238 3380 264244 3392
rect 250036 3352 264244 3380
rect 250036 3340 250042 3352
rect 264238 3340 264244 3352
rect 264296 3340 264302 3392
rect 266538 3340 266544 3392
rect 266596 3380 266602 3392
rect 283650 3380 283656 3392
rect 266596 3352 283656 3380
rect 266596 3340 266602 3352
rect 283650 3340 283656 3352
rect 283708 3340 283714 3392
rect 291378 3340 291384 3392
rect 291436 3380 291442 3392
rect 306668 3380 306696 3420
rect 306742 3408 306748 3460
rect 306800 3448 306806 3460
rect 311158 3448 311164 3460
rect 306800 3420 311164 3448
rect 306800 3408 306806 3420
rect 311158 3408 311164 3420
rect 311216 3408 311222 3460
rect 312630 3408 312636 3460
rect 312688 3448 312694 3460
rect 331306 3448 331312 3460
rect 312688 3420 331312 3448
rect 312688 3408 312694 3420
rect 331306 3408 331312 3420
rect 331364 3408 331370 3460
rect 337470 3408 337476 3460
rect 337528 3448 337534 3460
rect 338298 3448 338304 3460
rect 337528 3420 338304 3448
rect 337528 3408 337534 3420
rect 338298 3408 338304 3420
rect 338356 3408 338362 3460
rect 343634 3408 343640 3460
rect 343692 3448 343698 3460
rect 356330 3448 356336 3460
rect 343692 3420 356336 3448
rect 343692 3408 343698 3420
rect 356330 3408 356336 3420
rect 356388 3408 356394 3460
rect 359458 3408 359464 3460
rect 359516 3448 359522 3460
rect 367002 3448 367008 3460
rect 359516 3420 367008 3448
rect 359516 3408 359522 3420
rect 367002 3408 367008 3420
rect 367060 3408 367066 3460
rect 369486 3448 369492 3460
rect 367112 3420 369492 3448
rect 291436 3352 306512 3380
rect 306668 3352 307156 3380
rect 291436 3340 291442 3352
rect 106976 3284 113174 3312
rect 106976 3272 106982 3284
rect 118694 3272 118700 3324
rect 118752 3312 118758 3324
rect 119890 3312 119896 3324
rect 118752 3284 119896 3312
rect 118752 3272 118758 3284
rect 119890 3272 119896 3284
rect 119948 3272 119954 3324
rect 242158 3312 242164 3324
rect 122806 3284 242164 3312
rect 114002 3204 114008 3256
rect 114060 3244 114066 3256
rect 122806 3244 122834 3284
rect 242158 3272 242164 3284
rect 242216 3272 242222 3324
rect 253474 3272 253480 3324
rect 253532 3312 253538 3324
rect 265618 3312 265624 3324
rect 253532 3284 265624 3312
rect 253532 3272 253538 3284
rect 265618 3272 265624 3284
rect 265676 3272 265682 3324
rect 293678 3272 293684 3324
rect 293736 3312 293742 3324
rect 305638 3312 305644 3324
rect 293736 3284 305644 3312
rect 293736 3272 293742 3284
rect 305638 3272 305644 3284
rect 305696 3272 305702 3324
rect 114060 3216 122834 3244
rect 114060 3204 114066 3216
rect 124674 3204 124680 3256
rect 124732 3244 124738 3256
rect 244918 3244 244924 3256
rect 124732 3216 244924 3244
rect 124732 3204 124738 3216
rect 244918 3204 244924 3216
rect 244976 3204 244982 3256
rect 257062 3204 257068 3256
rect 257120 3244 257126 3256
rect 268378 3244 268384 3256
rect 257120 3216 268384 3244
rect 257120 3204 257126 3216
rect 268378 3204 268384 3216
rect 268436 3204 268442 3256
rect 281902 3204 281908 3256
rect 281960 3244 281966 3256
rect 294046 3244 294052 3256
rect 281960 3216 294052 3244
rect 281960 3204 281966 3216
rect 294046 3204 294052 3216
rect 294104 3204 294110 3256
rect 143534 3136 143540 3188
rect 143592 3176 143598 3188
rect 144730 3176 144736 3188
rect 143592 3148 144736 3176
rect 143592 3136 143598 3148
rect 144730 3136 144736 3148
rect 144788 3136 144794 3188
rect 259454 3136 259460 3188
rect 259512 3176 259518 3188
rect 268470 3176 268476 3188
rect 259512 3148 268476 3176
rect 259512 3136 259518 3148
rect 268470 3136 268476 3148
rect 268528 3136 268534 3188
rect 306484 3176 306512 3352
rect 307128 3244 307156 3352
rect 307938 3340 307944 3392
rect 307996 3380 308002 3392
rect 312722 3380 312728 3392
rect 307996 3352 312728 3380
rect 307996 3340 308002 3352
rect 312722 3340 312728 3352
rect 312780 3340 312786 3392
rect 319714 3340 319720 3392
rect 319772 3380 319778 3392
rect 332870 3380 332876 3392
rect 319772 3352 332876 3380
rect 319772 3340 319778 3352
rect 332870 3340 332876 3352
rect 332928 3340 332934 3392
rect 342530 3340 342536 3392
rect 342588 3380 342594 3392
rect 342588 3352 344784 3380
rect 342588 3340 342594 3352
rect 309042 3272 309048 3324
rect 309100 3312 309106 3324
rect 319438 3312 319444 3324
rect 309100 3284 319444 3312
rect 309100 3272 309106 3284
rect 319438 3272 319444 3284
rect 319496 3272 319502 3324
rect 323302 3272 323308 3324
rect 323360 3312 323366 3324
rect 333974 3312 333980 3324
rect 323360 3284 333980 3312
rect 323360 3272 323366 3284
rect 333974 3272 333980 3284
rect 334032 3272 334038 3324
rect 336274 3272 336280 3324
rect 336332 3312 336338 3324
rect 338206 3312 338212 3324
rect 336332 3284 338212 3312
rect 336332 3272 336338 3284
rect 338206 3272 338212 3284
rect 338264 3272 338270 3324
rect 338666 3272 338672 3324
rect 338724 3312 338730 3324
rect 339678 3312 339684 3324
rect 338724 3284 339684 3312
rect 338724 3272 338730 3284
rect 339678 3272 339684 3284
rect 339736 3272 339742 3324
rect 342254 3272 342260 3324
rect 342312 3312 342318 3324
rect 342312 3284 344692 3312
rect 342312 3272 342318 3284
rect 309134 3244 309140 3256
rect 307128 3216 309140 3244
rect 309134 3204 309140 3216
rect 309192 3204 309198 3256
rect 324406 3204 324412 3256
rect 324464 3244 324470 3256
rect 334250 3244 334256 3256
rect 324464 3216 334256 3244
rect 324464 3204 324470 3216
rect 334250 3204 334256 3216
rect 334308 3204 334314 3256
rect 312538 3176 312544 3188
rect 306484 3148 312544 3176
rect 312538 3136 312544 3148
rect 312596 3136 312602 3188
rect 327994 3136 328000 3188
rect 328052 3176 328058 3188
rect 335538 3176 335544 3188
rect 328052 3148 335544 3176
rect 328052 3136 328058 3148
rect 335538 3136 335544 3148
rect 335596 3136 335602 3188
rect 339586 3136 339592 3188
rect 339644 3176 339650 3188
rect 340966 3176 340972 3188
rect 339644 3148 340972 3176
rect 339644 3136 339650 3148
rect 340966 3136 340972 3148
rect 341024 3136 341030 3188
rect 341150 3136 341156 3188
rect 341208 3176 341214 3188
rect 344554 3176 344560 3188
rect 341208 3148 344560 3176
rect 341208 3136 341214 3148
rect 344554 3136 344560 3148
rect 344612 3136 344618 3188
rect 344664 3176 344692 3284
rect 344756 3244 344784 3352
rect 346394 3340 346400 3392
rect 346452 3380 346458 3392
rect 346452 3352 355272 3380
rect 346452 3340 346458 3352
rect 345014 3272 345020 3324
rect 345072 3312 345078 3324
rect 345072 3284 354674 3312
rect 345072 3272 345078 3284
rect 351638 3244 351644 3256
rect 344756 3216 351644 3244
rect 351638 3204 351644 3216
rect 351696 3204 351702 3256
rect 349246 3176 349252 3188
rect 344664 3148 349252 3176
rect 349246 3136 349252 3148
rect 349304 3136 349310 3188
rect 297266 3068 297272 3120
rect 297324 3108 297330 3120
rect 307018 3108 307024 3120
rect 297324 3080 307024 3108
rect 297324 3068 297330 3080
rect 307018 3068 307024 3080
rect 307076 3068 307082 3120
rect 322106 3068 322112 3120
rect 322164 3108 322170 3120
rect 334158 3108 334164 3120
rect 322164 3080 334164 3108
rect 322164 3068 322170 3080
rect 334158 3068 334164 3080
rect 334216 3068 334222 3120
rect 342438 3068 342444 3120
rect 342496 3108 342502 3120
rect 348050 3108 348056 3120
rect 342496 3080 348056 3108
rect 342496 3068 342502 3080
rect 348050 3068 348056 3080
rect 348108 3068 348114 3120
rect 329190 3000 329196 3052
rect 329248 3040 329254 3052
rect 335630 3040 335636 3052
rect 329248 3012 335636 3040
rect 329248 3000 329254 3012
rect 335630 3000 335636 3012
rect 335688 3000 335694 3052
rect 341242 3000 341248 3052
rect 341300 3040 341306 3052
rect 343358 3040 343364 3052
rect 341300 3012 343364 3040
rect 341300 3000 341306 3012
rect 343358 3000 343364 3012
rect 343416 3000 343422 3052
rect 350442 3040 350448 3052
rect 344986 3012 350448 3040
rect 342346 2932 342352 2984
rect 342404 2972 342410 2984
rect 344986 2972 345014 3012
rect 350442 3000 350448 3012
rect 350500 3000 350506 3052
rect 342404 2944 345014 2972
rect 354646 2972 354674 3284
rect 355244 3244 355272 3352
rect 355410 3340 355416 3392
rect 355468 3380 355474 3392
rect 357526 3380 357532 3392
rect 355468 3352 357532 3380
rect 355468 3340 355474 3352
rect 357526 3340 357532 3352
rect 357584 3340 357590 3392
rect 363598 3340 363604 3392
rect 363656 3380 363662 3392
rect 367112 3380 367140 3420
rect 369486 3408 369492 3420
rect 369544 3408 369550 3460
rect 370498 3408 370504 3460
rect 370556 3448 370562 3460
rect 371694 3448 371700 3460
rect 370556 3420 371700 3448
rect 370556 3408 370562 3420
rect 371694 3408 371700 3420
rect 371752 3408 371758 3460
rect 371786 3408 371792 3460
rect 371844 3448 371850 3460
rect 397730 3448 397736 3460
rect 371844 3420 397736 3448
rect 371844 3408 371850 3420
rect 397730 3408 397736 3420
rect 397788 3408 397794 3460
rect 411254 3408 411260 3460
rect 411312 3448 411318 3460
rect 571518 3448 571524 3460
rect 411312 3420 571524 3448
rect 411312 3408 411318 3420
rect 571518 3408 571524 3420
rect 571576 3408 571582 3460
rect 363656 3352 367140 3380
rect 363656 3340 363662 3352
rect 369210 3340 369216 3392
rect 369268 3380 369274 3392
rect 369268 3352 371924 3380
rect 369268 3340 369274 3352
rect 362218 3272 362224 3324
rect 362276 3312 362282 3324
rect 371896 3312 371924 3352
rect 371970 3340 371976 3392
rect 372028 3380 372034 3392
rect 388254 3380 388260 3392
rect 372028 3352 388260 3380
rect 372028 3340 372034 3352
rect 388254 3340 388260 3352
rect 388312 3340 388318 3392
rect 388438 3340 388444 3392
rect 388496 3380 388502 3392
rect 415486 3380 415492 3392
rect 388496 3352 415492 3380
rect 388496 3340 388502 3352
rect 415486 3340 415492 3352
rect 415544 3340 415550 3392
rect 423674 3340 423680 3392
rect 423732 3380 423738 3392
rect 424962 3380 424968 3392
rect 423732 3352 424968 3380
rect 423732 3340 423738 3352
rect 424962 3340 424968 3352
rect 425020 3340 425026 3392
rect 448606 3340 448612 3392
rect 448664 3380 448670 3392
rect 449802 3380 449808 3392
rect 448664 3352 449808 3380
rect 448664 3340 448670 3352
rect 449802 3340 449808 3352
rect 449860 3340 449866 3392
rect 468662 3380 468668 3392
rect 449912 3352 468668 3380
rect 395338 3312 395344 3324
rect 362276 3284 369854 3312
rect 371896 3284 395344 3312
rect 362276 3272 362282 3284
rect 362310 3244 362316 3256
rect 355244 3216 362316 3244
rect 362310 3204 362316 3216
rect 362368 3204 362374 3256
rect 369826 3244 369854 3284
rect 395338 3272 395344 3284
rect 395396 3272 395402 3324
rect 442718 3272 442724 3324
rect 442776 3312 442782 3324
rect 449912 3312 449940 3352
rect 468662 3340 468668 3352
rect 468720 3340 468726 3392
rect 489914 3340 489920 3392
rect 489972 3380 489978 3392
rect 490742 3380 490748 3392
rect 489972 3352 490748 3380
rect 489972 3340 489978 3352
rect 490742 3340 490748 3352
rect 490800 3340 490806 3392
rect 442776 3284 449940 3312
rect 442776 3272 442782 3284
rect 449986 3272 449992 3324
rect 450044 3312 450050 3324
rect 461578 3312 461584 3324
rect 450044 3284 461584 3312
rect 450044 3272 450050 3284
rect 461578 3272 461584 3284
rect 461636 3272 461642 3324
rect 384758 3244 384764 3256
rect 369826 3216 384764 3244
rect 384758 3204 384764 3216
rect 384816 3204 384822 3256
rect 439498 3204 439504 3256
rect 439556 3244 439562 3256
rect 458082 3244 458088 3256
rect 439556 3216 458088 3244
rect 439556 3204 439562 3216
rect 458082 3204 458088 3216
rect 458140 3204 458146 3256
rect 355318 3136 355324 3188
rect 355376 3176 355382 3188
rect 361482 3176 361488 3188
rect 355376 3148 361488 3176
rect 355376 3136 355382 3148
rect 361482 3136 361488 3148
rect 361540 3136 361546 3188
rect 371786 3176 371792 3188
rect 361592 3148 371792 3176
rect 357434 3068 357440 3120
rect 357492 3108 357498 3120
rect 361592 3108 361620 3148
rect 371786 3136 371792 3148
rect 371844 3136 371850 3188
rect 371878 3136 371884 3188
rect 371936 3176 371942 3188
rect 371936 3148 373028 3176
rect 371936 3136 371942 3148
rect 357492 3080 361620 3108
rect 357492 3068 357498 3080
rect 367830 3068 367836 3120
rect 367888 3108 367894 3120
rect 372890 3108 372896 3120
rect 367888 3080 372896 3108
rect 367888 3068 367894 3080
rect 372890 3068 372896 3080
rect 372948 3068 372954 3120
rect 373000 3108 373028 3148
rect 373350 3136 373356 3188
rect 373408 3176 373414 3188
rect 394234 3176 394240 3188
rect 373408 3148 394240 3176
rect 373408 3136 373414 3148
rect 394234 3136 394240 3148
rect 394292 3136 394298 3188
rect 422938 3136 422944 3188
rect 422996 3176 423002 3188
rect 429654 3176 429660 3188
rect 422996 3148 429660 3176
rect 422996 3136 423002 3148
rect 429654 3136 429660 3148
rect 429712 3136 429718 3188
rect 440878 3136 440884 3188
rect 440936 3176 440942 3188
rect 454494 3176 454500 3188
rect 440936 3148 454500 3176
rect 440936 3136 440942 3148
rect 454494 3136 454500 3148
rect 454552 3136 454558 3188
rect 379974 3108 379980 3120
rect 373000 3080 379980 3108
rect 379974 3068 379980 3080
rect 380032 3068 380038 3120
rect 436830 3068 436836 3120
rect 436888 3108 436894 3120
rect 447410 3108 447416 3120
rect 436888 3080 447416 3108
rect 436888 3068 436894 3080
rect 447410 3068 447416 3080
rect 447468 3068 447474 3120
rect 358078 3000 358084 3052
rect 358136 3040 358142 3052
rect 361114 3040 361120 3052
rect 358136 3012 361120 3040
rect 358136 3000 358142 3012
rect 361114 3000 361120 3012
rect 361172 3000 361178 3052
rect 425698 3000 425704 3052
rect 425756 3040 425762 3052
rect 433242 3040 433248 3052
rect 425756 3012 433248 3040
rect 425756 3000 425762 3012
rect 433242 3000 433248 3012
rect 433300 3000 433306 3052
rect 443638 3000 443644 3052
rect 443696 3040 443702 3052
rect 449986 3040 449992 3052
rect 443696 3012 449992 3040
rect 443696 3000 443702 3012
rect 449986 3000 449992 3012
rect 450044 3000 450050 3052
rect 359918 2972 359924 2984
rect 354646 2944 359924 2972
rect 342404 2932 342410 2944
rect 359918 2932 359924 2944
rect 359976 2932 359982 2984
rect 366358 2932 366364 2984
rect 366416 2972 366422 2984
rect 371970 2972 371976 2984
rect 366416 2944 371976 2972
rect 366416 2932 366422 2944
rect 371970 2932 371976 2944
rect 372028 2932 372034 2984
<< via1 >>
rect 331220 702992 331272 703044
rect 332508 702992 332560 703044
rect 318800 700952 318852 701004
rect 413652 700952 413704 701004
rect 218980 700884 219032 700936
rect 327908 700884 327960 700936
rect 314660 700816 314712 700868
rect 478512 700816 478564 700868
rect 154120 700748 154172 700800
rect 333244 700748 333296 700800
rect 137836 700680 137888 700732
rect 329104 700680 329156 700732
rect 202788 700612 202840 700664
rect 327724 700612 327776 700664
rect 327816 700612 327868 700664
rect 527180 700612 527232 700664
rect 309140 700544 309192 700596
rect 543464 700544 543516 700596
rect 89168 700476 89220 700528
rect 338764 700476 338816 700528
rect 72976 700408 73028 700460
rect 331864 700408 331916 700460
rect 24308 700340 24360 700392
rect 342904 700340 342956 700392
rect 8116 700272 8168 700324
rect 331956 700272 332008 700324
rect 317420 700204 317472 700256
rect 397460 700204 397512 700256
rect 267648 700136 267700 700188
rect 324964 700136 325016 700188
rect 322940 700068 322992 700120
rect 348792 700068 348844 700120
rect 303620 696940 303672 696992
rect 580172 696940 580224 696992
rect 305000 683204 305052 683256
rect 580172 683204 580224 683256
rect 3424 683136 3476 683188
rect 349160 683136 349212 683188
rect 300860 670760 300912 670812
rect 580172 670760 580224 670812
rect 3516 670692 3568 670744
rect 351920 670692 351972 670744
rect 3424 656888 3476 656940
rect 350540 656888 350592 656940
rect 298100 643084 298152 643136
rect 580172 643084 580224 643136
rect 3424 632068 3476 632120
rect 353300 632068 353352 632120
rect 299572 630640 299624 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 356060 618264 356112 618316
rect 296720 616836 296772 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 354680 605820 354732 605872
rect 293960 590656 294012 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 358820 579640 358872 579692
rect 295340 576852 295392 576904
rect 580172 576852 580224 576904
rect 3424 565836 3476 565888
rect 361580 565836 361632 565888
rect 292580 563048 292632 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 337384 553392 337436 553444
rect 288440 536800 288492 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 362960 527144 363012 527196
rect 289820 524424 289872 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 345664 514768 345716 514820
rect 287060 510620 287112 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 341524 500964 341576 501016
rect 284300 484372 284352 484424
rect 580172 484372 580224 484424
rect 252652 478864 252704 478916
rect 577596 478864 577648 478916
rect 3424 474716 3476 474768
rect 368020 474716 368072 474768
rect 285864 470568 285916 470620
rect 579988 470568 580040 470620
rect 3240 462340 3292 462392
rect 349068 462340 349120 462392
rect 299480 462204 299532 462256
rect 325700 462204 325752 462256
rect 321376 462136 321428 462188
rect 364340 462136 364392 462188
rect 234620 462068 234672 462120
rect 330208 462068 330260 462120
rect 316592 462000 316644 462052
rect 429200 462000 429252 462052
rect 313188 461932 313240 461984
rect 462320 461932 462372 461984
rect 169760 461864 169812 461916
rect 334900 461864 334952 461916
rect 311808 461796 311860 461848
rect 494060 461796 494112 461848
rect 104900 461728 104952 461780
rect 339684 461728 339736 461780
rect 307116 461660 307168 461712
rect 558920 461660 558972 461712
rect 40040 461592 40092 461644
rect 344376 461592 344428 461644
rect 272340 460912 272392 460964
rect 578884 460912 578936 460964
rect 3884 460640 3936 460692
rect 380900 460640 380952 460692
rect 3608 460572 3660 460624
rect 383936 460572 383988 460624
rect 324964 460504 325016 460556
rect 327080 460504 327132 460556
rect 329104 460504 329156 460556
rect 336740 460504 336792 460556
rect 342904 460504 342956 460556
rect 347780 460504 347832 460556
rect 308680 460436 308732 460488
rect 327816 460436 327868 460488
rect 333244 460436 333296 460488
rect 338120 460436 338172 460488
rect 345664 460436 345716 460488
rect 366456 460436 366508 460488
rect 282920 460368 282972 460420
rect 328552 460368 328604 460420
rect 331864 460368 331916 460420
rect 341248 460368 341300 460420
rect 341524 460368 341576 460420
rect 364892 460368 364944 460420
rect 255044 460300 255096 460352
rect 308956 460300 309008 460352
rect 322848 460300 322900 460352
rect 331220 460300 331272 460352
rect 331956 460300 332008 460352
rect 345940 460300 345992 460352
rect 349068 460300 349120 460352
rect 371240 460300 371292 460352
rect 250260 460232 250312 460284
rect 321560 460232 321612 460284
rect 337384 460232 337436 460284
rect 360200 460232 360252 460284
rect 277124 460164 277176 460216
rect 378048 460164 378100 460216
rect 281448 460096 281500 460148
rect 415032 460096 415084 460148
rect 280068 460028 280120 460080
rect 580080 460028 580132 460080
rect 269028 459960 269080 460012
rect 577412 459960 577464 460012
rect 234344 459892 234396 459944
rect 248052 459892 248104 459944
rect 264520 459892 264572 459944
rect 580632 459892 580684 459944
rect 4988 459824 5040 459876
rect 369860 459824 369912 459876
rect 3332 459756 3384 459808
rect 375932 459756 375984 459808
rect 3792 459688 3844 459740
rect 379152 459688 379204 459740
rect 234436 459620 234488 459672
rect 243268 459620 243320 459672
rect 327908 459620 327960 459672
rect 333336 459620 333388 459672
rect 234528 459552 234580 459604
rect 238852 459552 238904 459604
rect 327724 459552 327776 459604
rect 331772 459552 331824 459604
rect 338764 459552 338816 459604
rect 342812 459552 342864 459604
rect 360660 459552 360712 459604
rect 374368 459552 374420 459604
rect 231216 459144 231268 459196
rect 399668 459144 399720 459196
rect 231124 459076 231176 459128
rect 404360 459076 404412 459128
rect 378048 459008 378100 459060
rect 580816 459008 580868 459060
rect 321560 458940 321612 458992
rect 580264 458940 580316 458992
rect 283472 458872 283524 458924
rect 580172 458872 580224 458924
rect 270408 458804 270460 458856
rect 577320 458804 577372 458856
rect 267648 458736 267700 458788
rect 574836 458736 574888 458788
rect 262864 458668 262916 458720
rect 574744 458668 574796 458720
rect 257988 458600 258040 458652
rect 577780 458600 577832 458652
rect 3240 458532 3292 458584
rect 372804 458532 372856 458584
rect 3976 458464 4028 458516
rect 377588 458464 377640 458516
rect 3700 458396 3752 458448
rect 382280 458396 382332 458448
rect 3516 458328 3568 458380
rect 387064 458328 387116 458380
rect 3424 458260 3476 458312
rect 391940 458260 391992 458312
rect 4896 458192 4948 458244
rect 396862 458192 396914 458244
rect 4068 457444 4120 457496
rect 261300 457444 261352 457496
rect 266084 457444 266136 457496
rect 234160 457104 234212 457156
rect 273996 457444 274048 457496
rect 275560 457444 275612 457496
rect 278596 457444 278648 457496
rect 360660 457444 360712 457496
rect 388628 457444 388680 457496
rect 580172 457036 580224 457088
rect 580908 456968 580960 457020
rect 580724 456900 580776 456952
rect 578148 456832 578200 456884
rect 577964 456764 578016 456816
rect 2780 449828 2832 449880
rect 4988 449828 5040 449880
rect 415032 419432 415084 419484
rect 579988 419432 580040 419484
rect 341018 337764 341070 337816
rect 341248 337764 341300 337816
rect 252560 336744 252612 336796
rect 252836 336744 252888 336796
rect 265164 336744 265216 336796
rect 265348 336744 265400 336796
rect 306564 336744 306616 336796
rect 307208 336744 307260 336796
rect 309232 336744 309284 336796
rect 309508 336744 309560 336796
rect 361764 336744 361816 336796
rect 362316 336744 362368 336796
rect 390652 336744 390704 336796
rect 391204 336744 391256 336796
rect 177304 336676 177356 336728
rect 268844 336676 268896 336728
rect 305644 336676 305696 336728
rect 325424 336676 325476 336728
rect 340788 336676 340840 336728
rect 341340 336676 341392 336728
rect 361580 336676 361632 336728
rect 361948 336676 362000 336728
rect 365628 336676 365680 336728
rect 388536 336676 388588 336728
rect 390560 336676 390612 336728
rect 390836 336676 390888 336728
rect 396080 336676 396132 336728
rect 396356 336676 396408 336728
rect 401600 336676 401652 336728
rect 401876 336676 401928 336728
rect 414020 336676 414072 336728
rect 450544 336676 450596 336728
rect 173164 336608 173216 336660
rect 266636 336608 266688 336660
rect 290280 336608 290332 336660
rect 324320 336608 324372 336660
rect 346400 336608 346452 336660
rect 358084 336608 358136 336660
rect 360108 336608 360160 336660
rect 373080 336608 373132 336660
rect 376760 336608 376812 336660
rect 377036 336608 377088 336660
rect 378968 336608 379020 336660
rect 428464 336608 428516 336660
rect 163504 336540 163556 336592
rect 264428 336540 264480 336592
rect 284300 336540 284352 336592
rect 322480 336540 322532 336592
rect 355876 336540 355928 336592
rect 366456 336540 366508 336592
rect 367560 336540 367612 336592
rect 422944 336540 422996 336592
rect 153844 336472 153896 336524
rect 262220 336472 262272 336524
rect 268384 336472 268436 336524
rect 314108 336472 314160 336524
rect 315028 336472 315080 336524
rect 331956 336472 332008 336524
rect 353760 336472 353812 336524
rect 362132 336472 362184 336524
rect 371148 336472 371200 336524
rect 425796 336472 425848 336524
rect 149704 336404 149756 336456
rect 261116 336404 261168 336456
rect 273628 336404 273680 336456
rect 319260 336404 319312 336456
rect 331220 336404 331272 336456
rect 337108 336404 337160 336456
rect 355784 336404 355836 336456
rect 367652 336404 367704 336456
rect 368664 336404 368716 336456
rect 425704 336404 425756 336456
rect 145564 336336 145616 336388
rect 259000 336336 259052 336388
rect 265624 336336 265676 336388
rect 45560 336268 45612 336320
rect 249064 336268 249116 336320
rect 268568 336268 268620 336320
rect 309600 336268 309652 336320
rect 312544 336336 312596 336388
rect 324688 336336 324740 336388
rect 347688 336336 347740 336388
rect 362316 336336 362368 336388
rect 374184 336336 374236 336388
rect 378968 336336 379020 336388
rect 379612 336336 379664 336388
rect 442264 336336 442316 336388
rect 313004 336268 313056 336320
rect 316408 336268 316460 336320
rect 332692 336268 332744 336320
rect 348608 336268 348660 336320
rect 364984 336268 365036 336320
rect 373172 336268 373224 336320
rect 436744 336268 436796 336320
rect 31760 336200 31812 336252
rect 244740 336200 244792 336252
rect 264244 336200 264296 336252
rect 311900 336200 311952 336252
rect 312728 336200 312780 336252
rect 330576 336200 330628 336252
rect 345296 336200 345348 336252
rect 355416 336200 355468 336252
rect 356888 336200 356940 336252
rect 373356 336200 373408 336252
rect 376668 336200 376720 336252
rect 439504 336200 439556 336252
rect 24860 336132 24912 336184
rect 242532 336132 242584 336184
rect 262864 336132 262916 336184
rect 310796 336132 310848 336184
rect 313280 336132 313332 336184
rect 331588 336132 331640 336184
rect 350356 336132 350408 336184
rect 367836 336132 367888 336184
rect 381820 336132 381872 336184
rect 447784 336132 447836 336184
rect 15200 336064 15252 336116
rect 239588 336064 239640 336116
rect 5540 335996 5592 336048
rect 236644 335996 236696 336048
rect 239404 335996 239456 336048
rect 265532 336064 265584 336116
rect 269396 336064 269448 336116
rect 318156 336064 318208 336116
rect 352564 336064 352616 336116
rect 371884 336064 371936 336116
rect 377496 336064 377548 336116
rect 443644 336064 443696 336116
rect 262220 335996 262272 336048
rect 316040 335996 316092 336048
rect 319444 335996 319496 336048
rect 330208 335996 330260 336048
rect 349988 335996 350040 336048
rect 370504 335996 370556 336048
rect 375288 335996 375340 336048
rect 440884 335996 440936 336048
rect 185584 335928 185636 335980
rect 271052 335928 271104 335980
rect 307024 335928 307076 335980
rect 326528 335928 326580 335980
rect 363236 335928 363288 335980
rect 388444 335928 388496 335980
rect 388536 335928 388588 335980
rect 391204 335928 391256 335980
rect 412548 335928 412600 335980
rect 431224 335928 431276 335980
rect 188344 335860 188396 335912
rect 272156 335860 272208 335912
rect 311256 335860 311308 335912
rect 329472 335860 329524 335912
rect 358820 335860 358872 335912
rect 374644 335860 374696 335912
rect 408408 335860 408460 335912
rect 418896 335860 418948 335912
rect 261576 335792 261628 335844
rect 258816 335724 258868 335776
rect 290188 335724 290240 335776
rect 258724 335656 258776 335708
rect 288900 335656 288952 335708
rect 309600 335792 309652 335844
rect 314844 335792 314896 335844
rect 317420 335792 317472 335844
rect 333060 335792 333112 335844
rect 357164 335792 357216 335844
rect 369124 335792 369176 335844
rect 410340 335792 410392 335844
rect 418804 335792 418856 335844
rect 307116 335724 307168 335776
rect 322112 335724 322164 335776
rect 350816 335724 350868 335776
rect 363604 335724 363656 335776
rect 307484 335656 307536 335708
rect 315304 335656 315356 335708
rect 327080 335656 327132 335708
rect 244924 335588 244976 335640
rect 273260 335588 273312 335640
rect 307208 335588 307260 335640
rect 315212 335588 315264 335640
rect 354864 335588 354916 335640
rect 366272 335724 366324 335776
rect 242164 335520 242216 335572
rect 269948 335520 270000 335572
rect 236644 335452 236696 335504
rect 263324 335452 263376 335504
rect 352656 335452 352708 335504
rect 358176 335452 358228 335504
rect 242256 335384 242308 335436
rect 267832 335384 267884 335436
rect 351828 335384 351880 335436
rect 356704 335384 356756 335436
rect 330208 335316 330260 335368
rect 336740 335316 336792 335368
rect 350448 335316 350500 335368
rect 355324 335316 355376 335368
rect 371976 335316 372028 335368
rect 376024 335316 376076 335368
rect 278964 330760 279016 330812
rect 280252 330760 280304 330812
rect 339684 330760 339736 330812
rect 342444 330760 342496 330812
rect 386604 330760 386656 330812
rect 404452 330760 404504 330812
rect 234620 330624 234672 330676
rect 234804 330624 234856 330676
rect 278964 330556 279016 330608
rect 280252 330556 280304 330608
rect 285680 330556 285732 330608
rect 286048 330556 286100 330608
rect 302240 330556 302292 330608
rect 302608 330556 302660 330608
rect 305000 330556 305052 330608
rect 305368 330556 305420 330608
rect 339684 330556 339736 330608
rect 342444 330556 342496 330608
rect 386604 330556 386656 330608
rect 404452 330556 404504 330608
rect 405740 330556 405792 330608
rect 406844 330556 406896 330608
rect 236092 330488 236144 330540
rect 237012 330488 237064 330540
rect 237472 330488 237524 330540
rect 238484 330488 238536 330540
rect 240140 330488 240192 330540
rect 240692 330488 240744 330540
rect 254032 330488 254084 330540
rect 254952 330488 255004 330540
rect 255504 330488 255556 330540
rect 256424 330488 256476 330540
rect 256700 330488 256752 330540
rect 257160 330488 257212 330540
rect 258172 330488 258224 330540
rect 258632 330488 258684 330540
rect 259644 330488 259696 330540
rect 260380 330488 260432 330540
rect 261024 330488 261076 330540
rect 261852 330488 261904 330540
rect 262404 330488 262456 330540
rect 262956 330488 263008 330540
rect 266544 330488 266596 330540
rect 267372 330488 267424 330540
rect 271972 330488 272024 330540
rect 272800 330488 272852 330540
rect 273352 330488 273404 330540
rect 273904 330488 273956 330540
rect 274640 330488 274692 330540
rect 275744 330488 275796 330540
rect 276112 330488 276164 330540
rect 276848 330488 276900 330540
rect 277584 330488 277636 330540
rect 278320 330488 278372 330540
rect 278872 330488 278924 330540
rect 279424 330488 279476 330540
rect 280344 330488 280396 330540
rect 281264 330488 281316 330540
rect 283104 330488 283156 330540
rect 283748 330488 283800 330540
rect 284392 330488 284444 330540
rect 284852 330488 284904 330540
rect 285772 330488 285824 330540
rect 286324 330488 286376 330540
rect 287060 330488 287112 330540
rect 288164 330488 288216 330540
rect 289912 330488 289964 330540
rect 290372 330488 290424 330540
rect 291292 330488 291344 330540
rect 292212 330488 292264 330540
rect 302332 330488 302384 330540
rect 302792 330488 302844 330540
rect 303712 330488 303764 330540
rect 304632 330488 304684 330540
rect 305092 330488 305144 330540
rect 305736 330488 305788 330540
rect 306472 330488 306524 330540
rect 306840 330488 306892 330540
rect 307852 330488 307904 330540
rect 308588 330488 308640 330540
rect 309324 330488 309376 330540
rect 310060 330488 310112 330540
rect 314844 330488 314896 330540
rect 315580 330488 315632 330540
rect 318892 330488 318944 330540
rect 319904 330488 319956 330540
rect 333980 330488 334032 330540
rect 334532 330488 334584 330540
rect 336832 330488 336884 330540
rect 337844 330488 337896 330540
rect 339592 330488 339644 330540
rect 340052 330488 340104 330540
rect 341064 330488 341116 330540
rect 341524 330488 341576 330540
rect 342352 330488 342404 330540
rect 342996 330488 343048 330540
rect 343640 330488 343692 330540
rect 344744 330488 344796 330540
rect 345020 330488 345072 330540
rect 345848 330488 345900 330540
rect 351920 330488 351972 330540
rect 352840 330488 352892 330540
rect 356060 330488 356112 330540
rect 357256 330488 357308 330540
rect 357532 330488 357584 330540
rect 358268 330488 358320 330540
rect 363052 330488 363104 330540
rect 363788 330488 363840 330540
rect 365812 330488 365864 330540
rect 366364 330488 366416 330540
rect 367100 330488 367152 330540
rect 367744 330488 367796 330540
rect 368572 330488 368624 330540
rect 369216 330488 369268 330540
rect 371240 330488 371292 330540
rect 372160 330488 372212 330540
rect 372804 330488 372856 330540
rect 373264 330488 373316 330540
rect 374000 330488 374052 330540
rect 374736 330488 374788 330540
rect 376852 330488 376904 330540
rect 377680 330488 377732 330540
rect 378324 330488 378376 330540
rect 379152 330488 379204 330540
rect 379520 330488 379572 330540
rect 380532 330488 380584 330540
rect 382280 330488 382332 330540
rect 382740 330488 382792 330540
rect 383752 330488 383804 330540
rect 384580 330488 384632 330540
rect 385040 330488 385092 330540
rect 385684 330488 385736 330540
rect 386512 330488 386564 330540
rect 387524 330488 387576 330540
rect 387800 330488 387852 330540
rect 388628 330488 388680 330540
rect 389180 330488 389232 330540
rect 389732 330488 389784 330540
rect 390836 330488 390888 330540
rect 391480 330488 391532 330540
rect 391940 330488 391992 330540
rect 392952 330488 393004 330540
rect 393504 330488 393556 330540
rect 394424 330488 394476 330540
rect 394700 330488 394752 330540
rect 395160 330488 395212 330540
rect 396172 330488 396224 330540
rect 396632 330488 396684 330540
rect 397460 330488 397512 330540
rect 398472 330488 398524 330540
rect 399024 330488 399076 330540
rect 399944 330488 399996 330540
rect 400220 330488 400272 330540
rect 400680 330488 400732 330540
rect 401692 330488 401744 330540
rect 402152 330488 402204 330540
rect 403164 330488 403216 330540
rect 403900 330488 403952 330540
rect 404544 330488 404596 330540
rect 405372 330488 405424 330540
rect 405924 330488 405976 330540
rect 406108 330488 406160 330540
rect 408500 330488 408552 330540
rect 409420 330488 409472 330540
rect 409880 330488 409932 330540
rect 410524 330488 410576 330540
rect 240232 330420 240284 330472
rect 241060 330420 241112 330472
rect 255320 330420 255372 330472
rect 256056 330420 256108 330472
rect 256792 330420 256844 330472
rect 257528 330420 257580 330472
rect 259460 330420 259512 330472
rect 260012 330420 260064 330472
rect 273444 330420 273496 330472
rect 274272 330420 274324 330472
rect 277400 330420 277452 330472
rect 277952 330420 278004 330472
rect 282920 330420 282972 330472
rect 283380 330420 283432 330472
rect 284484 330420 284536 330472
rect 285220 330420 285272 330472
rect 285864 330420 285916 330472
rect 286692 330420 286744 330472
rect 290004 330420 290056 330472
rect 290740 330420 290792 330472
rect 302424 330420 302476 330472
rect 303160 330420 303212 330472
rect 305184 330420 305236 330472
rect 306104 330420 306156 330472
rect 309140 330420 309192 330472
rect 309692 330420 309744 330472
rect 340972 330420 341024 330472
rect 341892 330420 341944 330472
rect 365720 330420 365772 330472
rect 366732 330420 366784 330472
rect 368664 330420 368716 330472
rect 369584 330420 369636 330472
rect 372620 330420 372672 330472
rect 373632 330420 373684 330472
rect 378140 330420 378192 330472
rect 378784 330420 378836 330472
rect 385132 330420 385184 330472
rect 386052 330420 386104 330472
rect 389272 330420 389324 330472
rect 390100 330420 390152 330472
rect 405832 330420 405884 330472
rect 406476 330420 406528 330472
rect 409972 330420 410024 330472
rect 410892 330420 410944 330472
rect 310704 329944 310756 329996
rect 311532 329944 311584 329996
rect 281540 329808 281592 329860
rect 282368 329808 282420 329860
rect 234804 329400 234856 329452
rect 235540 329400 235592 329452
rect 367284 329400 367336 329452
rect 368112 329400 368164 329452
rect 237380 329264 237432 329316
rect 238116 329264 238168 329316
rect 243084 329128 243136 329180
rect 244004 329128 244056 329180
rect 317604 328924 317656 328976
rect 318524 328924 318576 328976
rect 265072 328788 265124 328840
rect 265900 328788 265952 328840
rect 375380 328720 375432 328772
rect 375840 328720 375892 328772
rect 316316 328584 316368 328636
rect 317052 328584 317104 328636
rect 393320 328448 393372 328500
rect 394056 328448 394108 328500
rect 398840 328448 398892 328500
rect 399576 328448 399628 328500
rect 263692 327496 263744 327548
rect 264060 327496 264112 327548
rect 380992 327428 381044 327480
rect 382004 327428 382056 327480
rect 245844 326816 245896 326868
rect 267832 326816 267884 326868
rect 268476 326816 268528 326868
rect 311992 326816 312044 326868
rect 312636 326816 312688 326868
rect 245844 326612 245896 326664
rect 292672 326408 292724 326460
rect 293684 326408 293736 326460
rect 294052 326408 294104 326460
rect 294788 326408 294840 326460
rect 298284 326408 298336 326460
rect 298468 326408 298520 326460
rect 299572 326408 299624 326460
rect 300584 326408 300636 326460
rect 245752 326340 245804 326392
rect 246212 326340 246264 326392
rect 247040 326340 247092 326392
rect 247960 326340 248012 326392
rect 249892 326340 249944 326392
rect 250904 326340 250956 326392
rect 251180 326340 251232 326392
rect 251640 326340 251692 326392
rect 292580 326340 292632 326392
rect 293316 326340 293368 326392
rect 293960 326340 294012 326392
rect 294420 326340 294472 326392
rect 298100 326340 298152 326392
rect 298744 326340 298796 326392
rect 299480 326340 299532 326392
rect 299848 326340 299900 326392
rect 300952 326340 301004 326392
rect 301688 326340 301740 326392
rect 321652 326340 321704 326392
rect 321836 326340 321888 326392
rect 322940 326340 322992 326392
rect 323584 326340 323636 326392
rect 327172 326340 327224 326392
rect 327632 326340 327684 326392
rect 329932 326340 329984 326392
rect 330944 326340 330996 326392
rect 294144 326272 294196 326324
rect 295156 326272 295208 326324
rect 296720 326136 296772 326188
rect 297640 326136 297692 326188
rect 394792 326068 394844 326120
rect 395528 326068 395580 326120
rect 400312 326068 400364 326120
rect 401048 326068 401100 326120
rect 252652 326000 252704 326052
rect 253112 326000 253164 326052
rect 242900 325728 242952 325780
rect 243636 325728 243688 325780
rect 577320 325456 577372 325508
rect 580724 325456 580776 325508
rect 249800 323824 249852 323876
rect 250536 323824 250588 323876
rect 325792 323552 325844 323604
rect 325976 323552 326028 323604
rect 323124 323212 323176 323264
rect 323952 323212 324004 323264
rect 251272 322192 251324 322244
rect 252008 322192 252060 322244
rect 328460 320832 328512 320884
rect 328644 320832 328696 320884
rect 245660 319200 245712 319252
rect 245936 319200 245988 319252
rect 3332 306280 3384 306332
rect 233608 306280 233660 306332
rect 577412 299412 577464 299464
rect 579620 299412 579672 299464
rect 578148 273164 578200 273216
rect 579620 273164 579672 273216
rect 574836 259360 574888 259412
rect 579804 259360 579856 259412
rect 3148 255212 3200 255264
rect 233792 255212 233844 255264
rect 3516 241408 3568 241460
rect 234160 241408 234212 241460
rect 577964 233180 578016 233232
rect 579620 233180 579672 233232
rect 574744 219376 574796 219428
rect 580172 219376 580224 219428
rect 3424 202784 3476 202836
rect 233976 202784 234028 202836
rect 578056 193128 578108 193180
rect 579620 193128 579672 193180
rect 3424 188980 3476 189032
rect 234252 188980 234304 189032
rect 577780 179324 577832 179376
rect 580080 179324 580132 179376
rect 2780 163752 2832 163804
rect 4896 163752 4948 163804
rect 3424 150356 3476 150408
rect 231216 150356 231268 150408
rect 577596 139340 577648 139392
rect 579620 139340 579672 139392
rect 3240 137912 3292 137964
rect 234068 137912 234120 137964
rect 577872 112956 577924 113008
rect 580540 112956 580592 113008
rect 234344 100648 234396 100700
rect 580172 100648 580224 100700
rect 3424 97928 3476 97980
rect 231124 97928 231176 97980
rect 3148 85484 3200 85536
rect 233884 85484 233936 85536
rect 577688 73108 577740 73160
rect 579712 73108 579764 73160
rect 2780 71612 2832 71664
rect 4804 71612 4856 71664
rect 234436 60664 234488 60716
rect 580172 60664 580224 60716
rect 577504 33056 577556 33108
rect 579620 33056 579672 33108
rect 3424 20612 3476 20664
rect 414940 20612 414992 20664
rect 234528 20544 234580 20596
rect 580172 20544 580224 20596
rect 74540 20272 74592 20324
rect 258264 20272 258316 20324
rect 70400 20204 70452 20256
rect 256884 20204 256936 20256
rect 67640 20136 67692 20188
rect 255596 20136 255648 20188
rect 63500 20068 63552 20120
rect 254216 20068 254268 20120
rect 60740 20000 60792 20052
rect 252836 20000 252888 20052
rect 234712 19932 234764 19984
rect 580264 19932 580316 19984
rect 149060 19252 149112 19304
rect 280436 19252 280488 19304
rect 144920 19184 144972 19236
rect 279056 19184 279108 19236
rect 62120 19116 62172 19168
rect 254124 19116 254176 19168
rect 59360 19048 59412 19100
rect 252652 19048 252704 19100
rect 55220 18980 55272 19032
rect 251272 18980 251324 19032
rect 56600 18912 56652 18964
rect 252744 18912 252796 18964
rect 52460 18844 52512 18896
rect 251364 18844 251416 18896
rect 49700 18776 49752 18828
rect 250076 18776 250128 18828
rect 44180 18708 44232 18760
rect 248604 18708 248656 18760
rect 41420 18640 41472 18692
rect 247224 18640 247276 18692
rect 37280 18572 37332 18624
rect 245936 18572 245988 18624
rect 151820 18504 151872 18556
rect 281724 18504 281776 18556
rect 198740 18436 198792 18488
rect 295524 18436 295576 18488
rect 201500 18368 201552 18420
rect 296996 18368 297048 18420
rect 204260 17892 204312 17944
rect 298284 17892 298336 17944
rect 201592 17824 201644 17876
rect 296904 17824 296956 17876
rect 194600 17756 194652 17808
rect 294144 17756 294196 17808
rect 191840 17688 191892 17740
rect 294236 17688 294288 17740
rect 153200 17620 153252 17672
rect 281540 17620 281592 17672
rect 151912 17552 151964 17604
rect 281632 17552 281684 17604
rect 150440 17484 150492 17536
rect 280344 17484 280396 17536
rect 147680 17416 147732 17468
rect 280160 17416 280212 17468
rect 146300 17348 146352 17400
rect 280252 17348 280304 17400
rect 143540 17280 143592 17332
rect 278872 17280 278924 17332
rect 142160 17212 142212 17264
rect 278964 17212 279016 17264
rect 208400 17144 208452 17196
rect 298376 17144 298428 17196
rect 211160 17076 211212 17128
rect 299756 17076 299808 17128
rect 215300 17008 215352 17060
rect 301044 17008 301096 17060
rect 171968 16532 172020 16584
rect 287336 16532 287388 16584
rect 168380 16464 168432 16516
rect 285864 16464 285916 16516
rect 164424 16396 164476 16448
rect 285956 16396 286008 16448
rect 161296 16328 161348 16380
rect 284668 16328 284720 16380
rect 125600 16260 125652 16312
rect 273536 16260 273588 16312
rect 123024 16192 123076 16244
rect 271972 16192 272024 16244
rect 118700 16124 118752 16176
rect 272064 16124 272116 16176
rect 116400 16056 116452 16108
rect 270684 16056 270736 16108
rect 34520 15988 34572 16040
rect 245844 15988 245896 16040
rect 368664 15988 368716 16040
rect 436744 15988 436796 16040
rect 30840 15920 30892 15972
rect 244372 15920 244424 15972
rect 378416 15920 378468 15972
rect 465172 15920 465224 15972
rect 27712 15852 27764 15904
rect 243176 15852 243228 15904
rect 412824 15852 412876 15904
rect 578608 15852 578660 15904
rect 218060 15784 218112 15836
rect 302516 15784 302568 15836
rect 221096 15716 221148 15768
rect 302424 15716 302476 15768
rect 225144 15648 225196 15700
rect 303896 15648 303948 15700
rect 102232 15104 102284 15156
rect 266452 15104 266504 15156
rect 394884 15104 394936 15156
rect 517888 15104 517940 15156
rect 98184 15036 98236 15088
rect 265164 15036 265216 15088
rect 396264 15036 396316 15088
rect 521660 15036 521712 15088
rect 93860 14968 93912 15020
rect 263692 14968 263744 15020
rect 396356 14968 396408 15020
rect 525432 14968 525484 15020
rect 91560 14900 91612 14952
rect 262404 14900 262456 14952
rect 397736 14900 397788 14952
rect 528560 14900 528612 14952
rect 87512 14832 87564 14884
rect 261024 14832 261076 14884
rect 399116 14832 399168 14884
rect 532056 14832 532108 14884
rect 84200 14764 84252 14816
rect 260932 14764 260984 14816
rect 400404 14764 400456 14816
rect 536104 14764 536156 14816
rect 80888 14696 80940 14748
rect 259736 14696 259788 14748
rect 401784 14696 401836 14748
rect 539600 14696 539652 14748
rect 77392 14628 77444 14680
rect 258172 14628 258224 14680
rect 401876 14628 401928 14680
rect 542728 14628 542780 14680
rect 73344 14560 73396 14612
rect 256792 14560 256844 14612
rect 403256 14560 403308 14612
rect 546500 14560 546552 14612
rect 69848 14492 69900 14544
rect 255504 14492 255556 14544
rect 406016 14492 406068 14544
rect 553768 14492 553820 14544
rect 66720 14424 66772 14476
rect 255412 14424 255464 14476
rect 408776 14424 408828 14476
rect 564440 14424 564492 14476
rect 105728 14356 105780 14408
rect 266544 14356 266596 14408
rect 393596 14356 393648 14408
rect 514760 14356 514812 14408
rect 109040 14288 109092 14340
rect 267832 14288 267884 14340
rect 390836 14288 390888 14340
rect 507216 14288 507268 14340
rect 112352 14220 112404 14272
rect 269304 14220 269356 14272
rect 367284 14220 367336 14272
rect 432052 14220 432104 14272
rect 118792 13744 118844 13796
rect 270776 13744 270828 13796
rect 367192 13744 367244 13796
rect 428464 13744 428516 13796
rect 114744 13676 114796 13728
rect 270592 13676 270644 13728
rect 372804 13676 372856 13728
rect 448520 13676 448572 13728
rect 110420 13608 110472 13660
rect 269212 13608 269264 13660
rect 374092 13608 374144 13660
rect 451648 13608 451700 13660
rect 108120 13540 108172 13592
rect 267924 13540 267976 13592
rect 375472 13540 375524 13592
rect 455696 13540 455748 13592
rect 104072 13472 104124 13524
rect 266636 13472 266688 13524
rect 376944 13472 376996 13524
rect 459192 13472 459244 13524
rect 100760 13404 100812 13456
rect 265072 13404 265124 13456
rect 376852 13404 376904 13456
rect 462320 13404 462372 13456
rect 97448 13336 97500 13388
rect 265256 13336 265308 13388
rect 393504 13336 393556 13388
rect 517152 13336 517204 13388
rect 93952 13268 94004 13320
rect 263784 13268 263836 13320
rect 394792 13268 394844 13320
rect 520280 13268 520332 13320
rect 52552 13200 52604 13252
rect 249892 13200 249944 13252
rect 396172 13200 396224 13252
rect 523776 13200 523828 13252
rect 48504 13132 48556 13184
rect 249984 13132 250036 13184
rect 397644 13132 397696 13184
rect 527824 13132 527876 13184
rect 44272 13064 44324 13116
rect 248512 13064 248564 13116
rect 405924 13064 405976 13116
rect 554780 13064 554832 13116
rect 122288 12996 122340 13048
rect 272156 12996 272208 13048
rect 365996 12996 366048 13048
rect 423680 12996 423732 13048
rect 156144 12928 156196 12980
rect 283196 12928 283248 12980
rect 364524 12928 364576 12980
rect 420920 12928 420972 12980
rect 160100 12860 160152 12912
rect 284576 12860 284628 12912
rect 363052 12860 363104 12912
rect 417424 12860 417476 12912
rect 223580 12384 223632 12436
rect 303804 12384 303856 12436
rect 385316 12384 385368 12436
rect 487160 12384 487212 12436
rect 219992 12316 220044 12368
rect 302332 12316 302384 12368
rect 386604 12316 386656 12368
rect 489920 12316 489972 12368
rect 216864 12248 216916 12300
rect 300952 12248 301004 12300
rect 385132 12248 385184 12300
rect 490012 12248 490064 12300
rect 213368 12180 213420 12232
rect 299572 12180 299624 12232
rect 386696 12180 386748 12232
rect 493048 12180 493100 12232
rect 209780 12112 209832 12164
rect 299664 12112 299716 12164
rect 386512 12112 386564 12164
rect 494704 12112 494756 12164
rect 206192 12044 206244 12096
rect 298192 12044 298244 12096
rect 387984 12044 388036 12096
rect 497096 12044 497148 12096
rect 138848 11976 138900 12028
rect 277676 11976 277728 12028
rect 389456 11976 389508 12028
rect 500592 11976 500644 12028
rect 135260 11908 135312 11960
rect 276296 11908 276348 11960
rect 390744 11908 390796 11960
rect 503720 11908 503772 11960
rect 36728 11840 36780 11892
rect 245752 11840 245804 11892
rect 392216 11840 392268 11892
rect 511264 11840 511316 11892
rect 17960 11772 18012 11824
rect 240416 11772 240468 11824
rect 403164 11772 403216 11824
rect 547880 11772 547932 11824
rect 13544 11704 13596 11756
rect 238852 11704 238904 11756
rect 276020 11704 276072 11756
rect 276756 11704 276808 11756
rect 404636 11704 404688 11756
rect 551008 11704 551060 11756
rect 201500 11636 201552 11688
rect 202696 11636 202748 11688
rect 226340 11636 226392 11688
rect 305276 11636 305328 11688
rect 385224 11636 385276 11688
rect 486424 11636 486476 11688
rect 231032 11568 231084 11620
rect 305184 11568 305236 11620
rect 383936 11568 383988 11620
rect 484032 11568 484084 11620
rect 234620 11500 234672 11552
rect 306564 11500 306616 11552
rect 382464 11500 382516 11552
rect 480536 11500 480588 11552
rect 176660 10956 176712 11008
rect 290096 10956 290148 11008
rect 372712 10956 372764 11008
rect 445760 10956 445812 11008
rect 173900 10888 173952 10940
rect 288532 10888 288584 10940
rect 372620 10888 372672 10940
rect 448612 10888 448664 10940
rect 170312 10820 170364 10872
rect 287244 10820 287296 10872
rect 374000 10820 374052 10872
rect 453304 10820 453356 10872
rect 167184 10752 167236 10804
rect 285772 10752 285824 10804
rect 375380 10752 375432 10804
rect 456892 10752 456944 10804
rect 163412 10684 163464 10736
rect 284484 10684 284536 10736
rect 376760 10684 376812 10736
rect 459928 10684 459980 10736
rect 158904 10616 158956 10668
rect 283104 10616 283156 10668
rect 378232 10616 378284 10668
rect 463976 10616 464028 10668
rect 155408 10548 155460 10600
rect 283012 10548 283064 10600
rect 378324 10548 378376 10600
rect 467472 10548 467524 10600
rect 126980 10480 127032 10532
rect 273444 10480 273496 10532
rect 379704 10480 379756 10532
rect 470600 10480 470652 10532
rect 89904 10412 89956 10464
rect 262312 10412 262364 10464
rect 381084 10412 381136 10464
rect 474096 10412 474148 10464
rect 86408 10344 86460 10396
rect 261116 10344 261168 10396
rect 382372 10344 382424 10396
rect 478144 10344 478196 10396
rect 83280 10276 83332 10328
rect 259644 10276 259696 10328
rect 383844 10276 383896 10328
rect 482376 10276 482428 10328
rect 180984 10208 181036 10260
rect 290004 10208 290056 10260
rect 371424 10208 371476 10260
rect 442172 10208 442224 10260
rect 184940 10140 184992 10192
rect 291476 10140 291528 10192
rect 369952 10140 370004 10192
rect 439136 10140 439188 10192
rect 188252 10072 188304 10124
rect 292856 10072 292908 10124
rect 368572 10072 368624 10124
rect 435088 10072 435140 10124
rect 151728 9596 151780 9648
rect 153016 9596 153068 9648
rect 222752 9596 222804 9648
rect 303620 9596 303672 9648
rect 400312 9596 400364 9648
rect 538404 9596 538456 9648
rect 219256 9528 219308 9580
rect 302240 9528 302292 9580
rect 401692 9528 401744 9580
rect 541992 9528 542044 9580
rect 141240 9460 141292 9512
rect 277584 9460 277636 9512
rect 403072 9460 403124 9512
rect 545488 9460 545540 9512
rect 137652 9392 137704 9444
rect 277492 9392 277544 9444
rect 404452 9392 404504 9444
rect 549076 9392 549128 9444
rect 76196 9324 76248 9376
rect 258356 9324 258408 9376
rect 404544 9324 404596 9376
rect 552664 9324 552716 9376
rect 72608 9256 72660 9308
rect 256700 9256 256752 9308
rect 405832 9256 405884 9308
rect 556160 9256 556212 9308
rect 33600 9188 33652 9240
rect 244464 9188 244516 9240
rect 407212 9188 407264 9240
rect 559748 9188 559800 9240
rect 30104 9120 30156 9172
rect 243084 9120 243136 9172
rect 408684 9120 408736 9172
rect 563244 9120 563296 9172
rect 26516 9052 26568 9104
rect 242992 9052 243044 9104
rect 410064 9052 410116 9104
rect 566832 9052 566884 9104
rect 21824 8984 21876 9036
rect 241612 8984 241664 9036
rect 409972 8984 410024 9036
rect 570328 8984 570380 9036
rect 4068 8916 4120 8968
rect 236184 8916 236236 8968
rect 238116 8916 238168 8968
rect 307944 8916 307996 8968
rect 411444 8916 411496 8968
rect 573916 8916 573968 8968
rect 226432 8848 226484 8900
rect 303712 8848 303764 8900
rect 399024 8848 399076 8900
rect 534908 8848 534960 8900
rect 229836 8780 229888 8832
rect 305092 8780 305144 8832
rect 398932 8780 398984 8832
rect 531320 8780 531372 8832
rect 233424 8712 233476 8764
rect 306472 8712 306524 8764
rect 361856 8712 361908 8764
rect 414296 8712 414348 8764
rect 187332 8236 187384 8288
rect 292764 8236 292816 8288
rect 380992 8236 381044 8288
rect 476948 8236 477000 8288
rect 183744 8168 183796 8220
rect 291384 8168 291436 8220
rect 383660 8168 383712 8220
rect 481732 8168 481784 8220
rect 180248 8100 180300 8152
rect 289912 8100 289964 8152
rect 383752 8100 383804 8152
rect 485228 8100 485280 8152
rect 176752 8032 176804 8084
rect 288624 8032 288676 8084
rect 385040 8032 385092 8084
rect 488816 8032 488868 8084
rect 173072 7964 173124 8016
rect 287060 7964 287112 8016
rect 386420 7964 386472 8016
rect 492312 7964 492364 8016
rect 169576 7896 169628 7948
rect 287152 7896 287204 7948
rect 387892 7896 387944 7948
rect 495900 7896 495952 7948
rect 166080 7828 166132 7880
rect 285680 7828 285732 7880
rect 389364 7828 389416 7880
rect 499396 7828 499448 7880
rect 157800 7760 157852 7812
rect 282920 7760 282972 7812
rect 283656 7760 283708 7812
rect 316316 7760 316368 7812
rect 389272 7760 389324 7812
rect 502984 7760 503036 7812
rect 134156 7692 134208 7744
rect 276204 7692 276256 7744
rect 277492 7692 277544 7744
rect 313464 7692 313516 7744
rect 390652 7692 390704 7744
rect 506480 7692 506532 7744
rect 130568 7624 130620 7676
rect 274824 7624 274876 7676
rect 275192 7624 275244 7676
rect 311992 7624 312044 7676
rect 392124 7624 392176 7676
rect 510068 7624 510120 7676
rect 127072 7556 127124 7608
rect 273352 7556 273404 7608
rect 274548 7556 274600 7608
rect 310704 7556 310756 7608
rect 393412 7556 393464 7608
rect 513564 7556 513616 7608
rect 190828 7488 190880 7540
rect 292672 7488 292724 7540
rect 380900 7488 380952 7540
rect 473452 7488 473504 7540
rect 194416 7420 194468 7472
rect 294052 7420 294104 7472
rect 379612 7420 379664 7472
rect 469864 7420 469916 7472
rect 197912 7352 197964 7404
rect 295432 7352 295484 7404
rect 378140 7352 378192 7404
rect 466276 7352 466328 7404
rect 69112 6808 69164 6860
rect 255320 6808 255372 6860
rect 279516 6808 279568 6860
rect 320272 6808 320324 6860
rect 365720 6808 365772 6860
rect 427268 6808 427320 6860
rect 65524 6740 65576 6792
rect 254032 6740 254084 6792
rect 276020 6740 276072 6792
rect 318892 6740 318944 6792
rect 367100 6740 367152 6792
rect 430856 6740 430908 6792
rect 62028 6672 62080 6724
rect 253940 6672 253992 6724
rect 272432 6672 272484 6724
rect 318984 6672 319036 6724
rect 368480 6672 368532 6724
rect 434444 6672 434496 6724
rect 58440 6604 58492 6656
rect 252560 6604 252612 6656
rect 268844 6604 268896 6656
rect 317696 6604 317748 6656
rect 369860 6604 369912 6656
rect 437940 6604 437992 6656
rect 54944 6536 54996 6588
rect 251180 6536 251232 6588
rect 265348 6536 265400 6588
rect 316224 6536 316276 6588
rect 371332 6536 371384 6588
rect 441528 6536 441580 6588
rect 51356 6468 51408 6520
rect 249800 6468 249852 6520
rect 261760 6468 261812 6520
rect 314844 6468 314896 6520
rect 371240 6468 371292 6520
rect 445024 6468 445076 6520
rect 47860 6400 47912 6452
rect 248696 6400 248748 6452
rect 258264 6400 258316 6452
rect 314752 6400 314804 6452
rect 407120 6400 407172 6452
rect 558552 6400 558604 6452
rect 12348 6332 12400 6384
rect 237472 6332 237524 6384
rect 254676 6332 254728 6384
rect 313372 6332 313424 6384
rect 408592 6332 408644 6384
rect 562048 6332 562100 6384
rect 7656 6264 7708 6316
rect 236092 6264 236144 6316
rect 239312 6264 239364 6316
rect 307852 6264 307904 6316
rect 365812 6264 365864 6316
rect 391848 6264 391900 6316
rect 408500 6264 408552 6316
rect 565636 6264 565688 6316
rect 2872 6196 2924 6248
rect 234804 6196 234856 6248
rect 240508 6196 240560 6248
rect 309416 6196 309468 6248
rect 360292 6196 360344 6248
rect 407212 6196 407264 6248
rect 409880 6196 409932 6248
rect 569132 6196 569184 6248
rect 1676 6128 1728 6180
rect 234896 6128 234948 6180
rect 237012 6128 237064 6180
rect 307760 6128 307812 6180
rect 360384 6128 360436 6180
rect 409604 6128 409656 6180
rect 412640 6128 412692 6180
rect 576308 6128 576360 6180
rect 140044 6060 140096 6112
rect 277400 6060 277452 6112
rect 286600 6060 286652 6112
rect 323216 6060 323268 6112
rect 365904 6060 365956 6112
rect 423772 6060 423824 6112
rect 143632 5992 143684 6044
rect 278780 5992 278832 6044
rect 299296 5992 299348 6044
rect 310612 5992 310664 6044
rect 364432 5992 364484 6044
rect 420184 5992 420236 6044
rect 232228 5924 232280 5976
rect 306656 5924 306708 5976
rect 362960 5924 363012 5976
rect 416688 5924 416740 5976
rect 235816 5856 235868 5908
rect 261484 5856 261536 5908
rect 361764 5856 361816 5908
rect 413100 5856 413152 5908
rect 361672 5788 361724 5840
rect 410800 5788 410852 5840
rect 85672 5448 85724 5500
rect 149704 5448 149756 5500
rect 210976 5448 211028 5500
rect 299480 5448 299532 5500
rect 364340 5448 364392 5500
rect 384948 5448 385000 5500
rect 390560 5448 390612 5500
rect 505376 5448 505428 5500
rect 89168 5380 89220 5432
rect 153844 5380 153896 5432
rect 207388 5380 207440 5432
rect 298100 5380 298152 5432
rect 301504 5380 301556 5432
rect 312084 5380 312136 5432
rect 361580 5380 361632 5432
rect 382280 5380 382332 5432
rect 392032 5380 392084 5432
rect 508872 5380 508924 5432
rect 110512 5312 110564 5364
rect 177304 5312 177356 5364
rect 203892 5312 203944 5364
rect 296720 5312 296772 5364
rect 297180 5312 297232 5364
rect 310796 5312 310848 5364
rect 352012 5312 352064 5364
rect 378876 5312 378928 5364
rect 391940 5312 391992 5364
rect 512460 5312 512512 5364
rect 78588 5244 78640 5296
rect 145564 5244 145616 5296
rect 196808 5244 196860 5296
rect 295340 5244 295392 5296
rect 303160 5244 303212 5296
rect 328644 5244 328696 5296
rect 351920 5244 351972 5296
rect 382372 5244 382424 5296
rect 393320 5244 393372 5296
rect 515956 5244 516008 5296
rect 117596 5176 117648 5228
rect 185584 5176 185636 5228
rect 193220 5176 193272 5228
rect 293960 5176 294012 5228
rect 294052 5176 294104 5228
rect 321652 5176 321704 5228
rect 353392 5176 353444 5228
rect 385960 5176 386012 5228
rect 394700 5176 394752 5228
rect 519544 5176 519596 5228
rect 121092 5108 121144 5160
rect 188344 5108 188396 5160
rect 189724 5108 189776 5160
rect 292580 5108 292632 5160
rect 299664 5108 299716 5160
rect 327264 5108 327316 5160
rect 353484 5108 353536 5160
rect 387156 5108 387208 5160
rect 396080 5108 396132 5160
rect 523040 5108 523092 5160
rect 96252 5040 96304 5092
rect 163504 5040 163556 5092
rect 186136 5040 186188 5092
rect 291292 5040 291344 5092
rect 296076 5040 296128 5092
rect 325792 5040 325844 5092
rect 354680 5040 354732 5092
rect 389456 5040 389508 5092
rect 397552 5040 397604 5092
rect 526628 5040 526680 5092
rect 103336 4972 103388 5024
rect 173164 4972 173216 5024
rect 182548 4972 182600 5024
rect 291200 4972 291252 5024
rect 292580 4972 292632 5024
rect 324504 4972 324556 5024
rect 356152 4972 356204 5024
rect 393044 4972 393096 5024
rect 398840 4972 398892 5024
rect 533712 4972 533764 5024
rect 146944 4904 146996 4956
rect 276112 4904 276164 4956
rect 285404 4904 285456 4956
rect 323032 4904 323084 4956
rect 356060 4904 356112 4956
rect 396540 4904 396592 4956
rect 400220 4904 400272 4956
rect 537208 4904 537260 4956
rect 132960 4836 133012 4888
rect 274640 4836 274692 4888
rect 278320 4836 278372 4888
rect 320180 4836 320232 4888
rect 357624 4836 357676 4888
rect 398932 4836 398984 4888
rect 401600 4836 401652 4888
rect 540796 4836 540848 4888
rect 129372 4768 129424 4820
rect 274732 4768 274784 4820
rect 274824 4768 274876 4820
rect 319076 4768 319128 4820
rect 357532 4768 357584 4820
rect 400128 4768 400180 4820
rect 402980 4768 403032 4820
rect 544384 4768 544436 4820
rect 136456 4700 136508 4752
rect 146944 4700 146996 4752
rect 214472 4700 214524 4752
rect 300860 4700 300912 4752
rect 389180 4700 389232 4752
rect 501788 4700 501840 4752
rect 175464 4632 175516 4684
rect 258724 4632 258776 4684
rect 264152 4632 264204 4684
rect 316132 4632 316184 4684
rect 387800 4632 387852 4684
rect 498200 4632 498252 4684
rect 179052 4564 179104 4616
rect 258816 4564 258868 4616
rect 288992 4564 289044 4616
rect 323124 4564 323176 4616
rect 360200 4564 360252 4616
rect 406016 4564 406068 4616
rect 291844 4496 291896 4548
rect 317604 4496 317656 4548
rect 358912 4496 358964 4548
rect 403624 4496 403676 4548
rect 291752 4428 291804 4480
rect 317512 4428 317564 4480
rect 358820 4428 358872 4480
rect 402520 4428 402572 4480
rect 126980 4156 127032 4208
rect 128176 4156 128228 4208
rect 176660 4156 176712 4208
rect 177856 4156 177908 4208
rect 226340 4156 226392 4208
rect 227536 4156 227588 4208
rect 361764 4156 361816 4208
rect 99840 4088 99892 4140
rect 239404 4088 239456 4140
rect 246396 4088 246448 4140
rect 262864 4088 262916 4140
rect 271236 4088 271288 4140
rect 291844 4088 291896 4140
rect 298468 4088 298520 4140
rect 315304 4088 315356 4140
rect 320916 4088 320968 4140
rect 92756 4020 92808 4072
rect 236644 4020 236696 4072
rect 255872 4020 255924 4072
rect 277492 4020 277544 4072
rect 283104 4020 283156 4072
rect 307116 4020 307168 4072
rect 316224 4020 316276 4072
rect 331404 4020 331456 4072
rect 333888 4088 333940 4140
rect 336832 4088 336884 4140
rect 346492 4088 346544 4140
rect 361856 4088 361908 4140
rect 334072 4020 334124 4072
rect 343824 4020 343876 4072
rect 354036 4020 354088 4072
rect 358176 4020 358228 4072
rect 362316 4088 362368 4140
rect 364340 4088 364392 4140
rect 364984 4088 365036 4140
rect 368204 4088 368256 4140
rect 382280 4088 382332 4140
rect 411904 4088 411956 4140
rect 418804 4088 418856 4140
rect 419080 4088 419132 4140
rect 425796 4088 425848 4140
rect 440332 4088 440384 4140
rect 442264 4088 442316 4140
rect 442724 4088 442776 4140
rect 447784 4088 447836 4140
rect 475752 4088 475804 4140
rect 82084 3952 82136 4004
rect 259460 3952 259512 4004
rect 267740 3952 267792 4004
rect 291752 3952 291804 4004
rect 294880 3952 294932 4004
rect 325884 3952 325936 4004
rect 345112 3952 345164 4004
rect 358728 3952 358780 4004
rect 377680 4020 377732 4072
rect 379520 4020 379572 4072
rect 472256 4020 472308 4072
rect 381176 3952 381228 4004
rect 382464 3952 382516 4004
rect 479340 3952 479392 4004
rect 43076 3884 43128 3936
rect 247040 3884 247092 3936
rect 252376 3884 252428 3936
rect 275192 3884 275244 3936
rect 287796 3884 287848 3936
rect 322940 3884 322992 3936
rect 325608 3884 325660 3936
rect 335360 3884 335412 3936
rect 340972 3884 341024 3936
rect 346952 3884 347004 3936
rect 347872 3884 347924 3936
rect 359464 3884 359516 3936
rect 35992 3816 36044 3868
rect 245660 3816 245712 3868
rect 248788 3816 248840 3868
rect 274548 3816 274600 3868
rect 280712 3816 280764 3868
rect 321744 3816 321796 3868
rect 326804 3816 326856 3868
rect 335452 3816 335504 3868
rect 343916 3816 343968 3868
rect 355232 3816 355284 3868
rect 356704 3816 356756 3868
rect 361764 3884 361816 3936
rect 361856 3884 361908 3936
rect 363512 3884 363564 3936
rect 367744 3884 367796 3936
rect 390652 3884 390704 3936
rect 391204 3884 391256 3936
rect 422576 3884 422628 3936
rect 428556 3884 428608 3936
rect 450912 3884 450964 3936
rect 454684 3884 454736 3936
rect 583392 3884 583444 3936
rect 361488 3816 361540 3868
rect 374092 3816 374144 3868
rect 376024 3816 376076 3868
rect 443828 3816 443880 3868
rect 450544 3816 450596 3868
rect 581000 3816 581052 3868
rect 28908 3748 28960 3800
rect 242900 3748 242952 3800
rect 260656 3748 260708 3800
rect 307208 3748 307260 3800
rect 311440 3748 311492 3800
rect 329932 3748 329984 3800
rect 347964 3748 348016 3800
rect 369400 3748 369452 3800
rect 369492 3748 369544 3800
rect 375288 3748 375340 3800
rect 377404 3748 377456 3800
rect 408408 3748 408460 3800
rect 418896 3748 418948 3800
rect 560852 3748 560904 3800
rect 24216 3680 24268 3732
rect 241796 3680 241848 3732
rect 247592 3680 247644 3732
rect 297180 3680 297232 3732
rect 310244 3680 310296 3732
rect 312636 3680 312688 3732
rect 312728 3680 312780 3732
rect 330024 3680 330076 3732
rect 335084 3680 335136 3732
rect 338120 3680 338172 3732
rect 341064 3680 341116 3732
rect 345756 3680 345808 3732
rect 347780 3680 347832 3732
rect 365812 3680 365864 3732
rect 366456 3680 366508 3732
rect 391848 3680 391900 3732
rect 391940 3680 391992 3732
rect 426164 3680 426216 3732
rect 431224 3680 431276 3732
rect 575112 3680 575164 3732
rect 19432 3612 19484 3664
rect 240140 3612 240192 3664
rect 251180 3612 251232 3664
rect 301504 3612 301556 3664
rect 305552 3612 305604 3664
rect 328736 3612 328788 3664
rect 349160 3612 349212 3664
rect 370596 3612 370648 3664
rect 374644 3612 374696 3664
rect 401324 3612 401376 3664
rect 404360 3612 404412 3664
rect 550272 3612 550324 3664
rect 20628 3544 20680 3596
rect 240232 3544 240284 3596
rect 244096 3544 244148 3596
rect 297732 3544 297784 3596
rect 304356 3544 304408 3596
rect 328552 3544 328604 3596
rect 332692 3544 332744 3596
rect 336924 3544 336976 3596
rect 350540 3544 350592 3596
rect 376484 3544 376536 3596
rect 384948 3544 385000 3596
rect 418988 3544 419040 3596
rect 419080 3544 419132 3596
rect 568028 3544 568080 3596
rect 14740 3476 14792 3528
rect 238944 3476 238996 3528
rect 245200 3476 245252 3528
rect 299296 3476 299348 3528
rect 301964 3476 302016 3528
rect 327356 3476 327408 3528
rect 343732 3476 343784 3528
rect 352840 3476 352892 3528
rect 353300 3476 353352 3528
rect 383568 3476 383620 3528
rect 405740 3476 405792 3528
rect 557356 3476 557408 3528
rect 11152 3408 11204 3460
rect 237380 3408 237432 3460
rect 242900 3408 242952 3460
rect 44180 3340 44232 3392
rect 45100 3340 45152 3392
rect 52460 3340 52512 3392
rect 53380 3340 53432 3392
rect 93860 3340 93912 3392
rect 94780 3340 94832 3392
rect 110420 3340 110472 3392
rect 111616 3340 111668 3392
rect 106924 3272 106976 3324
rect 242256 3340 242308 3392
rect 249984 3340 250036 3392
rect 264244 3340 264296 3392
rect 266544 3340 266596 3392
rect 283656 3340 283708 3392
rect 291384 3340 291436 3392
rect 306748 3408 306800 3460
rect 311164 3408 311216 3460
rect 312636 3408 312688 3460
rect 331312 3408 331364 3460
rect 337476 3408 337528 3460
rect 338304 3408 338356 3460
rect 343640 3408 343692 3460
rect 356336 3408 356388 3460
rect 359464 3408 359516 3460
rect 367008 3408 367060 3460
rect 118700 3272 118752 3324
rect 119896 3272 119948 3324
rect 114008 3204 114060 3256
rect 242164 3272 242216 3324
rect 253480 3272 253532 3324
rect 265624 3272 265676 3324
rect 293684 3272 293736 3324
rect 305644 3272 305696 3324
rect 124680 3204 124732 3256
rect 244924 3204 244976 3256
rect 257068 3204 257120 3256
rect 268384 3204 268436 3256
rect 281908 3204 281960 3256
rect 294052 3204 294104 3256
rect 143540 3136 143592 3188
rect 144736 3136 144788 3188
rect 259460 3136 259512 3188
rect 268476 3136 268528 3188
rect 307944 3340 307996 3392
rect 312728 3340 312780 3392
rect 319720 3340 319772 3392
rect 332876 3340 332928 3392
rect 342536 3340 342588 3392
rect 309048 3272 309100 3324
rect 319444 3272 319496 3324
rect 323308 3272 323360 3324
rect 333980 3272 334032 3324
rect 336280 3272 336332 3324
rect 338212 3272 338264 3324
rect 338672 3272 338724 3324
rect 339684 3272 339736 3324
rect 342260 3272 342312 3324
rect 309140 3204 309192 3256
rect 324412 3204 324464 3256
rect 334256 3204 334308 3256
rect 312544 3136 312596 3188
rect 328000 3136 328052 3188
rect 335544 3136 335596 3188
rect 339592 3136 339644 3188
rect 340972 3136 341024 3188
rect 341156 3136 341208 3188
rect 344560 3136 344612 3188
rect 346400 3340 346452 3392
rect 345020 3272 345072 3324
rect 351644 3204 351696 3256
rect 349252 3136 349304 3188
rect 297272 3068 297324 3120
rect 307024 3068 307076 3120
rect 322112 3068 322164 3120
rect 334164 3068 334216 3120
rect 342444 3068 342496 3120
rect 348056 3068 348108 3120
rect 329196 3000 329248 3052
rect 335636 3000 335688 3052
rect 341248 3000 341300 3052
rect 343364 3000 343416 3052
rect 342352 2932 342404 2984
rect 350448 3000 350500 3052
rect 355416 3340 355468 3392
rect 357532 3340 357584 3392
rect 363604 3340 363656 3392
rect 369492 3408 369544 3460
rect 370504 3408 370556 3460
rect 371700 3408 371752 3460
rect 371792 3408 371844 3460
rect 397736 3408 397788 3460
rect 411260 3408 411312 3460
rect 571524 3408 571576 3460
rect 369216 3340 369268 3392
rect 362224 3272 362276 3324
rect 371976 3340 372028 3392
rect 388260 3340 388312 3392
rect 388444 3340 388496 3392
rect 415492 3340 415544 3392
rect 423680 3340 423732 3392
rect 424968 3340 425020 3392
rect 448612 3340 448664 3392
rect 449808 3340 449860 3392
rect 362316 3204 362368 3256
rect 395344 3272 395396 3324
rect 442724 3272 442776 3324
rect 468668 3340 468720 3392
rect 489920 3340 489972 3392
rect 490748 3340 490800 3392
rect 449992 3272 450044 3324
rect 461584 3272 461636 3324
rect 384764 3204 384816 3256
rect 439504 3204 439556 3256
rect 458088 3204 458140 3256
rect 355324 3136 355376 3188
rect 361488 3136 361540 3188
rect 357440 3068 357492 3120
rect 371792 3136 371844 3188
rect 371884 3136 371936 3188
rect 367836 3068 367888 3120
rect 372896 3068 372948 3120
rect 373356 3136 373408 3188
rect 394240 3136 394292 3188
rect 422944 3136 422996 3188
rect 429660 3136 429712 3188
rect 440884 3136 440936 3188
rect 454500 3136 454552 3188
rect 379980 3068 380032 3120
rect 436836 3068 436888 3120
rect 447416 3068 447468 3120
rect 358084 3000 358136 3052
rect 361120 3000 361172 3052
rect 425704 3000 425756 3052
rect 433248 3000 433300 3052
rect 443644 3000 443696 3052
rect 449992 3000 450044 3052
rect 359924 2932 359976 2984
rect 366364 2932 366416 2984
rect 371976 2932 372028 2984
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40052 703582 40356 703610
rect 8128 700330 8156 703520
rect 24320 700398 24348 703520
rect 24308 700392 24360 700398
rect 24308 700334 24360 700340
rect 8116 700324 8168 700330
rect 8116 700266 8168 700272
rect 3422 684312 3478 684321
rect 3422 684247 3478 684256
rect 3436 683194 3464 684247
rect 3424 683188 3476 683194
rect 3424 683130 3476 683136
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 40052 461650 40080 703582
rect 40328 703474 40356 703582
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 104912 703582 105308 703610
rect 40512 703474 40540 703520
rect 40328 703446 40540 703474
rect 72988 700466 73016 703520
rect 89180 700534 89208 703520
rect 89168 700528 89220 700534
rect 89168 700470 89220 700476
rect 72976 700460 73028 700466
rect 72976 700402 73028 700408
rect 104912 461786 104940 703582
rect 105280 703474 105308 703582
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 234632 703582 235028 703610
rect 105464 703474 105492 703520
rect 105280 703446 105492 703474
rect 137848 700738 137876 703520
rect 154132 700806 154160 703520
rect 170324 702434 170352 703520
rect 169772 702406 170352 702434
rect 154120 700800 154172 700806
rect 154120 700742 154172 700748
rect 137836 700732 137888 700738
rect 137836 700674 137888 700680
rect 169772 461922 169800 702406
rect 202800 700670 202828 703520
rect 218992 700942 219020 703520
rect 218980 700936 219032 700942
rect 218980 700878 219032 700884
rect 202788 700664 202840 700670
rect 202788 700606 202840 700612
rect 234632 462126 234660 703582
rect 235000 703474 235028 703582
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 299492 703582 299980 703610
rect 235184 703474 235212 703520
rect 235000 703446 235212 703474
rect 267660 700194 267688 703520
rect 283852 702434 283880 703520
rect 282932 702406 283880 702434
rect 267648 700188 267700 700194
rect 267648 700130 267700 700136
rect 252652 478916 252704 478922
rect 252652 478858 252704 478864
rect 234620 462120 234672 462126
rect 234620 462062 234672 462068
rect 169760 461916 169812 461922
rect 169760 461858 169812 461864
rect 104900 461780 104952 461786
rect 104900 461722 104952 461728
rect 40040 461644 40092 461650
rect 40040 461586 40092 461592
rect 3884 460692 3936 460698
rect 3884 460634 3936 460640
rect 3608 460624 3660 460630
rect 3608 460566 3660 460572
rect 3332 459808 3384 459814
rect 3332 459750 3384 459756
rect 3240 458584 3292 458590
rect 3240 458526 3292 458532
rect 2780 449880 2832 449886
rect 2780 449822 2832 449828
rect 2792 449585 2820 449822
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 3252 423609 3280 458526
rect 3238 423600 3294 423609
rect 3238 423535 3294 423544
rect 3344 410553 3372 459750
rect 3516 458380 3568 458386
rect 3516 458322 3568 458328
rect 3424 458312 3476 458318
rect 3424 458254 3476 458260
rect 3330 410544 3386 410553
rect 3330 410479 3386 410488
rect 3332 306332 3384 306338
rect 3332 306274 3384 306280
rect 3344 306241 3372 306274
rect 3330 306232 3386 306241
rect 3330 306167 3386 306176
rect 3148 255264 3200 255270
rect 3148 255206 3200 255212
rect 3160 254153 3188 255206
rect 3146 254144 3202 254153
rect 3146 254079 3202 254088
rect 3436 214985 3464 458254
rect 3528 267209 3556 458322
rect 3620 293185 3648 460566
rect 3792 459740 3844 459746
rect 3792 459682 3844 459688
rect 3700 458448 3752 458454
rect 3700 458390 3752 458396
rect 3712 319297 3740 458390
rect 3804 345409 3832 459682
rect 3896 358465 3924 460634
rect 237286 460456 237342 460465
rect 237286 460391 237342 460400
rect 234344 459944 234396 459950
rect 234344 459886 234396 459892
rect 4988 459876 5040 459882
rect 4988 459818 5040 459824
rect 3976 458516 4028 458522
rect 3976 458458 4028 458464
rect 3988 371385 4016 458458
rect 4802 458280 4858 458289
rect 4802 458215 4858 458224
rect 4896 458244 4948 458250
rect 4068 457496 4120 457502
rect 4068 457438 4120 457444
rect 4080 397497 4108 457438
rect 4066 397488 4122 397497
rect 4066 397423 4122 397432
rect 3974 371376 4030 371385
rect 3974 371311 4030 371320
rect 3882 358456 3938 358465
rect 3882 358391 3938 358400
rect 3790 345400 3846 345409
rect 3790 345335 3846 345344
rect 3698 319288 3754 319297
rect 3698 319223 3754 319232
rect 3606 293176 3662 293185
rect 3606 293111 3662 293120
rect 3514 267200 3570 267209
rect 3514 267135 3570 267144
rect 3516 241460 3568 241466
rect 3516 241402 3568 241408
rect 3528 241097 3556 241402
rect 3514 241088 3570 241097
rect 3514 241023 3570 241032
rect 3422 214976 3478 214985
rect 3422 214911 3478 214920
rect 3424 202836 3476 202842
rect 3424 202778 3476 202784
rect 3436 201929 3464 202778
rect 3422 201920 3478 201929
rect 3422 201855 3478 201864
rect 3424 189032 3476 189038
rect 3424 188974 3476 188980
rect 3436 188873 3464 188974
rect 3422 188864 3478 188873
rect 3422 188799 3478 188808
rect 2780 163804 2832 163810
rect 2780 163746 2832 163752
rect 2792 162897 2820 163746
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 3424 150408 3476 150414
rect 3424 150350 3476 150356
rect 3436 149841 3464 150350
rect 3422 149832 3478 149841
rect 3422 149767 3478 149776
rect 3240 137964 3292 137970
rect 3240 137906 3292 137912
rect 3252 136785 3280 137906
rect 3238 136776 3294 136785
rect 3238 136711 3294 136720
rect 3424 97980 3476 97986
rect 3424 97922 3476 97928
rect 3436 97617 3464 97922
rect 3422 97608 3478 97617
rect 3422 97543 3478 97552
rect 3148 85536 3200 85542
rect 3148 85478 3200 85484
rect 3160 84697 3188 85478
rect 3146 84688 3202 84697
rect 3146 84623 3202 84632
rect 4816 71670 4844 458215
rect 4896 458186 4948 458192
rect 4908 163810 4936 458186
rect 5000 449886 5028 459818
rect 231216 459196 231268 459202
rect 231216 459138 231268 459144
rect 231124 459128 231176 459134
rect 231124 459070 231176 459076
rect 4988 449880 5040 449886
rect 4988 449822 5040 449828
rect 177304 336728 177356 336734
rect 177304 336670 177356 336676
rect 173164 336660 173216 336666
rect 173164 336602 173216 336608
rect 163504 336592 163556 336598
rect 163504 336534 163556 336540
rect 153844 336524 153896 336530
rect 153844 336466 153896 336472
rect 149704 336456 149756 336462
rect 149704 336398 149756 336404
rect 145564 336388 145616 336394
rect 145564 336330 145616 336336
rect 45560 336320 45612 336326
rect 45560 336262 45612 336268
rect 31760 336252 31812 336258
rect 31760 336194 31812 336200
rect 24860 336184 24912 336190
rect 24860 336126 24912 336132
rect 15200 336116 15252 336122
rect 15200 336058 15252 336064
rect 5540 336048 5592 336054
rect 5540 335990 5592 335996
rect 4896 163804 4948 163810
rect 4896 163746 4948 163752
rect 2780 71664 2832 71670
rect 2778 71632 2780 71641
rect 4804 71664 4856 71670
rect 2832 71632 2834 71641
rect 4804 71606 4856 71612
rect 2778 71567 2834 71576
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3514 19952 3570 19961
rect 3514 19887 3570 19896
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 110 15872 166 15881
rect 110 15807 166 15816
rect 124 354 152 15807
rect 3528 6914 3556 19887
rect 5552 16574 5580 335990
rect 9678 18592 9734 18601
rect 9678 18527 9734 18536
rect 5552 16546 6040 16574
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3436 6886 3556 6914
rect 3436 6497 3464 6886
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 6248 2924 6254
rect 2872 6190 2924 6196
rect 1676 6180 1728 6186
rect 1676 6122 1728 6128
rect 1688 480 1716 6122
rect 2884 480 2912 6190
rect 4080 480 4108 8910
rect 5262 3360 5318 3369
rect 5262 3295 5318 3304
rect 5276 480 5304 3295
rect 542 354 654 480
rect 124 326 654 354
rect 542 -960 654 326
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6012 354 6040 16546
rect 8758 11656 8814 11665
rect 8758 11591 8814 11600
rect 7656 6316 7708 6322
rect 7656 6258 7708 6264
rect 7668 480 7696 6258
rect 8772 480 8800 11591
rect 6430 354 6542 480
rect 6012 326 6542 354
rect 6430 -960 6542 326
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9692 354 9720 18527
rect 15212 16574 15240 336058
rect 24872 16574 24900 336126
rect 31772 16574 31800 336194
rect 38658 336016 38714 336025
rect 38658 335951 38714 335960
rect 37280 18624 37332 18630
rect 37280 18566 37332 18572
rect 37292 16574 37320 18566
rect 38672 16574 38700 335951
rect 44180 18760 44232 18766
rect 44180 18702 44232 18708
rect 41420 18692 41472 18698
rect 41420 18634 41472 18640
rect 41432 16574 41460 18634
rect 15212 16546 15976 16574
rect 24872 16546 25360 16574
rect 31772 16546 31984 16574
rect 37292 16546 38424 16574
rect 38672 16546 39160 16574
rect 41432 16546 41920 16574
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 11152 3460 11204 3466
rect 11152 3402 11204 3408
rect 11164 480 11192 3402
rect 12360 480 12388 6326
rect 13556 480 13584 11698
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14752 480 14780 3470
rect 15948 480 15976 16546
rect 22558 14512 22614 14521
rect 22558 14447 22614 14456
rect 17960 11824 18012 11830
rect 17960 11766 18012 11772
rect 17038 8936 17094 8945
rect 17038 8871 17094 8880
rect 17052 480 17080 8871
rect 9926 354 10038 480
rect 9692 326 10038 354
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 17972 354 18000 11766
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 19432 3664 19484 3670
rect 19432 3606 19484 3612
rect 19444 480 19472 3606
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20640 480 20668 3538
rect 21836 480 21864 8978
rect 18206 354 18318 480
rect 17972 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22572 354 22600 14447
rect 24216 3732 24268 3738
rect 24216 3674 24268 3680
rect 24228 480 24256 3674
rect 25332 480 25360 16546
rect 30840 15972 30892 15978
rect 30840 15914 30892 15920
rect 27712 15904 27764 15910
rect 27712 15846 27764 15852
rect 26516 9104 26568 9110
rect 26516 9046 26568 9052
rect 26528 480 26556 9046
rect 27724 480 27752 15846
rect 30104 9172 30156 9178
rect 30104 9114 30156 9120
rect 28908 3800 28960 3806
rect 28908 3742 28960 3748
rect 28920 480 28948 3742
rect 30116 480 30144 9114
rect 22990 354 23102 480
rect 22572 326 23102 354
rect 22990 -960 23102 326
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 30852 354 30880 15914
rect 31270 354 31382 480
rect 30852 326 31382 354
rect 31956 354 31984 16546
rect 34520 16040 34572 16046
rect 34520 15982 34572 15988
rect 33600 9240 33652 9246
rect 33600 9182 33652 9188
rect 33612 480 33640 9182
rect 32374 354 32486 480
rect 31956 326 32486 354
rect 31270 -960 31382 326
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34532 354 34560 15982
rect 36728 11892 36780 11898
rect 36728 11834 36780 11840
rect 35992 3868 36044 3874
rect 35992 3810 36044 3816
rect 36004 480 36032 3810
rect 34766 354 34878 480
rect 34532 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36740 354 36768 11834
rect 38396 480 38424 16546
rect 37158 354 37270 480
rect 36740 326 37270 354
rect 37158 -960 37270 326
rect 38354 -960 38466 480
rect 39132 354 39160 16546
rect 40222 13016 40278 13025
rect 40222 12951 40278 12960
rect 39550 354 39662 480
rect 39132 326 39662 354
rect 40236 354 40264 12951
rect 41892 480 41920 16546
rect 43076 3936 43128 3942
rect 43076 3878 43128 3884
rect 43088 480 43116 3878
rect 44192 3398 44220 18702
rect 45572 16574 45600 336262
rect 74540 20324 74592 20330
rect 74540 20266 74592 20272
rect 70400 20256 70452 20262
rect 70400 20198 70452 20204
rect 67640 20188 67692 20194
rect 67640 20130 67692 20136
rect 63500 20120 63552 20126
rect 63500 20062 63552 20068
rect 60740 20052 60792 20058
rect 60740 19994 60792 20000
rect 59360 19100 59412 19106
rect 59360 19042 59412 19048
rect 55220 19032 55272 19038
rect 55220 18974 55272 18980
rect 52460 18896 52512 18902
rect 52460 18838 52512 18844
rect 49700 18828 49752 18834
rect 49700 18770 49752 18776
rect 49712 16574 49740 18770
rect 45572 16546 46704 16574
rect 49712 16546 50200 16574
rect 44272 13116 44324 13122
rect 44272 13058 44324 13064
rect 44180 3392 44232 3398
rect 44180 3334 44232 3340
rect 44284 480 44312 13058
rect 45100 3392 45152 3398
rect 45100 3334 45152 3340
rect 40654 354 40766 480
rect 40236 326 40766 354
rect 39550 -960 39662 326
rect 40654 -960 40766 326
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45112 354 45140 3334
rect 46676 480 46704 16546
rect 48504 13184 48556 13190
rect 48504 13126 48556 13132
rect 47860 6452 47912 6458
rect 47860 6394 47912 6400
rect 47872 480 47900 6394
rect 45438 354 45550 480
rect 45112 326 45550 354
rect 45438 -960 45550 326
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48516 354 48544 13126
rect 50172 480 50200 16546
rect 51356 6520 51408 6526
rect 51356 6462 51408 6468
rect 51368 480 51396 6462
rect 52472 3398 52500 18838
rect 55232 16574 55260 18974
rect 56600 18964 56652 18970
rect 56600 18906 56652 18912
rect 56612 16574 56640 18906
rect 55232 16546 56088 16574
rect 56612 16546 56824 16574
rect 52552 13252 52604 13258
rect 52552 13194 52604 13200
rect 52460 3392 52512 3398
rect 52460 3334 52512 3340
rect 52564 480 52592 13194
rect 54944 6588 54996 6594
rect 54944 6530 54996 6536
rect 53380 3392 53432 3398
rect 53380 3334 53432 3340
rect 48934 354 49046 480
rect 48516 326 49046 354
rect 48934 -960 49046 326
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53392 354 53420 3334
rect 54956 480 54984 6530
rect 56060 480 56088 16546
rect 53718 354 53830 480
rect 53392 326 53830 354
rect 53718 -960 53830 326
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 56796 354 56824 16546
rect 58440 6656 58492 6662
rect 58440 6598 58492 6604
rect 58452 480 58480 6598
rect 57214 354 57326 480
rect 56796 326 57326 354
rect 57214 -960 57326 326
rect 58410 -960 58522 480
rect 59372 354 59400 19042
rect 60752 16574 60780 19994
rect 62120 19168 62172 19174
rect 62120 19110 62172 19116
rect 62132 16574 62160 19110
rect 63512 16574 63540 20062
rect 60752 16546 60872 16574
rect 62132 16546 63264 16574
rect 63512 16546 64368 16574
rect 60844 480 60872 16546
rect 62028 6724 62080 6730
rect 62028 6666 62080 6672
rect 62040 480 62068 6666
rect 63236 480 63264 16546
rect 64340 480 64368 16546
rect 66720 14476 66772 14482
rect 66720 14418 66772 14424
rect 65524 6792 65576 6798
rect 65524 6734 65576 6740
rect 65536 480 65564 6734
rect 66732 480 66760 14418
rect 59606 354 59718 480
rect 59372 326 59718 354
rect 59606 -960 59718 326
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67652 354 67680 20130
rect 70412 16574 70440 20198
rect 74552 16574 74580 20266
rect 144920 19236 144972 19242
rect 144920 19178 144972 19184
rect 143540 17332 143592 17338
rect 143540 17274 143592 17280
rect 142160 17264 142212 17270
rect 131118 17232 131174 17241
rect 142160 17206 142212 17212
rect 131118 17167 131174 17176
rect 131132 16574 131160 17167
rect 70412 16546 71544 16574
rect 74552 16546 75040 16574
rect 131132 16546 131344 16574
rect 69848 14544 69900 14550
rect 69848 14486 69900 14492
rect 69112 6860 69164 6866
rect 69112 6802 69164 6808
rect 69124 480 69152 6802
rect 67886 354 67998 480
rect 67652 326 67998 354
rect 67886 -960 67998 326
rect 69082 -960 69194 480
rect 69860 354 69888 14486
rect 71516 480 71544 16546
rect 73344 14612 73396 14618
rect 73344 14554 73396 14560
rect 72608 9308 72660 9314
rect 72608 9250 72660 9256
rect 72620 480 72648 9250
rect 70278 354 70390 480
rect 69860 326 70390 354
rect 70278 -960 70390 326
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73356 354 73384 14554
rect 75012 480 75040 16546
rect 125600 16312 125652 16318
rect 125600 16254 125652 16260
rect 123024 16244 123076 16250
rect 123024 16186 123076 16192
rect 118700 16176 118752 16182
rect 118700 16118 118752 16124
rect 116400 16108 116452 16114
rect 116400 16050 116452 16056
rect 102232 15156 102284 15162
rect 102232 15098 102284 15104
rect 98184 15088 98236 15094
rect 98184 15030 98236 15036
rect 93860 15020 93912 15026
rect 93860 14962 93912 14968
rect 91560 14952 91612 14958
rect 91560 14894 91612 14900
rect 87512 14884 87564 14890
rect 87512 14826 87564 14832
rect 84200 14816 84252 14822
rect 84200 14758 84252 14764
rect 80888 14748 80940 14754
rect 80888 14690 80940 14696
rect 77392 14680 77444 14686
rect 77392 14622 77444 14628
rect 76196 9376 76248 9382
rect 76196 9318 76248 9324
rect 76208 480 76236 9318
rect 77404 480 77432 14622
rect 79230 10296 79286 10305
rect 79230 10231 79286 10240
rect 78588 5296 78640 5302
rect 78588 5238 78640 5244
rect 78600 480 78628 5238
rect 73774 354 73886 480
rect 73356 326 73886 354
rect 73774 -960 73886 326
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79244 354 79272 10231
rect 80900 480 80928 14690
rect 83280 10328 83332 10334
rect 83280 10270 83332 10276
rect 82084 4004 82136 4010
rect 82084 3946 82136 3952
rect 82096 480 82124 3946
rect 83292 480 83320 10270
rect 79662 354 79774 480
rect 79244 326 79774 354
rect 79662 -960 79774 326
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84212 354 84240 14758
rect 86408 10396 86460 10402
rect 86408 10338 86460 10344
rect 85672 5500 85724 5506
rect 85672 5442 85724 5448
rect 85684 480 85712 5442
rect 84446 354 84558 480
rect 84212 326 84558 354
rect 84446 -960 84558 326
rect 85642 -960 85754 480
rect 86420 354 86448 10338
rect 86838 354 86950 480
rect 86420 326 86950 354
rect 87524 354 87552 14826
rect 89904 10464 89956 10470
rect 89904 10406 89956 10412
rect 89168 5432 89220 5438
rect 89168 5374 89220 5380
rect 89180 480 89208 5374
rect 87942 354 88054 480
rect 87524 326 88054 354
rect 86838 -960 86950 326
rect 87942 -960 88054 326
rect 89138 -960 89250 480
rect 89916 354 89944 10406
rect 91572 480 91600 14894
rect 92756 4072 92808 4078
rect 92756 4014 92808 4020
rect 92768 480 92796 4014
rect 93872 3398 93900 14962
rect 97448 13388 97500 13394
rect 97448 13330 97500 13336
rect 93952 13320 94004 13326
rect 93952 13262 94004 13268
rect 93860 3392 93912 3398
rect 93860 3334 93912 3340
rect 93964 480 93992 13262
rect 96252 5092 96304 5098
rect 96252 5034 96304 5040
rect 94780 3392 94832 3398
rect 94780 3334 94832 3340
rect 90334 354 90446 480
rect 89916 326 90446 354
rect 90334 -960 90446 326
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 94792 354 94820 3334
rect 96264 480 96292 5034
rect 97460 480 97488 13330
rect 95118 354 95230 480
rect 94792 326 95230 354
rect 95118 -960 95230 326
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98196 354 98224 15030
rect 100760 13456 100812 13462
rect 100760 13398 100812 13404
rect 99840 4140 99892 4146
rect 99840 4082 99892 4088
rect 99852 480 99880 4082
rect 98614 354 98726 480
rect 98196 326 98726 354
rect 98614 -960 98726 326
rect 99810 -960 99922 480
rect 100772 354 100800 13398
rect 102244 480 102272 15098
rect 105728 14408 105780 14414
rect 105728 14350 105780 14356
rect 104072 13524 104124 13530
rect 104072 13466 104124 13472
rect 103336 5024 103388 5030
rect 103336 4966 103388 4972
rect 103348 480 103376 4966
rect 101006 354 101118 480
rect 100772 326 101118 354
rect 101006 -960 101118 326
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104084 354 104112 13466
rect 105740 480 105768 14350
rect 109040 14340 109092 14346
rect 109040 14282 109092 14288
rect 108120 13592 108172 13598
rect 108120 13534 108172 13540
rect 106924 3324 106976 3330
rect 106924 3266 106976 3272
rect 106936 480 106964 3266
rect 108132 480 108160 13534
rect 104502 354 104614 480
rect 104084 326 104614 354
rect 104502 -960 104614 326
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109052 354 109080 14282
rect 112352 14272 112404 14278
rect 112352 14214 112404 14220
rect 110420 13660 110472 13666
rect 110420 13602 110472 13608
rect 110432 3398 110460 13602
rect 110512 5364 110564 5370
rect 110512 5306 110564 5312
rect 110420 3392 110472 3398
rect 110420 3334 110472 3340
rect 110524 480 110552 5306
rect 111616 3392 111668 3398
rect 111616 3334 111668 3340
rect 111628 480 111656 3334
rect 109286 354 109398 480
rect 109052 326 109398 354
rect 109286 -960 109398 326
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112364 354 112392 14214
rect 114744 13728 114796 13734
rect 114744 13670 114796 13676
rect 114008 3256 114060 3262
rect 114008 3198 114060 3204
rect 114020 480 114048 3198
rect 112782 354 112894 480
rect 112364 326 112894 354
rect 112782 -960 112894 326
rect 113978 -960 114090 480
rect 114756 354 114784 13670
rect 116412 480 116440 16050
rect 117596 5228 117648 5234
rect 117596 5170 117648 5176
rect 117608 480 117636 5170
rect 118712 3330 118740 16118
rect 118792 13796 118844 13802
rect 118792 13738 118844 13744
rect 118700 3324 118752 3330
rect 118700 3266 118752 3272
rect 118804 480 118832 13738
rect 122288 13048 122340 13054
rect 122288 12990 122340 12996
rect 121092 5160 121144 5166
rect 121092 5102 121144 5108
rect 119896 3324 119948 3330
rect 119896 3266 119948 3272
rect 119908 480 119936 3266
rect 121104 480 121132 5102
rect 122300 480 122328 12990
rect 115174 354 115286 480
rect 114756 326 115286 354
rect 115174 -960 115286 326
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123036 354 123064 16186
rect 124680 3256 124732 3262
rect 124680 3198 124732 3204
rect 124692 480 124720 3198
rect 123454 354 123566 480
rect 123036 326 123566 354
rect 123454 -960 123566 326
rect 124650 -960 124762 480
rect 125612 354 125640 16254
rect 126980 10532 127032 10538
rect 126980 10474 127032 10480
rect 126992 4214 127020 10474
rect 130568 7676 130620 7682
rect 130568 7618 130620 7624
rect 127072 7608 127124 7614
rect 127072 7550 127124 7556
rect 126980 4208 127032 4214
rect 126980 4150 127032 4156
rect 127084 3482 127112 7550
rect 129372 4820 129424 4826
rect 129372 4762 129424 4768
rect 128176 4208 128228 4214
rect 128176 4150 128228 4156
rect 126992 3454 127112 3482
rect 126992 480 127020 3454
rect 128188 480 128216 4150
rect 129384 480 129412 4762
rect 130580 480 130608 7618
rect 125846 354 125958 480
rect 125612 326 125958 354
rect 125846 -960 125958 326
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131316 354 131344 16546
rect 138848 12028 138900 12034
rect 138848 11970 138900 11976
rect 135260 11960 135312 11966
rect 135260 11902 135312 11908
rect 134156 7744 134208 7750
rect 134156 7686 134208 7692
rect 132960 4888 133012 4894
rect 132960 4830 133012 4836
rect 132972 480 133000 4830
rect 134168 480 134196 7686
rect 135272 480 135300 11902
rect 137652 9444 137704 9450
rect 137652 9386 137704 9392
rect 136456 4752 136508 4758
rect 136456 4694 136508 4700
rect 136468 480 136496 4694
rect 137664 480 137692 9386
rect 138860 480 138888 11970
rect 141240 9512 141292 9518
rect 141240 9454 141292 9460
rect 140044 6112 140096 6118
rect 140044 6054 140096 6060
rect 140056 480 140084 6054
rect 141252 480 141280 9454
rect 131734 354 131846 480
rect 131316 326 131846 354
rect 131734 -960 131846 326
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142172 354 142200 17206
rect 143552 3194 143580 17274
rect 144932 16574 144960 19178
rect 144932 16546 145512 16574
rect 143632 6044 143684 6050
rect 143632 5986 143684 5992
rect 143540 3188 143592 3194
rect 143540 3130 143592 3136
rect 143644 3074 143672 5986
rect 144736 3188 144788 3194
rect 144736 3130 144788 3136
rect 143552 3046 143672 3074
rect 143552 480 143580 3046
rect 144748 480 144776 3130
rect 142406 354 142518 480
rect 142172 326 142518 354
rect 142406 -960 142518 326
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145484 354 145512 16546
rect 145576 5302 145604 336330
rect 149060 19304 149112 19310
rect 149060 19246 149112 19252
rect 147680 17468 147732 17474
rect 147680 17410 147732 17416
rect 146300 17400 146352 17406
rect 146300 17342 146352 17348
rect 146312 16574 146340 17342
rect 147692 16574 147720 17410
rect 149072 16574 149100 19246
rect 146312 16546 147168 16574
rect 147692 16546 147904 16574
rect 149072 16546 149560 16574
rect 145564 5296 145616 5302
rect 145564 5238 145616 5244
rect 146944 4956 146996 4962
rect 146944 4898 146996 4904
rect 146956 4758 146984 4898
rect 146944 4752 146996 4758
rect 146944 4694 146996 4700
rect 147140 480 147168 16546
rect 145902 354 146014 480
rect 145484 326 146014 354
rect 145902 -960 146014 326
rect 147098 -960 147210 480
rect 147876 354 147904 16546
rect 149532 480 149560 16546
rect 149716 5506 149744 336398
rect 151820 18556 151872 18562
rect 151820 18498 151872 18504
rect 150440 17536 150492 17542
rect 150440 17478 150492 17484
rect 150452 16574 150480 17478
rect 150452 16546 150664 16574
rect 149704 5500 149756 5506
rect 149704 5442 149756 5448
rect 150636 480 150664 16546
rect 151832 9674 151860 18498
rect 153200 17672 153252 17678
rect 153200 17614 153252 17620
rect 151912 17604 151964 17610
rect 151912 17546 151964 17552
rect 151740 9654 151860 9674
rect 151728 9648 151860 9654
rect 151780 9646 151860 9648
rect 151728 9590 151780 9596
rect 151924 6914 151952 17546
rect 153212 16574 153240 17614
rect 153212 16546 153792 16574
rect 153016 9648 153068 9654
rect 153016 9590 153068 9596
rect 151832 6886 151952 6914
rect 151832 480 151860 6886
rect 153028 480 153056 9590
rect 148294 354 148406 480
rect 147876 326 148406 354
rect 148294 -960 148406 326
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 153764 354 153792 16546
rect 153856 5438 153884 336466
rect 161296 16380 161348 16386
rect 161296 16322 161348 16328
rect 156144 12980 156196 12986
rect 156144 12922 156196 12928
rect 155408 10600 155460 10606
rect 155408 10542 155460 10548
rect 153844 5432 153896 5438
rect 153844 5374 153896 5380
rect 155420 480 155448 10542
rect 154182 354 154294 480
rect 153764 326 154294 354
rect 154182 -960 154294 326
rect 155378 -960 155490 480
rect 156156 354 156184 12922
rect 160100 12912 160152 12918
rect 160100 12854 160152 12860
rect 158904 10668 158956 10674
rect 158904 10610 158956 10616
rect 157800 7812 157852 7818
rect 157800 7754 157852 7760
rect 157812 480 157840 7754
rect 158916 480 158944 10610
rect 160112 480 160140 12854
rect 161308 480 161336 16322
rect 163412 10736 163464 10742
rect 163412 10678 163464 10684
rect 162490 7576 162546 7585
rect 162490 7511 162546 7520
rect 162504 480 162532 7511
rect 163424 3482 163452 10678
rect 163516 5098 163544 336534
rect 171968 16584 172020 16590
rect 171968 16526 172020 16532
rect 168380 16516 168432 16522
rect 168380 16458 168432 16464
rect 164424 16448 164476 16454
rect 164424 16390 164476 16396
rect 163504 5092 163556 5098
rect 163504 5034 163556 5040
rect 163424 3454 163728 3482
rect 163700 480 163728 3454
rect 156574 354 156686 480
rect 156156 326 156686 354
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164436 354 164464 16390
rect 167184 10804 167236 10810
rect 167184 10746 167236 10752
rect 166080 7880 166132 7886
rect 166080 7822 166132 7828
rect 166092 480 166120 7822
rect 167196 480 167224 10746
rect 168392 480 168420 16458
rect 170312 10872 170364 10878
rect 170312 10814 170364 10820
rect 169576 7948 169628 7954
rect 169576 7890 169628 7896
rect 169588 480 169616 7890
rect 164854 354 164966 480
rect 164436 326 164966 354
rect 164854 -960 164966 326
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170324 354 170352 10814
rect 171980 480 172008 16526
rect 173072 8016 173124 8022
rect 173072 7958 173124 7964
rect 173084 3482 173112 7958
rect 173176 5030 173204 336602
rect 176660 11008 176712 11014
rect 176660 10950 176712 10956
rect 173900 10940 173952 10946
rect 173900 10882 173952 10888
rect 173164 5024 173216 5030
rect 173164 4966 173216 4972
rect 173084 3454 173204 3482
rect 173176 480 173204 3454
rect 170742 354 170854 480
rect 170324 326 170854 354
rect 170742 -960 170854 326
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173912 354 173940 10882
rect 175464 4684 175516 4690
rect 175464 4626 175516 4632
rect 175476 480 175504 4626
rect 176672 4214 176700 10950
rect 176752 8084 176804 8090
rect 176752 8026 176804 8032
rect 176660 4208 176712 4214
rect 176660 4150 176712 4156
rect 176764 3482 176792 8026
rect 177316 5370 177344 336670
rect 185584 335980 185636 335986
rect 185584 335922 185636 335928
rect 180984 10260 181036 10266
rect 180984 10202 181036 10208
rect 180248 8152 180300 8158
rect 180248 8094 180300 8100
rect 177304 5364 177356 5370
rect 177304 5306 177356 5312
rect 179052 4616 179104 4622
rect 179052 4558 179104 4564
rect 177856 4208 177908 4214
rect 177856 4150 177908 4156
rect 176672 3454 176792 3482
rect 176672 480 176700 3454
rect 177868 480 177896 4150
rect 179064 480 179092 4558
rect 180260 480 180288 8094
rect 174238 354 174350 480
rect 173912 326 174350 354
rect 174238 -960 174350 326
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 180996 354 181024 10202
rect 184940 10192 184992 10198
rect 184940 10134 184992 10140
rect 183744 8220 183796 8226
rect 183744 8162 183796 8168
rect 182548 5024 182600 5030
rect 182548 4966 182600 4972
rect 182560 480 182588 4966
rect 183756 480 183784 8162
rect 184952 480 184980 10134
rect 185596 5234 185624 335922
rect 188344 335912 188396 335918
rect 188344 335854 188396 335860
rect 188252 10124 188304 10130
rect 188252 10066 188304 10072
rect 187332 8288 187384 8294
rect 187332 8230 187384 8236
rect 185584 5228 185636 5234
rect 185584 5170 185636 5176
rect 186136 5092 186188 5098
rect 186136 5034 186188 5040
rect 186148 480 186176 5034
rect 187344 480 187372 8230
rect 188264 3482 188292 10066
rect 188356 5166 188384 335854
rect 231136 97986 231164 459070
rect 231228 150414 231256 459138
rect 234250 457328 234306 457337
rect 234250 457263 234306 457272
rect 234066 457192 234122 457201
rect 234066 457127 234122 457136
rect 234160 457156 234212 457162
rect 233882 457056 233938 457065
rect 233882 456991 233938 457000
rect 233606 456376 233662 456385
rect 233606 456311 233662 456320
rect 233620 306338 233648 456311
rect 233790 456240 233846 456249
rect 233790 456175 233846 456184
rect 233608 306332 233660 306338
rect 233608 306274 233660 306280
rect 233804 255270 233832 456175
rect 233792 255264 233844 255270
rect 233792 255206 233844 255212
rect 231216 150408 231268 150414
rect 231216 150350 231268 150356
rect 231124 97980 231176 97986
rect 231124 97922 231176 97928
rect 233896 85542 233924 456991
rect 233974 456104 234030 456113
rect 233974 456039 234030 456048
rect 233988 202842 234016 456039
rect 233976 202836 234028 202842
rect 233976 202778 234028 202784
rect 234080 137970 234108 457127
rect 234160 457098 234212 457104
rect 234172 241466 234200 457098
rect 234160 241460 234212 241466
rect 234160 241402 234212 241408
rect 234264 189038 234292 457263
rect 234252 189032 234304 189038
rect 234252 188974 234304 188980
rect 234068 137964 234120 137970
rect 234068 137906 234120 137912
rect 234356 100706 234384 459886
rect 234436 459672 234488 459678
rect 234436 459614 234488 459620
rect 234344 100700 234396 100706
rect 234344 100642 234396 100648
rect 233884 85536 233936 85542
rect 233884 85478 233936 85484
rect 234448 60722 234476 459614
rect 234528 459604 234580 459610
rect 234528 459546 234580 459552
rect 234436 60716 234488 60722
rect 234436 60658 234488 60664
rect 234540 20602 234568 459546
rect 237300 457994 237328 460391
rect 250260 460284 250312 460290
rect 250260 460226 250312 460232
rect 248052 459944 248104 459950
rect 246946 459912 247002 459921
rect 248052 459886 248104 459892
rect 246946 459847 247002 459856
rect 242346 459776 242402 459785
rect 242346 459711 242402 459720
rect 238852 459604 238904 459610
rect 238852 459546 238904 459552
rect 238864 457994 238892 459546
rect 240782 458552 240838 458561
rect 240782 458487 240838 458496
rect 240796 457994 240824 458487
rect 242360 457994 242388 459711
rect 243268 459672 243320 459678
rect 243268 459614 243320 459620
rect 237300 457966 237360 457994
rect 238864 457966 238924 457994
rect 240488 457966 240824 457994
rect 242052 457966 242388 457994
rect 243280 457994 243308 459614
rect 245566 458688 245622 458697
rect 245566 458623 245622 458632
rect 245580 457994 245608 458623
rect 246960 457994 246988 459847
rect 243280 457966 243616 457994
rect 245272 457966 245608 457994
rect 246836 457966 246988 457994
rect 248064 457994 248092 459886
rect 250272 457994 250300 460226
rect 251822 460048 251878 460057
rect 251822 459983 251878 459992
rect 251836 457994 251864 459983
rect 248064 457966 248400 457994
rect 249964 457966 250300 457994
rect 251528 457966 251864 457994
rect 252664 457994 252692 478858
rect 272340 460964 272392 460970
rect 272340 460906 272392 460912
rect 255044 460352 255096 460358
rect 255044 460294 255096 460300
rect 259366 460320 259422 460329
rect 255056 457994 255084 460294
rect 259366 460255 259422 460264
rect 256606 460184 256662 460193
rect 256606 460119 256662 460128
rect 256620 457994 256648 460119
rect 257988 458652 258040 458658
rect 257988 458594 258040 458600
rect 252664 457966 253092 457994
rect 254748 457966 255084 457994
rect 256312 457966 256648 457994
rect 258000 457858 258028 458594
rect 259380 457994 259408 460255
rect 269028 460012 269080 460018
rect 269028 459954 269080 459960
rect 264520 459944 264572 459950
rect 264520 459886 264572 459892
rect 262864 458720 262916 458726
rect 262864 458662 262916 458668
rect 262876 457994 262904 458662
rect 264532 457994 264560 459886
rect 267648 458788 267700 458794
rect 267648 458730 267700 458736
rect 267660 457994 267688 458730
rect 269040 457994 269068 459954
rect 270408 458856 270460 458862
rect 270408 458798 270460 458804
rect 259380 457966 259440 457994
rect 262568 457966 262904 457994
rect 264224 457966 264560 457994
rect 267352 457966 267688 457994
rect 268916 457966 269068 457994
rect 270420 457994 270448 458798
rect 272352 457994 272380 460906
rect 282932 460426 282960 702406
rect 298100 643136 298152 643142
rect 298100 643078 298152 643084
rect 296720 616888 296772 616894
rect 296720 616830 296772 616836
rect 293960 590708 294012 590714
rect 293960 590650 294012 590656
rect 292580 563100 292632 563106
rect 292580 563042 292632 563048
rect 288440 536852 288492 536858
rect 288440 536794 288492 536800
rect 287060 510672 287112 510678
rect 287060 510614 287112 510620
rect 284300 484424 284352 484430
rect 284300 484366 284352 484372
rect 282920 460420 282972 460426
rect 282920 460362 282972 460368
rect 277124 460216 277176 460222
rect 277124 460158 277176 460164
rect 277136 457994 277164 460158
rect 281448 460148 281500 460154
rect 281448 460090 281500 460096
rect 280068 460080 280120 460086
rect 280068 460022 280120 460028
rect 280080 457994 280108 460022
rect 270420 457966 270480 457994
rect 272044 457966 272380 457994
rect 276828 457966 277164 457994
rect 279956 457966 280108 457994
rect 281460 457994 281488 460090
rect 283472 458924 283524 458930
rect 283472 458866 283524 458872
rect 283484 457994 283512 458866
rect 281460 457966 281520 457994
rect 283176 457966 283512 457994
rect 284312 457994 284340 484366
rect 287072 480254 287100 510614
rect 288452 480254 288480 536794
rect 289820 524476 289872 524482
rect 289820 524418 289872 524424
rect 289832 480254 289860 524418
rect 287072 480226 287468 480254
rect 288452 480226 289032 480254
rect 289832 480226 290596 480254
rect 285864 470620 285916 470626
rect 285864 470562 285916 470568
rect 285876 457994 285904 470562
rect 287440 457994 287468 480226
rect 289004 457994 289032 480226
rect 290568 457994 290596 480226
rect 292592 457994 292620 563042
rect 293972 457994 294000 590650
rect 295340 576904 295392 576910
rect 295340 576846 295392 576852
rect 295352 457994 295380 576846
rect 296732 480254 296760 616830
rect 298112 480254 298140 643078
rect 296732 480226 296944 480254
rect 298112 480226 298508 480254
rect 296916 457994 296944 480226
rect 298480 457994 298508 480226
rect 299492 462262 299520 703582
rect 299952 703474 299980 703582
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 300136 703474 300164 703520
rect 299952 703446 300164 703474
rect 332520 703050 332548 703520
rect 331220 703044 331272 703050
rect 331220 702986 331272 702992
rect 332508 703044 332560 703050
rect 332508 702986 332560 702992
rect 318800 701004 318852 701010
rect 318800 700946 318852 700952
rect 314660 700868 314712 700874
rect 314660 700810 314712 700816
rect 309140 700596 309192 700602
rect 309140 700538 309192 700544
rect 303620 696992 303672 696998
rect 303620 696934 303672 696940
rect 300860 670812 300912 670818
rect 300860 670754 300912 670760
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299584 480254 299612 630634
rect 300872 480254 300900 670754
rect 299584 480226 300072 480254
rect 300872 480226 301728 480254
rect 299480 462256 299532 462262
rect 299480 462198 299532 462204
rect 300044 457994 300072 480226
rect 301700 457994 301728 480226
rect 303632 457994 303660 696934
rect 305000 683256 305052 683262
rect 305000 683198 305052 683204
rect 305012 457994 305040 683198
rect 309152 480254 309180 700538
rect 309152 480226 309548 480254
rect 307116 461712 307168 461718
rect 307116 461654 307168 461660
rect 307128 457994 307156 461654
rect 308680 460488 308732 460494
rect 308680 460430 308732 460436
rect 308692 457994 308720 460430
rect 308956 460352 309008 460358
rect 308956 460294 309008 460300
rect 284312 457966 284740 457994
rect 285876 457966 286304 457994
rect 287440 457966 287868 457994
rect 289004 457966 289432 457994
rect 290568 457966 290996 457994
rect 292592 457966 292652 457994
rect 293972 457966 294216 457994
rect 295352 457966 295780 457994
rect 296916 457966 297344 457994
rect 298480 457966 298908 457994
rect 300044 457966 300472 457994
rect 301700 457966 302128 457994
rect 303632 457966 303692 457994
rect 305012 457966 305256 457994
rect 306820 457966 307156 457994
rect 308384 457966 308720 457994
rect 257876 457830 258028 457858
rect 261300 457496 261352 457502
rect 234724 457422 235796 457450
rect 261004 457444 261300 457450
rect 266084 457496 266136 457502
rect 261004 457438 261352 457444
rect 265788 457444 266084 457450
rect 273996 457496 274048 457502
rect 265788 457438 266136 457444
rect 273700 457444 273996 457450
rect 275560 457496 275612 457502
rect 273700 457438 274048 457444
rect 275264 457444 275560 457450
rect 278596 457496 278648 457502
rect 275264 457438 275612 457444
rect 278392 457444 278596 457450
rect 308968 457473 308996 460294
rect 309520 457994 309548 480226
rect 313188 461984 313240 461990
rect 313188 461926 313240 461932
rect 311808 461848 311860 461854
rect 311808 461790 311860 461796
rect 311820 457994 311848 461790
rect 313200 458266 313228 461926
rect 309520 457966 309948 457994
rect 311604 457966 311848 457994
rect 313154 458238 313228 458266
rect 313154 457980 313182 458238
rect 314672 457994 314700 700810
rect 317420 700256 317472 700262
rect 317420 700198 317472 700204
rect 316592 462052 316644 462058
rect 316592 461994 316644 462000
rect 316604 457994 316632 461994
rect 314672 457966 314732 457994
rect 316296 457966 316632 457994
rect 317432 457994 317460 700198
rect 318812 480254 318840 700946
rect 327908 700936 327960 700942
rect 327908 700878 327960 700884
rect 327724 700664 327776 700670
rect 327724 700606 327776 700612
rect 327816 700664 327868 700670
rect 327816 700606 327868 700612
rect 324964 700188 325016 700194
rect 324964 700130 325016 700136
rect 322940 700120 322992 700126
rect 322940 700062 322992 700068
rect 322952 480254 322980 700062
rect 318812 480226 319024 480254
rect 322952 480226 323808 480254
rect 318996 457994 319024 480226
rect 321376 462188 321428 462194
rect 321376 462130 321428 462136
rect 321388 457994 321416 462130
rect 322848 460352 322900 460358
rect 322848 460294 322900 460300
rect 321560 460284 321612 460290
rect 321560 460226 321612 460232
rect 321572 458998 321600 460226
rect 321560 458992 321612 458998
rect 321560 458934 321612 458940
rect 322860 457994 322888 460294
rect 317432 457966 317860 457994
rect 318996 457966 319424 457994
rect 321080 457966 321416 457994
rect 322644 457966 322888 457994
rect 323780 457994 323808 480226
rect 324976 460562 325004 700130
rect 325700 462256 325752 462262
rect 325700 462198 325752 462204
rect 324964 460556 325016 460562
rect 324964 460498 325016 460504
rect 325712 457994 325740 462198
rect 327080 460556 327132 460562
rect 327080 460498 327132 460504
rect 327092 457994 327120 460498
rect 327736 459610 327764 700606
rect 327828 460494 327856 700606
rect 327816 460488 327868 460494
rect 327816 460430 327868 460436
rect 327920 459678 327948 700878
rect 329104 700732 329156 700738
rect 329104 700674 329156 700680
rect 329116 460562 329144 700674
rect 330208 462120 330260 462126
rect 330208 462062 330260 462068
rect 329104 460556 329156 460562
rect 329104 460498 329156 460504
rect 328552 460420 328604 460426
rect 328552 460362 328604 460368
rect 327908 459672 327960 459678
rect 327908 459614 327960 459620
rect 327724 459604 327776 459610
rect 327724 459546 327776 459552
rect 328564 457994 328592 460362
rect 330220 457994 330248 462062
rect 331232 460358 331260 702986
rect 333244 700800 333296 700806
rect 333244 700742 333296 700748
rect 331864 700460 331916 700466
rect 331864 700402 331916 700408
rect 331876 460426 331904 700402
rect 331956 700324 332008 700330
rect 331956 700266 332008 700272
rect 331864 460420 331916 460426
rect 331864 460362 331916 460368
rect 331968 460358 331996 700266
rect 333256 460494 333284 700742
rect 338764 700528 338816 700534
rect 338764 700470 338816 700476
rect 337384 553444 337436 553450
rect 337384 553386 337436 553392
rect 334900 461916 334952 461922
rect 334900 461858 334952 461864
rect 333244 460488 333296 460494
rect 333244 460430 333296 460436
rect 331220 460352 331272 460358
rect 331220 460294 331272 460300
rect 331956 460352 332008 460358
rect 331956 460294 332008 460300
rect 333336 459672 333388 459678
rect 333336 459614 333388 459620
rect 331772 459604 331824 459610
rect 331772 459546 331824 459552
rect 331784 457994 331812 459546
rect 333348 457994 333376 459614
rect 334912 457994 334940 461858
rect 336740 460556 336792 460562
rect 336740 460498 336792 460504
rect 336752 457994 336780 460498
rect 337396 460290 337424 553386
rect 338120 460488 338172 460494
rect 338120 460430 338172 460436
rect 337384 460284 337436 460290
rect 337384 460226 337436 460232
rect 338132 457994 338160 460430
rect 338776 459610 338804 700470
rect 342904 700392 342956 700398
rect 342904 700334 342956 700340
rect 341524 501016 341576 501022
rect 341524 500958 341576 500964
rect 339684 461780 339736 461786
rect 339684 461722 339736 461728
rect 338764 459604 338816 459610
rect 338764 459546 338816 459552
rect 339696 457994 339724 461722
rect 341536 460426 341564 500958
rect 342916 460562 342944 700334
rect 348804 700126 348832 703520
rect 364996 702434 365024 703520
rect 364352 702406 365024 702434
rect 348792 700120 348844 700126
rect 348792 700062 348844 700068
rect 349160 683188 349212 683194
rect 349160 683130 349212 683136
rect 345664 514820 345716 514826
rect 345664 514762 345716 514768
rect 344376 461644 344428 461650
rect 344376 461586 344428 461592
rect 342904 460556 342956 460562
rect 342904 460498 342956 460504
rect 341248 460420 341300 460426
rect 341248 460362 341300 460368
rect 341524 460420 341576 460426
rect 341524 460362 341576 460368
rect 341260 457994 341288 460362
rect 342812 459604 342864 459610
rect 342812 459546 342864 459552
rect 342824 457994 342852 459546
rect 344388 457994 344416 461586
rect 345676 460494 345704 514762
rect 349068 462392 349120 462398
rect 349068 462334 349120 462340
rect 347780 460556 347832 460562
rect 347780 460498 347832 460504
rect 345664 460488 345716 460494
rect 345664 460430 345716 460436
rect 345940 460352 345992 460358
rect 345940 460294 345992 460300
rect 345952 457994 345980 460294
rect 347792 457994 347820 460498
rect 349080 460358 349108 462334
rect 349068 460352 349120 460358
rect 349068 460294 349120 460300
rect 349172 457994 349200 683130
rect 351920 670744 351972 670750
rect 351920 670686 351972 670692
rect 350540 656940 350592 656946
rect 350540 656882 350592 656888
rect 350552 480254 350580 656882
rect 351932 480254 351960 670686
rect 353300 632120 353352 632126
rect 353300 632062 353352 632068
rect 353312 480254 353340 632062
rect 356060 618316 356112 618322
rect 356060 618258 356112 618264
rect 354680 605872 354732 605878
rect 354680 605814 354732 605820
rect 354692 480254 354720 605814
rect 356072 480254 356100 618258
rect 358820 579692 358872 579698
rect 358820 579634 358872 579640
rect 350552 480226 350672 480254
rect 351932 480226 352236 480254
rect 353312 480226 353800 480254
rect 354692 480226 355364 480254
rect 356072 480226 356928 480254
rect 350644 457994 350672 480226
rect 352208 457994 352236 480226
rect 353772 457994 353800 480226
rect 355336 457994 355364 480226
rect 356900 457994 356928 480226
rect 358832 457994 358860 579634
rect 361580 565888 361632 565894
rect 361580 565830 361632 565836
rect 361592 480254 361620 565830
rect 362960 527196 363012 527202
rect 362960 527138 363012 527144
rect 362972 480254 363000 527138
rect 361592 480226 361712 480254
rect 362972 480226 363276 480254
rect 360200 460284 360252 460290
rect 360200 460226 360252 460232
rect 360212 457994 360240 460226
rect 360660 459604 360712 459610
rect 360660 459546 360712 459552
rect 323780 457966 324208 457994
rect 325712 457966 325772 457994
rect 327092 457966 327336 457994
rect 328564 457966 328900 457994
rect 330220 457966 330556 457994
rect 331784 457966 332120 457994
rect 333348 457966 333684 457994
rect 334912 457966 335248 457994
rect 336752 457966 336812 457994
rect 338132 457966 338376 457994
rect 339696 457966 340032 457994
rect 341260 457966 341596 457994
rect 342824 457966 343160 457994
rect 344388 457966 344724 457994
rect 345952 457966 346288 457994
rect 347792 457966 347852 457994
rect 349172 457966 349508 457994
rect 350644 457966 351072 457994
rect 352208 457966 352636 457994
rect 353772 457966 354200 457994
rect 355336 457966 355764 457994
rect 356900 457966 357328 457994
rect 358832 457966 358984 457994
rect 360212 457966 360548 457994
rect 360672 457502 360700 459546
rect 361684 457994 361712 480226
rect 363248 457994 363276 480226
rect 364352 462194 364380 702406
rect 397472 700262 397500 703520
rect 413664 701010 413692 703520
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 397460 700256 397512 700262
rect 397460 700198 397512 700204
rect 368020 474768 368072 474774
rect 368020 474710 368072 474716
rect 364340 462188 364392 462194
rect 364340 462130 364392 462136
rect 366456 460488 366508 460494
rect 366456 460430 366508 460436
rect 364892 460420 364944 460426
rect 364892 460362 364944 460368
rect 364904 457994 364932 460362
rect 366468 457994 366496 460430
rect 368032 457994 368060 474710
rect 429212 462058 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494072 703582 494652 703610
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 429200 462052 429252 462058
rect 429200 461994 429252 462000
rect 462332 461990 462360 703520
rect 478524 700874 478552 703520
rect 478512 700868 478564 700874
rect 478512 700810 478564 700816
rect 462320 461984 462372 461990
rect 462320 461926 462372 461932
rect 494072 461854 494100 703582
rect 494624 703474 494652 703582
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 494808 703474 494836 703520
rect 494624 703446 494836 703474
rect 527192 700670 527220 703520
rect 527180 700664 527232 700670
rect 527180 700606 527232 700612
rect 543476 700602 543504 703520
rect 559668 702434 559696 703520
rect 558932 702406 559696 702434
rect 543464 700596 543516 700602
rect 543464 700538 543516 700544
rect 494060 461848 494112 461854
rect 494060 461790 494112 461796
rect 558932 461718 558960 702406
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683262 580212 683839
rect 580172 683256 580224 683262
rect 580172 683198 580224 683204
rect 580172 670812 580224 670818
rect 580172 670754 580224 670760
rect 580184 670721 580212 670754
rect 580170 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 577596 478916 577648 478922
rect 577596 478858 577648 478864
rect 558920 461712 558972 461718
rect 558920 461654 558972 461660
rect 380900 460692 380952 460698
rect 380900 460634 380952 460640
rect 371240 460352 371292 460358
rect 371240 460294 371292 460300
rect 369860 459876 369912 459882
rect 369860 459818 369912 459824
rect 369872 457994 369900 459818
rect 371252 457994 371280 460294
rect 378048 460216 378100 460222
rect 378048 460158 378100 460164
rect 375932 459808 375984 459814
rect 375932 459750 375984 459756
rect 374368 459604 374420 459610
rect 374368 459546 374420 459552
rect 372804 458584 372856 458590
rect 372804 458526 372856 458532
rect 372816 457994 372844 458526
rect 374380 457994 374408 459546
rect 375944 457994 375972 459750
rect 378060 459066 378088 460158
rect 379152 459740 379204 459746
rect 379152 459682 379204 459688
rect 378048 459060 378100 459066
rect 378048 459002 378100 459008
rect 377588 458516 377640 458522
rect 377588 458458 377640 458464
rect 377600 457994 377628 458458
rect 379164 457994 379192 459682
rect 380912 457994 380940 460634
rect 383936 460624 383988 460630
rect 383936 460566 383988 460572
rect 382280 458448 382332 458454
rect 382280 458390 382332 458396
rect 382292 457994 382320 458390
rect 383948 457994 383976 460566
rect 577502 460456 577558 460465
rect 577502 460391 577558 460400
rect 415032 460148 415084 460154
rect 415032 460090 415084 460096
rect 399668 459196 399720 459202
rect 399668 459138 399720 459144
rect 387064 458380 387116 458386
rect 387064 458322 387116 458328
rect 387076 457994 387104 458322
rect 391940 458312 391992 458318
rect 391940 458254 391992 458260
rect 391952 457994 391980 458254
rect 396862 458244 396914 458250
rect 396862 458186 396914 458192
rect 361684 457966 362112 457994
rect 363248 457966 363676 457994
rect 364904 457966 365240 457994
rect 366468 457966 366804 457994
rect 368032 457966 368460 457994
rect 369872 457966 370024 457994
rect 371252 457966 371588 457994
rect 372816 457966 373152 457994
rect 374380 457966 374716 457994
rect 375944 457966 376280 457994
rect 377600 457966 377936 457994
rect 379164 457966 379500 457994
rect 380912 457966 381064 457994
rect 382292 457966 382628 457994
rect 383948 457966 384192 457994
rect 387076 457966 387412 457994
rect 391952 457966 392104 457994
rect 396874 457980 396902 458186
rect 399680 457994 399708 459138
rect 404360 459128 404412 459134
rect 404360 459070 404412 459076
rect 401230 458416 401286 458425
rect 401230 458351 401286 458360
rect 401244 457994 401272 458351
rect 404372 457994 404400 459070
rect 406336 458280 406392 458289
rect 406336 458215 406392 458224
rect 399680 457966 400016 457994
rect 401244 457966 401580 457994
rect 404372 457966 404708 457994
rect 406350 457980 406378 458215
rect 360660 457496 360712 457502
rect 278392 457438 278648 457444
rect 308954 457464 309010 457473
rect 261004 457422 261340 457438
rect 265788 457422 266124 457438
rect 273700 457422 274036 457438
rect 275264 457422 275600 457438
rect 278392 457422 278636 457438
rect 234724 345014 234752 457422
rect 388628 457496 388680 457502
rect 360660 457438 360712 457444
rect 385406 457464 385462 457473
rect 308954 457399 309010 457408
rect 385462 457422 385756 457450
rect 390190 457464 390246 457473
rect 388680 457444 388976 457450
rect 388628 457438 388976 457444
rect 388640 457422 388976 457438
rect 385406 457399 385462 457408
rect 393502 457464 393558 457473
rect 390246 457422 390540 457450
rect 390190 457399 390246 457408
rect 394974 457464 395030 457473
rect 393558 457422 393668 457450
rect 393502 457399 393558 457408
rect 398102 457464 398158 457473
rect 395030 457422 395232 457450
rect 394974 457399 395030 457408
rect 402978 457464 403034 457473
rect 398158 457422 398452 457450
rect 398102 457399 398158 457408
rect 407578 457464 407634 457473
rect 403034 457422 403144 457450
rect 402978 457399 403034 457408
rect 409142 457464 409198 457473
rect 407634 457422 407928 457450
rect 407578 457399 407634 457408
rect 410706 457464 410762 457473
rect 409198 457422 409492 457450
rect 409142 457399 409198 457408
rect 412270 457464 412326 457473
rect 410762 457422 411056 457450
rect 410706 457399 410762 457408
rect 412326 457422 412620 457450
rect 414184 457422 414980 457450
rect 412270 457399 412326 457408
rect 234632 344986 234752 345014
rect 234632 330682 234660 344986
rect 265052 338150 265296 338178
rect 234724 338014 235152 338042
rect 235276 338014 235428 338042
rect 235552 338014 235796 338042
rect 234620 330676 234672 330682
rect 234620 330618 234672 330624
rect 234724 330562 234752 338014
rect 234804 330676 234856 330682
rect 234804 330618 234856 330624
rect 234632 330534 234752 330562
rect 234528 20596 234580 20602
rect 234528 20538 234580 20544
rect 198740 18488 198792 18494
rect 198740 18430 198792 18436
rect 194600 17808 194652 17814
rect 194600 17750 194652 17756
rect 191840 17740 191892 17746
rect 191840 17682 191892 17688
rect 191852 16574 191880 17682
rect 194612 16574 194640 17750
rect 191852 16546 192064 16574
rect 194612 16546 195192 16574
rect 190828 7540 190880 7546
rect 190828 7482 190880 7488
rect 188344 5160 188396 5166
rect 188344 5102 188396 5108
rect 189724 5160 189776 5166
rect 189724 5102 189776 5108
rect 188264 3454 188568 3482
rect 188540 480 188568 3454
rect 189736 480 189764 5102
rect 190840 480 190868 7482
rect 192036 480 192064 16546
rect 194416 7472 194468 7478
rect 194416 7414 194468 7420
rect 193220 5228 193272 5234
rect 193220 5170 193272 5176
rect 193232 480 193260 5170
rect 194428 480 194456 7414
rect 181414 354 181526 480
rect 180996 326 181526 354
rect 181414 -960 181526 326
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195164 354 195192 16546
rect 197912 7404 197964 7410
rect 197912 7346 197964 7352
rect 196808 5296 196860 5302
rect 196808 5238 196860 5244
rect 196820 480 196848 5238
rect 197924 480 197952 7346
rect 195582 354 195694 480
rect 195164 326 195694 354
rect 195582 -960 195694 326
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 198752 354 198780 18430
rect 201500 18420 201552 18426
rect 201500 18362 201552 18368
rect 201512 11694 201540 18362
rect 204260 17944 204312 17950
rect 204260 17886 204312 17892
rect 201592 17876 201644 17882
rect 201592 17818 201644 17824
rect 201500 11688 201552 11694
rect 201500 11630 201552 11636
rect 201604 6914 201632 17818
rect 204272 16574 204300 17886
rect 208400 17196 208452 17202
rect 208400 17138 208452 17144
rect 208412 16574 208440 17138
rect 211160 17128 211212 17134
rect 211160 17070 211212 17076
rect 211172 16574 211200 17070
rect 215300 17060 215352 17066
rect 215300 17002 215352 17008
rect 204272 16546 205128 16574
rect 208412 16546 208624 16574
rect 211172 16546 211752 16574
rect 202696 11688 202748 11694
rect 202696 11630 202748 11636
rect 201512 6886 201632 6914
rect 200302 4856 200358 4865
rect 200302 4791 200358 4800
rect 200316 480 200344 4791
rect 201512 480 201540 6886
rect 202708 480 202736 11630
rect 203892 5364 203944 5370
rect 203892 5306 203944 5312
rect 203904 480 203932 5306
rect 205100 480 205128 16546
rect 206192 12096 206244 12102
rect 206192 12038 206244 12044
rect 206204 480 206232 12038
rect 207388 5432 207440 5438
rect 207388 5374 207440 5380
rect 207400 480 207428 5374
rect 208596 480 208624 16546
rect 209780 12164 209832 12170
rect 209780 12106 209832 12112
rect 209792 480 209820 12106
rect 210976 5500 211028 5506
rect 210976 5442 211028 5448
rect 210988 480 211016 5442
rect 199078 354 199190 480
rect 198752 326 199190 354
rect 199078 -960 199190 326
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 211724 354 211752 16546
rect 213368 12232 213420 12238
rect 213368 12174 213420 12180
rect 213380 480 213408 12174
rect 214472 4752 214524 4758
rect 214472 4694 214524 4700
rect 214484 480 214512 4694
rect 212142 354 212254 480
rect 211724 326 212254 354
rect 212142 -960 212254 326
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215312 354 215340 17002
rect 234632 15881 234660 330534
rect 234816 330426 234844 330618
rect 234724 330398 234844 330426
rect 234724 19990 234752 330398
rect 234804 329452 234856 329458
rect 234804 329394 234856 329400
rect 234712 19984 234764 19990
rect 234712 19926 234764 19932
rect 234618 15872 234674 15881
rect 218060 15836 218112 15842
rect 234618 15807 234674 15816
rect 218060 15778 218112 15784
rect 216864 12300 216916 12306
rect 216864 12242 216916 12248
rect 216876 480 216904 12242
rect 218072 480 218100 15778
rect 221096 15768 221148 15774
rect 221096 15710 221148 15716
rect 219992 12368 220044 12374
rect 219992 12310 220044 12316
rect 219256 9580 219308 9586
rect 219256 9522 219308 9528
rect 219268 480 219296 9522
rect 215638 354 215750 480
rect 215312 326 215750 354
rect 215638 -960 215750 326
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220004 354 220032 12310
rect 220422 354 220534 480
rect 220004 326 220534 354
rect 221108 354 221136 15710
rect 225144 15700 225196 15706
rect 225144 15642 225196 15648
rect 223580 12436 223632 12442
rect 223580 12378 223632 12384
rect 222752 9648 222804 9654
rect 222752 9590 222804 9596
rect 222764 480 222792 9590
rect 221526 354 221638 480
rect 221108 326 221638 354
rect 220422 -960 220534 326
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223592 354 223620 12378
rect 225156 480 225184 15642
rect 226340 11688 226392 11694
rect 226340 11630 226392 11636
rect 226352 4214 226380 11630
rect 231032 11620 231084 11626
rect 231032 11562 231084 11568
rect 226432 8900 226484 8906
rect 226432 8842 226484 8848
rect 226340 4208 226392 4214
rect 226340 4150 226392 4156
rect 226444 3482 226472 8842
rect 229836 8832 229888 8838
rect 229836 8774 229888 8780
rect 228730 6216 228786 6225
rect 228730 6151 228786 6160
rect 227536 4208 227588 4214
rect 227536 4150 227588 4156
rect 226352 3454 226472 3482
rect 226352 480 226380 3454
rect 227548 480 227576 4150
rect 228744 480 228772 6151
rect 229848 480 229876 8774
rect 231044 480 231072 11562
rect 234620 11552 234672 11558
rect 234620 11494 234672 11500
rect 233424 8764 233476 8770
rect 233424 8706 233476 8712
rect 232228 5976 232280 5982
rect 232228 5918 232280 5924
rect 232240 480 232268 5918
rect 233436 480 233464 8706
rect 234632 480 234660 11494
rect 234816 6254 234844 329394
rect 235276 316034 235304 338014
rect 235552 329458 235580 338014
rect 236150 337770 236178 338028
rect 236288 338014 236532 338042
rect 236656 338014 236900 338042
rect 237024 338014 237268 338042
rect 237576 338014 237636 338042
rect 237760 338014 238004 338042
rect 238128 338014 238372 338042
rect 238496 338014 238740 338042
rect 238864 338014 239108 338042
rect 239232 338014 239476 338042
rect 239600 338014 239844 338042
rect 240212 338014 240364 338042
rect 236150 337742 236224 337770
rect 236092 330540 236144 330546
rect 236092 330482 236144 330488
rect 235540 329452 235592 329458
rect 235540 329394 235592 329400
rect 234908 316006 235304 316034
rect 234804 6248 234856 6254
rect 234804 6190 234856 6196
rect 234908 6186 234936 316006
rect 236104 6322 236132 330482
rect 236196 8974 236224 337742
rect 236184 8968 236236 8974
rect 236184 8910 236236 8916
rect 236092 6316 236144 6322
rect 236092 6258 236144 6264
rect 234896 6180 234948 6186
rect 234896 6122 234948 6128
rect 235816 5908 235868 5914
rect 235816 5850 235868 5856
rect 235828 480 235856 5850
rect 236288 3369 236316 338014
rect 236656 336054 236684 338014
rect 236644 336048 236696 336054
rect 236644 335990 236696 335996
rect 236644 335504 236696 335510
rect 236644 335446 236696 335452
rect 236656 4078 236684 335446
rect 237024 330546 237052 338014
rect 237012 330540 237064 330546
rect 237012 330482 237064 330488
rect 237472 330540 237524 330546
rect 237472 330482 237524 330488
rect 237380 329316 237432 329322
rect 237380 329258 237432 329264
rect 237012 6180 237064 6186
rect 237012 6122 237064 6128
rect 236644 4072 236696 4078
rect 236644 4014 236696 4020
rect 236274 3360 236330 3369
rect 236274 3295 236330 3304
rect 237024 480 237052 6122
rect 237392 3466 237420 329258
rect 237484 6390 237512 330482
rect 237576 11665 237604 338014
rect 237760 316034 237788 338014
rect 238128 329322 238156 338014
rect 238496 330546 238524 338014
rect 238484 330540 238536 330546
rect 238484 330482 238536 330488
rect 238116 329316 238168 329322
rect 238116 329258 238168 329264
rect 237668 316006 237788 316034
rect 237668 18601 237696 316006
rect 237654 18592 237710 18601
rect 237654 18527 237710 18536
rect 238864 11762 238892 338014
rect 239232 316034 239260 338014
rect 239600 336122 239628 338014
rect 239588 336116 239640 336122
rect 239588 336058 239640 336064
rect 239404 336048 239456 336054
rect 239404 335990 239456 335996
rect 238956 316006 239260 316034
rect 238852 11756 238904 11762
rect 238852 11698 238904 11704
rect 237562 11656 237618 11665
rect 237562 11591 237618 11600
rect 238116 8968 238168 8974
rect 238116 8910 238168 8916
rect 237472 6384 237524 6390
rect 237472 6326 237524 6332
rect 237380 3460 237432 3466
rect 237380 3402 237432 3408
rect 238128 480 238156 8910
rect 238956 3534 238984 316006
rect 239312 6316 239364 6322
rect 239312 6258 239364 6264
rect 238944 3528 238996 3534
rect 238944 3470 238996 3476
rect 239324 480 239352 6258
rect 239416 4146 239444 335990
rect 240140 330540 240192 330546
rect 240140 330482 240192 330488
rect 239404 4140 239456 4146
rect 239404 4082 239456 4088
rect 240152 3670 240180 330482
rect 240232 330472 240284 330478
rect 240232 330414 240284 330420
rect 240140 3664 240192 3670
rect 240140 3606 240192 3612
rect 240244 3602 240272 330414
rect 240336 8945 240364 338014
rect 240428 338014 240580 338042
rect 240704 338014 240948 338042
rect 241072 338014 241316 338042
rect 241624 338014 241684 338042
rect 241808 338014 242052 338042
rect 242176 338014 242420 338042
rect 242544 338014 242788 338042
rect 243004 338014 243156 338042
rect 243280 338014 243524 338042
rect 243648 338014 243892 338042
rect 244016 338014 244260 338042
rect 244384 338014 244628 338042
rect 244752 338014 244996 338042
rect 245120 338014 245364 338042
rect 245732 338014 245884 338042
rect 240428 11830 240456 338014
rect 240704 330546 240732 338014
rect 240692 330540 240744 330546
rect 240692 330482 240744 330488
rect 241072 330478 241100 338014
rect 241060 330472 241112 330478
rect 241060 330414 241112 330420
rect 240416 11824 240468 11830
rect 240416 11766 240468 11772
rect 241624 9042 241652 338014
rect 241808 335354 241836 338014
rect 242176 336682 242204 338014
rect 241716 335326 241836 335354
rect 241992 336654 242204 336682
rect 241716 14521 241744 335326
rect 241992 316034 242020 336654
rect 242544 336190 242572 338014
rect 242532 336184 242584 336190
rect 242532 336126 242584 336132
rect 242164 335572 242216 335578
rect 242164 335514 242216 335520
rect 241808 316006 242020 316034
rect 241702 14512 241758 14521
rect 241702 14447 241758 14456
rect 241612 9036 241664 9042
rect 241612 8978 241664 8984
rect 240322 8936 240378 8945
rect 240322 8871 240378 8880
rect 240508 6248 240560 6254
rect 240508 6190 240560 6196
rect 240232 3596 240284 3602
rect 240232 3538 240284 3544
rect 240520 480 240548 6190
rect 241808 3738 241836 316006
rect 241796 3732 241848 3738
rect 241796 3674 241848 3680
rect 241702 3360 241758 3369
rect 242176 3330 242204 335514
rect 242256 335436 242308 335442
rect 242256 335378 242308 335384
rect 242268 3398 242296 335378
rect 242900 325780 242952 325786
rect 242900 325722 242952 325728
rect 242912 3806 242940 325722
rect 243004 9110 243032 338014
rect 243084 329180 243136 329186
rect 243084 329122 243136 329128
rect 243096 9178 243124 329122
rect 243280 316034 243308 338014
rect 243648 325786 243676 338014
rect 244016 329186 244044 338014
rect 244004 329180 244056 329186
rect 244004 329122 244056 329128
rect 243636 325780 243688 325786
rect 243636 325722 243688 325728
rect 243188 316006 243308 316034
rect 243188 15910 243216 316006
rect 244384 15978 244412 338014
rect 244752 336258 244780 338014
rect 245120 336682 245148 338014
rect 244844 336654 245148 336682
rect 244740 336252 244792 336258
rect 244740 336194 244792 336200
rect 244844 316034 244872 336654
rect 244924 335640 244976 335646
rect 244924 335582 244976 335588
rect 244476 316006 244872 316034
rect 244372 15972 244424 15978
rect 244372 15914 244424 15920
rect 243176 15904 243228 15910
rect 243176 15846 243228 15852
rect 244476 9246 244504 316006
rect 244464 9240 244516 9246
rect 244464 9182 244516 9188
rect 243084 9172 243136 9178
rect 243084 9114 243136 9120
rect 242992 9104 243044 9110
rect 242992 9046 243044 9052
rect 242900 3800 242952 3806
rect 242900 3742 242952 3748
rect 244096 3596 244148 3602
rect 244096 3538 244148 3544
rect 242900 3460 242952 3466
rect 242900 3402 242952 3408
rect 242256 3392 242308 3398
rect 242256 3334 242308 3340
rect 241702 3295 241758 3304
rect 242164 3324 242216 3330
rect 241716 480 241744 3295
rect 242164 3266 242216 3272
rect 242912 480 242940 3402
rect 244108 480 244136 3538
rect 244936 3262 244964 335582
rect 245856 326874 245884 338014
rect 245948 338014 246100 338042
rect 246224 338014 246468 338042
rect 246592 338014 246836 338042
rect 247052 338014 247112 338042
rect 247236 338014 247480 338042
rect 247604 338014 247848 338042
rect 247972 338014 248216 338042
rect 248524 338014 248584 338042
rect 248708 338014 248952 338042
rect 249076 338014 249320 338042
rect 249444 338014 249688 338042
rect 249996 338014 250056 338042
rect 250180 338014 250424 338042
rect 250548 338014 250792 338042
rect 250916 338014 251160 338042
rect 251376 338014 251528 338042
rect 251652 338014 251896 338042
rect 252020 338014 252264 338042
rect 252632 338014 252784 338042
rect 245844 326868 245896 326874
rect 245844 326810 245896 326816
rect 245844 326664 245896 326670
rect 245844 326606 245896 326612
rect 245752 326392 245804 326398
rect 245752 326334 245804 326340
rect 245660 319252 245712 319258
rect 245660 319194 245712 319200
rect 245672 3874 245700 319194
rect 245764 11898 245792 326334
rect 245856 16046 245884 326606
rect 245948 319258 245976 338014
rect 246224 326398 246252 338014
rect 246212 326392 246264 326398
rect 246212 326334 246264 326340
rect 245936 319252 245988 319258
rect 245936 319194 245988 319200
rect 246592 316034 246620 338014
rect 247052 336025 247080 338014
rect 247038 336016 247094 336025
rect 247038 335951 247094 335960
rect 247236 335354 247264 338014
rect 247144 335326 247264 335354
rect 247040 326392 247092 326398
rect 247040 326334 247092 326340
rect 245948 316006 246620 316034
rect 245948 18630 245976 316006
rect 245936 18624 245988 18630
rect 245936 18566 245988 18572
rect 245844 16040 245896 16046
rect 245844 15982 245896 15988
rect 245752 11892 245804 11898
rect 245752 11834 245804 11840
rect 246396 4140 246448 4146
rect 246396 4082 246448 4088
rect 245660 3868 245712 3874
rect 245660 3810 245712 3816
rect 245200 3528 245252 3534
rect 245200 3470 245252 3476
rect 244924 3256 244976 3262
rect 244924 3198 244976 3204
rect 245212 480 245240 3470
rect 246408 480 246436 4082
rect 247052 3942 247080 326334
rect 247144 13025 247172 335326
rect 247604 316034 247632 338014
rect 247972 326398 248000 338014
rect 247960 326392 248012 326398
rect 247960 326334 248012 326340
rect 247236 316006 247632 316034
rect 247236 18698 247264 316006
rect 247224 18692 247276 18698
rect 247224 18634 247276 18640
rect 248524 13122 248552 338014
rect 248708 335354 248736 338014
rect 249076 336326 249104 338014
rect 249064 336320 249116 336326
rect 249064 336262 249116 336268
rect 248616 335326 248736 335354
rect 248616 18766 248644 335326
rect 249444 316034 249472 338014
rect 249892 326392 249944 326398
rect 249892 326334 249944 326340
rect 249800 323876 249852 323882
rect 249800 323818 249852 323824
rect 248708 316006 249472 316034
rect 248604 18760 248656 18766
rect 248604 18702 248656 18708
rect 248512 13116 248564 13122
rect 248512 13058 248564 13064
rect 247130 13016 247186 13025
rect 247130 12951 247186 12960
rect 248708 6458 248736 316006
rect 249812 6526 249840 323818
rect 249904 13258 249932 326334
rect 249892 13252 249944 13258
rect 249892 13194 249944 13200
rect 249996 13190 250024 338014
rect 250180 316034 250208 338014
rect 250548 323882 250576 338014
rect 250916 326398 250944 338014
rect 250904 326392 250956 326398
rect 250904 326334 250956 326340
rect 251180 326392 251232 326398
rect 251180 326334 251232 326340
rect 250536 323876 250588 323882
rect 250536 323818 250588 323824
rect 250088 316006 250208 316034
rect 250088 18834 250116 316006
rect 250076 18828 250128 18834
rect 250076 18770 250128 18776
rect 249984 13184 250036 13190
rect 249984 13126 250036 13132
rect 251192 6594 251220 326334
rect 251272 322244 251324 322250
rect 251272 322186 251324 322192
rect 251284 19038 251312 322186
rect 251272 19032 251324 19038
rect 251272 18974 251324 18980
rect 251376 18902 251404 338014
rect 251652 326398 251680 338014
rect 251640 326392 251692 326398
rect 251640 326334 251692 326340
rect 252020 322250 252048 338014
rect 252560 336796 252612 336802
rect 252560 336738 252612 336744
rect 252008 322244 252060 322250
rect 252008 322186 252060 322192
rect 251364 18896 251416 18902
rect 251364 18838 251416 18844
rect 252572 6662 252600 336738
rect 252652 326052 252704 326058
rect 252652 325994 252704 326000
rect 252664 19106 252692 325994
rect 252652 19100 252704 19106
rect 252652 19042 252704 19048
rect 252756 18970 252784 338014
rect 252848 338014 253000 338042
rect 253124 338014 253368 338042
rect 253492 338014 253736 338042
rect 253952 338014 254104 338042
rect 254228 338014 254472 338042
rect 254596 338014 254840 338042
rect 254964 338014 255208 338042
rect 255424 338014 255576 338042
rect 255700 338014 255944 338042
rect 256068 338014 256312 338042
rect 256436 338014 256680 338042
rect 256896 338014 257048 338042
rect 257172 338014 257416 338042
rect 257540 338014 257784 338042
rect 258152 338014 258304 338042
rect 252848 336802 252876 338014
rect 252836 336796 252888 336802
rect 252836 336738 252888 336744
rect 253124 326058 253152 338014
rect 253112 326052 253164 326058
rect 253112 325994 253164 326000
rect 253492 316034 253520 338014
rect 252848 316006 253520 316034
rect 252848 20058 252876 316006
rect 252836 20052 252888 20058
rect 252836 19994 252888 20000
rect 252744 18964 252796 18970
rect 252744 18906 252796 18912
rect 253952 6730 253980 338014
rect 254228 335354 254256 338014
rect 254136 335326 254256 335354
rect 254032 330540 254084 330546
rect 254032 330482 254084 330488
rect 254044 6798 254072 330482
rect 254136 19174 254164 335326
rect 254596 316034 254624 338014
rect 254964 330546 254992 338014
rect 254952 330540 255004 330546
rect 254952 330482 255004 330488
rect 255320 330472 255372 330478
rect 255320 330414 255372 330420
rect 254228 316006 254624 316034
rect 254228 20126 254256 316006
rect 254216 20120 254268 20126
rect 254216 20062 254268 20068
rect 254124 19168 254176 19174
rect 254124 19110 254176 19116
rect 255332 6866 255360 330414
rect 255424 14482 255452 338014
rect 255504 330540 255556 330546
rect 255504 330482 255556 330488
rect 255516 14550 255544 330482
rect 255700 316034 255728 338014
rect 256068 330478 256096 338014
rect 256436 330546 256464 338014
rect 256424 330540 256476 330546
rect 256424 330482 256476 330488
rect 256700 330540 256752 330546
rect 256700 330482 256752 330488
rect 256056 330472 256108 330478
rect 256056 330414 256108 330420
rect 255608 316006 255728 316034
rect 255608 20194 255636 316006
rect 255596 20188 255648 20194
rect 255596 20130 255648 20136
rect 255504 14544 255556 14550
rect 255504 14486 255556 14492
rect 255412 14476 255464 14482
rect 255412 14418 255464 14424
rect 256712 9314 256740 330482
rect 256792 330472 256844 330478
rect 256792 330414 256844 330420
rect 256804 14618 256832 330414
rect 256896 20262 256924 338014
rect 257172 330546 257200 338014
rect 257160 330540 257212 330546
rect 257160 330482 257212 330488
rect 257540 330478 257568 338014
rect 258172 330540 258224 330546
rect 258172 330482 258224 330488
rect 257528 330472 257580 330478
rect 257528 330414 257580 330420
rect 256884 20256 256936 20262
rect 256884 20198 256936 20204
rect 258184 14686 258212 330482
rect 258276 20330 258304 338014
rect 258368 338014 258520 338042
rect 258644 338014 258888 338042
rect 259012 338014 259164 338042
rect 258264 20324 258316 20330
rect 258264 20266 258316 20272
rect 258172 14680 258224 14686
rect 258172 14622 258224 14628
rect 256792 14612 256844 14618
rect 256792 14554 256844 14560
rect 258368 9382 258396 338014
rect 258644 330546 258672 338014
rect 259012 336394 259040 338014
rect 259518 337770 259546 338028
rect 259748 338014 259900 338042
rect 260024 338014 260268 338042
rect 260392 338014 260636 338042
rect 260944 338014 261004 338042
rect 261128 338014 261372 338042
rect 261496 338014 261740 338042
rect 261864 338014 262108 338042
rect 262232 338014 262476 338042
rect 262600 338014 262844 338042
rect 262968 338014 263212 338042
rect 263336 338014 263580 338042
rect 263796 338014 263948 338042
rect 264072 338014 264316 338042
rect 264440 338014 264684 338042
rect 259518 337742 259592 337770
rect 259000 336388 259052 336394
rect 259000 336330 259052 336336
rect 258816 335776 258868 335782
rect 258816 335718 258868 335724
rect 258724 335708 258776 335714
rect 258724 335650 258776 335656
rect 258632 330540 258684 330546
rect 258632 330482 258684 330488
rect 258356 9376 258408 9382
rect 258356 9318 258408 9324
rect 256700 9308 256752 9314
rect 256700 9250 256752 9256
rect 255320 6860 255372 6866
rect 255320 6802 255372 6808
rect 254032 6792 254084 6798
rect 254032 6734 254084 6740
rect 253940 6724 253992 6730
rect 253940 6666 253992 6672
rect 252560 6656 252612 6662
rect 252560 6598 252612 6604
rect 251180 6588 251232 6594
rect 251180 6530 251232 6536
rect 249800 6520 249852 6526
rect 249800 6462 249852 6468
rect 248696 6452 248748 6458
rect 248696 6394 248748 6400
rect 258264 6452 258316 6458
rect 258264 6394 258316 6400
rect 254676 6384 254728 6390
rect 254676 6326 254728 6332
rect 247040 3936 247092 3942
rect 247040 3878 247092 3884
rect 252376 3936 252428 3942
rect 252376 3878 252428 3884
rect 248788 3868 248840 3874
rect 248788 3810 248840 3816
rect 247592 3732 247644 3738
rect 247592 3674 247644 3680
rect 247604 480 247632 3674
rect 248800 480 248828 3810
rect 251180 3664 251232 3670
rect 251180 3606 251232 3612
rect 249984 3392 250036 3398
rect 249984 3334 250036 3340
rect 249996 480 250024 3334
rect 251192 480 251220 3606
rect 252388 480 252416 3878
rect 253480 3324 253532 3330
rect 253480 3266 253532 3272
rect 253492 480 253520 3266
rect 254688 480 254716 6326
rect 255872 4072 255924 4078
rect 255872 4014 255924 4020
rect 255884 480 255912 4014
rect 257068 3256 257120 3262
rect 257068 3198 257120 3204
rect 257080 480 257108 3198
rect 258276 480 258304 6394
rect 258736 4690 258764 335650
rect 258724 4684 258776 4690
rect 258724 4626 258776 4632
rect 258828 4622 258856 335718
rect 259460 330472 259512 330478
rect 259460 330414 259512 330420
rect 258816 4616 258868 4622
rect 258816 4558 258868 4564
rect 259472 4010 259500 330414
rect 259564 10305 259592 337742
rect 259644 330540 259696 330546
rect 259644 330482 259696 330488
rect 259656 10334 259684 330482
rect 259748 14754 259776 338014
rect 260024 330478 260052 338014
rect 260392 330546 260420 338014
rect 260380 330540 260432 330546
rect 260380 330482 260432 330488
rect 260012 330472 260064 330478
rect 260012 330414 260064 330420
rect 260944 14822 260972 338014
rect 261128 336462 261156 338014
rect 261116 336456 261168 336462
rect 261116 336398 261168 336404
rect 261496 335354 261524 338014
rect 261576 335844 261628 335850
rect 261576 335786 261628 335792
rect 261404 335326 261524 335354
rect 261024 330540 261076 330546
rect 261024 330482 261076 330488
rect 261036 14890 261064 330482
rect 261404 316034 261432 335326
rect 261588 316034 261616 335786
rect 261864 330546 261892 338014
rect 262232 336530 262260 338014
rect 262220 336524 262272 336530
rect 262220 336466 262272 336472
rect 262220 336048 262272 336054
rect 262220 335990 262272 335996
rect 261852 330540 261904 330546
rect 261852 330482 261904 330488
rect 261128 316006 261432 316034
rect 261496 316006 261616 316034
rect 261024 14884 261076 14890
rect 261024 14826 261076 14832
rect 260932 14816 260984 14822
rect 260932 14758 260984 14764
rect 259736 14748 259788 14754
rect 259736 14690 259788 14696
rect 261128 10402 261156 316006
rect 261116 10396 261168 10402
rect 261116 10338 261168 10344
rect 259644 10328 259696 10334
rect 259550 10296 259606 10305
rect 259644 10270 259696 10276
rect 259550 10231 259606 10240
rect 261496 5914 261524 316006
rect 262232 6914 262260 335990
rect 262600 335354 262628 338014
rect 262864 336184 262916 336190
rect 262864 336126 262916 336132
rect 262324 335326 262628 335354
rect 262324 10470 262352 335326
rect 262404 330540 262456 330546
rect 262404 330482 262456 330488
rect 262416 14958 262444 330482
rect 262404 14952 262456 14958
rect 262404 14894 262456 14900
rect 262312 10464 262364 10470
rect 262312 10406 262364 10412
rect 262232 6886 262536 6914
rect 261760 6520 261812 6526
rect 261760 6462 261812 6468
rect 261484 5908 261536 5914
rect 261484 5850 261536 5856
rect 259460 4004 259512 4010
rect 259460 3946 259512 3952
rect 260656 3800 260708 3806
rect 260656 3742 260708 3748
rect 259460 3188 259512 3194
rect 259460 3130 259512 3136
rect 259472 480 259500 3130
rect 260668 480 260696 3742
rect 261772 480 261800 6462
rect 223918 354 224030 480
rect 223592 326 224030 354
rect 223918 -960 224030 326
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262508 354 262536 6886
rect 262876 4146 262904 336126
rect 262968 330546 262996 338014
rect 263336 335510 263364 338014
rect 263324 335504 263376 335510
rect 263324 335446 263376 335452
rect 262956 330540 263008 330546
rect 262956 330482 263008 330488
rect 263692 327548 263744 327554
rect 263692 327490 263744 327496
rect 263704 15026 263732 327490
rect 263692 15020 263744 15026
rect 263692 14962 263744 14968
rect 263796 13326 263824 338014
rect 264072 327554 264100 338014
rect 264440 336598 264468 338014
rect 265164 336796 265216 336802
rect 265164 336738 265216 336744
rect 264428 336592 264480 336598
rect 264428 336534 264480 336540
rect 264244 336252 264296 336258
rect 264244 336194 264296 336200
rect 264060 327548 264112 327554
rect 264060 327490 264112 327496
rect 263784 13320 263836 13326
rect 263784 13262 263836 13268
rect 264152 4684 264204 4690
rect 264152 4626 264204 4632
rect 262864 4140 262916 4146
rect 262864 4082 262916 4088
rect 264164 480 264192 4626
rect 264256 3398 264284 336194
rect 265072 328840 265124 328846
rect 265072 328782 265124 328788
rect 265084 13462 265112 328782
rect 265176 15094 265204 336738
rect 265164 15088 265216 15094
rect 265164 15030 265216 15036
rect 265072 13456 265124 13462
rect 265072 13398 265124 13404
rect 265268 13394 265296 338150
rect 341168 338150 341412 338178
rect 265360 338014 265420 338042
rect 265544 338014 265788 338042
rect 265912 338014 266156 338042
rect 266464 338014 266524 338042
rect 266648 338014 266892 338042
rect 267016 338014 267260 338042
rect 267384 338014 267628 338042
rect 267844 338014 267996 338042
rect 268120 338014 268364 338042
rect 268488 338014 268732 338042
rect 268856 338014 269100 338042
rect 269224 338014 269468 338042
rect 269592 338014 269836 338042
rect 269960 338014 270204 338042
rect 265360 336802 265388 338014
rect 265348 336796 265400 336802
rect 265348 336738 265400 336744
rect 265544 336122 265572 338014
rect 265624 336388 265676 336394
rect 265624 336330 265676 336336
rect 265532 336116 265584 336122
rect 265532 336058 265584 336064
rect 265256 13388 265308 13394
rect 265256 13330 265308 13336
rect 265348 6588 265400 6594
rect 265348 6530 265400 6536
rect 264244 3392 264296 3398
rect 264244 3334 264296 3340
rect 265360 480 265388 6530
rect 265636 3330 265664 336330
rect 265912 328846 265940 338014
rect 265900 328840 265952 328846
rect 265900 328782 265952 328788
rect 266464 15162 266492 338014
rect 266648 336666 266676 338014
rect 266636 336660 266688 336666
rect 266636 336602 266688 336608
rect 266544 330540 266596 330546
rect 266544 330482 266596 330488
rect 266452 15156 266504 15162
rect 266452 15098 266504 15104
rect 266556 14414 266584 330482
rect 267016 316034 267044 338014
rect 267384 330546 267412 338014
rect 267844 335442 267872 338014
rect 267832 335436 267884 335442
rect 267832 335378 267884 335384
rect 267372 330540 267424 330546
rect 267372 330482 267424 330488
rect 267832 326868 267884 326874
rect 267832 326810 267884 326816
rect 266648 316006 267044 316034
rect 266544 14408 266596 14414
rect 266544 14350 266596 14356
rect 266648 13530 266676 316006
rect 267844 14346 267872 326810
rect 268120 316034 268148 338014
rect 268384 336524 268436 336530
rect 268384 336466 268436 336472
rect 267936 316006 268148 316034
rect 267832 14340 267884 14346
rect 267832 14282 267884 14288
rect 267936 13598 267964 316006
rect 267924 13592 267976 13598
rect 267924 13534 267976 13540
rect 266636 13524 266688 13530
rect 266636 13466 266688 13472
rect 267740 4004 267792 4010
rect 267740 3946 267792 3952
rect 266544 3392 266596 3398
rect 266544 3334 266596 3340
rect 265624 3324 265676 3330
rect 265624 3266 265676 3272
rect 266556 480 266584 3334
rect 267752 480 267780 3946
rect 268396 3262 268424 336466
rect 268488 326874 268516 338014
rect 268856 336734 268884 338014
rect 268844 336728 268896 336734
rect 268844 336670 268896 336676
rect 268568 336320 268620 336326
rect 268568 336262 268620 336268
rect 268476 326868 268528 326874
rect 268476 326810 268528 326816
rect 268580 316034 268608 336262
rect 268488 316006 268608 316034
rect 268384 3256 268436 3262
rect 268384 3198 268436 3204
rect 268488 3194 268516 316006
rect 269224 13666 269252 338014
rect 269592 336682 269620 338014
rect 269316 336654 269620 336682
rect 269316 14278 269344 336654
rect 269396 336116 269448 336122
rect 269396 336058 269448 336064
rect 269408 16574 269436 336058
rect 269960 335578 269988 338014
rect 270558 337770 270586 338028
rect 270696 338014 270940 338042
rect 271064 338014 271216 338042
rect 271340 338014 271584 338042
rect 271952 338014 272104 338042
rect 270558 337742 270632 337770
rect 269948 335572 270000 335578
rect 269948 335514 270000 335520
rect 269408 16546 270080 16574
rect 269304 14272 269356 14278
rect 269304 14214 269356 14220
rect 269212 13660 269264 13666
rect 269212 13602 269264 13608
rect 268844 6656 268896 6662
rect 268844 6598 268896 6604
rect 268476 3188 268528 3194
rect 268476 3130 268528 3136
rect 268856 480 268884 6598
rect 270052 480 270080 16546
rect 270604 13734 270632 337742
rect 270696 16114 270724 338014
rect 271064 335986 271092 338014
rect 271052 335980 271104 335986
rect 271052 335922 271104 335928
rect 271340 316034 271368 338014
rect 271972 330540 272024 330546
rect 271972 330482 272024 330488
rect 270788 316006 271368 316034
rect 270684 16108 270736 16114
rect 270684 16050 270736 16056
rect 270788 13802 270816 316006
rect 271984 16250 272012 330482
rect 271972 16244 272024 16250
rect 271972 16186 272024 16192
rect 272076 16182 272104 338014
rect 272168 338014 272320 338042
rect 272444 338014 272688 338042
rect 272812 338014 273056 338042
rect 273272 338014 273424 338042
rect 273548 338014 273792 338042
rect 273916 338014 274160 338042
rect 274284 338014 274528 338042
rect 274744 338014 274896 338042
rect 275020 338014 275264 338042
rect 275388 338014 275632 338042
rect 275756 338014 276000 338042
rect 276216 338014 276368 338042
rect 276492 338014 276736 338042
rect 276860 338014 277104 338042
rect 272168 335918 272196 338014
rect 272156 335912 272208 335918
rect 272156 335854 272208 335860
rect 272444 316034 272472 338014
rect 272812 330546 272840 338014
rect 273272 335646 273300 338014
rect 273260 335640 273312 335646
rect 273260 335582 273312 335588
rect 272800 330540 272852 330546
rect 272800 330482 272852 330488
rect 273352 330540 273404 330546
rect 273352 330482 273404 330488
rect 272168 316006 272472 316034
rect 272064 16176 272116 16182
rect 272064 16118 272116 16124
rect 270776 13796 270828 13802
rect 270776 13738 270828 13744
rect 270592 13728 270644 13734
rect 270592 13670 270644 13676
rect 272168 13054 272196 316006
rect 272156 13048 272208 13054
rect 272156 12990 272208 12996
rect 273364 7614 273392 330482
rect 273444 330472 273496 330478
rect 273444 330414 273496 330420
rect 273456 10538 273484 330414
rect 273548 16318 273576 338014
rect 273628 336456 273680 336462
rect 273628 336398 273680 336404
rect 273536 16312 273588 16318
rect 273536 16254 273588 16260
rect 273444 10532 273496 10538
rect 273444 10474 273496 10480
rect 273352 7608 273404 7614
rect 273352 7550 273404 7556
rect 272432 6724 272484 6730
rect 272432 6666 272484 6672
rect 271236 4140 271288 4146
rect 271236 4082 271288 4088
rect 271248 480 271276 4082
rect 272444 480 272472 6666
rect 273640 480 273668 336398
rect 273916 330546 273944 338014
rect 273904 330540 273956 330546
rect 273904 330482 273956 330488
rect 274284 330478 274312 338014
rect 274640 330540 274692 330546
rect 274640 330482 274692 330488
rect 274272 330472 274324 330478
rect 274272 330414 274324 330420
rect 274548 7608 274600 7614
rect 274548 7550 274600 7556
rect 274560 3874 274588 7550
rect 274652 4894 274680 330482
rect 274640 4888 274692 4894
rect 274640 4830 274692 4836
rect 274744 4826 274772 338014
rect 275020 335354 275048 338014
rect 274836 335326 275048 335354
rect 274836 7682 274864 335326
rect 275388 316034 275416 338014
rect 275756 330546 275784 338014
rect 276018 336016 276074 336025
rect 276018 335951 276074 335960
rect 275744 330540 275796 330546
rect 275744 330482 275796 330488
rect 274928 316006 275416 316034
rect 274928 17241 274956 316006
rect 274914 17232 274970 17241
rect 274914 17167 274970 17176
rect 276032 11762 276060 335951
rect 276112 330540 276164 330546
rect 276112 330482 276164 330488
rect 276020 11756 276072 11762
rect 276020 11698 276072 11704
rect 274824 7676 274876 7682
rect 274824 7618 274876 7624
rect 275192 7676 275244 7682
rect 275192 7618 275244 7624
rect 274732 4820 274784 4826
rect 274732 4762 274784 4768
rect 274824 4820 274876 4826
rect 274824 4762 274876 4768
rect 274548 3868 274600 3874
rect 274548 3810 274600 3816
rect 274836 480 274864 4762
rect 275204 3942 275232 7618
rect 276020 6792 276072 6798
rect 276020 6734 276072 6740
rect 275192 3936 275244 3942
rect 275192 3878 275244 3884
rect 276032 480 276060 6734
rect 276124 4962 276152 330482
rect 276216 7750 276244 338014
rect 276492 316034 276520 338014
rect 276860 330546 276888 338014
rect 277458 337770 277486 338028
rect 277688 338014 277840 338042
rect 277964 338014 278208 338042
rect 278332 338014 278576 338042
rect 277458 337742 277532 337770
rect 276848 330540 276900 330546
rect 276848 330482 276900 330488
rect 277400 330472 277452 330478
rect 277400 330414 277452 330420
rect 276308 316006 276520 316034
rect 276308 11966 276336 316006
rect 276296 11960 276348 11966
rect 276296 11902 276348 11908
rect 276756 11756 276808 11762
rect 276756 11698 276808 11704
rect 276204 7744 276256 7750
rect 276204 7686 276256 7692
rect 276112 4956 276164 4962
rect 276112 4898 276164 4904
rect 262926 354 263038 480
rect 262508 326 263038 354
rect 262926 -960 263038 326
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 276768 354 276796 11698
rect 277412 6118 277440 330414
rect 277504 9450 277532 337742
rect 277584 330540 277636 330546
rect 277584 330482 277636 330488
rect 277596 9518 277624 330482
rect 277688 12034 277716 338014
rect 277964 330478 277992 338014
rect 278332 330546 278360 338014
rect 278930 337770 278958 338028
rect 279068 338014 279312 338042
rect 279436 338014 279680 338042
rect 279804 338014 280048 338042
rect 280264 338014 280416 338042
rect 280540 338014 280784 338042
rect 280908 338014 281152 338042
rect 281276 338014 281520 338042
rect 281644 338014 281888 338042
rect 282012 338014 282256 338042
rect 282380 338014 282624 338042
rect 278930 337742 279004 337770
rect 278976 330818 279004 337742
rect 278964 330812 279016 330818
rect 278964 330754 279016 330760
rect 279068 330698 279096 338014
rect 278792 330670 279096 330698
rect 278320 330540 278372 330546
rect 278320 330482 278372 330488
rect 277952 330472 278004 330478
rect 277952 330414 278004 330420
rect 277676 12028 277728 12034
rect 277676 11970 277728 11976
rect 277584 9512 277636 9518
rect 277584 9454 277636 9460
rect 277492 9444 277544 9450
rect 277492 9386 277544 9392
rect 277492 7744 277544 7750
rect 277492 7686 277544 7692
rect 277400 6112 277452 6118
rect 277400 6054 277452 6060
rect 277504 4078 277532 7686
rect 278792 6050 278820 330670
rect 278964 330608 279016 330614
rect 278964 330550 279016 330556
rect 278872 330540 278924 330546
rect 278872 330482 278924 330488
rect 278884 17338 278912 330482
rect 278872 17332 278924 17338
rect 278872 17274 278924 17280
rect 278976 17270 279004 330550
rect 279436 330546 279464 338014
rect 279424 330540 279476 330546
rect 279424 330482 279476 330488
rect 279804 316034 279832 338014
rect 280264 330818 280292 338014
rect 280540 335354 280568 338014
rect 280356 335326 280568 335354
rect 280252 330812 280304 330818
rect 280252 330754 280304 330760
rect 280356 330698 280384 335326
rect 279068 316006 279832 316034
rect 280172 330670 280384 330698
rect 279068 19242 279096 316006
rect 279056 19236 279108 19242
rect 279056 19178 279108 19184
rect 280172 17474 280200 330670
rect 280252 330608 280304 330614
rect 280252 330550 280304 330556
rect 280160 17468 280212 17474
rect 280160 17410 280212 17416
rect 280264 17406 280292 330550
rect 280344 330540 280396 330546
rect 280344 330482 280396 330488
rect 280356 17542 280384 330482
rect 280908 316034 280936 338014
rect 281276 330546 281304 338014
rect 281264 330540 281316 330546
rect 281264 330482 281316 330488
rect 281540 329860 281592 329866
rect 281540 329802 281592 329808
rect 280448 316006 280936 316034
rect 280448 19310 280476 316006
rect 280436 19304 280488 19310
rect 280436 19246 280488 19252
rect 281552 17678 281580 329802
rect 281540 17672 281592 17678
rect 281540 17614 281592 17620
rect 281644 17610 281672 338014
rect 282012 316034 282040 338014
rect 282380 329866 282408 338014
rect 282978 337770 283006 338028
rect 283208 338014 283268 338042
rect 283392 338014 283636 338042
rect 283760 338014 284004 338042
rect 284372 338014 284616 338042
rect 282978 337742 283052 337770
rect 282920 330472 282972 330478
rect 282920 330414 282972 330420
rect 282368 329860 282420 329866
rect 282368 329802 282420 329808
rect 281736 316006 282040 316034
rect 281736 18562 281764 316006
rect 281724 18556 281776 18562
rect 281724 18498 281776 18504
rect 281632 17604 281684 17610
rect 281632 17546 281684 17552
rect 280344 17536 280396 17542
rect 280344 17478 280396 17484
rect 280252 17400 280304 17406
rect 280252 17342 280304 17348
rect 278964 17264 279016 17270
rect 278964 17206 279016 17212
rect 282932 7818 282960 330414
rect 283024 10606 283052 337742
rect 283104 330540 283156 330546
rect 283104 330482 283156 330488
rect 283116 10674 283144 330482
rect 283208 12986 283236 338014
rect 283392 330478 283420 338014
rect 283760 330546 283788 338014
rect 284300 336592 284352 336598
rect 284300 336534 284352 336540
rect 283748 330540 283800 330546
rect 283748 330482 283800 330488
rect 283380 330472 283432 330478
rect 283380 330414 283432 330420
rect 283196 12980 283248 12986
rect 283196 12922 283248 12928
rect 283104 10668 283156 10674
rect 283104 10610 283156 10616
rect 283012 10600 283064 10606
rect 283012 10542 283064 10548
rect 282920 7812 282972 7818
rect 282920 7754 282972 7760
rect 283656 7812 283708 7818
rect 283656 7754 283708 7760
rect 279516 6860 279568 6866
rect 279516 6802 279568 6808
rect 278780 6044 278832 6050
rect 278780 5986 278832 5992
rect 278320 4888 278372 4894
rect 278320 4830 278372 4836
rect 277492 4072 277544 4078
rect 277492 4014 277544 4020
rect 278332 480 278360 4830
rect 279528 480 279556 6802
rect 283104 4072 283156 4078
rect 283104 4014 283156 4020
rect 280712 3868 280764 3874
rect 280712 3810 280764 3816
rect 280724 480 280752 3810
rect 281908 3256 281960 3262
rect 281908 3198 281960 3204
rect 281920 480 281948 3198
rect 283116 480 283144 4014
rect 283668 3398 283696 7754
rect 283656 3392 283708 3398
rect 283656 3334 283708 3340
rect 284312 480 284340 336534
rect 284392 330540 284444 330546
rect 284392 330482 284444 330488
rect 284404 7585 284432 330482
rect 284484 330472 284536 330478
rect 284484 330414 284536 330420
rect 284496 10742 284524 330414
rect 284588 12918 284616 338014
rect 284680 338014 284740 338042
rect 284864 338014 285108 338042
rect 285232 338014 285476 338042
rect 284680 16386 284708 338014
rect 284864 330546 284892 338014
rect 284852 330540 284904 330546
rect 284852 330482 284904 330488
rect 285232 330478 285260 338014
rect 285830 337770 285858 338028
rect 286060 338014 286212 338042
rect 286336 338014 286580 338042
rect 286704 338014 286948 338042
rect 287164 338014 287316 338042
rect 287440 338014 287684 338042
rect 287808 338014 288052 338042
rect 288176 338014 288420 338042
rect 288544 338014 288788 338042
rect 288912 338014 289156 338042
rect 289280 338014 289524 338042
rect 289892 338014 290136 338042
rect 285830 337742 285904 337770
rect 285680 330608 285732 330614
rect 285680 330550 285732 330556
rect 285876 330562 285904 337742
rect 286060 330614 286088 338014
rect 286048 330608 286100 330614
rect 285220 330472 285272 330478
rect 285220 330414 285272 330420
rect 284668 16380 284720 16386
rect 284668 16322 284720 16328
rect 284576 12912 284628 12918
rect 284576 12854 284628 12860
rect 284484 10736 284536 10742
rect 284484 10678 284536 10684
rect 285692 7886 285720 330550
rect 285772 330540 285824 330546
rect 285876 330534 285996 330562
rect 286048 330550 286100 330556
rect 286336 330546 286364 338014
rect 285772 330482 285824 330488
rect 285784 10810 285812 330482
rect 285864 330472 285916 330478
rect 285864 330414 285916 330420
rect 285876 16522 285904 330414
rect 285864 16516 285916 16522
rect 285864 16458 285916 16464
rect 285968 16454 285996 330534
rect 286324 330540 286376 330546
rect 286324 330482 286376 330488
rect 286704 330478 286732 338014
rect 287060 330540 287112 330546
rect 287060 330482 287112 330488
rect 286692 330472 286744 330478
rect 286692 330414 286744 330420
rect 285956 16448 286008 16454
rect 285956 16390 286008 16396
rect 285772 10804 285824 10810
rect 285772 10746 285824 10752
rect 287072 8022 287100 330482
rect 287060 8016 287112 8022
rect 287060 7958 287112 7964
rect 287164 7954 287192 338014
rect 287440 335354 287468 338014
rect 287256 335326 287468 335354
rect 287256 10878 287284 335326
rect 287808 316034 287836 338014
rect 288176 330546 288204 338014
rect 288164 330540 288216 330546
rect 288164 330482 288216 330488
rect 287348 316006 287836 316034
rect 287348 16590 287376 316006
rect 287336 16584 287388 16590
rect 287336 16526 287388 16532
rect 288544 10946 288572 338014
rect 288912 335714 288940 338014
rect 288900 335708 288952 335714
rect 288900 335650 288952 335656
rect 289280 316034 289308 338014
rect 289912 330540 289964 330546
rect 289912 330482 289964 330488
rect 288636 316006 289308 316034
rect 288532 10940 288584 10946
rect 288532 10882 288584 10888
rect 287244 10872 287296 10878
rect 287244 10814 287296 10820
rect 288636 8090 288664 316006
rect 289924 8158 289952 330482
rect 290004 330472 290056 330478
rect 290004 330414 290056 330420
rect 290016 10266 290044 330414
rect 290108 11014 290136 338014
rect 290200 338014 290260 338042
rect 290384 338014 290628 338042
rect 290752 338014 290996 338042
rect 291212 338014 291364 338042
rect 291488 338014 291732 338042
rect 291856 338014 292100 338042
rect 292224 338014 292468 338042
rect 292776 338014 292836 338042
rect 292960 338014 293204 338042
rect 293328 338014 293572 338042
rect 293696 338014 293940 338042
rect 294248 338014 294308 338042
rect 294432 338014 294676 338042
rect 294800 338014 295044 338042
rect 295168 338014 295320 338042
rect 295444 338014 295688 338042
rect 295812 338014 296056 338042
rect 296180 338014 296424 338042
rect 290200 335782 290228 338014
rect 290280 336660 290332 336666
rect 290280 336602 290332 336608
rect 290188 335776 290240 335782
rect 290188 335718 290240 335724
rect 290292 316034 290320 336602
rect 290384 330546 290412 338014
rect 290372 330540 290424 330546
rect 290372 330482 290424 330488
rect 290752 330478 290780 338014
rect 290740 330472 290792 330478
rect 290740 330414 290792 330420
rect 290200 316006 290320 316034
rect 290096 11008 290148 11014
rect 290096 10950 290148 10956
rect 290004 10260 290056 10266
rect 290004 10202 290056 10208
rect 289912 8152 289964 8158
rect 289912 8094 289964 8100
rect 288624 8084 288676 8090
rect 288624 8026 288676 8032
rect 287152 7948 287204 7954
rect 287152 7890 287204 7896
rect 285680 7880 285732 7886
rect 285680 7822 285732 7828
rect 284390 7576 284446 7585
rect 284390 7511 284446 7520
rect 286600 6112 286652 6118
rect 286600 6054 286652 6060
rect 285404 4956 285456 4962
rect 285404 4898 285456 4904
rect 285416 480 285444 4898
rect 286612 480 286640 6054
rect 288992 4616 289044 4622
rect 288992 4558 289044 4564
rect 287796 3936 287848 3942
rect 287796 3878 287848 3884
rect 287808 480 287836 3878
rect 289004 480 289032 4558
rect 290200 480 290228 316006
rect 291212 5030 291240 338014
rect 291488 335354 291516 338014
rect 291396 335326 291516 335354
rect 291292 330540 291344 330546
rect 291292 330482 291344 330488
rect 291304 5098 291332 330482
rect 291396 8226 291424 335326
rect 291856 316034 291884 338014
rect 292224 330546 292252 338014
rect 292212 330540 292264 330546
rect 292212 330482 292264 330488
rect 292672 326460 292724 326466
rect 292672 326402 292724 326408
rect 292580 326392 292632 326398
rect 292580 326334 292632 326340
rect 291488 316006 291884 316034
rect 291488 10198 291516 316006
rect 291476 10192 291528 10198
rect 291476 10134 291528 10140
rect 291384 8220 291436 8226
rect 291384 8162 291436 8168
rect 292592 5166 292620 326334
rect 292684 7546 292712 326402
rect 292776 8294 292804 338014
rect 292960 316034 292988 338014
rect 293328 326398 293356 338014
rect 293696 326466 293724 338014
rect 293684 326460 293736 326466
rect 293684 326402 293736 326408
rect 294052 326460 294104 326466
rect 294052 326402 294104 326408
rect 293316 326392 293368 326398
rect 293316 326334 293368 326340
rect 293960 326392 294012 326398
rect 293960 326334 294012 326340
rect 292868 316006 292988 316034
rect 292868 10130 292896 316006
rect 292856 10124 292908 10130
rect 292856 10066 292908 10072
rect 292764 8288 292816 8294
rect 292764 8230 292816 8236
rect 292672 7540 292724 7546
rect 292672 7482 292724 7488
rect 293972 5234 294000 326334
rect 294064 7478 294092 326402
rect 294144 326324 294196 326330
rect 294144 326266 294196 326272
rect 294156 17814 294184 326266
rect 294144 17808 294196 17814
rect 294144 17750 294196 17756
rect 294248 17746 294276 338014
rect 294432 326398 294460 338014
rect 294800 326466 294828 338014
rect 294788 326460 294840 326466
rect 294788 326402 294840 326408
rect 294420 326392 294472 326398
rect 294420 326334 294472 326340
rect 295168 326330 295196 338014
rect 295444 336682 295472 338014
rect 295352 336654 295472 336682
rect 295156 326324 295208 326330
rect 295156 326266 295208 326272
rect 294236 17740 294288 17746
rect 294236 17682 294288 17688
rect 294052 7472 294104 7478
rect 294052 7414 294104 7420
rect 295352 5302 295380 336654
rect 295812 335354 295840 338014
rect 295444 335326 295840 335354
rect 295444 7410 295472 335326
rect 296180 316034 296208 338014
rect 296778 337770 296806 338028
rect 296916 338014 297160 338042
rect 297284 338014 297528 338042
rect 297652 338014 297896 338042
rect 296778 337742 296852 337770
rect 296720 326188 296772 326194
rect 296720 326130 296772 326136
rect 295536 316006 296208 316034
rect 295536 18494 295564 316006
rect 295524 18488 295576 18494
rect 295524 18430 295576 18436
rect 295432 7404 295484 7410
rect 295432 7346 295484 7352
rect 296732 5370 296760 326130
rect 296824 16574 296852 337742
rect 296916 17882 296944 338014
rect 297284 316034 297312 338014
rect 297652 326194 297680 338014
rect 298250 337770 298278 338028
rect 298388 338014 298632 338042
rect 298756 338014 299000 338042
rect 299124 338014 299368 338042
rect 299676 338014 299736 338042
rect 299860 338014 300104 338042
rect 300228 338014 300472 338042
rect 300596 338014 300840 338042
rect 300964 338014 301208 338042
rect 301332 338014 301576 338042
rect 301700 338014 301944 338042
rect 302312 338014 302464 338042
rect 298250 337742 298324 337770
rect 298296 326466 298324 337742
rect 298284 326460 298336 326466
rect 298284 326402 298336 326408
rect 298100 326392 298152 326398
rect 298100 326334 298152 326340
rect 297640 326188 297692 326194
rect 297640 326130 297692 326136
rect 297008 316006 297312 316034
rect 297008 18426 297036 316006
rect 296996 18420 297048 18426
rect 296996 18362 297048 18368
rect 296904 17876 296956 17882
rect 296904 17818 296956 17824
rect 296824 16546 296944 16574
rect 296720 5364 296772 5370
rect 296720 5306 296772 5312
rect 295340 5296 295392 5302
rect 295340 5238 295392 5244
rect 293960 5228 294012 5234
rect 293960 5170 294012 5176
rect 294052 5228 294104 5234
rect 294052 5170 294104 5176
rect 292580 5160 292632 5166
rect 292580 5102 292632 5108
rect 291292 5092 291344 5098
rect 291292 5034 291344 5040
rect 291200 5024 291252 5030
rect 291200 4966 291252 4972
rect 292580 5024 292632 5030
rect 292580 4966 292632 4972
rect 291844 4548 291896 4554
rect 291844 4490 291896 4496
rect 291752 4480 291804 4486
rect 291752 4422 291804 4428
rect 291764 4010 291792 4422
rect 291856 4146 291884 4490
rect 291844 4140 291896 4146
rect 291844 4082 291896 4088
rect 291752 4004 291804 4010
rect 291752 3946 291804 3952
rect 291384 3392 291436 3398
rect 291384 3334 291436 3340
rect 291396 480 291424 3334
rect 292592 480 292620 4966
rect 293684 3324 293736 3330
rect 293684 3266 293736 3272
rect 293696 480 293724 3266
rect 294064 3262 294092 5170
rect 296076 5092 296128 5098
rect 296076 5034 296128 5040
rect 294880 4004 294932 4010
rect 294880 3946 294932 3952
rect 294052 3256 294104 3262
rect 294052 3198 294104 3204
rect 294892 480 294920 3946
rect 296088 480 296116 5034
rect 296916 5001 296944 16546
rect 298112 5438 298140 326334
rect 298388 323626 298416 338014
rect 298468 326460 298520 326466
rect 298468 326402 298520 326408
rect 298204 323598 298416 323626
rect 298204 12102 298232 323598
rect 298480 318794 298508 326402
rect 298756 326398 298784 338014
rect 298744 326392 298796 326398
rect 298744 326334 298796 326340
rect 298296 318766 298508 318794
rect 298296 17950 298324 318766
rect 299124 316034 299152 338014
rect 299572 326460 299624 326466
rect 299572 326402 299624 326408
rect 299480 326392 299532 326398
rect 299480 326334 299532 326340
rect 298388 316006 299152 316034
rect 298284 17944 298336 17950
rect 298284 17886 298336 17892
rect 298388 17202 298416 316006
rect 298376 17196 298428 17202
rect 298376 17138 298428 17144
rect 298192 12096 298244 12102
rect 298192 12038 298244 12044
rect 299296 6044 299348 6050
rect 299296 5986 299348 5992
rect 298100 5432 298152 5438
rect 298100 5374 298152 5380
rect 297180 5364 297232 5370
rect 297180 5306 297232 5312
rect 296902 4992 296958 5001
rect 296902 4927 296958 4936
rect 297192 3738 297220 5306
rect 297730 4856 297786 4865
rect 297730 4791 297786 4800
rect 297180 3732 297232 3738
rect 297180 3674 297232 3680
rect 297744 3602 297772 4791
rect 298468 4140 298520 4146
rect 298468 4082 298520 4088
rect 297732 3596 297784 3602
rect 297732 3538 297784 3544
rect 297272 3120 297324 3126
rect 297272 3062 297324 3068
rect 297284 480 297312 3062
rect 298480 480 298508 4082
rect 299308 3534 299336 5986
rect 299492 5506 299520 326334
rect 299584 12238 299612 326402
rect 299572 12232 299624 12238
rect 299572 12174 299624 12180
rect 299676 12170 299704 338014
rect 299860 326398 299888 338014
rect 299848 326392 299900 326398
rect 299848 326334 299900 326340
rect 300228 316034 300256 338014
rect 300596 326466 300624 338014
rect 300964 335354 300992 338014
rect 300872 335326 300992 335354
rect 300584 326460 300636 326466
rect 300584 326402 300636 326408
rect 299768 316006 300256 316034
rect 299768 17134 299796 316006
rect 299756 17128 299808 17134
rect 299756 17070 299808 17076
rect 299664 12164 299716 12170
rect 299664 12106 299716 12112
rect 299480 5500 299532 5506
rect 299480 5442 299532 5448
rect 299664 5160 299716 5166
rect 299664 5102 299716 5108
rect 299296 3528 299348 3534
rect 299296 3470 299348 3476
rect 299676 480 299704 5102
rect 300872 4758 300900 335326
rect 300952 326392 301004 326398
rect 300952 326334 301004 326340
rect 300964 12306 300992 326334
rect 301332 316034 301360 338014
rect 301700 326398 301728 338014
rect 302240 330608 302292 330614
rect 302240 330550 302292 330556
rect 302436 330562 302464 338014
rect 302620 338014 302680 338042
rect 302804 338014 303048 338042
rect 303172 338014 303416 338042
rect 303632 338014 303784 338042
rect 303908 338014 304152 338042
rect 304276 338014 304520 338042
rect 304644 338014 304888 338042
rect 305196 338014 305256 338042
rect 305380 338014 305624 338042
rect 305748 338014 305992 338042
rect 306116 338014 306360 338042
rect 306668 338014 306728 338042
rect 306852 338014 307096 338042
rect 307220 338014 307372 338042
rect 307496 338014 307740 338042
rect 307864 338014 308108 338042
rect 308232 338014 308476 338042
rect 308600 338014 308844 338042
rect 309212 338014 309456 338042
rect 302620 330614 302648 338014
rect 302608 330608 302660 330614
rect 301688 326392 301740 326398
rect 301688 326334 301740 326340
rect 301056 316006 301360 316034
rect 301056 17066 301084 316006
rect 301044 17060 301096 17066
rect 301044 17002 301096 17008
rect 300952 12300 301004 12306
rect 300952 12242 301004 12248
rect 302252 9586 302280 330550
rect 302332 330540 302384 330546
rect 302436 330534 302556 330562
rect 302608 330550 302660 330556
rect 302804 330546 302832 338014
rect 302332 330482 302384 330488
rect 302344 12374 302372 330482
rect 302424 330472 302476 330478
rect 302424 330414 302476 330420
rect 302436 15774 302464 330414
rect 302528 15842 302556 330534
rect 302792 330540 302844 330546
rect 302792 330482 302844 330488
rect 303172 330478 303200 338014
rect 303160 330472 303212 330478
rect 303160 330414 303212 330420
rect 302516 15836 302568 15842
rect 302516 15778 302568 15784
rect 302424 15768 302476 15774
rect 302424 15710 302476 15716
rect 302332 12368 302384 12374
rect 302332 12310 302384 12316
rect 303632 9654 303660 338014
rect 303908 335354 303936 338014
rect 303816 335326 303936 335354
rect 303712 330540 303764 330546
rect 303712 330482 303764 330488
rect 303620 9648 303672 9654
rect 303620 9590 303672 9596
rect 302240 9580 302292 9586
rect 302240 9522 302292 9528
rect 303724 8906 303752 330482
rect 303816 12442 303844 335326
rect 304276 316034 304304 338014
rect 304644 330546 304672 338014
rect 305000 330608 305052 330614
rect 305000 330550 305052 330556
rect 305196 330562 305224 338014
rect 305380 330614 305408 338014
rect 305644 336728 305696 336734
rect 305644 336670 305696 336676
rect 305368 330608 305420 330614
rect 304632 330540 304684 330546
rect 304632 330482 304684 330488
rect 303908 316006 304304 316034
rect 303908 15706 303936 316006
rect 303896 15700 303948 15706
rect 303896 15642 303948 15648
rect 303804 12436 303856 12442
rect 303804 12378 303856 12384
rect 303712 8900 303764 8906
rect 303712 8842 303764 8848
rect 305012 6225 305040 330550
rect 305092 330540 305144 330546
rect 305196 330534 305316 330562
rect 305368 330550 305420 330556
rect 305092 330482 305144 330488
rect 305104 8838 305132 330482
rect 305184 330472 305236 330478
rect 305184 330414 305236 330420
rect 305196 11626 305224 330414
rect 305288 11694 305316 330534
rect 305276 11688 305328 11694
rect 305276 11630 305328 11636
rect 305184 11620 305236 11626
rect 305184 11562 305236 11568
rect 305092 8832 305144 8838
rect 305092 8774 305144 8780
rect 304998 6216 305054 6225
rect 304998 6151 305054 6160
rect 301504 5432 301556 5438
rect 301504 5374 301556 5380
rect 300860 4752 300912 4758
rect 300860 4694 300912 4700
rect 301516 3670 301544 5374
rect 303160 5296 303212 5302
rect 303160 5238 303212 5244
rect 301504 3664 301556 3670
rect 301504 3606 301556 3612
rect 301964 3528 302016 3534
rect 300766 3496 300822 3505
rect 301964 3470 302016 3476
rect 300766 3431 300822 3440
rect 300780 480 300808 3431
rect 301976 480 302004 3470
rect 303172 480 303200 5238
rect 305552 3664 305604 3670
rect 305552 3606 305604 3612
rect 304356 3596 304408 3602
rect 304356 3538 304408 3544
rect 304368 480 304396 3538
rect 305564 480 305592 3606
rect 305656 3330 305684 336670
rect 305748 330546 305776 338014
rect 305736 330540 305788 330546
rect 305736 330482 305788 330488
rect 306116 330478 306144 338014
rect 306564 336796 306616 336802
rect 306564 336738 306616 336744
rect 306472 330540 306524 330546
rect 306472 330482 306524 330488
rect 306104 330472 306156 330478
rect 306104 330414 306156 330420
rect 306484 8770 306512 330482
rect 306576 11558 306604 336738
rect 306564 11552 306616 11558
rect 306564 11494 306616 11500
rect 306472 8764 306524 8770
rect 306472 8706 306524 8712
rect 306668 5982 306696 338014
rect 306852 330546 306880 338014
rect 307220 336802 307248 338014
rect 307208 336796 307260 336802
rect 307208 336738 307260 336744
rect 307024 335980 307076 335986
rect 307024 335922 307076 335928
rect 306840 330540 306892 330546
rect 306840 330482 306892 330488
rect 306656 5976 306708 5982
rect 306656 5918 306708 5924
rect 306748 3460 306800 3466
rect 306748 3402 306800 3408
rect 305644 3324 305696 3330
rect 305644 3266 305696 3272
rect 306760 480 306788 3402
rect 307036 3126 307064 335922
rect 307116 335776 307168 335782
rect 307116 335718 307168 335724
rect 307128 4078 307156 335718
rect 307496 335714 307524 338014
rect 307484 335708 307536 335714
rect 307484 335650 307536 335656
rect 307208 335640 307260 335646
rect 307208 335582 307260 335588
rect 307116 4072 307168 4078
rect 307116 4014 307168 4020
rect 307220 3806 307248 335582
rect 307864 335354 307892 338014
rect 307772 335326 307892 335354
rect 307772 6186 307800 335326
rect 307852 330540 307904 330546
rect 307852 330482 307904 330488
rect 307864 6322 307892 330482
rect 308232 316034 308260 338014
rect 308600 330546 308628 338014
rect 309232 336796 309284 336802
rect 309232 336738 309284 336744
rect 308588 330540 308640 330546
rect 308588 330482 308640 330488
rect 309140 330472 309192 330478
rect 309140 330414 309192 330420
rect 307956 316006 308260 316034
rect 307956 8974 307984 316006
rect 307944 8968 307996 8974
rect 307944 8910 307996 8916
rect 307852 6316 307904 6322
rect 307852 6258 307904 6264
rect 307760 6180 307812 6186
rect 307760 6122 307812 6128
rect 307208 3800 307260 3806
rect 307208 3742 307260 3748
rect 307944 3392 307996 3398
rect 307944 3334 307996 3340
rect 307024 3120 307076 3126
rect 307024 3062 307076 3068
rect 307956 480 307984 3334
rect 309048 3324 309100 3330
rect 309048 3266 309100 3272
rect 309060 480 309088 3266
rect 309152 3262 309180 330414
rect 309244 3369 309272 336738
rect 309324 330540 309376 330546
rect 309324 330482 309376 330488
rect 309336 4865 309364 330482
rect 309428 6254 309456 338014
rect 309520 338014 309580 338042
rect 309704 338014 309948 338042
rect 310072 338014 310316 338042
rect 310624 338014 310684 338042
rect 310808 338014 311052 338042
rect 311176 338014 311420 338042
rect 311544 338014 311788 338042
rect 311912 338014 312156 338042
rect 312280 338014 312524 338042
rect 312648 338014 312892 338042
rect 313016 338014 313260 338042
rect 313384 338014 313628 338042
rect 313752 338014 313996 338042
rect 314120 338014 314364 338042
rect 309520 336802 309548 338014
rect 309508 336796 309560 336802
rect 309508 336738 309560 336744
rect 309600 336320 309652 336326
rect 309600 336262 309652 336268
rect 309612 335850 309640 336262
rect 309600 335844 309652 335850
rect 309600 335786 309652 335792
rect 309704 330478 309732 338014
rect 310072 330546 310100 338014
rect 310060 330540 310112 330546
rect 310060 330482 310112 330488
rect 309692 330472 309744 330478
rect 309692 330414 309744 330420
rect 309416 6248 309468 6254
rect 309416 6190 309468 6196
rect 310624 6050 310652 338014
rect 310808 336190 310836 338014
rect 310796 336184 310848 336190
rect 310796 336126 310848 336132
rect 311176 335354 311204 338014
rect 311256 335912 311308 335918
rect 311256 335854 311308 335860
rect 311084 335326 311204 335354
rect 310704 329996 310756 330002
rect 310704 329938 310756 329944
rect 310716 7614 310744 329938
rect 311084 316034 311112 335326
rect 311268 316034 311296 335854
rect 311544 330002 311572 338014
rect 311912 336258 311940 338014
rect 311900 336252 311952 336258
rect 311900 336194 311952 336200
rect 311532 329996 311584 330002
rect 311532 329938 311584 329944
rect 311992 326868 312044 326874
rect 311992 326810 312044 326816
rect 310808 316006 311112 316034
rect 311176 316006 311296 316034
rect 310704 7608 310756 7614
rect 310704 7550 310756 7556
rect 310612 6044 310664 6050
rect 310612 5986 310664 5992
rect 310808 5370 310836 316006
rect 310796 5364 310848 5370
rect 310796 5306 310848 5312
rect 309322 4856 309378 4865
rect 309322 4791 309378 4800
rect 310244 3732 310296 3738
rect 310244 3674 310296 3680
rect 309230 3360 309286 3369
rect 309230 3295 309286 3304
rect 309140 3256 309192 3262
rect 309140 3198 309192 3204
rect 310256 480 310284 3674
rect 311176 3466 311204 316006
rect 312004 7682 312032 326810
rect 312280 316034 312308 338014
rect 312544 336388 312596 336394
rect 312544 336330 312596 336336
rect 312096 316006 312308 316034
rect 311992 7676 312044 7682
rect 311992 7618 312044 7624
rect 312096 5438 312124 316006
rect 312084 5432 312136 5438
rect 312084 5374 312136 5380
rect 311440 3800 311492 3806
rect 311440 3742 311492 3748
rect 311164 3460 311216 3466
rect 311164 3402 311216 3408
rect 311452 480 311480 3742
rect 312556 3194 312584 336330
rect 312648 326874 312676 338014
rect 313016 336326 313044 338014
rect 313004 336320 313056 336326
rect 313004 336262 313056 336268
rect 312728 336252 312780 336258
rect 312728 336194 312780 336200
rect 312636 326868 312688 326874
rect 312636 326810 312688 326816
rect 312740 316034 312768 336194
rect 313280 336184 313332 336190
rect 313280 336126 313332 336132
rect 312648 316006 312768 316034
rect 312648 3738 312676 316006
rect 312636 3732 312688 3738
rect 312636 3674 312688 3680
rect 312728 3732 312780 3738
rect 312728 3674 312780 3680
rect 312636 3460 312688 3466
rect 312636 3402 312688 3408
rect 312544 3188 312596 3194
rect 312544 3130 312596 3136
rect 312648 480 312676 3402
rect 312740 3398 312768 3674
rect 313292 3482 313320 336126
rect 313384 6390 313412 338014
rect 313752 316034 313780 338014
rect 314120 336530 314148 338014
rect 314718 337770 314746 338028
rect 314856 338014 315100 338042
rect 315224 338014 315468 338042
rect 315592 338014 315836 338042
rect 316052 338014 316204 338042
rect 316328 338014 316572 338042
rect 316696 338014 316940 338042
rect 317064 338014 317308 338042
rect 317524 338014 317676 338042
rect 317800 338014 318044 338042
rect 318168 338014 318412 338042
rect 318536 338014 318780 338042
rect 318996 338014 319148 338042
rect 319272 338014 319424 338042
rect 319548 338014 319792 338042
rect 319916 338014 320160 338042
rect 320284 338014 320528 338042
rect 320652 338014 320896 338042
rect 321020 338014 321264 338042
rect 321632 338014 321784 338042
rect 314718 337742 314792 337770
rect 314108 336524 314160 336530
rect 314108 336466 314160 336472
rect 313476 316006 313780 316034
rect 313476 7750 313504 316006
rect 313464 7744 313516 7750
rect 313464 7686 313516 7692
rect 314764 6458 314792 337742
rect 314856 335850 314884 338014
rect 315028 336524 315080 336530
rect 315028 336466 315080 336472
rect 314844 335844 314896 335850
rect 314844 335786 314896 335792
rect 314844 330540 314896 330546
rect 314844 330482 314896 330488
rect 314856 6526 314884 330482
rect 314844 6520 314896 6526
rect 314844 6462 314896 6468
rect 314752 6452 314804 6458
rect 314752 6394 314804 6400
rect 313372 6384 313424 6390
rect 313372 6326 313424 6332
rect 313292 3454 313872 3482
rect 312728 3392 312780 3398
rect 312728 3334 312780 3340
rect 313844 480 313872 3454
rect 315040 480 315068 336466
rect 315224 335646 315252 338014
rect 315304 335708 315356 335714
rect 315304 335650 315356 335656
rect 315212 335640 315264 335646
rect 315212 335582 315264 335588
rect 315316 4146 315344 335650
rect 315592 330546 315620 338014
rect 316052 336054 316080 338014
rect 316328 336818 316356 338014
rect 316144 336790 316356 336818
rect 316040 336048 316092 336054
rect 316040 335990 316092 335996
rect 315580 330540 315632 330546
rect 315580 330482 315632 330488
rect 316144 4690 316172 336790
rect 316696 336682 316724 338014
rect 316236 336654 316724 336682
rect 316236 6594 316264 336654
rect 316408 336320 316460 336326
rect 316408 336262 316460 336268
rect 316316 328636 316368 328642
rect 316316 328578 316368 328584
rect 316328 7818 316356 328578
rect 316420 16574 316448 336262
rect 317064 328642 317092 338014
rect 317420 335844 317472 335850
rect 317420 335786 317472 335792
rect 317052 328636 317104 328642
rect 317052 328578 317104 328584
rect 316420 16546 317368 16574
rect 316316 7812 316368 7818
rect 316316 7754 316368 7760
rect 316224 6588 316276 6594
rect 316224 6530 316276 6536
rect 316132 4684 316184 4690
rect 316132 4626 316184 4632
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 316224 4072 316276 4078
rect 316224 4014 316276 4020
rect 316236 480 316264 4014
rect 317340 480 317368 16546
rect 317432 1170 317460 335786
rect 317524 4486 317552 338014
rect 317604 328976 317656 328982
rect 317604 328918 317656 328924
rect 317616 4554 317644 328918
rect 317800 316034 317828 338014
rect 318168 336122 318196 338014
rect 318156 336116 318208 336122
rect 318156 336058 318208 336064
rect 318536 328982 318564 338014
rect 318892 330540 318944 330546
rect 318892 330482 318944 330488
rect 318524 328976 318576 328982
rect 318524 328918 318576 328924
rect 317708 316006 317828 316034
rect 317708 6662 317736 316006
rect 318904 6798 318932 330482
rect 318892 6792 318944 6798
rect 318892 6734 318944 6740
rect 318996 6730 319024 338014
rect 319272 336462 319300 338014
rect 319548 336682 319576 338014
rect 319364 336654 319576 336682
rect 319260 336456 319312 336462
rect 319260 336398 319312 336404
rect 319364 316034 319392 336654
rect 319444 336048 319496 336054
rect 319444 335990 319496 335996
rect 319088 316006 319392 316034
rect 318984 6724 319036 6730
rect 318984 6666 319036 6672
rect 317696 6656 317748 6662
rect 317696 6598 317748 6604
rect 319088 4826 319116 316006
rect 319076 4820 319128 4826
rect 319076 4762 319128 4768
rect 317604 4548 317656 4554
rect 317604 4490 317656 4496
rect 317512 4480 317564 4486
rect 317512 4422 317564 4428
rect 319456 3330 319484 335990
rect 319916 330546 319944 338014
rect 320284 336025 320312 338014
rect 320270 336016 320326 336025
rect 320270 335951 320326 335960
rect 320652 335354 320680 338014
rect 320192 335326 320680 335354
rect 319904 330540 319956 330546
rect 319904 330482 319956 330488
rect 320192 4894 320220 335326
rect 321020 316034 321048 338014
rect 321652 326392 321704 326398
rect 321652 326334 321704 326340
rect 320284 316006 321048 316034
rect 320284 6866 320312 316006
rect 320272 6860 320324 6866
rect 320272 6802 320324 6808
rect 321664 5234 321692 326334
rect 321652 5228 321704 5234
rect 321652 5170 321704 5176
rect 320180 4888 320232 4894
rect 320180 4830 320232 4836
rect 320916 4140 320968 4146
rect 320916 4082 320968 4088
rect 319720 3392 319772 3398
rect 319720 3334 319772 3340
rect 319444 3324 319496 3330
rect 319444 3266 319496 3272
rect 317432 1142 318104 1170
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 277094 -960 277206 326
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318076 354 318104 1142
rect 319732 480 319760 3334
rect 320928 480 320956 4082
rect 321756 3874 321784 338014
rect 321848 338014 322000 338042
rect 322124 338014 322368 338042
rect 322492 338014 322736 338042
rect 323044 338014 323104 338042
rect 323228 338014 323472 338042
rect 323596 338014 323840 338042
rect 323964 338014 324208 338042
rect 324332 338014 324576 338042
rect 324700 338014 324944 338042
rect 325068 338014 325312 338042
rect 325436 338014 325680 338042
rect 325896 338014 326048 338042
rect 326172 338014 326416 338042
rect 326540 338014 326784 338042
rect 327092 338014 327152 338042
rect 327276 338014 327520 338042
rect 327644 338014 327888 338042
rect 328012 338014 328256 338042
rect 328472 338014 328624 338042
rect 328748 338014 328992 338042
rect 329116 338014 329360 338042
rect 329484 338014 329728 338042
rect 330036 338014 330096 338042
rect 330220 338014 330464 338042
rect 330588 338014 330832 338042
rect 330956 338014 331108 338042
rect 331324 338014 331476 338042
rect 331600 338014 331844 338042
rect 331968 338014 332212 338042
rect 332336 338014 332580 338042
rect 332704 338014 332948 338042
rect 333072 338014 333316 338042
rect 333440 338014 333684 338042
rect 321848 326398 321876 338014
rect 322124 335782 322152 338014
rect 322492 336598 322520 338014
rect 322480 336592 322532 336598
rect 322480 336534 322532 336540
rect 322112 335776 322164 335782
rect 322112 335718 322164 335724
rect 321836 326392 321888 326398
rect 321836 326334 321888 326340
rect 322940 326392 322992 326398
rect 322940 326334 322992 326340
rect 322952 3942 322980 326334
rect 323044 4962 323072 338014
rect 323124 323264 323176 323270
rect 323124 323206 323176 323212
rect 323032 4956 323084 4962
rect 323032 4898 323084 4904
rect 323136 4622 323164 323206
rect 323228 6118 323256 338014
rect 323596 326398 323624 338014
rect 323584 326392 323636 326398
rect 323584 326334 323636 326340
rect 323964 323270 323992 338014
rect 324332 336666 324360 338014
rect 324320 336660 324372 336666
rect 324320 336602 324372 336608
rect 324700 336394 324728 338014
rect 324688 336388 324740 336394
rect 324688 336330 324740 336336
rect 323952 323264 324004 323270
rect 323952 323206 324004 323212
rect 325068 316034 325096 338014
rect 325436 336734 325464 338014
rect 325424 336728 325476 336734
rect 325424 336670 325476 336676
rect 325896 328454 325924 338014
rect 326172 335354 326200 338014
rect 326540 335986 326568 338014
rect 326528 335980 326580 335986
rect 326528 335922 326580 335928
rect 327092 335714 327120 338014
rect 327080 335708 327132 335714
rect 327080 335650 327132 335656
rect 325804 328426 325924 328454
rect 325988 335326 326200 335354
rect 325804 323762 325832 328426
rect 325804 323734 325924 323762
rect 325792 323604 325844 323610
rect 325792 323546 325844 323552
rect 324516 316006 325096 316034
rect 323216 6112 323268 6118
rect 323216 6054 323268 6060
rect 324516 5030 324544 316006
rect 325804 5098 325832 323546
rect 325792 5092 325844 5098
rect 325792 5034 325844 5040
rect 324504 5024 324556 5030
rect 324504 4966 324556 4972
rect 323124 4616 323176 4622
rect 323124 4558 323176 4564
rect 325896 4010 325924 323734
rect 325988 323610 326016 335326
rect 327172 326392 327224 326398
rect 327172 326334 327224 326340
rect 325976 323604 326028 323610
rect 325976 323546 326028 323552
rect 325884 4004 325936 4010
rect 325884 3946 325936 3952
rect 322940 3936 322992 3942
rect 322940 3878 322992 3884
rect 325608 3936 325660 3942
rect 325608 3878 325660 3884
rect 321744 3868 321796 3874
rect 321744 3810 321796 3816
rect 323308 3324 323360 3330
rect 323308 3266 323360 3272
rect 322112 3120 322164 3126
rect 322112 3062 322164 3068
rect 322124 480 322152 3062
rect 323320 480 323348 3266
rect 324412 3256 324464 3262
rect 324412 3198 324464 3204
rect 324424 480 324452 3198
rect 325620 480 325648 3878
rect 326804 3868 326856 3874
rect 326804 3810 326856 3816
rect 326816 480 326844 3810
rect 327184 3505 327212 326334
rect 327276 5166 327304 338014
rect 327644 326398 327672 338014
rect 327632 326392 327684 326398
rect 327632 326334 327684 326340
rect 328012 316034 328040 338014
rect 328472 320890 328500 338014
rect 328748 321554 328776 338014
rect 328564 321526 328776 321554
rect 328460 320884 328512 320890
rect 328460 320826 328512 320832
rect 327368 316006 328040 316034
rect 327264 5160 327316 5166
rect 327264 5102 327316 5108
rect 327368 3534 327396 316006
rect 328564 3602 328592 321526
rect 328644 320884 328696 320890
rect 328644 320826 328696 320832
rect 328656 5302 328684 320826
rect 329116 316034 329144 338014
rect 329484 335918 329512 338014
rect 329472 335912 329524 335918
rect 329472 335854 329524 335860
rect 329932 326392 329984 326398
rect 329932 326334 329984 326340
rect 328748 316006 329144 316034
rect 328644 5296 328696 5302
rect 328644 5238 328696 5244
rect 328748 3670 328776 316006
rect 329944 3806 329972 326334
rect 329932 3800 329984 3806
rect 329932 3742 329984 3748
rect 330036 3738 330064 338014
rect 330220 336054 330248 338014
rect 330588 336258 330616 338014
rect 330576 336252 330628 336258
rect 330576 336194 330628 336200
rect 330208 336048 330260 336054
rect 330208 335990 330260 335996
rect 330208 335368 330260 335374
rect 330208 335310 330260 335316
rect 330220 16574 330248 335310
rect 330956 326398 330984 338014
rect 331220 336456 331272 336462
rect 331220 336398 331272 336404
rect 330944 326392 330996 326398
rect 330944 326334 330996 326340
rect 330220 16546 330432 16574
rect 330024 3732 330076 3738
rect 330024 3674 330076 3680
rect 328736 3664 328788 3670
rect 328736 3606 328788 3612
rect 328552 3596 328604 3602
rect 328552 3538 328604 3544
rect 327356 3528 327408 3534
rect 327170 3496 327226 3505
rect 327356 3470 327408 3476
rect 327170 3431 327226 3440
rect 328000 3188 328052 3194
rect 328000 3130 328052 3136
rect 328012 480 328040 3130
rect 329196 3052 329248 3058
rect 329196 2994 329248 3000
rect 329208 480 329236 2994
rect 330404 480 330432 16546
rect 318494 354 318606 480
rect 318076 326 318606 354
rect 318494 -960 318606 326
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331232 354 331260 336398
rect 331324 3466 331352 338014
rect 331600 336190 331628 338014
rect 331968 336530 331996 338014
rect 331956 336524 332008 336530
rect 331956 336466 332008 336472
rect 331588 336184 331640 336190
rect 331588 336126 331640 336132
rect 332336 316034 332364 338014
rect 332704 336326 332732 338014
rect 332692 336320 332744 336326
rect 332692 336262 332744 336268
rect 333072 335850 333100 338014
rect 333060 335844 333112 335850
rect 333060 335786 333112 335792
rect 333440 316034 333468 338014
rect 334038 337770 334066 338028
rect 334176 338014 334420 338042
rect 334544 338014 334788 338042
rect 334912 338014 335156 338042
rect 335372 338014 335524 338042
rect 335648 338014 335892 338042
rect 336016 338014 336260 338042
rect 336384 338014 336628 338042
rect 336752 338014 336996 338042
rect 337120 338014 337364 338042
rect 337488 338014 337732 338042
rect 337856 338014 338100 338042
rect 338224 338014 338468 338042
rect 338592 338014 338836 338042
rect 338960 338014 339204 338042
rect 339572 338014 339724 338042
rect 334038 337742 334112 337770
rect 333980 330540 334032 330546
rect 333980 330482 334032 330488
rect 331416 316006 332364 316034
rect 332888 316006 333468 316034
rect 331416 4078 331444 316006
rect 331404 4072 331456 4078
rect 331404 4014 331456 4020
rect 332692 3596 332744 3602
rect 332692 3538 332744 3544
rect 331312 3460 331364 3466
rect 331312 3402 331364 3408
rect 332704 480 332732 3538
rect 332888 3398 332916 316006
rect 333888 4140 333940 4146
rect 333888 4082 333940 4088
rect 332876 3392 332928 3398
rect 332876 3334 332928 3340
rect 333900 480 333928 4082
rect 333992 3330 334020 330482
rect 334084 4078 334112 337742
rect 334072 4072 334124 4078
rect 334072 4014 334124 4020
rect 333980 3324 334032 3330
rect 333980 3266 334032 3272
rect 334176 3126 334204 338014
rect 334544 330546 334572 338014
rect 334532 330540 334584 330546
rect 334532 330482 334584 330488
rect 334912 316034 334940 338014
rect 334268 316006 334940 316034
rect 334268 3262 334296 316006
rect 335372 3942 335400 338014
rect 335648 336682 335676 338014
rect 335464 336654 335676 336682
rect 335360 3936 335412 3942
rect 335360 3878 335412 3884
rect 335464 3874 335492 336654
rect 336016 335354 336044 338014
rect 335556 335326 336044 335354
rect 335452 3868 335504 3874
rect 335452 3810 335504 3816
rect 335084 3732 335136 3738
rect 335084 3674 335136 3680
rect 334256 3256 334308 3262
rect 334256 3198 334308 3204
rect 334164 3120 334216 3126
rect 334164 3062 334216 3068
rect 335096 480 335124 3674
rect 335556 3194 335584 335326
rect 336384 316034 336412 338014
rect 336752 335374 336780 338014
rect 337120 336462 337148 338014
rect 337108 336456 337160 336462
rect 337108 336398 337160 336404
rect 336740 335368 336792 335374
rect 336740 335310 336792 335316
rect 336832 330540 336884 330546
rect 336832 330482 336884 330488
rect 335648 316006 336412 316034
rect 335544 3188 335596 3194
rect 335544 3130 335596 3136
rect 335648 3058 335676 316006
rect 336844 4146 336872 330482
rect 337488 316034 337516 338014
rect 337856 330546 337884 338014
rect 338224 336682 338252 338014
rect 338132 336654 338252 336682
rect 337844 330540 337896 330546
rect 337844 330482 337896 330488
rect 336936 316006 337516 316034
rect 336832 4140 336884 4146
rect 336832 4082 336884 4088
rect 336936 3602 336964 316006
rect 338132 3738 338160 336654
rect 338592 335354 338620 338014
rect 338224 335326 338620 335354
rect 338120 3732 338172 3738
rect 338120 3674 338172 3680
rect 336924 3596 336976 3602
rect 336924 3538 336976 3544
rect 337476 3460 337528 3466
rect 337476 3402 337528 3408
rect 336280 3324 336332 3330
rect 336280 3266 336332 3272
rect 335636 3052 335688 3058
rect 335636 2994 335688 3000
rect 336292 480 336320 3266
rect 337488 480 337516 3402
rect 338224 3330 338252 335326
rect 338960 316034 338988 338014
rect 339696 330818 339724 338014
rect 339788 338014 339940 338042
rect 340064 338014 340308 338042
rect 340676 338014 340828 338042
rect 339684 330812 339736 330818
rect 339684 330754 339736 330760
rect 339788 330698 339816 338014
rect 338316 316006 338988 316034
rect 339512 330670 339816 330698
rect 338316 3466 338344 316006
rect 338304 3460 338356 3466
rect 338304 3402 338356 3408
rect 338212 3324 338264 3330
rect 338212 3266 338264 3272
rect 338672 3324 338724 3330
rect 338672 3266 338724 3272
rect 338684 480 338712 3266
rect 331558 354 331670 480
rect 331232 326 331670 354
rect 331558 -960 331670 326
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339512 354 339540 330670
rect 339684 330608 339736 330614
rect 339684 330550 339736 330556
rect 339592 330540 339644 330546
rect 339592 330482 339644 330488
rect 339604 3194 339632 330482
rect 339696 3330 339724 330550
rect 340064 330546 340092 338014
rect 340800 336734 340828 338014
rect 341030 337822 341058 338028
rect 341018 337816 341070 337822
rect 341018 337758 341070 337764
rect 340788 336728 340840 336734
rect 340788 336670 340840 336676
rect 340052 330540 340104 330546
rect 340052 330482 340104 330488
rect 341064 330540 341116 330546
rect 341064 330482 341116 330488
rect 340972 330472 341024 330478
rect 340972 330414 341024 330420
rect 340984 3942 341012 330414
rect 340972 3936 341024 3942
rect 340972 3878 341024 3884
rect 341076 3738 341104 330482
rect 341064 3732 341116 3738
rect 341064 3674 341116 3680
rect 339684 3324 339736 3330
rect 339684 3266 339736 3272
rect 341168 3194 341196 338150
rect 341536 338014 341780 338042
rect 341904 338014 342148 338042
rect 342456 338014 342516 338042
rect 342640 338014 342884 338042
rect 343008 338014 343160 338042
rect 343284 338014 343528 338042
rect 343744 338014 343896 338042
rect 344020 338014 344264 338042
rect 344388 338014 344632 338042
rect 344756 338014 345000 338042
rect 345308 338014 345368 338042
rect 345492 338014 345736 338042
rect 345860 338014 346104 338042
rect 346412 338014 346472 338042
rect 346596 338014 346840 338042
rect 346964 338014 347208 338042
rect 347576 338014 347728 338042
rect 341248 337816 341300 337822
rect 341248 337758 341300 337764
rect 339592 3188 339644 3194
rect 339592 3130 339644 3136
rect 340972 3188 341024 3194
rect 340972 3130 341024 3136
rect 341156 3188 341208 3194
rect 341156 3130 341208 3136
rect 340984 480 341012 3130
rect 341260 3058 341288 337758
rect 341340 336728 341392 336734
rect 341340 336670 341392 336676
rect 341352 16574 341380 336670
rect 341536 330546 341564 338014
rect 341524 330540 341576 330546
rect 341524 330482 341576 330488
rect 341904 330478 341932 338014
rect 342456 330818 342484 338014
rect 342640 335354 342668 338014
rect 342548 335326 342668 335354
rect 342444 330812 342496 330818
rect 342444 330754 342496 330760
rect 342548 330698 342576 335326
rect 342272 330670 342576 330698
rect 341892 330472 341944 330478
rect 341892 330414 341944 330420
rect 341352 16546 342208 16574
rect 341248 3052 341300 3058
rect 341248 2994 341300 3000
rect 342180 480 342208 16546
rect 342272 3330 342300 330670
rect 342444 330608 342496 330614
rect 342444 330550 342496 330556
rect 342352 330540 342404 330546
rect 342352 330482 342404 330488
rect 342260 3324 342312 3330
rect 342260 3266 342312 3272
rect 342364 2990 342392 330482
rect 342456 3126 342484 330550
rect 343008 330546 343036 338014
rect 342996 330540 343048 330546
rect 342996 330482 343048 330488
rect 343284 316034 343312 338014
rect 343640 330540 343692 330546
rect 343640 330482 343692 330488
rect 342548 316006 343312 316034
rect 342548 3398 342576 316006
rect 343652 3466 343680 330482
rect 343744 3534 343772 338014
rect 344020 335354 344048 338014
rect 343836 335326 344048 335354
rect 343836 4078 343864 335326
rect 344388 316034 344416 338014
rect 344756 330546 344784 338014
rect 345308 336258 345336 338014
rect 345296 336252 345348 336258
rect 345296 336194 345348 336200
rect 344744 330540 344796 330546
rect 344744 330482 344796 330488
rect 345020 330540 345072 330546
rect 345020 330482 345072 330488
rect 343928 316006 344416 316034
rect 343824 4072 343876 4078
rect 343824 4014 343876 4020
rect 343928 3874 343956 316006
rect 343916 3868 343968 3874
rect 343916 3810 343968 3816
rect 343732 3528 343784 3534
rect 343732 3470 343784 3476
rect 343640 3460 343692 3466
rect 343640 3402 343692 3408
rect 342536 3392 342588 3398
rect 342536 3334 342588 3340
rect 345032 3330 345060 330482
rect 345492 316034 345520 338014
rect 345860 330546 345888 338014
rect 346412 336666 346440 338014
rect 346400 336660 346452 336666
rect 346400 336602 346452 336608
rect 346596 335354 346624 338014
rect 346412 335326 346624 335354
rect 345848 330540 345900 330546
rect 345848 330482 345900 330488
rect 345124 316006 345520 316034
rect 345124 4010 345152 316006
rect 345112 4004 345164 4010
rect 345112 3946 345164 3952
rect 345756 3732 345808 3738
rect 345756 3674 345808 3680
rect 345020 3324 345072 3330
rect 345020 3266 345072 3272
rect 344560 3188 344612 3194
rect 344560 3130 344612 3136
rect 342444 3120 342496 3126
rect 342444 3062 342496 3068
rect 343364 3052 343416 3058
rect 343364 2994 343416 3000
rect 342352 2984 342404 2990
rect 342352 2926 342404 2932
rect 343376 480 343404 2994
rect 344572 480 344600 3130
rect 345768 480 345796 3674
rect 346412 3398 346440 335326
rect 346964 316034 346992 338014
rect 347700 336394 347728 338014
rect 347792 338014 347944 338042
rect 348068 338014 348312 338042
rect 348620 338014 348680 338042
rect 348804 338014 349048 338042
rect 349172 338014 349416 338042
rect 349784 338014 350028 338042
rect 350152 338014 350396 338042
rect 347688 336388 347740 336394
rect 347688 336330 347740 336336
rect 346504 316006 346992 316034
rect 346504 4146 346532 316006
rect 346492 4140 346544 4146
rect 346492 4082 346544 4088
rect 346952 3936 347004 3942
rect 346952 3878 347004 3884
rect 346400 3392 346452 3398
rect 346400 3334 346452 3340
rect 346964 480 346992 3878
rect 347792 3738 347820 338014
rect 348068 335354 348096 338014
rect 348620 336326 348648 338014
rect 348608 336320 348660 336326
rect 348608 336262 348660 336268
rect 347884 335326 348096 335354
rect 347884 3942 347912 335326
rect 348804 316034 348832 338014
rect 347976 316006 348832 316034
rect 347872 3936 347924 3942
rect 347872 3878 347924 3884
rect 347976 3806 348004 316006
rect 347964 3800 348016 3806
rect 347964 3742 348016 3748
rect 347780 3732 347832 3738
rect 347780 3674 347832 3680
rect 349172 3670 349200 338014
rect 350000 336054 350028 338014
rect 350368 336190 350396 338014
rect 350460 338014 350520 338042
rect 350828 338014 350888 338042
rect 351012 338014 351256 338042
rect 351624 338014 351868 338042
rect 350356 336184 350408 336190
rect 350356 336126 350408 336132
rect 349988 336048 350040 336054
rect 349988 335990 350040 335996
rect 350460 335374 350488 338014
rect 350828 335782 350856 338014
rect 350816 335776 350868 335782
rect 350816 335718 350868 335724
rect 350448 335368 350500 335374
rect 350448 335310 350500 335316
rect 351012 316034 351040 338014
rect 351840 335442 351868 338014
rect 351978 337770 352006 338028
rect 352360 338014 352604 338042
rect 351978 337742 352052 337770
rect 351828 335436 351880 335442
rect 351828 335378 351880 335384
rect 351920 330540 351972 330546
rect 351920 330482 351972 330488
rect 350552 316006 351040 316034
rect 349160 3664 349212 3670
rect 349160 3606 349212 3612
rect 350552 3602 350580 316006
rect 351932 5302 351960 330482
rect 352024 5370 352052 337742
rect 352576 336122 352604 338014
rect 352668 338014 352728 338042
rect 352852 338014 353096 338042
rect 353312 338014 353464 338042
rect 353772 338014 353832 338042
rect 353956 338014 354200 338042
rect 354324 338014 354568 338042
rect 354876 338014 354936 338042
rect 355060 338014 355212 338042
rect 355580 338014 355824 338042
rect 352564 336116 352616 336122
rect 352564 336058 352616 336064
rect 352668 335510 352696 338014
rect 352656 335504 352708 335510
rect 352656 335446 352708 335452
rect 352852 330546 352880 338014
rect 352840 330540 352892 330546
rect 352840 330482 352892 330488
rect 352012 5364 352064 5370
rect 352012 5306 352064 5312
rect 351920 5296 351972 5302
rect 351920 5238 351972 5244
rect 350540 3596 350592 3602
rect 350540 3538 350592 3544
rect 353312 3534 353340 338014
rect 353772 336530 353800 338014
rect 353760 336524 353812 336530
rect 353760 336466 353812 336472
rect 353956 331214 353984 338014
rect 353404 331186 353984 331214
rect 353404 5234 353432 331186
rect 354324 316034 354352 338014
rect 354876 335646 354904 338014
rect 354864 335640 354916 335646
rect 354864 335582 354916 335588
rect 355060 316034 355088 338014
rect 355796 336462 355824 338014
rect 355888 338014 355948 338042
rect 356164 338014 356316 338042
rect 356684 338014 356928 338042
rect 357052 338014 357204 338042
rect 355888 336598 355916 338014
rect 355876 336592 355928 336598
rect 355876 336534 355928 336540
rect 355784 336456 355836 336462
rect 355784 336398 355836 336404
rect 355416 336252 355468 336258
rect 355416 336194 355468 336200
rect 355324 335368 355376 335374
rect 355324 335310 355376 335316
rect 353496 316006 354352 316034
rect 354692 316006 355088 316034
rect 353392 5228 353444 5234
rect 353392 5170 353444 5176
rect 353496 5166 353524 316006
rect 353484 5160 353536 5166
rect 353484 5102 353536 5108
rect 354692 5098 354720 316006
rect 354680 5092 354732 5098
rect 354680 5034 354732 5040
rect 354036 4072 354088 4078
rect 354036 4014 354088 4020
rect 352840 3528 352892 3534
rect 352840 3470 352892 3476
rect 353300 3528 353352 3534
rect 353300 3470 353352 3476
rect 351644 3256 351696 3262
rect 351644 3198 351696 3204
rect 349252 3188 349304 3194
rect 349252 3130 349304 3136
rect 348056 3120 348108 3126
rect 348056 3062 348108 3068
rect 348068 480 348096 3062
rect 349264 480 349292 3130
rect 350448 3052 350500 3058
rect 350448 2994 350500 3000
rect 350460 480 350488 2994
rect 351656 480 351684 3198
rect 352852 480 352880 3470
rect 354048 480 354076 4014
rect 355232 3868 355284 3874
rect 355232 3810 355284 3816
rect 355244 480 355272 3810
rect 355336 3194 355364 335310
rect 355428 3398 355456 336194
rect 356060 330540 356112 330546
rect 356060 330482 356112 330488
rect 356072 4962 356100 330482
rect 356164 5030 356192 338014
rect 356900 336258 356928 338014
rect 356888 336252 356940 336258
rect 356888 336194 356940 336200
rect 357176 335850 357204 338014
rect 357268 338014 357420 338042
rect 357544 338014 357788 338042
rect 357912 338014 358156 338042
rect 358280 338014 358524 338042
rect 358832 338014 358892 338042
rect 359016 338014 359260 338042
rect 359384 338014 359628 338042
rect 359996 338014 360148 338042
rect 357164 335844 357216 335850
rect 357164 335786 357216 335792
rect 356704 335436 356756 335442
rect 356704 335378 356756 335384
rect 356152 5024 356204 5030
rect 356152 4966 356204 4972
rect 356060 4956 356112 4962
rect 356060 4898 356112 4904
rect 356716 3874 356744 335378
rect 357268 330546 357296 338014
rect 357544 331214 357572 338014
rect 357452 331186 357572 331214
rect 357256 330540 357308 330546
rect 357256 330482 357308 330488
rect 356704 3868 356756 3874
rect 356704 3810 356756 3816
rect 356336 3460 356388 3466
rect 356336 3402 356388 3408
rect 355416 3392 355468 3398
rect 355416 3334 355468 3340
rect 355324 3188 355376 3194
rect 355324 3130 355376 3136
rect 356348 480 356376 3402
rect 357452 3126 357480 331186
rect 357532 330540 357584 330546
rect 357532 330482 357584 330488
rect 357544 4826 357572 330482
rect 357912 316034 357940 338014
rect 358084 336660 358136 336666
rect 358084 336602 358136 336608
rect 357636 316006 357940 316034
rect 357636 4894 357664 316006
rect 357624 4888 357676 4894
rect 357624 4830 357676 4836
rect 357532 4820 357584 4826
rect 357532 4762 357584 4768
rect 357532 3392 357584 3398
rect 357532 3334 357584 3340
rect 357440 3120 357492 3126
rect 357440 3062 357492 3068
rect 357544 480 357572 3334
rect 358096 3058 358124 336602
rect 358176 335504 358228 335510
rect 358176 335446 358228 335452
rect 358188 4078 358216 335446
rect 358280 330546 358308 338014
rect 358832 335918 358860 338014
rect 358820 335912 358872 335918
rect 358820 335854 358872 335860
rect 359016 331214 359044 338014
rect 358832 331186 359044 331214
rect 358268 330540 358320 330546
rect 358268 330482 358320 330488
rect 358832 4486 358860 331186
rect 359384 316034 359412 338014
rect 360120 336666 360148 338014
rect 360212 338014 360364 338042
rect 360488 338014 360732 338042
rect 361040 338014 361100 338042
rect 361224 338014 361468 338042
rect 361684 338014 361836 338042
rect 361960 338014 362204 338042
rect 362328 338014 362572 338042
rect 362696 338014 362940 338042
rect 363248 338014 363308 338042
rect 363432 338014 363676 338042
rect 363800 338014 364044 338042
rect 364352 338014 364412 338042
rect 364536 338014 364780 338042
rect 364904 338014 365148 338042
rect 365516 338014 365668 338042
rect 360108 336660 360160 336666
rect 360108 336602 360160 336608
rect 358924 316006 359412 316034
rect 358924 4554 358952 316006
rect 360212 4622 360240 338014
rect 360488 335354 360516 338014
rect 361040 336025 361068 338014
rect 361026 336016 361082 336025
rect 361026 335951 361082 335960
rect 360304 335326 360516 335354
rect 360304 6254 360332 335326
rect 361224 316034 361252 338014
rect 361580 336728 361632 336734
rect 361580 336670 361632 336676
rect 360396 316006 361252 316034
rect 360292 6248 360344 6254
rect 360292 6190 360344 6196
rect 360396 6186 360424 316006
rect 360384 6180 360436 6186
rect 360384 6122 360436 6128
rect 361592 5438 361620 336670
rect 361684 5846 361712 338014
rect 361764 336796 361816 336802
rect 361764 336738 361816 336744
rect 361776 5914 361804 336738
rect 361960 336734 361988 338014
rect 362328 336802 362356 338014
rect 362316 336796 362368 336802
rect 362316 336738 362368 336744
rect 361948 336728 362000 336734
rect 362696 336682 362724 338014
rect 361948 336670 362000 336676
rect 362052 336654 362724 336682
rect 362052 316034 362080 336654
rect 362132 336524 362184 336530
rect 362132 336466 362184 336472
rect 362144 325694 362172 336466
rect 362316 336388 362368 336394
rect 362316 336330 362368 336336
rect 362144 325666 362264 325694
rect 361868 316006 362080 316034
rect 361868 8770 361896 316006
rect 361856 8764 361908 8770
rect 361856 8706 361908 8712
rect 361764 5908 361816 5914
rect 361764 5850 361816 5856
rect 361672 5840 361724 5846
rect 361672 5782 361724 5788
rect 361580 5432 361632 5438
rect 361580 5374 361632 5380
rect 360200 4616 360252 4622
rect 360200 4558 360252 4564
rect 358912 4548 358964 4554
rect 358912 4490 358964 4496
rect 358820 4480 358872 4486
rect 358820 4422 358872 4428
rect 361764 4208 361816 4214
rect 361764 4150 361816 4156
rect 358176 4072 358228 4078
rect 358176 4014 358228 4020
rect 358728 4004 358780 4010
rect 358728 3946 358780 3952
rect 358084 3052 358136 3058
rect 358084 2994 358136 3000
rect 358740 480 358768 3946
rect 361776 3942 361804 4150
rect 361856 4140 361908 4146
rect 361856 4082 361908 4088
rect 361868 3942 361896 4082
rect 359464 3936 359516 3942
rect 359464 3878 359516 3884
rect 361764 3936 361816 3942
rect 361764 3878 361816 3884
rect 361856 3936 361908 3942
rect 361856 3878 361908 3884
rect 359476 3466 359504 3878
rect 361488 3868 361540 3874
rect 361488 3810 361540 3816
rect 359464 3460 359516 3466
rect 359464 3402 359516 3408
rect 361500 3194 361528 3810
rect 362236 3330 362264 325666
rect 362328 4146 362356 336330
rect 363248 335986 363276 338014
rect 363236 335980 363288 335986
rect 363236 335922 363288 335928
rect 363432 335354 363460 338014
rect 363604 335776 363656 335782
rect 363604 335718 363656 335724
rect 362972 335326 363460 335354
rect 362972 5982 363000 335326
rect 363052 330540 363104 330546
rect 363052 330482 363104 330488
rect 363064 12918 363092 330482
rect 363052 12912 363104 12918
rect 363052 12854 363104 12860
rect 362960 5976 363012 5982
rect 362960 5918 363012 5924
rect 362316 4140 362368 4146
rect 362316 4082 362368 4088
rect 363512 3936 363564 3942
rect 363512 3878 363564 3884
rect 362224 3324 362276 3330
rect 362224 3266 362276 3272
rect 362316 3256 362368 3262
rect 362316 3198 362368 3204
rect 361488 3188 361540 3194
rect 361488 3130 361540 3136
rect 361120 3052 361172 3058
rect 361120 2994 361172 3000
rect 359924 2984 359976 2990
rect 359924 2926 359976 2932
rect 359936 480 359964 2926
rect 361132 480 361160 2994
rect 362328 480 362356 3198
rect 363524 480 363552 3878
rect 363616 3398 363644 335718
rect 363800 330546 363828 338014
rect 363788 330540 363840 330546
rect 363788 330482 363840 330488
rect 364352 5506 364380 338014
rect 364536 335354 364564 338014
rect 364444 335326 364564 335354
rect 364444 6050 364472 335326
rect 364904 316034 364932 338014
rect 365640 336734 365668 338014
rect 365870 337770 365898 338028
rect 366008 338014 366252 338042
rect 366376 338014 366620 338042
rect 366744 338014 366988 338042
rect 367204 338014 367264 338042
rect 367572 338014 367632 338042
rect 367756 338014 368000 338042
rect 368124 338014 368368 338042
rect 368676 338014 368736 338042
rect 368860 338014 369104 338042
rect 369228 338014 369472 338042
rect 369596 338014 369840 338042
rect 369964 338014 370208 338042
rect 370332 338014 370576 338042
rect 370944 338014 371188 338042
rect 365870 337742 365944 337770
rect 365628 336728 365680 336734
rect 365628 336670 365680 336676
rect 364984 336320 365036 336326
rect 364984 336262 365036 336268
rect 364536 316006 364932 316034
rect 364536 12986 364564 316006
rect 364524 12980 364576 12986
rect 364524 12922 364576 12928
rect 364432 6044 364484 6050
rect 364432 5986 364484 5992
rect 364340 5500 364392 5506
rect 364340 5442 364392 5448
rect 364996 4146 365024 336262
rect 365812 330540 365864 330546
rect 365812 330482 365864 330488
rect 365720 330472 365772 330478
rect 365720 330414 365772 330420
rect 365732 6866 365760 330414
rect 365720 6860 365772 6866
rect 365720 6802 365772 6808
rect 365824 6322 365852 330482
rect 365812 6316 365864 6322
rect 365812 6258 365864 6264
rect 365916 6118 365944 337742
rect 366008 13054 366036 338014
rect 366272 335776 366324 335782
rect 366272 335718 366324 335724
rect 366284 325694 366312 335718
rect 366376 330546 366404 338014
rect 366456 336592 366508 336598
rect 366456 336534 366508 336540
rect 366364 330540 366416 330546
rect 366364 330482 366416 330488
rect 366284 325666 366404 325694
rect 365996 13048 366048 13054
rect 365996 12990 366048 12996
rect 365904 6112 365956 6118
rect 365904 6054 365956 6060
rect 364340 4140 364392 4146
rect 364340 4082 364392 4088
rect 364984 4140 365036 4146
rect 364984 4082 365036 4088
rect 363604 3392 363656 3398
rect 363604 3334 363656 3340
rect 364352 2122 364380 4082
rect 365812 3732 365864 3738
rect 365812 3674 365864 3680
rect 364352 2094 364656 2122
rect 364628 480 364656 2094
rect 365824 480 365852 3674
rect 366376 2990 366404 325666
rect 366468 3738 366496 336534
rect 366744 330478 366772 338014
rect 367100 330540 367152 330546
rect 367100 330482 367152 330488
rect 366732 330472 366784 330478
rect 366732 330414 366784 330420
rect 367112 6798 367140 330482
rect 367204 13802 367232 338014
rect 367572 336598 367600 338014
rect 367560 336592 367612 336598
rect 367560 336534 367612 336540
rect 367652 336456 367704 336462
rect 367652 336398 367704 336404
rect 367284 329452 367336 329458
rect 367284 329394 367336 329400
rect 367296 14278 367324 329394
rect 367664 325694 367692 336398
rect 367756 330546 367784 338014
rect 367836 336184 367888 336190
rect 367836 336126 367888 336132
rect 367744 330540 367796 330546
rect 367744 330482 367796 330488
rect 367664 325666 367784 325694
rect 367284 14272 367336 14278
rect 367284 14214 367336 14220
rect 367192 13796 367244 13802
rect 367192 13738 367244 13744
rect 367100 6792 367152 6798
rect 367100 6734 367152 6740
rect 367756 3942 367784 325666
rect 367744 3936 367796 3942
rect 367744 3878 367796 3884
rect 366456 3732 366508 3738
rect 366456 3674 366508 3680
rect 367008 3460 367060 3466
rect 367008 3402 367060 3408
rect 366364 2984 366416 2990
rect 366364 2926 366416 2932
rect 367020 480 367048 3402
rect 367848 3126 367876 336126
rect 368124 329458 368152 338014
rect 368676 336462 368704 338014
rect 368664 336456 368716 336462
rect 368664 336398 368716 336404
rect 368860 335354 368888 338014
rect 369124 335844 369176 335850
rect 369124 335786 369176 335792
rect 368492 335326 368888 335354
rect 368112 329452 368164 329458
rect 368112 329394 368164 329400
rect 368492 6730 368520 335326
rect 368572 330540 368624 330546
rect 368572 330482 368624 330488
rect 368584 10130 368612 330482
rect 368664 330472 368716 330478
rect 368664 330414 368716 330420
rect 368676 16046 368704 330414
rect 369136 16574 369164 335786
rect 369228 330546 369256 338014
rect 369216 330540 369268 330546
rect 369216 330482 369268 330488
rect 369596 330478 369624 338014
rect 369964 335354 369992 338014
rect 369872 335326 369992 335354
rect 369584 330472 369636 330478
rect 369584 330414 369636 330420
rect 369136 16546 369256 16574
rect 368664 16040 368716 16046
rect 368664 15982 368716 15988
rect 368572 10124 368624 10130
rect 368572 10066 368624 10072
rect 368480 6724 368532 6730
rect 368480 6666 368532 6672
rect 368204 4140 368256 4146
rect 368204 4082 368256 4088
rect 367836 3120 367888 3126
rect 367836 3062 367888 3068
rect 368216 480 368244 4082
rect 369228 3398 369256 16546
rect 369872 6662 369900 335326
rect 370332 316034 370360 338014
rect 371160 336530 371188 338014
rect 371298 337770 371326 338028
rect 371436 338014 371680 338042
rect 371988 338014 372048 338042
rect 372172 338014 372416 338042
rect 372724 338014 372784 338042
rect 371298 337742 371372 337770
rect 371148 336524 371200 336530
rect 371148 336466 371200 336472
rect 370504 336048 370556 336054
rect 370504 335990 370556 335996
rect 369964 316006 370360 316034
rect 369964 10198 369992 316006
rect 369952 10192 370004 10198
rect 369952 10134 370004 10140
rect 369860 6656 369912 6662
rect 369860 6598 369912 6604
rect 369400 3800 369452 3806
rect 369400 3742 369452 3748
rect 369492 3800 369544 3806
rect 369492 3742 369544 3748
rect 369216 3392 369268 3398
rect 369216 3334 369268 3340
rect 369412 480 369440 3742
rect 369504 3466 369532 3742
rect 370516 3466 370544 335990
rect 371240 330540 371292 330546
rect 371240 330482 371292 330488
rect 371252 6526 371280 330482
rect 371344 6594 371372 337742
rect 371436 10266 371464 338014
rect 371884 336116 371936 336122
rect 371884 336058 371936 336064
rect 371424 10260 371476 10266
rect 371424 10202 371476 10208
rect 371332 6588 371384 6594
rect 371332 6530 371384 6536
rect 371240 6520 371292 6526
rect 371240 6462 371292 6468
rect 370596 3664 370648 3670
rect 370596 3606 370648 3612
rect 369492 3460 369544 3466
rect 369492 3402 369544 3408
rect 370504 3460 370556 3466
rect 370504 3402 370556 3408
rect 370608 480 370636 3606
rect 371700 3460 371752 3466
rect 371700 3402 371752 3408
rect 371792 3460 371844 3466
rect 371792 3402 371844 3408
rect 371712 480 371740 3402
rect 371804 3194 371832 3402
rect 371896 3194 371924 336058
rect 371988 335374 372016 338014
rect 371976 335368 372028 335374
rect 371976 335310 372028 335316
rect 372172 330546 372200 338014
rect 372160 330540 372212 330546
rect 372160 330482 372212 330488
rect 372620 330472 372672 330478
rect 372620 330414 372672 330420
rect 372632 10946 372660 330414
rect 372724 11014 372752 338014
rect 373138 337770 373166 338028
rect 373276 338014 373520 338042
rect 373644 338014 373888 338042
rect 374196 338014 374256 338042
rect 374380 338014 374624 338042
rect 374748 338014 374992 338042
rect 375300 338014 375360 338042
rect 375484 338014 375728 338042
rect 375852 338014 376096 338042
rect 376464 338014 376708 338042
rect 376832 338014 376984 338042
rect 373138 337742 373212 337770
rect 373080 336660 373132 336666
rect 373080 336602 373132 336608
rect 372804 330540 372856 330546
rect 372804 330482 372856 330488
rect 372816 13734 372844 330482
rect 373092 325694 373120 336602
rect 373184 336326 373212 337742
rect 373172 336320 373224 336326
rect 373172 336262 373224 336268
rect 373276 330546 373304 338014
rect 373356 336252 373408 336258
rect 373356 336194 373408 336200
rect 373264 330540 373316 330546
rect 373264 330482 373316 330488
rect 373092 325666 373304 325694
rect 372804 13728 372856 13734
rect 372804 13670 372856 13676
rect 372712 11008 372764 11014
rect 372712 10950 372764 10956
rect 372620 10940 372672 10946
rect 372620 10882 372672 10888
rect 371976 3392 372028 3398
rect 373276 3369 373304 325666
rect 371976 3334 372028 3340
rect 373262 3360 373318 3369
rect 371792 3188 371844 3194
rect 371792 3130 371844 3136
rect 371884 3188 371936 3194
rect 371884 3130 371936 3136
rect 371988 2990 372016 3334
rect 373262 3295 373318 3304
rect 373368 3194 373396 336194
rect 373644 330478 373672 338014
rect 374196 336394 374224 338014
rect 374184 336388 374236 336394
rect 374184 336330 374236 336336
rect 374000 330540 374052 330546
rect 374000 330482 374052 330488
rect 373632 330472 373684 330478
rect 373632 330414 373684 330420
rect 374012 10878 374040 330482
rect 374380 316034 374408 338014
rect 374644 335912 374696 335918
rect 374644 335854 374696 335860
rect 374104 316006 374408 316034
rect 374104 13666 374132 316006
rect 374092 13660 374144 13666
rect 374092 13602 374144 13608
rect 374000 10872 374052 10878
rect 374000 10814 374052 10820
rect 374092 3868 374144 3874
rect 374092 3810 374144 3816
rect 373356 3188 373408 3194
rect 373356 3130 373408 3136
rect 372896 3120 372948 3126
rect 372896 3062 372948 3068
rect 371976 2984 372028 2990
rect 371976 2926 372028 2932
rect 372908 480 372936 3062
rect 374104 480 374132 3810
rect 374656 3670 374684 335854
rect 374748 330546 374776 338014
rect 375300 336054 375328 338014
rect 375288 336048 375340 336054
rect 375288 335990 375340 335996
rect 374736 330540 374788 330546
rect 374736 330482 374788 330488
rect 375380 328772 375432 328778
rect 375380 328714 375432 328720
rect 375392 10810 375420 328714
rect 375484 13598 375512 338014
rect 375852 328778 375880 338014
rect 376680 336258 376708 338014
rect 376760 336660 376812 336666
rect 376760 336602 376812 336608
rect 376668 336252 376720 336258
rect 376668 336194 376720 336200
rect 376024 335368 376076 335374
rect 376024 335310 376076 335316
rect 375840 328772 375892 328778
rect 375840 328714 375892 328720
rect 375472 13592 375524 13598
rect 375472 13534 375524 13540
rect 375380 10804 375432 10810
rect 375380 10746 375432 10752
rect 376036 3874 376064 335310
rect 376772 10742 376800 336602
rect 376852 330540 376904 330546
rect 376852 330482 376904 330488
rect 376864 13462 376892 330482
rect 376956 13530 376984 338014
rect 377048 338014 377200 338042
rect 377508 338014 377568 338042
rect 377692 338014 377936 338042
rect 378244 338014 378304 338042
rect 378428 338014 378672 338042
rect 378796 338014 379040 338042
rect 379164 338014 379316 338042
rect 379624 338014 379684 338042
rect 379808 338014 380052 338042
rect 380176 338014 380420 338042
rect 380544 338014 380788 338042
rect 380912 338014 381156 338042
rect 381280 338014 381524 338042
rect 381832 338014 381892 338042
rect 382016 338014 382260 338042
rect 382384 338014 382628 338042
rect 382752 338014 382996 338042
rect 383120 338014 383364 338042
rect 383672 338014 383732 338042
rect 383856 338014 384100 338042
rect 384224 338014 384468 338042
rect 384592 338014 384836 338042
rect 377048 336666 377076 338014
rect 377036 336660 377088 336666
rect 377036 336602 377088 336608
rect 377508 336122 377536 338014
rect 377496 336116 377548 336122
rect 377496 336058 377548 336064
rect 377402 336016 377458 336025
rect 377402 335951 377458 335960
rect 376944 13524 376996 13530
rect 376944 13466 376996 13472
rect 376852 13456 376904 13462
rect 376852 13398 376904 13404
rect 376760 10736 376812 10742
rect 376760 10678 376812 10684
rect 376024 3868 376076 3874
rect 376024 3810 376076 3816
rect 377416 3806 377444 335951
rect 377692 330546 377720 338014
rect 377680 330540 377732 330546
rect 377680 330482 377732 330488
rect 378140 330472 378192 330478
rect 378140 330414 378192 330420
rect 378152 7410 378180 330414
rect 378244 10674 378272 338014
rect 378324 330540 378376 330546
rect 378324 330482 378376 330488
rect 378232 10668 378284 10674
rect 378232 10610 378284 10616
rect 378336 10606 378364 330482
rect 378428 15978 378456 338014
rect 378796 330478 378824 338014
rect 378968 336660 379020 336666
rect 378968 336602 379020 336608
rect 378980 336394 379008 336602
rect 378968 336388 379020 336394
rect 378968 336330 379020 336336
rect 379164 330546 379192 338014
rect 379624 336394 379652 338014
rect 379612 336388 379664 336394
rect 379612 336330 379664 336336
rect 379808 335354 379836 338014
rect 379624 335326 379836 335354
rect 379152 330540 379204 330546
rect 379152 330482 379204 330488
rect 379520 330540 379572 330546
rect 379520 330482 379572 330488
rect 378784 330472 378836 330478
rect 378784 330414 378836 330420
rect 378416 15972 378468 15978
rect 378416 15914 378468 15920
rect 378324 10600 378376 10606
rect 378324 10542 378376 10548
rect 378140 7404 378192 7410
rect 378140 7346 378192 7352
rect 378876 5364 378928 5370
rect 378876 5306 378928 5312
rect 377680 4072 377732 4078
rect 377680 4014 377732 4020
rect 375288 3800 375340 3806
rect 375288 3742 375340 3748
rect 377404 3800 377456 3806
rect 377404 3742 377456 3748
rect 374644 3664 374696 3670
rect 374644 3606 374696 3612
rect 375300 480 375328 3742
rect 376484 3596 376536 3602
rect 376484 3538 376536 3544
rect 376496 480 376524 3538
rect 377692 480 377720 4014
rect 378888 480 378916 5306
rect 379532 4078 379560 330482
rect 379624 7478 379652 335326
rect 380176 316034 380204 338014
rect 380544 330546 380572 338014
rect 380532 330540 380584 330546
rect 380532 330482 380584 330488
rect 379716 316006 380204 316034
rect 379716 10538 379744 316006
rect 379704 10532 379756 10538
rect 379704 10474 379756 10480
rect 380912 7546 380940 338014
rect 380992 327480 381044 327486
rect 380992 327422 381044 327428
rect 381004 8294 381032 327422
rect 381280 316034 381308 338014
rect 381832 336190 381860 338014
rect 381820 336184 381872 336190
rect 381820 336126 381872 336132
rect 382016 327486 382044 338014
rect 382280 330540 382332 330546
rect 382280 330482 382332 330488
rect 382004 327480 382056 327486
rect 382004 327422 382056 327428
rect 381096 316006 381308 316034
rect 381096 10470 381124 316006
rect 381084 10464 381136 10470
rect 381084 10406 381136 10412
rect 380992 8288 381044 8294
rect 380992 8230 381044 8236
rect 380900 7540 380952 7546
rect 380900 7482 380952 7488
rect 379612 7472 379664 7478
rect 379612 7414 379664 7420
rect 382292 6914 382320 330482
rect 382384 10402 382412 338014
rect 382752 330546 382780 338014
rect 382740 330540 382792 330546
rect 382740 330482 382792 330488
rect 383120 316034 383148 338014
rect 382476 316006 383148 316034
rect 382476 11558 382504 316006
rect 382464 11552 382516 11558
rect 382464 11494 382516 11500
rect 382372 10396 382424 10402
rect 382372 10338 382424 10344
rect 383672 8226 383700 338014
rect 383752 330540 383804 330546
rect 383752 330482 383804 330488
rect 383660 8220 383712 8226
rect 383660 8162 383712 8168
rect 383764 8158 383792 330482
rect 383856 10334 383884 338014
rect 384224 316034 384252 338014
rect 384592 330546 384620 338014
rect 385190 337770 385218 338028
rect 385328 338014 385572 338042
rect 385696 338014 385940 338042
rect 386064 338014 386308 338042
rect 386616 338014 386676 338042
rect 386800 338014 387044 338042
rect 387168 338014 387412 338042
rect 387536 338014 387780 338042
rect 387904 338014 388148 338042
rect 388272 338014 388516 338042
rect 388640 338014 388884 338042
rect 389252 338014 389404 338042
rect 385190 337742 385264 337770
rect 384580 330540 384632 330546
rect 384580 330482 384632 330488
rect 385040 330540 385092 330546
rect 385040 330482 385092 330488
rect 383948 316006 384252 316034
rect 383948 11626 383976 316006
rect 383936 11620 383988 11626
rect 383936 11562 383988 11568
rect 383844 10328 383896 10334
rect 383844 10270 383896 10276
rect 383752 8152 383804 8158
rect 383752 8094 383804 8100
rect 385052 8090 385080 330482
rect 385132 330472 385184 330478
rect 385132 330414 385184 330420
rect 385144 12306 385172 330414
rect 385132 12300 385184 12306
rect 385132 12242 385184 12248
rect 385236 11694 385264 337742
rect 385328 12442 385356 338014
rect 385696 330546 385724 338014
rect 385684 330540 385736 330546
rect 385684 330482 385736 330488
rect 386064 330478 386092 338014
rect 386616 330818 386644 338014
rect 386800 335354 386828 338014
rect 386708 335326 386828 335354
rect 386604 330812 386656 330818
rect 386604 330754 386656 330760
rect 386708 330698 386736 335326
rect 386432 330670 386736 330698
rect 386052 330472 386104 330478
rect 386052 330414 386104 330420
rect 385316 12436 385368 12442
rect 385316 12378 385368 12384
rect 385224 11688 385276 11694
rect 385224 11630 385276 11636
rect 385040 8084 385092 8090
rect 385040 8026 385092 8032
rect 386432 8022 386460 330670
rect 386604 330608 386656 330614
rect 386604 330550 386656 330556
rect 386512 330540 386564 330546
rect 386512 330482 386564 330488
rect 386524 12170 386552 330482
rect 386616 12374 386644 330550
rect 387168 316034 387196 338014
rect 387536 330546 387564 338014
rect 387524 330540 387576 330546
rect 387524 330482 387576 330488
rect 387800 330540 387852 330546
rect 387800 330482 387852 330488
rect 386708 316006 387196 316034
rect 386604 12368 386656 12374
rect 386604 12310 386656 12316
rect 386708 12238 386736 316006
rect 386696 12232 386748 12238
rect 386696 12174 386748 12180
rect 386512 12164 386564 12170
rect 386512 12106 386564 12112
rect 386420 8016 386472 8022
rect 386420 7958 386472 7964
rect 382292 6886 382504 6914
rect 382280 5432 382332 5438
rect 382280 5374 382332 5380
rect 382292 4146 382320 5374
rect 382372 5296 382424 5302
rect 382372 5238 382424 5244
rect 382280 4140 382332 4146
rect 382280 4082 382332 4088
rect 379520 4072 379572 4078
rect 379520 4014 379572 4020
rect 381176 4004 381228 4010
rect 381176 3946 381228 3952
rect 379980 3120 380032 3126
rect 379980 3062 380032 3068
rect 379992 480 380020 3062
rect 381188 480 381216 3946
rect 382384 480 382412 5238
rect 382476 4010 382504 6886
rect 384948 5500 385000 5506
rect 384948 5442 385000 5448
rect 382464 4004 382516 4010
rect 382464 3946 382516 3952
rect 384960 3602 384988 5442
rect 385960 5228 386012 5234
rect 385960 5170 386012 5176
rect 384948 3596 385000 3602
rect 384948 3538 385000 3544
rect 383568 3528 383620 3534
rect 383568 3470 383620 3476
rect 383580 480 383608 3470
rect 384764 3256 384816 3262
rect 384764 3198 384816 3204
rect 384776 480 384804 3198
rect 385972 480 386000 5170
rect 387156 5160 387208 5166
rect 387156 5102 387208 5108
rect 387168 480 387196 5102
rect 387812 4690 387840 330482
rect 387904 7954 387932 338014
rect 388272 316034 388300 338014
rect 388536 336728 388588 336734
rect 388536 336670 388588 336676
rect 388548 335986 388576 336670
rect 388444 335980 388496 335986
rect 388444 335922 388496 335928
rect 388536 335980 388588 335986
rect 388536 335922 388588 335928
rect 387996 316006 388300 316034
rect 387996 12102 388024 316006
rect 387984 12096 388036 12102
rect 387984 12038 388036 12044
rect 387892 7948 387944 7954
rect 387892 7890 387944 7896
rect 387800 4684 387852 4690
rect 387800 4626 387852 4632
rect 388456 3398 388484 335922
rect 388640 330546 388668 338014
rect 388628 330540 388680 330546
rect 388628 330482 388680 330488
rect 389180 330540 389232 330546
rect 389180 330482 389232 330488
rect 389192 4758 389220 330482
rect 389272 330472 389324 330478
rect 389272 330414 389324 330420
rect 389284 7818 389312 330414
rect 389376 7886 389404 338014
rect 389468 338014 389620 338042
rect 389744 338014 389988 338042
rect 390112 338014 390356 338042
rect 389468 12034 389496 338014
rect 389744 330546 389772 338014
rect 389732 330540 389784 330546
rect 389732 330482 389784 330488
rect 390112 330478 390140 338014
rect 390710 337770 390738 338028
rect 390848 338014 391092 338042
rect 391216 338014 391368 338042
rect 391492 338014 391736 338042
rect 392044 338014 392104 338042
rect 392228 338014 392472 338042
rect 392596 338014 392840 338042
rect 392964 338014 393208 338042
rect 393424 338014 393576 338042
rect 393700 338014 393944 338042
rect 394068 338014 394312 338042
rect 394436 338014 394680 338042
rect 394896 338014 395048 338042
rect 395172 338014 395416 338042
rect 395540 338014 395784 338042
rect 396152 338014 396304 338042
rect 390710 337742 390784 337770
rect 390652 336796 390704 336802
rect 390652 336738 390704 336744
rect 390560 336728 390612 336734
rect 390560 336670 390612 336676
rect 390100 330472 390152 330478
rect 390100 330414 390152 330420
rect 389456 12028 389508 12034
rect 389456 11970 389508 11976
rect 389364 7880 389416 7886
rect 389364 7822 389416 7828
rect 389272 7812 389324 7818
rect 389272 7754 389324 7760
rect 390572 5506 390600 336670
rect 390664 7750 390692 336738
rect 390756 11966 390784 337742
rect 390848 336734 390876 338014
rect 391216 336802 391244 338014
rect 391204 336796 391256 336802
rect 391204 336738 391256 336744
rect 390836 336728 390888 336734
rect 390836 336670 390888 336676
rect 391204 335980 391256 335986
rect 391204 335922 391256 335928
rect 390836 330540 390888 330546
rect 390836 330482 390888 330488
rect 390848 14346 390876 330482
rect 390836 14340 390888 14346
rect 390836 14282 390888 14288
rect 390744 11960 390796 11966
rect 390744 11902 390796 11908
rect 390652 7744 390704 7750
rect 390652 7686 390704 7692
rect 390560 5500 390612 5506
rect 390560 5442 390612 5448
rect 389456 5092 389508 5098
rect 389456 5034 389508 5040
rect 389180 4752 389232 4758
rect 389180 4694 389232 4700
rect 388260 3392 388312 3398
rect 388260 3334 388312 3340
rect 388444 3392 388496 3398
rect 388444 3334 388496 3340
rect 388272 480 388300 3334
rect 389468 480 389496 5034
rect 391216 3942 391244 335922
rect 391492 330546 391520 338014
rect 391480 330540 391532 330546
rect 391480 330482 391532 330488
rect 391940 330540 391992 330546
rect 391940 330482 391992 330488
rect 391848 6316 391900 6322
rect 391848 6258 391900 6264
rect 390652 3936 390704 3942
rect 390652 3878 390704 3884
rect 391204 3936 391256 3942
rect 391204 3878 391256 3884
rect 391860 3890 391888 6258
rect 391952 5370 391980 330482
rect 392044 5438 392072 338014
rect 392228 335354 392256 338014
rect 392136 335326 392256 335354
rect 392136 7682 392164 335326
rect 392596 316034 392624 338014
rect 392964 330546 392992 338014
rect 392952 330540 393004 330546
rect 392952 330482 393004 330488
rect 393320 328500 393372 328506
rect 393320 328442 393372 328448
rect 392228 316006 392624 316034
rect 392228 11898 392256 316006
rect 392216 11892 392268 11898
rect 392216 11834 392268 11840
rect 392124 7676 392176 7682
rect 392124 7618 392176 7624
rect 392032 5432 392084 5438
rect 392032 5374 392084 5380
rect 391940 5364 391992 5370
rect 391940 5306 391992 5312
rect 393332 5302 393360 328442
rect 393424 7614 393452 338014
rect 393504 330540 393556 330546
rect 393504 330482 393556 330488
rect 393516 13394 393544 330482
rect 393700 316034 393728 338014
rect 394068 328506 394096 338014
rect 394436 330546 394464 338014
rect 394424 330540 394476 330546
rect 394424 330482 394476 330488
rect 394700 330540 394752 330546
rect 394700 330482 394752 330488
rect 394056 328500 394108 328506
rect 394056 328442 394108 328448
rect 393608 316006 393728 316034
rect 393608 14414 393636 316006
rect 393596 14408 393648 14414
rect 393596 14350 393648 14356
rect 393504 13388 393556 13394
rect 393504 13330 393556 13336
rect 393412 7608 393464 7614
rect 393412 7550 393464 7556
rect 393320 5296 393372 5302
rect 393320 5238 393372 5244
rect 394712 5234 394740 330482
rect 394792 326120 394844 326126
rect 394792 326062 394844 326068
rect 394804 13326 394832 326062
rect 394896 15162 394924 338014
rect 395172 330546 395200 338014
rect 395160 330540 395212 330546
rect 395160 330482 395212 330488
rect 395540 326126 395568 338014
rect 396080 336728 396132 336734
rect 396080 336670 396132 336676
rect 395528 326120 395580 326126
rect 395528 326062 395580 326068
rect 394884 15156 394936 15162
rect 394884 15098 394936 15104
rect 394792 13320 394844 13326
rect 394792 13262 394844 13268
rect 394700 5228 394752 5234
rect 394700 5170 394752 5176
rect 396092 5166 396120 336670
rect 396172 330540 396224 330546
rect 396172 330482 396224 330488
rect 396184 13258 396212 330482
rect 396276 15094 396304 338014
rect 396368 338014 396520 338042
rect 396644 338014 396888 338042
rect 397012 338014 397256 338042
rect 397564 338014 397624 338042
rect 397748 338014 397992 338042
rect 398116 338014 398360 338042
rect 398484 338014 398728 338042
rect 398944 338014 399096 338042
rect 399220 338014 399464 338042
rect 399588 338014 399832 338042
rect 399956 338014 400200 338042
rect 400416 338014 400568 338042
rect 400692 338014 400936 338042
rect 401060 338014 401304 338042
rect 401672 338014 401824 338042
rect 396368 336734 396396 338014
rect 396356 336728 396408 336734
rect 396356 336670 396408 336676
rect 396644 330546 396672 338014
rect 396632 330540 396684 330546
rect 396632 330482 396684 330488
rect 397012 316034 397040 338014
rect 397460 330540 397512 330546
rect 397460 330482 397512 330488
rect 396368 316006 397040 316034
rect 396264 15088 396316 15094
rect 396264 15030 396316 15036
rect 396368 15026 396396 316006
rect 396356 15020 396408 15026
rect 396356 14962 396408 14968
rect 396172 13252 396224 13258
rect 396172 13194 396224 13200
rect 396080 5160 396132 5166
rect 396080 5102 396132 5108
rect 393044 5024 393096 5030
rect 393044 4966 393096 4972
rect 390664 480 390692 3878
rect 391860 3862 391980 3890
rect 391952 3738 391980 3862
rect 391848 3732 391900 3738
rect 391848 3674 391900 3680
rect 391940 3732 391992 3738
rect 391940 3674 391992 3680
rect 391860 480 391888 3674
rect 393056 480 393084 4966
rect 396540 4956 396592 4962
rect 396540 4898 396592 4904
rect 395344 3324 395396 3330
rect 395344 3266 395396 3272
rect 394240 3188 394292 3194
rect 394240 3130 394292 3136
rect 394252 480 394280 3130
rect 395356 480 395384 3266
rect 396552 480 396580 4898
rect 397472 4865 397500 330482
rect 397564 5098 397592 338014
rect 397748 335354 397776 338014
rect 397656 335326 397776 335354
rect 397656 13190 397684 335326
rect 398116 316034 398144 338014
rect 398484 330546 398512 338014
rect 398472 330540 398524 330546
rect 398472 330482 398524 330488
rect 398840 328500 398892 328506
rect 398840 328442 398892 328448
rect 397748 316006 398144 316034
rect 397748 14958 397776 316006
rect 397736 14952 397788 14958
rect 397736 14894 397788 14900
rect 397644 13184 397696 13190
rect 397644 13126 397696 13132
rect 397552 5092 397604 5098
rect 397552 5034 397604 5040
rect 398852 5030 398880 328442
rect 398944 8838 398972 338014
rect 399024 330540 399076 330546
rect 399024 330482 399076 330488
rect 399036 8906 399064 330482
rect 399220 316034 399248 338014
rect 399588 328506 399616 338014
rect 399956 330546 399984 338014
rect 399944 330540 399996 330546
rect 399944 330482 399996 330488
rect 400220 330540 400272 330546
rect 400220 330482 400272 330488
rect 399576 328500 399628 328506
rect 399576 328442 399628 328448
rect 399128 316006 399248 316034
rect 399128 14890 399156 316006
rect 399116 14884 399168 14890
rect 399116 14826 399168 14832
rect 399024 8900 399076 8906
rect 399024 8842 399076 8848
rect 398932 8832 398984 8838
rect 398932 8774 398984 8780
rect 398840 5024 398892 5030
rect 398840 4966 398892 4972
rect 400232 4962 400260 330482
rect 400312 326120 400364 326126
rect 400312 326062 400364 326068
rect 400324 9654 400352 326062
rect 400416 14822 400444 338014
rect 400692 330546 400720 338014
rect 400680 330540 400732 330546
rect 400680 330482 400732 330488
rect 401060 326126 401088 338014
rect 401600 336728 401652 336734
rect 401600 336670 401652 336676
rect 401048 326120 401100 326126
rect 401048 326062 401100 326068
rect 400404 14816 400456 14822
rect 400404 14758 400456 14764
rect 400312 9648 400364 9654
rect 400312 9590 400364 9596
rect 400220 4956 400272 4962
rect 400220 4898 400272 4904
rect 401612 4894 401640 336670
rect 401692 330540 401744 330546
rect 401692 330482 401744 330488
rect 401704 9586 401732 330482
rect 401796 14754 401824 338014
rect 401888 338014 402040 338042
rect 402164 338014 402408 338042
rect 402532 338014 402776 338042
rect 402992 338014 403144 338042
rect 403268 338014 403420 338042
rect 403544 338014 403788 338042
rect 403912 338014 404156 338042
rect 404464 338014 404524 338042
rect 404648 338014 404892 338042
rect 405016 338014 405260 338042
rect 405384 338014 405628 338042
rect 401888 336734 401916 338014
rect 401876 336728 401928 336734
rect 401876 336670 401928 336676
rect 402164 330546 402192 338014
rect 402152 330540 402204 330546
rect 402152 330482 402204 330488
rect 402532 316034 402560 338014
rect 401888 316006 402560 316034
rect 401784 14748 401836 14754
rect 401784 14690 401836 14696
rect 401888 14686 401916 316006
rect 401876 14680 401928 14686
rect 401876 14622 401928 14628
rect 401692 9580 401744 9586
rect 401692 9522 401744 9528
rect 398932 4888 398984 4894
rect 397458 4856 397514 4865
rect 398932 4830 398984 4836
rect 401600 4888 401652 4894
rect 401600 4830 401652 4836
rect 397458 4791 397514 4800
rect 397736 3460 397788 3466
rect 397736 3402 397788 3408
rect 397748 480 397776 3402
rect 398944 480 398972 4830
rect 402992 4826 403020 338014
rect 403268 335354 403296 338014
rect 403084 335326 403296 335354
rect 403084 9518 403112 335326
rect 403164 330540 403216 330546
rect 403164 330482 403216 330488
rect 403176 11830 403204 330482
rect 403544 316034 403572 338014
rect 403912 330546 403940 338014
rect 404464 330818 404492 338014
rect 404648 335354 404676 338014
rect 404556 335326 404676 335354
rect 404452 330812 404504 330818
rect 404452 330754 404504 330760
rect 404556 330698 404584 335326
rect 404372 330670 404584 330698
rect 403900 330540 403952 330546
rect 403900 330482 403952 330488
rect 403268 316006 403572 316034
rect 403268 14618 403296 316006
rect 403256 14612 403308 14618
rect 403256 14554 403308 14560
rect 403164 11824 403216 11830
rect 403164 11766 403216 11772
rect 403072 9512 403124 9518
rect 403072 9454 403124 9460
rect 400128 4820 400180 4826
rect 400128 4762 400180 4768
rect 402980 4820 403032 4826
rect 402980 4762 403032 4768
rect 400140 480 400168 4762
rect 403624 4548 403676 4554
rect 403624 4490 403676 4496
rect 402520 4480 402572 4486
rect 402520 4422 402572 4428
rect 401324 3664 401376 3670
rect 401324 3606 401376 3612
rect 401336 480 401364 3606
rect 402532 480 402560 4422
rect 403636 480 403664 4490
rect 404372 3670 404400 330670
rect 404452 330608 404504 330614
rect 404452 330550 404504 330556
rect 404464 9450 404492 330550
rect 404544 330540 404596 330546
rect 404544 330482 404596 330488
rect 404452 9444 404504 9450
rect 404452 9386 404504 9392
rect 404556 9382 404584 330482
rect 405016 316034 405044 338014
rect 405384 330546 405412 338014
rect 405982 337770 406010 338028
rect 406120 338014 406364 338042
rect 406488 338014 406732 338042
rect 406856 338014 407100 338042
rect 407224 338014 407468 338042
rect 407592 338014 407836 338042
rect 408204 338014 408448 338042
rect 405982 337742 406056 337770
rect 405740 330608 405792 330614
rect 405740 330550 405792 330556
rect 405372 330540 405424 330546
rect 405372 330482 405424 330488
rect 404648 316006 405044 316034
rect 404648 11762 404676 316006
rect 404636 11756 404688 11762
rect 404636 11698 404688 11704
rect 404544 9376 404596 9382
rect 404544 9318 404596 9324
rect 404360 3664 404412 3670
rect 404360 3606 404412 3612
rect 405752 3534 405780 330550
rect 405924 330540 405976 330546
rect 405924 330482 405976 330488
rect 405832 330472 405884 330478
rect 405832 330414 405884 330420
rect 405844 9314 405872 330414
rect 405936 13122 405964 330482
rect 406028 14550 406056 337742
rect 406120 330546 406148 338014
rect 406108 330540 406160 330546
rect 406108 330482 406160 330488
rect 406488 330478 406516 338014
rect 406856 330614 406884 338014
rect 407224 335354 407252 338014
rect 407132 335326 407252 335354
rect 406844 330608 406896 330614
rect 406844 330550 406896 330556
rect 406476 330472 406528 330478
rect 406476 330414 406528 330420
rect 406016 14544 406068 14550
rect 406016 14486 406068 14492
rect 405924 13116 405976 13122
rect 405924 13058 405976 13064
rect 405832 9308 405884 9314
rect 405832 9250 405884 9256
rect 407132 6458 407160 335326
rect 407592 316034 407620 338014
rect 408420 335918 408448 338014
rect 408558 337770 408586 338028
rect 408696 338014 408940 338042
rect 409064 338014 409308 338042
rect 409432 338014 409676 338042
rect 408558 337742 408632 337770
rect 408408 335912 408460 335918
rect 408408 335854 408460 335860
rect 408500 330540 408552 330546
rect 408500 330482 408552 330488
rect 407224 316006 407620 316034
rect 407224 9246 407252 316006
rect 407212 9240 407264 9246
rect 407212 9182 407264 9188
rect 407120 6452 407172 6458
rect 407120 6394 407172 6400
rect 408512 6322 408540 330482
rect 408604 6390 408632 337742
rect 408696 9178 408724 338014
rect 409064 316034 409092 338014
rect 409432 330546 409460 338014
rect 410030 337770 410058 338028
rect 410352 338014 410412 338042
rect 410536 338014 410780 338042
rect 410904 338014 411148 338042
rect 411272 338014 411516 338042
rect 411640 338014 411884 338042
rect 412008 338014 412252 338042
rect 412560 338014 412620 338042
rect 412744 338014 412988 338042
rect 413112 338014 413356 338042
rect 413480 338014 413724 338042
rect 414032 338014 414092 338042
rect 414216 338014 414460 338042
rect 414768 338014 414828 338042
rect 410030 337742 410104 337770
rect 409420 330540 409472 330546
rect 409420 330482 409472 330488
rect 409880 330540 409932 330546
rect 409880 330482 409932 330488
rect 408788 316006 409092 316034
rect 408788 14482 408816 316006
rect 408776 14476 408828 14482
rect 408776 14418 408828 14424
rect 408684 9172 408736 9178
rect 408684 9114 408736 9120
rect 408592 6384 408644 6390
rect 408592 6326 408644 6332
rect 408500 6316 408552 6322
rect 408500 6258 408552 6264
rect 409892 6254 409920 330482
rect 409972 330472 410024 330478
rect 409972 330414 410024 330420
rect 409984 9042 410012 330414
rect 410076 9110 410104 337742
rect 410352 335850 410380 338014
rect 410340 335844 410392 335850
rect 410340 335786 410392 335792
rect 410536 330546 410564 338014
rect 410524 330540 410576 330546
rect 410524 330482 410576 330488
rect 410904 330478 410932 338014
rect 410892 330472 410944 330478
rect 410892 330414 410944 330420
rect 410064 9104 410116 9110
rect 410064 9046 410116 9052
rect 409972 9036 410024 9042
rect 409972 8978 410024 8984
rect 407212 6248 407264 6254
rect 407212 6190 407264 6196
rect 409880 6248 409932 6254
rect 409880 6190 409932 6196
rect 406016 4616 406068 4622
rect 406016 4558 406068 4564
rect 405740 3528 405792 3534
rect 405740 3470 405792 3476
rect 404818 3360 404874 3369
rect 404818 3295 404874 3304
rect 404832 480 404860 3295
rect 406028 480 406056 4558
rect 407224 480 407252 6190
rect 409604 6180 409656 6186
rect 409604 6122 409656 6128
rect 408408 3800 408460 3806
rect 408408 3742 408460 3748
rect 408420 480 408448 3742
rect 409616 480 409644 6122
rect 410800 5840 410852 5846
rect 410800 5782 410852 5788
rect 410812 480 410840 5782
rect 411272 3466 411300 338014
rect 411640 335354 411668 338014
rect 411364 335326 411668 335354
rect 411364 6225 411392 335326
rect 412008 316034 412036 338014
rect 412560 335986 412588 338014
rect 412744 336682 412772 338014
rect 412652 336654 412772 336682
rect 412548 335980 412600 335986
rect 412548 335922 412600 335928
rect 411456 316006 412036 316034
rect 411456 8974 411484 316006
rect 411444 8968 411496 8974
rect 411444 8910 411496 8916
rect 411350 6216 411406 6225
rect 412652 6186 412680 336654
rect 413112 335354 413140 338014
rect 412744 335326 413140 335354
rect 412744 8945 412772 335326
rect 413480 316034 413508 338014
rect 414032 336734 414060 338014
rect 414020 336728 414072 336734
rect 414020 336670 414072 336676
rect 414216 316034 414244 338014
rect 414768 336025 414796 338014
rect 414754 336016 414810 336025
rect 414754 335951 414810 335960
rect 412836 316006 413508 316034
rect 414032 316006 414244 316034
rect 412836 15910 412864 316006
rect 412824 15904 412876 15910
rect 412824 15846 412876 15852
rect 412730 8936 412786 8945
rect 412730 8871 412786 8880
rect 411350 6151 411406 6160
rect 412640 6180 412692 6186
rect 412640 6122 412692 6128
rect 413100 5908 413152 5914
rect 413100 5850 413152 5856
rect 411904 4140 411956 4146
rect 411904 4082 411956 4088
rect 411260 3460 411312 3466
rect 411260 3402 411312 3408
rect 411916 480 411944 4082
rect 413112 480 413140 5850
rect 414032 3369 414060 316006
rect 414952 20670 414980 457422
rect 415044 419490 415072 460090
rect 577412 460012 577464 460018
rect 577412 459954 577464 459960
rect 577320 458856 577372 458862
rect 577320 458798 577372 458804
rect 574836 458788 574888 458794
rect 574836 458730 574888 458736
rect 574744 458720 574796 458726
rect 574744 458662 574796 458668
rect 415032 419484 415084 419490
rect 415032 419426 415084 419432
rect 450544 336728 450596 336734
rect 450544 336670 450596 336676
rect 428464 336660 428516 336666
rect 428464 336602 428516 336608
rect 422944 336592 422996 336598
rect 422944 336534 422996 336540
rect 418896 335912 418948 335918
rect 418896 335854 418948 335860
rect 418804 335844 418856 335850
rect 418804 335786 418856 335792
rect 414940 20664 414992 20670
rect 414940 20606 414992 20612
rect 417424 12912 417476 12918
rect 417424 12854 417476 12860
rect 414296 8764 414348 8770
rect 414296 8706 414348 8712
rect 414018 3360 414074 3369
rect 414018 3295 414074 3304
rect 414308 480 414336 8706
rect 416688 5976 416740 5982
rect 416688 5918 416740 5924
rect 415492 3392 415544 3398
rect 415492 3334 415544 3340
rect 415504 480 415532 3334
rect 416700 480 416728 5918
rect 339838 354 339950 480
rect 339512 326 339950 354
rect 339838 -960 339950 326
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417436 354 417464 12854
rect 418816 4146 418844 335786
rect 418804 4140 418856 4146
rect 418804 4082 418856 4088
rect 418908 3806 418936 335854
rect 420920 12980 420972 12986
rect 420920 12922 420972 12928
rect 420184 6044 420236 6050
rect 420184 5986 420236 5992
rect 419080 4140 419132 4146
rect 419080 4082 419132 4088
rect 418896 3800 418948 3806
rect 418896 3742 418948 3748
rect 419092 3602 419120 4082
rect 418988 3596 419040 3602
rect 418988 3538 419040 3544
rect 419080 3596 419132 3602
rect 419080 3538 419132 3544
rect 419000 480 419028 3538
rect 420196 480 420224 5986
rect 417854 354 417966 480
rect 417436 326 417966 354
rect 417854 -960 417966 326
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 420932 354 420960 12922
rect 422576 3936 422628 3942
rect 422576 3878 422628 3884
rect 422588 480 422616 3878
rect 422956 3194 422984 336534
rect 425796 336524 425848 336530
rect 425796 336466 425848 336472
rect 425704 336456 425756 336462
rect 425704 336398 425756 336404
rect 423680 13048 423732 13054
rect 423680 12990 423732 12996
rect 423692 3398 423720 12990
rect 423772 6112 423824 6118
rect 423772 6054 423824 6060
rect 423680 3392 423732 3398
rect 423680 3334 423732 3340
rect 422944 3188 422996 3194
rect 422944 3130 422996 3136
rect 423784 480 423812 6054
rect 424968 3392 425020 3398
rect 424968 3334 425020 3340
rect 424980 480 425008 3334
rect 425716 3058 425744 336398
rect 425808 4146 425836 336466
rect 428476 16574 428504 336602
rect 442264 336388 442316 336394
rect 442264 336330 442316 336336
rect 436744 336320 436796 336326
rect 436744 336262 436796 336268
rect 431224 335980 431276 335986
rect 431224 335922 431276 335928
rect 428476 16546 428596 16574
rect 428464 13796 428516 13802
rect 428464 13738 428516 13744
rect 427268 6860 427320 6866
rect 427268 6802 427320 6808
rect 425796 4140 425848 4146
rect 425796 4082 425848 4088
rect 426164 3732 426216 3738
rect 426164 3674 426216 3680
rect 425704 3052 425756 3058
rect 425704 2994 425756 3000
rect 426176 480 426204 3674
rect 427280 480 427308 6802
rect 428476 480 428504 13738
rect 428568 3942 428596 16546
rect 430856 6792 430908 6798
rect 430856 6734 430908 6740
rect 428556 3936 428608 3942
rect 428556 3878 428608 3884
rect 429660 3188 429712 3194
rect 429660 3130 429712 3136
rect 429672 480 429700 3130
rect 430868 480 430896 6734
rect 431236 3738 431264 335922
rect 436756 16574 436784 336262
rect 439504 336252 439556 336258
rect 439504 336194 439556 336200
rect 436756 16546 436876 16574
rect 436744 16040 436796 16046
rect 436744 15982 436796 15988
rect 432052 14272 432104 14278
rect 432052 14214 432104 14220
rect 431224 3732 431276 3738
rect 431224 3674 431276 3680
rect 432064 480 432092 14214
rect 435088 10124 435140 10130
rect 435088 10066 435140 10072
rect 434444 6724 434496 6730
rect 434444 6666 434496 6672
rect 433248 3052 433300 3058
rect 433248 2994 433300 3000
rect 433260 480 433288 2994
rect 434456 480 434484 6666
rect 421350 354 421462 480
rect 420932 326 421462 354
rect 421350 -960 421462 326
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435100 354 435128 10066
rect 436756 480 436784 15982
rect 436848 3126 436876 16546
rect 439136 10192 439188 10198
rect 439136 10134 439188 10140
rect 437940 6656 437992 6662
rect 437940 6598 437992 6604
rect 436836 3120 436888 3126
rect 436836 3062 436888 3068
rect 437952 480 437980 6598
rect 439148 480 439176 10134
rect 439516 3262 439544 336194
rect 440884 336048 440936 336054
rect 440884 335990 440936 335996
rect 440332 4140 440384 4146
rect 440332 4082 440384 4088
rect 439504 3256 439556 3262
rect 439504 3198 439556 3204
rect 440344 480 440372 4082
rect 440896 3194 440924 335990
rect 442172 10260 442224 10266
rect 442172 10202 442224 10208
rect 441528 6588 441580 6594
rect 441528 6530 441580 6536
rect 440884 3188 440936 3194
rect 440884 3130 440936 3136
rect 441540 480 441568 6530
rect 442184 3482 442212 10202
rect 442276 4146 442304 336330
rect 447784 336184 447836 336190
rect 447784 336126 447836 336132
rect 443644 336116 443696 336122
rect 443644 336058 443696 336064
rect 442264 4140 442316 4146
rect 442264 4082 442316 4088
rect 442724 4140 442776 4146
rect 442724 4082 442776 4088
rect 442184 3454 442672 3482
rect 442644 480 442672 3454
rect 442736 3330 442764 4082
rect 442724 3324 442776 3330
rect 442724 3266 442776 3272
rect 443656 3058 443684 336058
rect 445760 11008 445812 11014
rect 445760 10950 445812 10956
rect 445024 6520 445076 6526
rect 445024 6462 445076 6468
rect 443828 3868 443880 3874
rect 443828 3810 443880 3816
rect 443644 3052 443696 3058
rect 443644 2994 443696 3000
rect 443840 480 443868 3810
rect 445036 480 445064 6462
rect 435518 354 435630 480
rect 435100 326 435630 354
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 445772 354 445800 10950
rect 447796 4146 447824 336126
rect 448520 13728 448572 13734
rect 448520 13670 448572 13676
rect 447784 4140 447836 4146
rect 447784 4082 447836 4088
rect 448532 3210 448560 13670
rect 448612 10940 448664 10946
rect 448612 10882 448664 10888
rect 448624 3398 448652 10882
rect 450556 3874 450584 336670
rect 454682 336016 454738 336025
rect 454682 335951 454738 335960
rect 451648 13660 451700 13666
rect 451648 13602 451700 13608
rect 450912 3936 450964 3942
rect 450912 3878 450964 3884
rect 450544 3868 450596 3874
rect 450544 3810 450596 3816
rect 448612 3392 448664 3398
rect 448612 3334 448664 3340
rect 449808 3392 449860 3398
rect 449808 3334 449860 3340
rect 448532 3182 448652 3210
rect 447416 3120 447468 3126
rect 447416 3062 447468 3068
rect 447428 480 447456 3062
rect 448624 480 448652 3182
rect 449820 480 449848 3334
rect 449992 3324 450044 3330
rect 449992 3266 450044 3272
rect 450004 3058 450032 3266
rect 449992 3052 450044 3058
rect 449992 2994 450044 3000
rect 450924 480 450952 3878
rect 446190 354 446302 480
rect 445772 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451660 354 451688 13602
rect 453304 10872 453356 10878
rect 453304 10814 453356 10820
rect 453316 480 453344 10814
rect 454696 3942 454724 335951
rect 574756 219434 574784 458662
rect 574848 259418 574876 458730
rect 577332 325514 577360 458798
rect 577320 325508 577372 325514
rect 577320 325450 577372 325456
rect 577424 299470 577452 459954
rect 577412 299464 577464 299470
rect 577412 299406 577464 299412
rect 574836 259412 574888 259418
rect 574836 259354 574888 259360
rect 574744 219428 574796 219434
rect 574744 219370 574796 219376
rect 577516 33114 577544 460391
rect 577608 139398 577636 478858
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 578884 460964 578936 460970
rect 578884 460906 578936 460912
rect 578054 460184 578110 460193
rect 578054 460119 578110 460128
rect 577870 459912 577926 459921
rect 577870 459847 577926 459856
rect 577686 459776 577742 459785
rect 577686 459711 577742 459720
rect 577596 139392 577648 139398
rect 577596 139334 577648 139340
rect 577700 73166 577728 459711
rect 577780 458652 577832 458658
rect 577780 458594 577832 458600
rect 577792 179382 577820 458594
rect 577780 179376 577832 179382
rect 577780 179318 577832 179324
rect 577884 113014 577912 459847
rect 577964 456816 578016 456822
rect 577964 456758 578016 456764
rect 577976 233238 578004 456758
rect 577964 233232 578016 233238
rect 577964 233174 578016 233180
rect 578068 193186 578096 460119
rect 578148 456884 578200 456890
rect 578148 456826 578200 456832
rect 578160 273222 578188 456826
rect 578896 312089 578924 460906
rect 580538 460320 580594 460329
rect 580538 460255 580594 460264
rect 580080 460080 580132 460086
rect 580080 460022 580132 460028
rect 580354 460048 580410 460057
rect 580092 431633 580120 460022
rect 580354 459983 580410 459992
rect 580264 458992 580316 458998
rect 580264 458934 580316 458940
rect 580172 458924 580224 458930
rect 580172 458866 580224 458872
rect 580184 458153 580212 458866
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580172 457088 580224 457094
rect 580172 457030 580224 457036
rect 580078 431624 580134 431633
rect 580078 431559 580134 431568
rect 579988 419484 580040 419490
rect 579988 419426 580040 419432
rect 580000 418305 580028 419426
rect 579986 418296 580042 418305
rect 579986 418231 580042 418240
rect 580184 404977 580212 457030
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 578882 312080 578938 312089
rect 578882 312015 578938 312024
rect 579620 299464 579672 299470
rect 579620 299406 579672 299412
rect 579632 298761 579660 299406
rect 579618 298752 579674 298761
rect 579618 298687 579674 298696
rect 578148 273216 578200 273222
rect 578148 273158 578200 273164
rect 579620 273216 579672 273222
rect 579620 273158 579672 273164
rect 579632 272241 579660 273158
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 579804 259412 579856 259418
rect 579804 259354 579856 259360
rect 579816 258913 579844 259354
rect 579802 258904 579858 258913
rect 579802 258839 579858 258848
rect 579620 233232 579672 233238
rect 579620 233174 579672 233180
rect 579632 232393 579660 233174
rect 579618 232384 579674 232393
rect 579618 232319 579674 232328
rect 580172 219428 580224 219434
rect 580172 219370 580224 219376
rect 580184 219065 580212 219370
rect 580170 219056 580226 219065
rect 580170 218991 580226 219000
rect 578056 193180 578108 193186
rect 578056 193122 578108 193128
rect 579620 193180 579672 193186
rect 579620 193122 579672 193128
rect 579632 192545 579660 193122
rect 579618 192536 579674 192545
rect 579618 192471 579674 192480
rect 580080 179376 580132 179382
rect 580080 179318 580132 179324
rect 580092 179217 580120 179318
rect 580078 179208 580134 179217
rect 580078 179143 580134 179152
rect 579620 139392 579672 139398
rect 579618 139360 579620 139369
rect 579672 139360 579674 139369
rect 579618 139295 579674 139304
rect 580276 126041 580304 458934
rect 580368 152697 580396 459983
rect 580446 457464 580502 457473
rect 580446 457399 580502 457408
rect 580460 165889 580488 457399
rect 580552 205737 580580 460255
rect 580632 459944 580684 459950
rect 580632 459886 580684 459892
rect 580644 245585 580672 459886
rect 580816 459060 580868 459066
rect 580816 459002 580868 459008
rect 580724 456952 580776 456958
rect 580724 456894 580776 456900
rect 580736 351937 580764 456894
rect 580828 365129 580856 459002
rect 580908 457020 580960 457026
rect 580908 456962 580960 456968
rect 580920 378457 580948 456962
rect 580906 378448 580962 378457
rect 580906 378383 580962 378392
rect 580814 365120 580870 365129
rect 580814 365055 580870 365064
rect 580722 351928 580778 351937
rect 580722 351863 580778 351872
rect 580724 325508 580776 325514
rect 580724 325450 580776 325456
rect 580736 325281 580764 325450
rect 580722 325272 580778 325281
rect 580722 325207 580778 325216
rect 580630 245576 580686 245585
rect 580630 245511 580686 245520
rect 580538 205728 580594 205737
rect 580538 205663 580594 205672
rect 580446 165880 580502 165889
rect 580446 165815 580502 165824
rect 580354 152688 580410 152697
rect 580354 152623 580410 152632
rect 580262 126032 580318 126041
rect 580262 125967 580318 125976
rect 577872 113008 577924 113014
rect 577872 112950 577924 112956
rect 580540 113008 580592 113014
rect 580540 112950 580592 112956
rect 580552 112849 580580 112950
rect 580538 112840 580594 112849
rect 580538 112775 580594 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 577688 73160 577740 73166
rect 577688 73102 577740 73108
rect 579712 73160 579764 73166
rect 579712 73102 579764 73108
rect 579724 73001 579752 73102
rect 579710 72992 579766 73001
rect 579710 72927 579766 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 579618 33144 579674 33153
rect 577504 33108 577556 33114
rect 579618 33079 579620 33088
rect 577504 33050 577556 33056
rect 579672 33079 579674 33088
rect 579620 33050 579672 33056
rect 580172 20596 580224 20602
rect 580172 20538 580224 20544
rect 580184 19825 580212 20538
rect 580264 19984 580316 19990
rect 580264 19926 580316 19932
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 465172 15972 465224 15978
rect 465172 15914 465224 15920
rect 455696 13592 455748 13598
rect 455696 13534 455748 13540
rect 454684 3936 454736 3942
rect 454684 3878 454736 3884
rect 454500 3188 454552 3194
rect 454500 3130 454552 3136
rect 454512 480 454540 3130
rect 455708 480 455736 13534
rect 459192 13524 459244 13530
rect 459192 13466 459244 13472
rect 456892 10804 456944 10810
rect 456892 10746 456944 10752
rect 456904 480 456932 10746
rect 458088 3256 458140 3262
rect 458088 3198 458140 3204
rect 458100 480 458128 3198
rect 459204 480 459232 13466
rect 462320 13456 462372 13462
rect 462320 13398 462372 13404
rect 459928 10736 459980 10742
rect 459928 10678 459980 10684
rect 452078 354 452190 480
rect 451660 326 452190 354
rect 452078 -960 452190 326
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459940 354 459968 10678
rect 461584 3324 461636 3330
rect 461584 3266 461636 3272
rect 461596 480 461624 3266
rect 460358 354 460470 480
rect 459940 326 460470 354
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462332 354 462360 13398
rect 463976 10668 464028 10674
rect 463976 10610 464028 10616
rect 463988 480 464016 10610
rect 465184 480 465212 15914
rect 578608 15904 578660 15910
rect 578608 15846 578660 15852
rect 517888 15156 517940 15162
rect 517888 15098 517940 15104
rect 514760 14408 514812 14414
rect 514760 14350 514812 14356
rect 507216 14340 507268 14346
rect 507216 14282 507268 14288
rect 487160 12436 487212 12442
rect 487160 12378 487212 12384
rect 486424 11688 486476 11694
rect 486424 11630 486476 11636
rect 484032 11620 484084 11626
rect 484032 11562 484084 11568
rect 480536 11552 480588 11558
rect 480536 11494 480588 11500
rect 467472 10600 467524 10606
rect 467472 10542 467524 10548
rect 466276 7404 466328 7410
rect 466276 7346 466328 7352
rect 466288 480 466316 7346
rect 467484 480 467512 10542
rect 470600 10532 470652 10538
rect 470600 10474 470652 10480
rect 469864 7472 469916 7478
rect 469864 7414 469916 7420
rect 468668 3392 468720 3398
rect 468668 3334 468720 3340
rect 468680 480 468708 3334
rect 469876 480 469904 7414
rect 462750 354 462862 480
rect 462332 326 462862 354
rect 462750 -960 462862 326
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 470612 354 470640 10474
rect 474096 10464 474148 10470
rect 474096 10406 474148 10412
rect 473452 7540 473504 7546
rect 473452 7482 473504 7488
rect 472256 4072 472308 4078
rect 472256 4014 472308 4020
rect 472268 480 472296 4014
rect 473464 480 473492 7482
rect 471030 354 471142 480
rect 470612 326 471142 354
rect 471030 -960 471142 326
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474108 354 474136 10406
rect 478144 10396 478196 10402
rect 478144 10338 478196 10344
rect 476948 8288 477000 8294
rect 476948 8230 477000 8236
rect 475752 4140 475804 4146
rect 475752 4082 475804 4088
rect 475764 480 475792 4082
rect 476960 480 476988 8230
rect 478156 480 478184 10338
rect 479340 4004 479392 4010
rect 479340 3946 479392 3952
rect 479352 480 479380 3946
rect 480548 480 480576 11494
rect 482376 10328 482428 10334
rect 482376 10270 482428 10276
rect 481732 8220 481784 8226
rect 481732 8162 481784 8168
rect 481744 480 481772 8162
rect 474526 354 474638 480
rect 474108 326 474638 354
rect 474526 -960 474638 326
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482388 354 482416 10270
rect 484044 480 484072 11562
rect 485228 8152 485280 8158
rect 485228 8094 485280 8100
rect 485240 480 485268 8094
rect 486436 480 486464 11630
rect 482806 354 482918 480
rect 482388 326 482918 354
rect 482806 -960 482918 326
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487172 354 487200 12378
rect 489920 12368 489972 12374
rect 489920 12310 489972 12316
rect 488816 8084 488868 8090
rect 488816 8026 488868 8032
rect 488828 480 488856 8026
rect 489932 3398 489960 12310
rect 490012 12300 490064 12306
rect 490012 12242 490064 12248
rect 489920 3392 489972 3398
rect 489920 3334 489972 3340
rect 490024 3210 490052 12242
rect 493048 12232 493100 12238
rect 493048 12174 493100 12180
rect 492312 8016 492364 8022
rect 492312 7958 492364 7964
rect 490748 3392 490800 3398
rect 490748 3334 490800 3340
rect 489932 3182 490052 3210
rect 489932 480 489960 3182
rect 487590 354 487702 480
rect 487172 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 490760 354 490788 3334
rect 492324 480 492352 7958
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 491086 -960 491198 326
rect 492282 -960 492394 480
rect 493060 354 493088 12174
rect 494704 12164 494756 12170
rect 494704 12106 494756 12112
rect 494716 480 494744 12106
rect 497096 12096 497148 12102
rect 497096 12038 497148 12044
rect 495900 7948 495952 7954
rect 495900 7890 495952 7896
rect 495912 480 495940 7890
rect 497108 480 497136 12038
rect 500592 12028 500644 12034
rect 500592 11970 500644 11976
rect 499396 7880 499448 7886
rect 499396 7822 499448 7828
rect 498200 4684 498252 4690
rect 498200 4626 498252 4632
rect 498212 480 498240 4626
rect 499408 480 499436 7822
rect 500604 480 500632 11970
rect 503720 11960 503772 11966
rect 503720 11902 503772 11908
rect 502984 7812 503036 7818
rect 502984 7754 503036 7760
rect 501788 4752 501840 4758
rect 501788 4694 501840 4700
rect 501800 480 501828 4694
rect 502996 480 503024 7754
rect 493478 354 493590 480
rect 493060 326 493590 354
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 503732 354 503760 11902
rect 506480 7744 506532 7750
rect 506480 7686 506532 7692
rect 505376 5500 505428 5506
rect 505376 5442 505428 5448
rect 505388 480 505416 5442
rect 506492 480 506520 7686
rect 504150 354 504262 480
rect 503732 326 504262 354
rect 504150 -960 504262 326
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507228 354 507256 14282
rect 511264 11892 511316 11898
rect 511264 11834 511316 11840
rect 510068 7676 510120 7682
rect 510068 7618 510120 7624
rect 508872 5432 508924 5438
rect 508872 5374 508924 5380
rect 508884 480 508912 5374
rect 510080 480 510108 7618
rect 511276 480 511304 11834
rect 513564 7608 513616 7614
rect 513564 7550 513616 7556
rect 512460 5364 512512 5370
rect 512460 5306 512512 5312
rect 512472 480 512500 5306
rect 513576 480 513604 7550
rect 514772 480 514800 14350
rect 517152 13388 517204 13394
rect 517152 13330 517204 13336
rect 515956 5296 516008 5302
rect 515956 5238 516008 5244
rect 515968 480 515996 5238
rect 517164 480 517192 13330
rect 507646 354 507758 480
rect 507228 326 507758 354
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 517900 354 517928 15098
rect 521660 15088 521712 15094
rect 521660 15030 521712 15036
rect 520280 13320 520332 13326
rect 520280 13262 520332 13268
rect 519544 5228 519596 5234
rect 519544 5170 519596 5176
rect 519556 480 519584 5170
rect 518318 354 518430 480
rect 517900 326 518430 354
rect 518318 -960 518430 326
rect 519514 -960 519626 480
rect 520292 354 520320 13262
rect 520710 354 520822 480
rect 520292 326 520822 354
rect 521672 354 521700 15030
rect 525432 15020 525484 15026
rect 525432 14962 525484 14968
rect 523776 13252 523828 13258
rect 523776 13194 523828 13200
rect 523040 5160 523092 5166
rect 523040 5102 523092 5108
rect 523052 480 523080 5102
rect 521814 354 521926 480
rect 521672 326 521926 354
rect 520710 -960 520822 326
rect 521814 -960 521926 326
rect 523010 -960 523122 480
rect 523788 354 523816 13194
rect 525444 480 525472 14962
rect 528560 14952 528612 14958
rect 528560 14894 528612 14900
rect 527824 13184 527876 13190
rect 527824 13126 527876 13132
rect 526628 5092 526680 5098
rect 526628 5034 526680 5040
rect 526640 480 526668 5034
rect 527836 480 527864 13126
rect 524206 354 524318 480
rect 523788 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528572 354 528600 14894
rect 532056 14884 532108 14890
rect 532056 14826 532108 14832
rect 531320 8832 531372 8838
rect 531320 8774 531372 8780
rect 530122 4856 530178 4865
rect 530122 4791 530178 4800
rect 530136 480 530164 4791
rect 531332 480 531360 8774
rect 528990 354 529102 480
rect 528572 326 529102 354
rect 528990 -960 529102 326
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532068 354 532096 14826
rect 536104 14816 536156 14822
rect 536104 14758 536156 14764
rect 534908 8900 534960 8906
rect 534908 8842 534960 8848
rect 533712 5024 533764 5030
rect 533712 4966 533764 4972
rect 533724 480 533752 4966
rect 534920 480 534948 8842
rect 536116 480 536144 14758
rect 539600 14748 539652 14754
rect 539600 14690 539652 14696
rect 538404 9648 538456 9654
rect 538404 9590 538456 9596
rect 537208 4956 537260 4962
rect 537208 4898 537260 4904
rect 537220 480 537248 4898
rect 538416 480 538444 9590
rect 539612 480 539640 14690
rect 542728 14680 542780 14686
rect 542728 14622 542780 14628
rect 541992 9580 542044 9586
rect 541992 9522 542044 9528
rect 540796 4888 540848 4894
rect 540796 4830 540848 4836
rect 540808 480 540836 4830
rect 542004 480 542032 9522
rect 532486 354 532598 480
rect 532068 326 532598 354
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542740 354 542768 14622
rect 546500 14612 546552 14618
rect 546500 14554 546552 14560
rect 545488 9512 545540 9518
rect 545488 9454 545540 9460
rect 544384 4820 544436 4826
rect 544384 4762 544436 4768
rect 544396 480 544424 4762
rect 545500 480 545528 9454
rect 543158 354 543270 480
rect 542740 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546512 354 546540 14554
rect 553768 14544 553820 14550
rect 553768 14486 553820 14492
rect 547880 11824 547932 11830
rect 547880 11766 547932 11772
rect 547892 480 547920 11766
rect 551008 11756 551060 11762
rect 551008 11698 551060 11704
rect 549076 9444 549128 9450
rect 549076 9386 549128 9392
rect 549088 480 549116 9386
rect 550272 3664 550324 3670
rect 550272 3606 550324 3612
rect 550284 480 550312 3606
rect 546654 354 546766 480
rect 546512 326 546766 354
rect 546654 -960 546766 326
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551020 354 551048 11698
rect 552664 9376 552716 9382
rect 552664 9318 552716 9324
rect 552676 480 552704 9318
rect 553780 480 553808 14486
rect 564440 14476 564492 14482
rect 564440 14418 564492 14424
rect 554780 13116 554832 13122
rect 554780 13058 554832 13064
rect 551438 354 551550 480
rect 551020 326 551550 354
rect 551438 -960 551550 326
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554792 354 554820 13058
rect 556160 9308 556212 9314
rect 556160 9250 556212 9256
rect 556172 480 556200 9250
rect 559748 9240 559800 9246
rect 559748 9182 559800 9188
rect 558552 6452 558604 6458
rect 558552 6394 558604 6400
rect 557356 3528 557408 3534
rect 557356 3470 557408 3476
rect 557368 480 557396 3470
rect 558564 480 558592 6394
rect 559760 480 559788 9182
rect 563244 9172 563296 9178
rect 563244 9114 563296 9120
rect 562048 6384 562100 6390
rect 562048 6326 562100 6332
rect 560852 3800 560904 3806
rect 560852 3742 560904 3748
rect 560864 480 560892 3742
rect 562060 480 562088 6326
rect 563256 480 563284 9114
rect 564452 480 564480 14418
rect 566832 9104 566884 9110
rect 566832 9046 566884 9052
rect 565636 6316 565688 6322
rect 565636 6258 565688 6264
rect 565648 480 565676 6258
rect 566844 480 566872 9046
rect 570328 9036 570380 9042
rect 570328 8978 570380 8984
rect 569132 6248 569184 6254
rect 569132 6190 569184 6196
rect 568028 3596 568080 3602
rect 568028 3538 568080 3544
rect 568040 480 568068 3538
rect 569144 480 569172 6190
rect 570340 480 570368 8978
rect 573916 8968 573968 8974
rect 573916 8910 573968 8916
rect 577410 8936 577466 8945
rect 572718 6216 572774 6225
rect 572718 6151 572774 6160
rect 571524 3460 571576 3466
rect 571524 3402 571576 3408
rect 571536 480 571564 3402
rect 572732 480 572760 6151
rect 573928 480 573956 8910
rect 577410 8871 577466 8880
rect 576308 6180 576360 6186
rect 576308 6122 576360 6128
rect 575112 3732 575164 3738
rect 575112 3674 575164 3680
rect 575124 480 575152 3674
rect 576320 480 576348 6122
rect 577424 480 577452 8871
rect 578620 480 578648 15846
rect 580276 6633 580304 19926
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 583392 3936 583444 3942
rect 583392 3878 583444 3884
rect 581000 3868 581052 3874
rect 581000 3810 581052 3816
rect 581012 480 581040 3810
rect 582194 3360 582250 3369
rect 582194 3295 582250 3304
rect 582208 480 582236 3295
rect 583404 480 583432 3878
rect 554934 354 555046 480
rect 554792 326 555046 354
rect 554934 -960 555046 326
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 684256 3478 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 2778 449520 2834 449576
rect 3238 423544 3294 423600
rect 3330 410488 3386 410544
rect 3330 306176 3386 306232
rect 3146 254088 3202 254144
rect 237286 460400 237342 460456
rect 4802 458224 4858 458280
rect 4066 397432 4122 397488
rect 3974 371320 4030 371376
rect 3882 358400 3938 358456
rect 3790 345344 3846 345400
rect 3698 319232 3754 319288
rect 3606 293120 3662 293176
rect 3514 267144 3570 267200
rect 3514 241032 3570 241088
rect 3422 214920 3478 214976
rect 3422 201864 3478 201920
rect 3422 188808 3478 188864
rect 2778 162832 2834 162888
rect 3422 149776 3478 149832
rect 3238 136720 3294 136776
rect 3422 97552 3478 97608
rect 3146 84632 3202 84688
rect 2778 71612 2780 71632
rect 2780 71612 2832 71632
rect 2832 71612 2834 71632
rect 2778 71576 2834 71612
rect 3514 19896 3570 19952
rect 3422 19352 3478 19408
rect 110 15816 166 15872
rect 9678 18536 9734 18592
rect 3422 6432 3478 6488
rect 5262 3304 5318 3360
rect 8758 11600 8814 11656
rect 38658 335960 38714 336016
rect 22558 14456 22614 14512
rect 17038 8880 17094 8936
rect 40222 12960 40278 13016
rect 131118 17176 131174 17232
rect 79230 10240 79286 10296
rect 162490 7520 162546 7576
rect 234250 457272 234306 457328
rect 234066 457136 234122 457192
rect 233882 457000 233938 457056
rect 233606 456320 233662 456376
rect 233790 456184 233846 456240
rect 233974 456048 234030 456104
rect 246946 459856 247002 459912
rect 242346 459720 242402 459776
rect 240782 458496 240838 458552
rect 245566 458632 245622 458688
rect 251822 459992 251878 460048
rect 259366 460264 259422 460320
rect 256606 460128 256662 460184
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670656 580226 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 577502 460400 577558 460456
rect 401230 458360 401286 458416
rect 406336 458224 406392 458280
rect 308954 457408 309010 457464
rect 385406 457408 385462 457464
rect 390190 457408 390246 457464
rect 393502 457408 393558 457464
rect 394974 457408 395030 457464
rect 398102 457408 398158 457464
rect 402978 457408 403034 457464
rect 407578 457408 407634 457464
rect 409142 457408 409198 457464
rect 410706 457408 410762 457464
rect 412270 457408 412326 457464
rect 200302 4800 200358 4856
rect 234618 15816 234674 15872
rect 228730 6160 228786 6216
rect 236274 3304 236330 3360
rect 237654 18536 237710 18592
rect 237562 11600 237618 11656
rect 241702 14456 241758 14512
rect 240322 8880 240378 8936
rect 241702 3304 241758 3360
rect 247038 335960 247094 336016
rect 247130 12960 247186 13016
rect 259550 10240 259606 10296
rect 276018 335960 276074 336016
rect 274914 17176 274970 17232
rect 284390 7520 284446 7576
rect 296902 4936 296958 4992
rect 297730 4800 297786 4856
rect 304998 6160 305054 6216
rect 300766 3440 300822 3496
rect 309322 4800 309378 4856
rect 309230 3304 309286 3360
rect 320270 335960 320326 336016
rect 327170 3440 327226 3496
rect 361026 335960 361082 336016
rect 373262 3304 373318 3360
rect 377402 335960 377458 336016
rect 397458 4800 397514 4856
rect 404818 3304 404874 3360
rect 411350 6160 411406 6216
rect 414754 335960 414810 336016
rect 412730 8880 412786 8936
rect 414018 3304 414074 3360
rect 454682 335960 454738 336016
rect 579986 471416 580042 471472
rect 578054 460128 578110 460184
rect 577870 459856 577926 459912
rect 577686 459720 577742 459776
rect 580538 460264 580594 460320
rect 580354 459992 580410 460048
rect 580170 458088 580226 458144
rect 580078 431568 580134 431624
rect 579986 418240 580042 418296
rect 580170 404912 580226 404968
rect 578882 312024 578938 312080
rect 579618 298696 579674 298752
rect 579618 272176 579674 272232
rect 579802 258848 579858 258904
rect 579618 232328 579674 232384
rect 580170 219000 580226 219056
rect 579618 192480 579674 192536
rect 580078 179152 580134 179208
rect 579618 139340 579620 139360
rect 579620 139340 579672 139360
rect 579672 139340 579674 139360
rect 579618 139304 579674 139340
rect 580446 457408 580502 457464
rect 580906 378392 580962 378448
rect 580814 365064 580870 365120
rect 580722 351872 580778 351928
rect 580722 325216 580778 325272
rect 580630 245520 580686 245576
rect 580538 205672 580594 205728
rect 580446 165824 580502 165880
rect 580354 152632 580410 152688
rect 580262 125976 580318 126032
rect 580538 112784 580594 112840
rect 580170 99456 580226 99512
rect 579710 72936 579766 72992
rect 580170 59608 580226 59664
rect 579618 33108 579674 33144
rect 579618 33088 579620 33108
rect 579620 33088 579672 33108
rect 579672 33088 579674 33108
rect 580170 19760 580226 19816
rect 530122 4800 530178 4856
rect 572718 6160 572774 6216
rect 577410 8880 577466 8936
rect 580262 6568 580318 6624
rect 582194 3304 582250 3360
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 3417 684314 3483 684317
rect -960 684312 3483 684314
rect -960 684256 3422 684312
rect 3478 684256 3483 684312
rect -960 684254 3483 684256
rect -960 684164 480 684254
rect 3417 684251 3483 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 237281 460458 237347 460461
rect 577497 460458 577563 460461
rect 237281 460456 577563 460458
rect 237281 460400 237286 460456
rect 237342 460400 577502 460456
rect 577558 460400 577563 460456
rect 237281 460398 577563 460400
rect 237281 460395 237347 460398
rect 577497 460395 577563 460398
rect 259361 460322 259427 460325
rect 580533 460322 580599 460325
rect 259361 460320 580599 460322
rect 259361 460264 259366 460320
rect 259422 460264 580538 460320
rect 580594 460264 580599 460320
rect 259361 460262 580599 460264
rect 259361 460259 259427 460262
rect 580533 460259 580599 460262
rect 256601 460186 256667 460189
rect 578049 460186 578115 460189
rect 256601 460184 578115 460186
rect 256601 460128 256606 460184
rect 256662 460128 578054 460184
rect 578110 460128 578115 460184
rect 256601 460126 578115 460128
rect 256601 460123 256667 460126
rect 578049 460123 578115 460126
rect 251817 460050 251883 460053
rect 580349 460050 580415 460053
rect 251817 460048 580415 460050
rect 251817 459992 251822 460048
rect 251878 459992 580354 460048
rect 580410 459992 580415 460048
rect 251817 459990 580415 459992
rect 251817 459987 251883 459990
rect 580349 459987 580415 459990
rect 246941 459914 247007 459917
rect 577865 459914 577931 459917
rect 246941 459912 577931 459914
rect 246941 459856 246946 459912
rect 247002 459856 577870 459912
rect 577926 459856 577931 459912
rect 246941 459854 577931 459856
rect 246941 459851 247007 459854
rect 577865 459851 577931 459854
rect 242341 459778 242407 459781
rect 577681 459778 577747 459781
rect 242341 459776 577747 459778
rect 242341 459720 242346 459776
rect 242402 459720 577686 459776
rect 577742 459720 577747 459776
rect 242341 459718 577747 459720
rect 242341 459715 242407 459718
rect 577681 459715 577747 459718
rect 245561 458690 245627 458693
rect 580390 458690 580396 458692
rect 245561 458688 580396 458690
rect 245561 458632 245566 458688
rect 245622 458632 580396 458688
rect 245561 458630 580396 458632
rect 245561 458627 245627 458630
rect 580390 458628 580396 458630
rect 580460 458628 580466 458692
rect 240777 458554 240843 458557
rect 580206 458554 580212 458556
rect 240777 458552 580212 458554
rect 240777 458496 240782 458552
rect 240838 458496 580212 458552
rect 240777 458494 580212 458496
rect 240777 458491 240843 458494
rect 580206 458492 580212 458494
rect 580276 458492 580282 458556
rect 3366 458356 3372 458420
rect 3436 458418 3442 458420
rect 401225 458418 401291 458421
rect 3436 458416 401291 458418
rect 3436 458360 401230 458416
rect 401286 458360 401291 458416
rect 3436 458358 401291 458360
rect 3436 458356 3442 458358
rect 401225 458355 401291 458358
rect 4797 458282 4863 458285
rect 406331 458282 406397 458285
rect 4797 458280 406397 458282
rect 4797 458224 4802 458280
rect 4858 458224 406336 458280
rect 406392 458224 406397 458280
rect 4797 458222 406397 458224
rect 4797 458219 4863 458222
rect 406331 458219 406397 458222
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 373950 457542 412650 457602
rect 308949 457466 309015 457469
rect 373950 457466 374010 457542
rect 385401 457468 385467 457469
rect 390185 457468 390251 457469
rect 385350 457466 385356 457468
rect 308949 457464 374010 457466
rect 308949 457408 308954 457464
rect 309010 457408 374010 457464
rect 308949 457406 374010 457408
rect 385310 457406 385356 457466
rect 385420 457464 385467 457468
rect 390134 457466 390140 457468
rect 385462 457408 385467 457464
rect 308949 457403 309015 457406
rect 385350 457404 385356 457406
rect 385420 457404 385467 457408
rect 390094 457406 390140 457466
rect 390204 457464 390251 457468
rect 393497 457466 393563 457469
rect 394969 457468 395035 457469
rect 394918 457466 394924 457468
rect 390246 457408 390251 457464
rect 390134 457404 390140 457406
rect 390204 457404 390251 457408
rect 385401 457403 385467 457404
rect 390185 457403 390251 457404
rect 393270 457464 393563 457466
rect 393270 457408 393502 457464
rect 393558 457408 393563 457464
rect 393270 457406 393563 457408
rect 394878 457406 394924 457466
rect 394988 457464 395035 457468
rect 398097 457466 398163 457469
rect 402973 457466 403039 457469
rect 407573 457466 407639 457469
rect 395030 457408 395035 457464
rect 234245 457330 234311 457333
rect 393270 457330 393330 457406
rect 393497 457403 393563 457406
rect 394918 457404 394924 457406
rect 394988 457404 395035 457408
rect 394969 457403 395035 457404
rect 395846 457464 398163 457466
rect 395846 457408 398102 457464
rect 398158 457408 398163 457464
rect 395846 457406 398163 457408
rect 234245 457328 393330 457330
rect 234245 457272 234250 457328
rect 234306 457272 393330 457328
rect 234245 457270 393330 457272
rect 234245 457267 234311 457270
rect 234061 457194 234127 457197
rect 395846 457194 395906 457406
rect 398097 457403 398163 457406
rect 402930 457464 403039 457466
rect 402930 457408 402978 457464
rect 403034 457408 403039 457464
rect 402930 457403 403039 457408
rect 405414 457464 407639 457466
rect 405414 457408 407578 457464
rect 407634 457408 407639 457464
rect 405414 457406 407639 457408
rect 234061 457192 395906 457194
rect 234061 457136 234066 457192
rect 234122 457136 395906 457192
rect 234061 457134 395906 457136
rect 234061 457131 234127 457134
rect 233877 457058 233943 457061
rect 402930 457058 402990 457403
rect 233877 457056 402990 457058
rect 233877 457000 233882 457056
rect 233938 457000 402990 457056
rect 233877 456998 402990 457000
rect 233877 456995 233943 456998
rect 233734 456860 233740 456924
rect 233804 456922 233810 456924
rect 405414 456922 405474 457406
rect 407573 457403 407639 457406
rect 408718 457404 408724 457468
rect 408788 457466 408794 457468
rect 409137 457466 409203 457469
rect 408788 457464 409203 457466
rect 408788 457408 409142 457464
rect 409198 457408 409203 457464
rect 408788 457406 409203 457408
rect 408788 457404 408794 457406
rect 409137 457403 409203 457406
rect 409822 457404 409828 457468
rect 409892 457466 409898 457468
rect 410701 457466 410767 457469
rect 409892 457464 410767 457466
rect 409892 457408 410706 457464
rect 410762 457408 410767 457464
rect 409892 457406 410767 457408
rect 409892 457404 409898 457406
rect 410701 457403 410767 457406
rect 411294 457404 411300 457468
rect 411364 457466 411370 457468
rect 412265 457466 412331 457469
rect 411364 457464 412331 457466
rect 411364 457408 412270 457464
rect 412326 457408 412331 457464
rect 411364 457406 412331 457408
rect 412590 457466 412650 457542
rect 580441 457466 580507 457469
rect 412590 457464 580507 457466
rect 412590 457408 580446 457464
rect 580502 457408 580507 457464
rect 412590 457406 580507 457408
rect 411364 457404 411370 457406
rect 412265 457403 412331 457406
rect 580441 457403 580507 457406
rect 233804 456862 405474 456922
rect 233804 456860 233810 456862
rect 233601 456378 233667 456381
rect 385350 456378 385356 456380
rect 233601 456376 385356 456378
rect 233601 456320 233606 456376
rect 233662 456320 385356 456376
rect 233601 456318 385356 456320
rect 233601 456315 233667 456318
rect 385350 456316 385356 456318
rect 385420 456316 385426 456380
rect 233785 456242 233851 456245
rect 390134 456242 390140 456244
rect 233785 456240 390140 456242
rect 233785 456184 233790 456240
rect 233846 456184 390140 456240
rect 233785 456182 390140 456184
rect 233785 456179 233851 456182
rect 390134 456180 390140 456182
rect 390204 456180 390210 456244
rect 233969 456106 234035 456109
rect 394918 456106 394924 456108
rect 233969 456104 394924 456106
rect 233969 456048 233974 456104
rect 234030 456048 394924 456104
rect 233969 456046 394924 456048
rect 233969 456043 234035 456046
rect 394918 456044 394924 456046
rect 394988 456044 394994 456108
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 580073 431626 580139 431629
rect 583520 431626 584960 431716
rect 580073 431624 584960 431626
rect 580073 431568 580078 431624
rect 580134 431568 584960 431624
rect 580073 431566 584960 431568
rect 580073 431563 580139 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 3233 423602 3299 423605
rect -960 423600 3299 423602
rect -960 423544 3238 423600
rect 3294 423544 3299 423600
rect -960 423542 3299 423544
rect -960 423452 480 423542
rect 3233 423539 3299 423542
rect 579981 418298 580047 418301
rect 583520 418298 584960 418388
rect 579981 418296 584960 418298
rect 579981 418240 579986 418296
rect 580042 418240 584960 418296
rect 579981 418238 584960 418240
rect 579981 418235 580047 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3325 410546 3391 410549
rect -960 410544 3391 410546
rect -960 410488 3330 410544
rect 3386 410488 3391 410544
rect -960 410486 3391 410488
rect -960 410396 480 410486
rect 3325 410483 3391 410486
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 4061 397490 4127 397493
rect -960 397488 4127 397490
rect -960 397432 4066 397488
rect 4122 397432 4127 397488
rect -960 397430 4127 397432
rect -960 397340 480 397430
rect 4061 397427 4127 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580901 378450 580967 378453
rect 583520 378450 584960 378540
rect 580901 378448 584960 378450
rect 580901 378392 580906 378448
rect 580962 378392 584960 378448
rect 580901 378390 584960 378392
rect 580901 378387 580967 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3969 371378 4035 371381
rect -960 371376 4035 371378
rect -960 371320 3974 371376
rect 4030 371320 4035 371376
rect -960 371318 4035 371320
rect -960 371228 480 371318
rect 3969 371315 4035 371318
rect 580809 365122 580875 365125
rect 583520 365122 584960 365212
rect 580809 365120 584960 365122
rect 580809 365064 580814 365120
rect 580870 365064 584960 365120
rect 580809 365062 584960 365064
rect 580809 365059 580875 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3877 358458 3943 358461
rect -960 358456 3943 358458
rect -960 358400 3882 358456
rect 3938 358400 3943 358456
rect -960 358398 3943 358400
rect -960 358308 480 358398
rect 3877 358395 3943 358398
rect 580717 351930 580783 351933
rect 583520 351930 584960 352020
rect 580717 351928 584960 351930
rect 580717 351872 580722 351928
rect 580778 351872 584960 351928
rect 580717 351870 584960 351872
rect 580717 351867 580783 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3785 345402 3851 345405
rect -960 345400 3851 345402
rect -960 345344 3790 345400
rect 3846 345344 3851 345400
rect -960 345342 3851 345344
rect -960 345252 480 345342
rect 3785 345339 3851 345342
rect 583520 338452 584960 338692
rect 38653 336018 38719 336021
rect 247033 336018 247099 336021
rect 38653 336016 247099 336018
rect 38653 335960 38658 336016
rect 38714 335960 247038 336016
rect 247094 335960 247099 336016
rect 38653 335958 247099 335960
rect 38653 335955 38719 335958
rect 247033 335955 247099 335958
rect 276013 336018 276079 336021
rect 320265 336018 320331 336021
rect 276013 336016 320331 336018
rect 276013 335960 276018 336016
rect 276074 335960 320270 336016
rect 320326 335960 320331 336016
rect 276013 335958 320331 335960
rect 276013 335955 276079 335958
rect 320265 335955 320331 335958
rect 361021 336018 361087 336021
rect 377397 336018 377463 336021
rect 361021 336016 377463 336018
rect 361021 335960 361026 336016
rect 361082 335960 377402 336016
rect 377458 335960 377463 336016
rect 361021 335958 377463 335960
rect 361021 335955 361087 335958
rect 377397 335955 377463 335958
rect 414749 336018 414815 336021
rect 454677 336018 454743 336021
rect 414749 336016 454743 336018
rect 414749 335960 414754 336016
rect 414810 335960 454682 336016
rect 454738 335960 454743 336016
rect 414749 335958 454743 335960
rect 414749 335955 414815 335958
rect 454677 335955 454743 335958
rect -960 332196 480 332436
rect 580717 325274 580783 325277
rect 583520 325274 584960 325364
rect 580717 325272 584960 325274
rect 580717 325216 580722 325272
rect 580778 325216 584960 325272
rect 580717 325214 584960 325216
rect 580717 325211 580783 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3693 319290 3759 319293
rect -960 319288 3759 319290
rect -960 319232 3698 319288
rect 3754 319232 3759 319288
rect -960 319230 3759 319232
rect -960 319140 480 319230
rect 3693 319227 3759 319230
rect 578877 312082 578943 312085
rect 583520 312082 584960 312172
rect 578877 312080 584960 312082
rect 578877 312024 578882 312080
rect 578938 312024 584960 312080
rect 578877 312022 584960 312024
rect 578877 312019 578943 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3325 306234 3391 306237
rect -960 306232 3391 306234
rect -960 306176 3330 306232
rect 3386 306176 3391 306232
rect -960 306174 3391 306176
rect -960 306084 480 306174
rect 3325 306171 3391 306174
rect 579613 298754 579679 298757
rect 583520 298754 584960 298844
rect 579613 298752 584960 298754
rect 579613 298696 579618 298752
rect 579674 298696 584960 298752
rect 579613 298694 584960 298696
rect 579613 298691 579679 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3601 293178 3667 293181
rect -960 293176 3667 293178
rect -960 293120 3606 293176
rect 3662 293120 3667 293176
rect -960 293118 3667 293120
rect -960 293028 480 293118
rect 3601 293115 3667 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3509 267202 3575 267205
rect -960 267200 3575 267202
rect -960 267144 3514 267200
rect 3570 267144 3575 267200
rect -960 267142 3575 267144
rect -960 267052 480 267142
rect 3509 267139 3575 267142
rect 579797 258906 579863 258909
rect 583520 258906 584960 258996
rect 579797 258904 584960 258906
rect 579797 258848 579802 258904
rect 579858 258848 584960 258904
rect 579797 258846 584960 258848
rect 579797 258843 579863 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 3141 254146 3207 254149
rect -960 254144 3207 254146
rect -960 254088 3146 254144
rect 3202 254088 3207 254144
rect -960 254086 3207 254088
rect -960 253996 480 254086
rect 3141 254083 3207 254086
rect 580625 245578 580691 245581
rect 583520 245578 584960 245668
rect 580625 245576 584960 245578
rect 580625 245520 580630 245576
rect 580686 245520 584960 245576
rect 580625 245518 584960 245520
rect 580625 245515 580691 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 3509 241090 3575 241093
rect -960 241088 3575 241090
rect -960 241032 3514 241088
rect 3570 241032 3575 241088
rect -960 241030 3575 241032
rect -960 240940 480 241030
rect 3509 241027 3575 241030
rect 579613 232386 579679 232389
rect 583520 232386 584960 232476
rect 579613 232384 584960 232386
rect 579613 232328 579618 232384
rect 579674 232328 584960 232384
rect 579613 232326 584960 232328
rect 579613 232323 579679 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580165 219058 580231 219061
rect 583520 219058 584960 219148
rect 580165 219056 584960 219058
rect 580165 219000 580170 219056
rect 580226 219000 584960 219056
rect 580165 218998 584960 219000
rect 580165 218995 580231 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 3417 214978 3483 214981
rect -960 214976 3483 214978
rect -960 214920 3422 214976
rect 3478 214920 3483 214976
rect -960 214918 3483 214920
rect -960 214828 480 214918
rect 3417 214915 3483 214918
rect 580533 205730 580599 205733
rect 583520 205730 584960 205820
rect 580533 205728 584960 205730
rect 580533 205672 580538 205728
rect 580594 205672 584960 205728
rect 580533 205670 584960 205672
rect 580533 205667 580599 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 3417 201922 3483 201925
rect -960 201920 3483 201922
rect -960 201864 3422 201920
rect 3478 201864 3483 201920
rect -960 201862 3483 201864
rect -960 201772 480 201862
rect 3417 201859 3483 201862
rect 579613 192538 579679 192541
rect 583520 192538 584960 192628
rect 579613 192536 584960 192538
rect 579613 192480 579618 192536
rect 579674 192480 584960 192536
rect 579613 192478 584960 192480
rect 579613 192475 579679 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 3417 188866 3483 188869
rect -960 188864 3483 188866
rect -960 188808 3422 188864
rect 3478 188808 3483 188864
rect -960 188806 3483 188808
rect -960 188716 480 188806
rect 3417 188803 3483 188806
rect 580073 179210 580139 179213
rect 583520 179210 584960 179300
rect 580073 179208 584960 179210
rect 580073 179152 580078 179208
rect 580134 179152 584960 179208
rect 580073 179150 584960 179152
rect 580073 179147 580139 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580441 165882 580507 165885
rect 583520 165882 584960 165972
rect 580441 165880 584960 165882
rect 580441 165824 580446 165880
rect 580502 165824 584960 165880
rect 580441 165822 584960 165824
rect 580441 165819 580507 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 580349 152690 580415 152693
rect 583520 152690 584960 152780
rect 580349 152688 584960 152690
rect 580349 152632 580354 152688
rect 580410 152632 584960 152688
rect 580349 152630 584960 152632
rect 580349 152627 580415 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3417 149834 3483 149837
rect -960 149832 3483 149834
rect -960 149776 3422 149832
rect 3478 149776 3483 149832
rect -960 149774 3483 149776
rect -960 149684 480 149774
rect 3417 149771 3483 149774
rect 579613 139362 579679 139365
rect 583520 139362 584960 139452
rect 579613 139360 584960 139362
rect 579613 139304 579618 139360
rect 579674 139304 584960 139360
rect 579613 139302 584960 139304
rect 579613 139299 579679 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3233 136778 3299 136781
rect -960 136776 3299 136778
rect -960 136720 3238 136776
rect 3294 136720 3299 136776
rect -960 136718 3299 136720
rect -960 136628 480 136718
rect 3233 136715 3299 136718
rect 580257 126034 580323 126037
rect 583520 126034 584960 126124
rect 580257 126032 584960 126034
rect 580257 125976 580262 126032
rect 580318 125976 584960 126032
rect 580257 125974 584960 125976
rect 580257 125971 580323 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580533 112842 580599 112845
rect 583520 112842 584960 112932
rect 580533 112840 584960 112842
rect 580533 112784 580538 112840
rect 580594 112784 584960 112840
rect 580533 112782 584960 112784
rect 580533 112779 580599 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 3366 110666 3372 110668
rect -960 110606 3372 110666
rect -960 110516 480 110606
rect 3366 110604 3372 110606
rect 3436 110604 3442 110668
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 3417 97610 3483 97613
rect -960 97608 3483 97610
rect -960 97552 3422 97608
rect 3478 97552 3483 97608
rect -960 97550 3483 97552
rect -960 97460 480 97550
rect 3417 97547 3483 97550
rect 580390 86124 580396 86188
rect 580460 86186 580466 86188
rect 583520 86186 584960 86276
rect 580460 86126 584960 86186
rect 580460 86124 580466 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3141 84690 3207 84693
rect -960 84688 3207 84690
rect -960 84632 3146 84688
rect 3202 84632 3207 84688
rect -960 84630 3207 84632
rect -960 84540 480 84630
rect 3141 84627 3207 84630
rect 579705 72994 579771 72997
rect 583520 72994 584960 73084
rect 579705 72992 584960 72994
rect 579705 72936 579710 72992
rect 579766 72936 584960 72992
rect 579705 72934 584960 72936
rect 579705 72931 579771 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 2773 71634 2839 71637
rect -960 71632 2839 71634
rect -960 71576 2778 71632
rect 2834 71576 2839 71632
rect -960 71574 2839 71576
rect -960 71484 480 71574
rect 2773 71571 2839 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect -960 58518 674 58578
rect -960 58442 480 58518
rect 614 58442 674 58518
rect -960 58428 674 58442
rect 246 58382 674 58428
rect 246 58034 306 58382
rect 408718 58034 408724 58036
rect 246 57974 408724 58034
rect 408718 57972 408724 57974
rect 408788 57972 408794 58036
rect 580206 46276 580212 46340
rect 580276 46338 580282 46340
rect 583520 46338 584960 46428
rect 580276 46278 584960 46338
rect 580276 46276 580282 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect -960 45462 674 45522
rect -960 45386 480 45462
rect 614 45386 674 45462
rect -960 45372 674 45386
rect 246 45326 674 45372
rect 246 44842 306 45326
rect 246 44782 6930 44842
rect 6870 44298 6930 44782
rect 233734 44298 233740 44300
rect 6870 44238 233740 44298
rect 233734 44236 233740 44238
rect 233804 44236 233810 44300
rect 579613 33146 579679 33149
rect 583520 33146 584960 33236
rect 579613 33144 584960 33146
rect 579613 33088 579618 33144
rect 579674 33088 584960 33144
rect 579613 33086 584960 33088
rect 579613 33083 579679 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect -960 32406 674 32466
rect -960 32330 480 32406
rect 614 32330 674 32406
rect -960 32316 674 32330
rect 246 32270 674 32316
rect 246 31786 306 32270
rect 409822 31786 409828 31788
rect 246 31726 409828 31786
rect 409822 31724 409828 31726
rect 409892 31724 409898 31788
rect 3509 19954 3575 19957
rect 411294 19954 411300 19956
rect 3509 19952 411300 19954
rect 3509 19896 3514 19952
rect 3570 19896 411300 19952
rect 3509 19894 411300 19896
rect 3509 19891 3575 19894
rect 411294 19892 411300 19894
rect 411364 19892 411370 19956
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 9673 18594 9739 18597
rect 237649 18594 237715 18597
rect 9673 18592 237715 18594
rect 9673 18536 9678 18592
rect 9734 18536 237654 18592
rect 237710 18536 237715 18592
rect 9673 18534 237715 18536
rect 9673 18531 9739 18534
rect 237649 18531 237715 18534
rect 131113 17234 131179 17237
rect 274909 17234 274975 17237
rect 131113 17232 274975 17234
rect 131113 17176 131118 17232
rect 131174 17176 274914 17232
rect 274970 17176 274975 17232
rect 131113 17174 274975 17176
rect 131113 17171 131179 17174
rect 274909 17171 274975 17174
rect 105 15874 171 15877
rect 234613 15874 234679 15877
rect 105 15872 234679 15874
rect 105 15816 110 15872
rect 166 15816 234618 15872
rect 234674 15816 234679 15872
rect 105 15814 234679 15816
rect 105 15811 171 15814
rect 234613 15811 234679 15814
rect 22553 14514 22619 14517
rect 241697 14514 241763 14517
rect 22553 14512 241763 14514
rect 22553 14456 22558 14512
rect 22614 14456 241702 14512
rect 241758 14456 241763 14512
rect 22553 14454 241763 14456
rect 22553 14451 22619 14454
rect 241697 14451 241763 14454
rect 40217 13018 40283 13021
rect 247125 13018 247191 13021
rect 40217 13016 247191 13018
rect 40217 12960 40222 13016
rect 40278 12960 247130 13016
rect 247186 12960 247191 13016
rect 40217 12958 247191 12960
rect 40217 12955 40283 12958
rect 247125 12955 247191 12958
rect 8753 11658 8819 11661
rect 237557 11658 237623 11661
rect 8753 11656 237623 11658
rect 8753 11600 8758 11656
rect 8814 11600 237562 11656
rect 237618 11600 237623 11656
rect 8753 11598 237623 11600
rect 8753 11595 8819 11598
rect 237557 11595 237623 11598
rect 79225 10298 79291 10301
rect 259545 10298 259611 10301
rect 79225 10296 259611 10298
rect 79225 10240 79230 10296
rect 79286 10240 259550 10296
rect 259606 10240 259611 10296
rect 79225 10238 259611 10240
rect 79225 10235 79291 10238
rect 259545 10235 259611 10238
rect 17033 8938 17099 8941
rect 240317 8938 240383 8941
rect 17033 8936 240383 8938
rect 17033 8880 17038 8936
rect 17094 8880 240322 8936
rect 240378 8880 240383 8936
rect 17033 8878 240383 8880
rect 17033 8875 17099 8878
rect 240317 8875 240383 8878
rect 412725 8938 412791 8941
rect 577405 8938 577471 8941
rect 412725 8936 577471 8938
rect 412725 8880 412730 8936
rect 412786 8880 577410 8936
rect 577466 8880 577471 8936
rect 412725 8878 577471 8880
rect 412725 8875 412791 8878
rect 577405 8875 577471 8878
rect 162485 7578 162551 7581
rect 284385 7578 284451 7581
rect 162485 7576 284451 7578
rect 162485 7520 162490 7576
rect 162546 7520 284390 7576
rect 284446 7520 284451 7576
rect 162485 7518 284451 7520
rect 162485 7515 162551 7518
rect 284385 7515 284451 7518
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect 583520 6476 584960 6566
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 228725 6218 228791 6221
rect 304993 6218 305059 6221
rect 228725 6216 305059 6218
rect 228725 6160 228730 6216
rect 228786 6160 304998 6216
rect 305054 6160 305059 6216
rect 228725 6158 305059 6160
rect 228725 6155 228791 6158
rect 304993 6155 305059 6158
rect 411345 6218 411411 6221
rect 572713 6218 572779 6221
rect 411345 6216 572779 6218
rect 411345 6160 411350 6216
rect 411406 6160 572718 6216
rect 572774 6160 572779 6216
rect 411345 6158 572779 6160
rect 411345 6155 411411 6158
rect 572713 6155 572779 6158
rect 296897 4994 296963 4997
rect 277350 4992 296963 4994
rect 277350 4936 296902 4992
rect 296958 4936 296963 4992
rect 277350 4934 296963 4936
rect 200297 4858 200363 4861
rect 277350 4858 277410 4934
rect 296897 4931 296963 4934
rect 200297 4856 277410 4858
rect 200297 4800 200302 4856
rect 200358 4800 277410 4856
rect 200297 4798 277410 4800
rect 297725 4858 297791 4861
rect 309317 4858 309383 4861
rect 297725 4856 309383 4858
rect 297725 4800 297730 4856
rect 297786 4800 309322 4856
rect 309378 4800 309383 4856
rect 297725 4798 309383 4800
rect 200297 4795 200363 4798
rect 297725 4795 297791 4798
rect 309317 4795 309383 4798
rect 397453 4858 397519 4861
rect 530117 4858 530183 4861
rect 397453 4856 530183 4858
rect 397453 4800 397458 4856
rect 397514 4800 530122 4856
rect 530178 4800 530183 4856
rect 397453 4798 530183 4800
rect 397453 4795 397519 4798
rect 530117 4795 530183 4798
rect 300761 3498 300827 3501
rect 327165 3498 327231 3501
rect 300761 3496 327231 3498
rect 300761 3440 300766 3496
rect 300822 3440 327170 3496
rect 327226 3440 327231 3496
rect 300761 3438 327231 3440
rect 300761 3435 300827 3438
rect 327165 3435 327231 3438
rect 5257 3362 5323 3365
rect 236269 3362 236335 3365
rect 5257 3360 236335 3362
rect 5257 3304 5262 3360
rect 5318 3304 236274 3360
rect 236330 3304 236335 3360
rect 5257 3302 236335 3304
rect 5257 3299 5323 3302
rect 236269 3299 236335 3302
rect 241697 3362 241763 3365
rect 309225 3362 309291 3365
rect 241697 3360 309291 3362
rect 241697 3304 241702 3360
rect 241758 3304 309230 3360
rect 309286 3304 309291 3360
rect 241697 3302 309291 3304
rect 241697 3299 241763 3302
rect 309225 3299 309291 3302
rect 373257 3362 373323 3365
rect 404813 3362 404879 3365
rect 373257 3360 404879 3362
rect 373257 3304 373262 3360
rect 373318 3304 404818 3360
rect 404874 3304 404879 3360
rect 373257 3302 404879 3304
rect 373257 3299 373323 3302
rect 404813 3299 404879 3302
rect 414013 3362 414079 3365
rect 582189 3362 582255 3365
rect 414013 3360 582255 3362
rect 414013 3304 414018 3360
rect 414074 3304 582194 3360
rect 582250 3304 582255 3360
rect 414013 3302 582255 3304
rect 414013 3299 414079 3302
rect 582189 3299 582255 3302
<< via3 >>
rect 580396 458628 580460 458692
rect 580212 458492 580276 458556
rect 3372 458356 3436 458420
rect 385356 457464 385420 457468
rect 385356 457408 385406 457464
rect 385406 457408 385420 457464
rect 385356 457404 385420 457408
rect 390140 457464 390204 457468
rect 390140 457408 390190 457464
rect 390190 457408 390204 457464
rect 390140 457404 390204 457408
rect 394924 457464 394988 457468
rect 394924 457408 394974 457464
rect 394974 457408 394988 457464
rect 394924 457404 394988 457408
rect 233740 456860 233804 456924
rect 408724 457404 408788 457468
rect 409828 457404 409892 457468
rect 411300 457404 411364 457468
rect 385356 456316 385420 456380
rect 390140 456180 390204 456244
rect 394924 456044 394988 456108
rect 3372 110604 3436 110668
rect 580396 86124 580460 86188
rect 408724 57972 408788 58036
rect 580212 46276 580276 46340
rect 233740 44236 233804 44300
rect 409828 31724 409892 31788
rect 411300 19892 411364 19956
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711002 -8694 711558
rect -8138 711002 -8106 711558
rect -8726 680614 -8106 711002
rect -8726 680058 -8694 680614
rect -8138 680058 -8106 680614
rect -8726 644614 -8106 680058
rect -8726 644058 -8694 644614
rect -8138 644058 -8106 644614
rect -8726 608614 -8106 644058
rect -8726 608058 -8694 608614
rect -8138 608058 -8106 608614
rect -8726 572614 -8106 608058
rect -8726 572058 -8694 572614
rect -8138 572058 -8106 572614
rect -8726 536614 -8106 572058
rect -8726 536058 -8694 536614
rect -8138 536058 -8106 536614
rect -8726 500614 -8106 536058
rect -8726 500058 -8694 500614
rect -8138 500058 -8106 500614
rect -8726 464614 -8106 500058
rect -8726 464058 -8694 464614
rect -8138 464058 -8106 464614
rect -8726 428614 -8106 464058
rect -8726 428058 -8694 428614
rect -8138 428058 -8106 428614
rect -8726 392614 -8106 428058
rect -8726 392058 -8694 392614
rect -8138 392058 -8106 392614
rect -8726 356614 -8106 392058
rect -8726 356058 -8694 356614
rect -8138 356058 -8106 356614
rect -8726 320614 -8106 356058
rect -8726 320058 -8694 320614
rect -8138 320058 -8106 320614
rect -8726 284614 -8106 320058
rect -8726 284058 -8694 284614
rect -8138 284058 -8106 284614
rect -8726 248614 -8106 284058
rect -8726 248058 -8694 248614
rect -8138 248058 -8106 248614
rect -8726 212614 -8106 248058
rect -8726 212058 -8694 212614
rect -8138 212058 -8106 212614
rect -8726 176614 -8106 212058
rect -8726 176058 -8694 176614
rect -8138 176058 -8106 176614
rect -8726 140614 -8106 176058
rect -8726 140058 -8694 140614
rect -8138 140058 -8106 140614
rect -8726 104614 -8106 140058
rect -8726 104058 -8694 104614
rect -8138 104058 -8106 104614
rect -8726 68614 -8106 104058
rect -8726 68058 -8694 68614
rect -8138 68058 -8106 68614
rect -8726 32614 -8106 68058
rect -8726 32058 -8694 32614
rect -8138 32058 -8106 32614
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710042 -7734 710598
rect -7178 710042 -7146 710598
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710042 12986 710598
rect 13542 710042 13574 710598
rect -7766 698058 -7734 698614
rect -7178 698058 -7146 698614
rect -7766 662614 -7146 698058
rect -7766 662058 -7734 662614
rect -7178 662058 -7146 662614
rect -7766 626614 -7146 662058
rect -7766 626058 -7734 626614
rect -7178 626058 -7146 626614
rect -7766 590614 -7146 626058
rect -7766 590058 -7734 590614
rect -7178 590058 -7146 590614
rect -7766 554614 -7146 590058
rect -7766 554058 -7734 554614
rect -7178 554058 -7146 554614
rect -7766 518614 -7146 554058
rect -7766 518058 -7734 518614
rect -7178 518058 -7146 518614
rect -7766 482614 -7146 518058
rect -7766 482058 -7734 482614
rect -7178 482058 -7146 482614
rect -7766 446614 -7146 482058
rect -7766 446058 -7734 446614
rect -7178 446058 -7146 446614
rect -7766 410614 -7146 446058
rect -7766 410058 -7734 410614
rect -7178 410058 -7146 410614
rect -7766 374614 -7146 410058
rect -7766 374058 -7734 374614
rect -7178 374058 -7146 374614
rect -7766 338614 -7146 374058
rect -7766 338058 -7734 338614
rect -7178 338058 -7146 338614
rect -7766 302614 -7146 338058
rect -7766 302058 -7734 302614
rect -7178 302058 -7146 302614
rect -7766 266614 -7146 302058
rect -7766 266058 -7734 266614
rect -7178 266058 -7146 266614
rect -7766 230614 -7146 266058
rect -7766 230058 -7734 230614
rect -7178 230058 -7146 230614
rect -7766 194614 -7146 230058
rect -7766 194058 -7734 194614
rect -7178 194058 -7146 194614
rect -7766 158614 -7146 194058
rect -7766 158058 -7734 158614
rect -7178 158058 -7146 158614
rect -7766 122614 -7146 158058
rect -7766 122058 -7734 122614
rect -7178 122058 -7146 122614
rect -7766 86614 -7146 122058
rect -7766 86058 -7734 86614
rect -7178 86058 -7146 86614
rect -7766 50614 -7146 86058
rect -7766 50058 -7734 50614
rect -7178 50058 -7146 50614
rect -7766 14614 -7146 50058
rect -7766 14058 -7734 14614
rect -7178 14058 -7146 14614
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709082 -6774 709638
rect -6218 709082 -6186 709638
rect -6806 676894 -6186 709082
rect -6806 676338 -6774 676894
rect -6218 676338 -6186 676894
rect -6806 640894 -6186 676338
rect -6806 640338 -6774 640894
rect -6218 640338 -6186 640894
rect -6806 604894 -6186 640338
rect -6806 604338 -6774 604894
rect -6218 604338 -6186 604894
rect -6806 568894 -6186 604338
rect -6806 568338 -6774 568894
rect -6218 568338 -6186 568894
rect -6806 532894 -6186 568338
rect -6806 532338 -6774 532894
rect -6218 532338 -6186 532894
rect -6806 496894 -6186 532338
rect -6806 496338 -6774 496894
rect -6218 496338 -6186 496894
rect -6806 460894 -6186 496338
rect -6806 460338 -6774 460894
rect -6218 460338 -6186 460894
rect -6806 424894 -6186 460338
rect -6806 424338 -6774 424894
rect -6218 424338 -6186 424894
rect -6806 388894 -6186 424338
rect -6806 388338 -6774 388894
rect -6218 388338 -6186 388894
rect -6806 352894 -6186 388338
rect -6806 352338 -6774 352894
rect -6218 352338 -6186 352894
rect -6806 316894 -6186 352338
rect -6806 316338 -6774 316894
rect -6218 316338 -6186 316894
rect -6806 280894 -6186 316338
rect -6806 280338 -6774 280894
rect -6218 280338 -6186 280894
rect -6806 244894 -6186 280338
rect -6806 244338 -6774 244894
rect -6218 244338 -6186 244894
rect -6806 208894 -6186 244338
rect -6806 208338 -6774 208894
rect -6218 208338 -6186 208894
rect -6806 172894 -6186 208338
rect -6806 172338 -6774 172894
rect -6218 172338 -6186 172894
rect -6806 136894 -6186 172338
rect -6806 136338 -6774 136894
rect -6218 136338 -6186 136894
rect -6806 100894 -6186 136338
rect -6806 100338 -6774 100894
rect -6218 100338 -6186 100894
rect -6806 64894 -6186 100338
rect -6806 64338 -6774 64894
rect -6218 64338 -6186 64894
rect -6806 28894 -6186 64338
rect -6806 28338 -6774 28894
rect -6218 28338 -6186 28894
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708122 -5814 708678
rect -5258 708122 -5226 708678
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708122 9266 708678
rect 9822 708122 9854 708678
rect -5846 694338 -5814 694894
rect -5258 694338 -5226 694894
rect -5846 658894 -5226 694338
rect -5846 658338 -5814 658894
rect -5258 658338 -5226 658894
rect -5846 622894 -5226 658338
rect -5846 622338 -5814 622894
rect -5258 622338 -5226 622894
rect -5846 586894 -5226 622338
rect -5846 586338 -5814 586894
rect -5258 586338 -5226 586894
rect -5846 550894 -5226 586338
rect -5846 550338 -5814 550894
rect -5258 550338 -5226 550894
rect -5846 514894 -5226 550338
rect -5846 514338 -5814 514894
rect -5258 514338 -5226 514894
rect -5846 478894 -5226 514338
rect -5846 478338 -5814 478894
rect -5258 478338 -5226 478894
rect -5846 442894 -5226 478338
rect -5846 442338 -5814 442894
rect -5258 442338 -5226 442894
rect -5846 406894 -5226 442338
rect -5846 406338 -5814 406894
rect -5258 406338 -5226 406894
rect -5846 370894 -5226 406338
rect -5846 370338 -5814 370894
rect -5258 370338 -5226 370894
rect -5846 334894 -5226 370338
rect -5846 334338 -5814 334894
rect -5258 334338 -5226 334894
rect -5846 298894 -5226 334338
rect -5846 298338 -5814 298894
rect -5258 298338 -5226 298894
rect -5846 262894 -5226 298338
rect -5846 262338 -5814 262894
rect -5258 262338 -5226 262894
rect -5846 226894 -5226 262338
rect -5846 226338 -5814 226894
rect -5258 226338 -5226 226894
rect -5846 190894 -5226 226338
rect -5846 190338 -5814 190894
rect -5258 190338 -5226 190894
rect -5846 154894 -5226 190338
rect -5846 154338 -5814 154894
rect -5258 154338 -5226 154894
rect -5846 118894 -5226 154338
rect -5846 118338 -5814 118894
rect -5258 118338 -5226 118894
rect -5846 82894 -5226 118338
rect -5846 82338 -5814 82894
rect -5258 82338 -5226 82894
rect -5846 46894 -5226 82338
rect -5846 46338 -5814 46894
rect -5258 46338 -5226 46894
rect -5846 10894 -5226 46338
rect -5846 10338 -5814 10894
rect -5258 10338 -5226 10894
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707162 -4854 707718
rect -4298 707162 -4266 707718
rect -4886 673174 -4266 707162
rect -4886 672618 -4854 673174
rect -4298 672618 -4266 673174
rect -4886 637174 -4266 672618
rect -4886 636618 -4854 637174
rect -4298 636618 -4266 637174
rect -4886 601174 -4266 636618
rect -4886 600618 -4854 601174
rect -4298 600618 -4266 601174
rect -4886 565174 -4266 600618
rect -4886 564618 -4854 565174
rect -4298 564618 -4266 565174
rect -4886 529174 -4266 564618
rect -4886 528618 -4854 529174
rect -4298 528618 -4266 529174
rect -4886 493174 -4266 528618
rect -4886 492618 -4854 493174
rect -4298 492618 -4266 493174
rect -4886 457174 -4266 492618
rect -4886 456618 -4854 457174
rect -4298 456618 -4266 457174
rect -4886 421174 -4266 456618
rect -4886 420618 -4854 421174
rect -4298 420618 -4266 421174
rect -4886 385174 -4266 420618
rect -4886 384618 -4854 385174
rect -4298 384618 -4266 385174
rect -4886 349174 -4266 384618
rect -4886 348618 -4854 349174
rect -4298 348618 -4266 349174
rect -4886 313174 -4266 348618
rect -4886 312618 -4854 313174
rect -4298 312618 -4266 313174
rect -4886 277174 -4266 312618
rect -4886 276618 -4854 277174
rect -4298 276618 -4266 277174
rect -4886 241174 -4266 276618
rect -4886 240618 -4854 241174
rect -4298 240618 -4266 241174
rect -4886 205174 -4266 240618
rect -4886 204618 -4854 205174
rect -4298 204618 -4266 205174
rect -4886 169174 -4266 204618
rect -4886 168618 -4854 169174
rect -4298 168618 -4266 169174
rect -4886 133174 -4266 168618
rect -4886 132618 -4854 133174
rect -4298 132618 -4266 133174
rect -4886 97174 -4266 132618
rect -4886 96618 -4854 97174
rect -4298 96618 -4266 97174
rect -4886 61174 -4266 96618
rect -4886 60618 -4854 61174
rect -4298 60618 -4266 61174
rect -4886 25174 -4266 60618
rect -4886 24618 -4854 25174
rect -4298 24618 -4266 25174
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706202 -3894 706758
rect -3338 706202 -3306 706758
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706202 5546 706758
rect 6102 706202 6134 706758
rect -3926 690618 -3894 691174
rect -3338 690618 -3306 691174
rect -3926 655174 -3306 690618
rect -3926 654618 -3894 655174
rect -3338 654618 -3306 655174
rect -3926 619174 -3306 654618
rect -3926 618618 -3894 619174
rect -3338 618618 -3306 619174
rect -3926 583174 -3306 618618
rect -3926 582618 -3894 583174
rect -3338 582618 -3306 583174
rect -3926 547174 -3306 582618
rect -3926 546618 -3894 547174
rect -3338 546618 -3306 547174
rect -3926 511174 -3306 546618
rect -3926 510618 -3894 511174
rect -3338 510618 -3306 511174
rect -3926 475174 -3306 510618
rect -3926 474618 -3894 475174
rect -3338 474618 -3306 475174
rect -3926 439174 -3306 474618
rect -3926 438618 -3894 439174
rect -3338 438618 -3306 439174
rect -3926 403174 -3306 438618
rect -3926 402618 -3894 403174
rect -3338 402618 -3306 403174
rect -3926 367174 -3306 402618
rect -3926 366618 -3894 367174
rect -3338 366618 -3306 367174
rect -3926 331174 -3306 366618
rect -3926 330618 -3894 331174
rect -3338 330618 -3306 331174
rect -3926 295174 -3306 330618
rect -3926 294618 -3894 295174
rect -3338 294618 -3306 295174
rect -3926 259174 -3306 294618
rect -3926 258618 -3894 259174
rect -3338 258618 -3306 259174
rect -3926 223174 -3306 258618
rect -3926 222618 -3894 223174
rect -3338 222618 -3306 223174
rect -3926 187174 -3306 222618
rect -3926 186618 -3894 187174
rect -3338 186618 -3306 187174
rect -3926 151174 -3306 186618
rect -3926 150618 -3894 151174
rect -3338 150618 -3306 151174
rect -3926 115174 -3306 150618
rect -3926 114618 -3894 115174
rect -3338 114618 -3306 115174
rect -3926 79174 -3306 114618
rect -3926 78618 -3894 79174
rect -3338 78618 -3306 79174
rect -3926 43174 -3306 78618
rect -3926 42618 -3894 43174
rect -3338 42618 -3306 43174
rect -3926 7174 -3306 42618
rect -3926 6618 -3894 7174
rect -3338 6618 -3306 7174
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705242 -2934 705798
rect -2378 705242 -2346 705798
rect -2966 669454 -2346 705242
rect -2966 668898 -2934 669454
rect -2378 668898 -2346 669454
rect -2966 633454 -2346 668898
rect -2966 632898 -2934 633454
rect -2378 632898 -2346 633454
rect -2966 597454 -2346 632898
rect -2966 596898 -2934 597454
rect -2378 596898 -2346 597454
rect -2966 561454 -2346 596898
rect -2966 560898 -2934 561454
rect -2378 560898 -2346 561454
rect -2966 525454 -2346 560898
rect -2966 524898 -2934 525454
rect -2378 524898 -2346 525454
rect -2966 489454 -2346 524898
rect -2966 488898 -2934 489454
rect -2378 488898 -2346 489454
rect -2966 453454 -2346 488898
rect -2966 452898 -2934 453454
rect -2378 452898 -2346 453454
rect -2966 417454 -2346 452898
rect -2966 416898 -2934 417454
rect -2378 416898 -2346 417454
rect -2966 381454 -2346 416898
rect -2966 380898 -2934 381454
rect -2378 380898 -2346 381454
rect -2966 345454 -2346 380898
rect -2966 344898 -2934 345454
rect -2378 344898 -2346 345454
rect -2966 309454 -2346 344898
rect -2966 308898 -2934 309454
rect -2378 308898 -2346 309454
rect -2966 273454 -2346 308898
rect -2966 272898 -2934 273454
rect -2378 272898 -2346 273454
rect -2966 237454 -2346 272898
rect -2966 236898 -2934 237454
rect -2378 236898 -2346 237454
rect -2966 201454 -2346 236898
rect -2966 200898 -2934 201454
rect -2378 200898 -2346 201454
rect -2966 165454 -2346 200898
rect -2966 164898 -2934 165454
rect -2378 164898 -2346 165454
rect -2966 129454 -2346 164898
rect -2966 128898 -2934 129454
rect -2378 128898 -2346 129454
rect -2966 93454 -2346 128898
rect -2966 92898 -2934 93454
rect -2378 92898 -2346 93454
rect -2966 57454 -2346 92898
rect -2966 56898 -2934 57454
rect -2378 56898 -2346 57454
rect -2966 21454 -2346 56898
rect -2966 20898 -2934 21454
rect -2378 20898 -2346 21454
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704282 -1974 704838
rect -1418 704282 -1386 704838
rect -2006 687454 -1386 704282
rect -2006 686898 -1974 687454
rect -1418 686898 -1386 687454
rect -2006 651454 -1386 686898
rect -2006 650898 -1974 651454
rect -1418 650898 -1386 651454
rect -2006 615454 -1386 650898
rect -2006 614898 -1974 615454
rect -1418 614898 -1386 615454
rect -2006 579454 -1386 614898
rect -2006 578898 -1974 579454
rect -1418 578898 -1386 579454
rect -2006 543454 -1386 578898
rect -2006 542898 -1974 543454
rect -1418 542898 -1386 543454
rect -2006 507454 -1386 542898
rect -2006 506898 -1974 507454
rect -1418 506898 -1386 507454
rect -2006 471454 -1386 506898
rect -2006 470898 -1974 471454
rect -1418 470898 -1386 471454
rect -2006 435454 -1386 470898
rect -2006 434898 -1974 435454
rect -1418 434898 -1386 435454
rect -2006 399454 -1386 434898
rect -2006 398898 -1974 399454
rect -1418 398898 -1386 399454
rect -2006 363454 -1386 398898
rect -2006 362898 -1974 363454
rect -1418 362898 -1386 363454
rect -2006 327454 -1386 362898
rect -2006 326898 -1974 327454
rect -1418 326898 -1386 327454
rect -2006 291454 -1386 326898
rect -2006 290898 -1974 291454
rect -1418 290898 -1386 291454
rect -2006 255454 -1386 290898
rect -2006 254898 -1974 255454
rect -1418 254898 -1386 255454
rect -2006 219454 -1386 254898
rect -2006 218898 -1974 219454
rect -1418 218898 -1386 219454
rect -2006 183454 -1386 218898
rect -2006 182898 -1974 183454
rect -1418 182898 -1386 183454
rect -2006 147454 -1386 182898
rect -2006 146898 -1974 147454
rect -1418 146898 -1386 147454
rect -2006 111454 -1386 146898
rect -2006 110898 -1974 111454
rect -1418 110898 -1386 111454
rect -2006 75454 -1386 110898
rect -2006 74898 -1974 75454
rect -1418 74898 -1386 75454
rect -2006 39454 -1386 74898
rect -2006 38898 -1974 39454
rect -1418 38898 -1386 39454
rect -2006 3454 -1386 38898
rect -2006 2898 -1974 3454
rect -1418 2898 -1386 3454
rect -2006 -346 -1386 2898
rect -2006 -902 -1974 -346
rect -1418 -902 -1386 -346
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704282 1826 704838
rect 2382 704282 2414 704838
rect 1794 687454 2414 704282
rect 1794 686898 1826 687454
rect 2382 686898 2414 687454
rect 1794 651454 2414 686898
rect 1794 650898 1826 651454
rect 2382 650898 2414 651454
rect 1794 615454 2414 650898
rect 1794 614898 1826 615454
rect 2382 614898 2414 615454
rect 1794 579454 2414 614898
rect 1794 578898 1826 579454
rect 2382 578898 2414 579454
rect 1794 543454 2414 578898
rect 1794 542898 1826 543454
rect 2382 542898 2414 543454
rect 1794 507454 2414 542898
rect 1794 506898 1826 507454
rect 2382 506898 2414 507454
rect 1794 471454 2414 506898
rect 1794 470898 1826 471454
rect 2382 470898 2414 471454
rect 1794 435454 2414 470898
rect 5514 691174 6134 706202
rect 5514 690618 5546 691174
rect 6102 690618 6134 691174
rect 5514 655174 6134 690618
rect 5514 654618 5546 655174
rect 6102 654618 6134 655174
rect 5514 619174 6134 654618
rect 5514 618618 5546 619174
rect 6102 618618 6134 619174
rect 5514 583174 6134 618618
rect 5514 582618 5546 583174
rect 6102 582618 6134 583174
rect 5514 547174 6134 582618
rect 5514 546618 5546 547174
rect 6102 546618 6134 547174
rect 5514 511174 6134 546618
rect 5514 510618 5546 511174
rect 6102 510618 6134 511174
rect 5514 475174 6134 510618
rect 5514 474618 5546 475174
rect 6102 474618 6134 475174
rect 3371 458420 3437 458421
rect 3371 458356 3372 458420
rect 3436 458356 3437 458420
rect 3371 458355 3437 458356
rect 1794 434898 1826 435454
rect 2382 434898 2414 435454
rect 1794 399454 2414 434898
rect 1794 398898 1826 399454
rect 2382 398898 2414 399454
rect 1794 363454 2414 398898
rect 1794 362898 1826 363454
rect 2382 362898 2414 363454
rect 1794 327454 2414 362898
rect 1794 326898 1826 327454
rect 2382 326898 2414 327454
rect 1794 291454 2414 326898
rect 1794 290898 1826 291454
rect 2382 290898 2414 291454
rect 1794 255454 2414 290898
rect 1794 254898 1826 255454
rect 2382 254898 2414 255454
rect 1794 219454 2414 254898
rect 1794 218898 1826 219454
rect 2382 218898 2414 219454
rect 1794 183454 2414 218898
rect 1794 182898 1826 183454
rect 2382 182898 2414 183454
rect 1794 147454 2414 182898
rect 1794 146898 1826 147454
rect 2382 146898 2414 147454
rect 1794 111454 2414 146898
rect 1794 110898 1826 111454
rect 2382 110898 2414 111454
rect 1794 75454 2414 110898
rect 3374 110669 3434 458355
rect 5514 439174 6134 474618
rect 5514 438618 5546 439174
rect 6102 438618 6134 439174
rect 5514 403174 6134 438618
rect 5514 402618 5546 403174
rect 6102 402618 6134 403174
rect 5514 367174 6134 402618
rect 5514 366618 5546 367174
rect 6102 366618 6134 367174
rect 5514 331174 6134 366618
rect 5514 330618 5546 331174
rect 6102 330618 6134 331174
rect 5514 295174 6134 330618
rect 5514 294618 5546 295174
rect 6102 294618 6134 295174
rect 5514 259174 6134 294618
rect 5514 258618 5546 259174
rect 6102 258618 6134 259174
rect 5514 223174 6134 258618
rect 5514 222618 5546 223174
rect 6102 222618 6134 223174
rect 5514 187174 6134 222618
rect 5514 186618 5546 187174
rect 6102 186618 6134 187174
rect 5514 151174 6134 186618
rect 5514 150618 5546 151174
rect 6102 150618 6134 151174
rect 5514 115174 6134 150618
rect 5514 114618 5546 115174
rect 6102 114618 6134 115174
rect 3371 110668 3437 110669
rect 3371 110604 3372 110668
rect 3436 110604 3437 110668
rect 3371 110603 3437 110604
rect 1794 74898 1826 75454
rect 2382 74898 2414 75454
rect 1794 39454 2414 74898
rect 1794 38898 1826 39454
rect 2382 38898 2414 39454
rect 1794 3454 2414 38898
rect 1794 2898 1826 3454
rect 2382 2898 2414 3454
rect 1794 -346 2414 2898
rect 1794 -902 1826 -346
rect 2382 -902 2414 -346
rect -2966 -1862 -2934 -1306
rect -2378 -1862 -2346 -1306
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 79174 6134 114618
rect 5514 78618 5546 79174
rect 6102 78618 6134 79174
rect 5514 43174 6134 78618
rect 5514 42618 5546 43174
rect 6102 42618 6134 43174
rect 5514 7174 6134 42618
rect 5514 6618 5546 7174
rect 6102 6618 6134 7174
rect -3926 -2822 -3894 -2266
rect -3338 -2822 -3306 -2266
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2822 5546 -2266
rect 6102 -2822 6134 -2266
rect -4886 -3782 -4854 -3226
rect -4298 -3782 -4266 -3226
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694338 9266 694894
rect 9822 694338 9854 694894
rect 9234 658894 9854 694338
rect 9234 658338 9266 658894
rect 9822 658338 9854 658894
rect 9234 622894 9854 658338
rect 9234 622338 9266 622894
rect 9822 622338 9854 622894
rect 9234 586894 9854 622338
rect 9234 586338 9266 586894
rect 9822 586338 9854 586894
rect 9234 550894 9854 586338
rect 9234 550338 9266 550894
rect 9822 550338 9854 550894
rect 9234 514894 9854 550338
rect 9234 514338 9266 514894
rect 9822 514338 9854 514894
rect 9234 478894 9854 514338
rect 9234 478338 9266 478894
rect 9822 478338 9854 478894
rect 9234 442894 9854 478338
rect 9234 442338 9266 442894
rect 9822 442338 9854 442894
rect 9234 406894 9854 442338
rect 9234 406338 9266 406894
rect 9822 406338 9854 406894
rect 9234 370894 9854 406338
rect 9234 370338 9266 370894
rect 9822 370338 9854 370894
rect 9234 334894 9854 370338
rect 9234 334338 9266 334894
rect 9822 334338 9854 334894
rect 9234 298894 9854 334338
rect 9234 298338 9266 298894
rect 9822 298338 9854 298894
rect 9234 262894 9854 298338
rect 9234 262338 9266 262894
rect 9822 262338 9854 262894
rect 9234 226894 9854 262338
rect 9234 226338 9266 226894
rect 9822 226338 9854 226894
rect 9234 190894 9854 226338
rect 9234 190338 9266 190894
rect 9822 190338 9854 190894
rect 9234 154894 9854 190338
rect 9234 154338 9266 154894
rect 9822 154338 9854 154894
rect 9234 118894 9854 154338
rect 9234 118338 9266 118894
rect 9822 118338 9854 118894
rect 9234 82894 9854 118338
rect 9234 82338 9266 82894
rect 9822 82338 9854 82894
rect 9234 46894 9854 82338
rect 9234 46338 9266 46894
rect 9822 46338 9854 46894
rect 9234 10894 9854 46338
rect 9234 10338 9266 10894
rect 9822 10338 9854 10894
rect -5846 -4742 -5814 -4186
rect -5258 -4742 -5226 -4186
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4742 9266 -4186
rect 9822 -4742 9854 -4186
rect -6806 -5702 -6774 -5146
rect -6218 -5702 -6186 -5146
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711002 30986 711558
rect 31542 711002 31574 711558
rect 27234 709638 27854 709670
rect 27234 709082 27266 709638
rect 27822 709082 27854 709638
rect 23514 707718 24134 707750
rect 23514 707162 23546 707718
rect 24102 707162 24134 707718
rect 12954 698058 12986 698614
rect 13542 698058 13574 698614
rect 12954 662614 13574 698058
rect 12954 662058 12986 662614
rect 13542 662058 13574 662614
rect 12954 626614 13574 662058
rect 12954 626058 12986 626614
rect 13542 626058 13574 626614
rect 12954 590614 13574 626058
rect 12954 590058 12986 590614
rect 13542 590058 13574 590614
rect 12954 554614 13574 590058
rect 12954 554058 12986 554614
rect 13542 554058 13574 554614
rect 12954 518614 13574 554058
rect 12954 518058 12986 518614
rect 13542 518058 13574 518614
rect 12954 482614 13574 518058
rect 12954 482058 12986 482614
rect 13542 482058 13574 482614
rect 12954 446614 13574 482058
rect 12954 446058 12986 446614
rect 13542 446058 13574 446614
rect 12954 410614 13574 446058
rect 12954 410058 12986 410614
rect 13542 410058 13574 410614
rect 12954 374614 13574 410058
rect 12954 374058 12986 374614
rect 13542 374058 13574 374614
rect 12954 338614 13574 374058
rect 12954 338058 12986 338614
rect 13542 338058 13574 338614
rect 12954 302614 13574 338058
rect 12954 302058 12986 302614
rect 13542 302058 13574 302614
rect 12954 266614 13574 302058
rect 12954 266058 12986 266614
rect 13542 266058 13574 266614
rect 12954 230614 13574 266058
rect 12954 230058 12986 230614
rect 13542 230058 13574 230614
rect 12954 194614 13574 230058
rect 12954 194058 12986 194614
rect 13542 194058 13574 194614
rect 12954 158614 13574 194058
rect 12954 158058 12986 158614
rect 13542 158058 13574 158614
rect 12954 122614 13574 158058
rect 12954 122058 12986 122614
rect 13542 122058 13574 122614
rect 12954 86614 13574 122058
rect 12954 86058 12986 86614
rect 13542 86058 13574 86614
rect 12954 50614 13574 86058
rect 12954 50058 12986 50614
rect 13542 50058 13574 50614
rect 12954 14614 13574 50058
rect 12954 14058 12986 14614
rect 13542 14058 13574 14614
rect -7766 -6662 -7734 -6106
rect -7178 -6662 -7146 -6106
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705242 19826 705798
rect 20382 705242 20414 705798
rect 19794 669454 20414 705242
rect 19794 668898 19826 669454
rect 20382 668898 20414 669454
rect 19794 633454 20414 668898
rect 19794 632898 19826 633454
rect 20382 632898 20414 633454
rect 19794 597454 20414 632898
rect 19794 596898 19826 597454
rect 20382 596898 20414 597454
rect 19794 561454 20414 596898
rect 19794 560898 19826 561454
rect 20382 560898 20414 561454
rect 19794 525454 20414 560898
rect 19794 524898 19826 525454
rect 20382 524898 20414 525454
rect 19794 489454 20414 524898
rect 19794 488898 19826 489454
rect 20382 488898 20414 489454
rect 19794 453454 20414 488898
rect 19794 452898 19826 453454
rect 20382 452898 20414 453454
rect 19794 417454 20414 452898
rect 19794 416898 19826 417454
rect 20382 416898 20414 417454
rect 19794 381454 20414 416898
rect 19794 380898 19826 381454
rect 20382 380898 20414 381454
rect 19794 345454 20414 380898
rect 19794 344898 19826 345454
rect 20382 344898 20414 345454
rect 19794 309454 20414 344898
rect 19794 308898 19826 309454
rect 20382 308898 20414 309454
rect 19794 273454 20414 308898
rect 19794 272898 19826 273454
rect 20382 272898 20414 273454
rect 19794 237454 20414 272898
rect 19794 236898 19826 237454
rect 20382 236898 20414 237454
rect 19794 201454 20414 236898
rect 19794 200898 19826 201454
rect 20382 200898 20414 201454
rect 19794 165454 20414 200898
rect 19794 164898 19826 165454
rect 20382 164898 20414 165454
rect 19794 129454 20414 164898
rect 19794 128898 19826 129454
rect 20382 128898 20414 129454
rect 19794 93454 20414 128898
rect 19794 92898 19826 93454
rect 20382 92898 20414 93454
rect 19794 57454 20414 92898
rect 19794 56898 19826 57454
rect 20382 56898 20414 57454
rect 19794 21454 20414 56898
rect 19794 20898 19826 21454
rect 20382 20898 20414 21454
rect 19794 -1306 20414 20898
rect 19794 -1862 19826 -1306
rect 20382 -1862 20414 -1306
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672618 23546 673174
rect 24102 672618 24134 673174
rect 23514 637174 24134 672618
rect 23514 636618 23546 637174
rect 24102 636618 24134 637174
rect 23514 601174 24134 636618
rect 23514 600618 23546 601174
rect 24102 600618 24134 601174
rect 23514 565174 24134 600618
rect 23514 564618 23546 565174
rect 24102 564618 24134 565174
rect 23514 529174 24134 564618
rect 23514 528618 23546 529174
rect 24102 528618 24134 529174
rect 23514 493174 24134 528618
rect 23514 492618 23546 493174
rect 24102 492618 24134 493174
rect 23514 457174 24134 492618
rect 23514 456618 23546 457174
rect 24102 456618 24134 457174
rect 23514 421174 24134 456618
rect 23514 420618 23546 421174
rect 24102 420618 24134 421174
rect 23514 385174 24134 420618
rect 23514 384618 23546 385174
rect 24102 384618 24134 385174
rect 23514 349174 24134 384618
rect 23514 348618 23546 349174
rect 24102 348618 24134 349174
rect 23514 313174 24134 348618
rect 23514 312618 23546 313174
rect 24102 312618 24134 313174
rect 23514 277174 24134 312618
rect 23514 276618 23546 277174
rect 24102 276618 24134 277174
rect 23514 241174 24134 276618
rect 23514 240618 23546 241174
rect 24102 240618 24134 241174
rect 23514 205174 24134 240618
rect 23514 204618 23546 205174
rect 24102 204618 24134 205174
rect 23514 169174 24134 204618
rect 23514 168618 23546 169174
rect 24102 168618 24134 169174
rect 23514 133174 24134 168618
rect 23514 132618 23546 133174
rect 24102 132618 24134 133174
rect 23514 97174 24134 132618
rect 23514 96618 23546 97174
rect 24102 96618 24134 97174
rect 23514 61174 24134 96618
rect 23514 60618 23546 61174
rect 24102 60618 24134 61174
rect 23514 25174 24134 60618
rect 23514 24618 23546 25174
rect 24102 24618 24134 25174
rect 23514 -3226 24134 24618
rect 23514 -3782 23546 -3226
rect 24102 -3782 24134 -3226
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676338 27266 676894
rect 27822 676338 27854 676894
rect 27234 640894 27854 676338
rect 27234 640338 27266 640894
rect 27822 640338 27854 640894
rect 27234 604894 27854 640338
rect 27234 604338 27266 604894
rect 27822 604338 27854 604894
rect 27234 568894 27854 604338
rect 27234 568338 27266 568894
rect 27822 568338 27854 568894
rect 27234 532894 27854 568338
rect 27234 532338 27266 532894
rect 27822 532338 27854 532894
rect 27234 496894 27854 532338
rect 27234 496338 27266 496894
rect 27822 496338 27854 496894
rect 27234 460894 27854 496338
rect 27234 460338 27266 460894
rect 27822 460338 27854 460894
rect 27234 424894 27854 460338
rect 27234 424338 27266 424894
rect 27822 424338 27854 424894
rect 27234 388894 27854 424338
rect 27234 388338 27266 388894
rect 27822 388338 27854 388894
rect 27234 352894 27854 388338
rect 27234 352338 27266 352894
rect 27822 352338 27854 352894
rect 27234 316894 27854 352338
rect 27234 316338 27266 316894
rect 27822 316338 27854 316894
rect 27234 280894 27854 316338
rect 27234 280338 27266 280894
rect 27822 280338 27854 280894
rect 27234 244894 27854 280338
rect 27234 244338 27266 244894
rect 27822 244338 27854 244894
rect 27234 208894 27854 244338
rect 27234 208338 27266 208894
rect 27822 208338 27854 208894
rect 27234 172894 27854 208338
rect 27234 172338 27266 172894
rect 27822 172338 27854 172894
rect 27234 136894 27854 172338
rect 27234 136338 27266 136894
rect 27822 136338 27854 136894
rect 27234 100894 27854 136338
rect 27234 100338 27266 100894
rect 27822 100338 27854 100894
rect 27234 64894 27854 100338
rect 27234 64338 27266 64894
rect 27822 64338 27854 64894
rect 27234 28894 27854 64338
rect 27234 28338 27266 28894
rect 27822 28338 27854 28894
rect 27234 -5146 27854 28338
rect 27234 -5702 27266 -5146
rect 27822 -5702 27854 -5146
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710042 48986 710598
rect 49542 710042 49574 710598
rect 45234 708678 45854 709670
rect 45234 708122 45266 708678
rect 45822 708122 45854 708678
rect 41514 706758 42134 707750
rect 41514 706202 41546 706758
rect 42102 706202 42134 706758
rect 30954 680058 30986 680614
rect 31542 680058 31574 680614
rect 30954 644614 31574 680058
rect 30954 644058 30986 644614
rect 31542 644058 31574 644614
rect 30954 608614 31574 644058
rect 30954 608058 30986 608614
rect 31542 608058 31574 608614
rect 30954 572614 31574 608058
rect 30954 572058 30986 572614
rect 31542 572058 31574 572614
rect 30954 536614 31574 572058
rect 30954 536058 30986 536614
rect 31542 536058 31574 536614
rect 30954 500614 31574 536058
rect 30954 500058 30986 500614
rect 31542 500058 31574 500614
rect 30954 464614 31574 500058
rect 30954 464058 30986 464614
rect 31542 464058 31574 464614
rect 30954 428614 31574 464058
rect 30954 428058 30986 428614
rect 31542 428058 31574 428614
rect 30954 392614 31574 428058
rect 30954 392058 30986 392614
rect 31542 392058 31574 392614
rect 30954 356614 31574 392058
rect 30954 356058 30986 356614
rect 31542 356058 31574 356614
rect 30954 320614 31574 356058
rect 30954 320058 30986 320614
rect 31542 320058 31574 320614
rect 30954 284614 31574 320058
rect 30954 284058 30986 284614
rect 31542 284058 31574 284614
rect 30954 248614 31574 284058
rect 30954 248058 30986 248614
rect 31542 248058 31574 248614
rect 30954 212614 31574 248058
rect 30954 212058 30986 212614
rect 31542 212058 31574 212614
rect 30954 176614 31574 212058
rect 30954 176058 30986 176614
rect 31542 176058 31574 176614
rect 30954 140614 31574 176058
rect 30954 140058 30986 140614
rect 31542 140058 31574 140614
rect 30954 104614 31574 140058
rect 30954 104058 30986 104614
rect 31542 104058 31574 104614
rect 30954 68614 31574 104058
rect 30954 68058 30986 68614
rect 31542 68058 31574 68614
rect 30954 32614 31574 68058
rect 30954 32058 30986 32614
rect 31542 32058 31574 32614
rect 12954 -6662 12986 -6106
rect 13542 -6662 13574 -6106
rect -8726 -7622 -8694 -7066
rect -8138 -7622 -8106 -7066
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704282 37826 704838
rect 38382 704282 38414 704838
rect 37794 687454 38414 704282
rect 37794 686898 37826 687454
rect 38382 686898 38414 687454
rect 37794 651454 38414 686898
rect 37794 650898 37826 651454
rect 38382 650898 38414 651454
rect 37794 615454 38414 650898
rect 37794 614898 37826 615454
rect 38382 614898 38414 615454
rect 37794 579454 38414 614898
rect 37794 578898 37826 579454
rect 38382 578898 38414 579454
rect 37794 543454 38414 578898
rect 37794 542898 37826 543454
rect 38382 542898 38414 543454
rect 37794 507454 38414 542898
rect 37794 506898 37826 507454
rect 38382 506898 38414 507454
rect 37794 471454 38414 506898
rect 37794 470898 37826 471454
rect 38382 470898 38414 471454
rect 37794 435454 38414 470898
rect 37794 434898 37826 435454
rect 38382 434898 38414 435454
rect 37794 399454 38414 434898
rect 37794 398898 37826 399454
rect 38382 398898 38414 399454
rect 37794 363454 38414 398898
rect 37794 362898 37826 363454
rect 38382 362898 38414 363454
rect 37794 327454 38414 362898
rect 37794 326898 37826 327454
rect 38382 326898 38414 327454
rect 37794 291454 38414 326898
rect 37794 290898 37826 291454
rect 38382 290898 38414 291454
rect 37794 255454 38414 290898
rect 37794 254898 37826 255454
rect 38382 254898 38414 255454
rect 37794 219454 38414 254898
rect 37794 218898 37826 219454
rect 38382 218898 38414 219454
rect 37794 183454 38414 218898
rect 37794 182898 37826 183454
rect 38382 182898 38414 183454
rect 37794 147454 38414 182898
rect 37794 146898 37826 147454
rect 38382 146898 38414 147454
rect 37794 111454 38414 146898
rect 37794 110898 37826 111454
rect 38382 110898 38414 111454
rect 37794 75454 38414 110898
rect 37794 74898 37826 75454
rect 38382 74898 38414 75454
rect 37794 39454 38414 74898
rect 37794 38898 37826 39454
rect 38382 38898 38414 39454
rect 37794 3454 38414 38898
rect 37794 2898 37826 3454
rect 38382 2898 38414 3454
rect 37794 -346 38414 2898
rect 37794 -902 37826 -346
rect 38382 -902 38414 -346
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690618 41546 691174
rect 42102 690618 42134 691174
rect 41514 655174 42134 690618
rect 41514 654618 41546 655174
rect 42102 654618 42134 655174
rect 41514 619174 42134 654618
rect 41514 618618 41546 619174
rect 42102 618618 42134 619174
rect 41514 583174 42134 618618
rect 41514 582618 41546 583174
rect 42102 582618 42134 583174
rect 41514 547174 42134 582618
rect 41514 546618 41546 547174
rect 42102 546618 42134 547174
rect 41514 511174 42134 546618
rect 41514 510618 41546 511174
rect 42102 510618 42134 511174
rect 41514 475174 42134 510618
rect 41514 474618 41546 475174
rect 42102 474618 42134 475174
rect 41514 439174 42134 474618
rect 41514 438618 41546 439174
rect 42102 438618 42134 439174
rect 41514 403174 42134 438618
rect 41514 402618 41546 403174
rect 42102 402618 42134 403174
rect 41514 367174 42134 402618
rect 41514 366618 41546 367174
rect 42102 366618 42134 367174
rect 41514 331174 42134 366618
rect 41514 330618 41546 331174
rect 42102 330618 42134 331174
rect 41514 295174 42134 330618
rect 41514 294618 41546 295174
rect 42102 294618 42134 295174
rect 41514 259174 42134 294618
rect 41514 258618 41546 259174
rect 42102 258618 42134 259174
rect 41514 223174 42134 258618
rect 41514 222618 41546 223174
rect 42102 222618 42134 223174
rect 41514 187174 42134 222618
rect 41514 186618 41546 187174
rect 42102 186618 42134 187174
rect 41514 151174 42134 186618
rect 41514 150618 41546 151174
rect 42102 150618 42134 151174
rect 41514 115174 42134 150618
rect 41514 114618 41546 115174
rect 42102 114618 42134 115174
rect 41514 79174 42134 114618
rect 41514 78618 41546 79174
rect 42102 78618 42134 79174
rect 41514 43174 42134 78618
rect 41514 42618 41546 43174
rect 42102 42618 42134 43174
rect 41514 7174 42134 42618
rect 41514 6618 41546 7174
rect 42102 6618 42134 7174
rect 41514 -2266 42134 6618
rect 41514 -2822 41546 -2266
rect 42102 -2822 42134 -2266
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694338 45266 694894
rect 45822 694338 45854 694894
rect 45234 658894 45854 694338
rect 45234 658338 45266 658894
rect 45822 658338 45854 658894
rect 45234 622894 45854 658338
rect 45234 622338 45266 622894
rect 45822 622338 45854 622894
rect 45234 586894 45854 622338
rect 45234 586338 45266 586894
rect 45822 586338 45854 586894
rect 45234 550894 45854 586338
rect 45234 550338 45266 550894
rect 45822 550338 45854 550894
rect 45234 514894 45854 550338
rect 45234 514338 45266 514894
rect 45822 514338 45854 514894
rect 45234 478894 45854 514338
rect 45234 478338 45266 478894
rect 45822 478338 45854 478894
rect 45234 442894 45854 478338
rect 45234 442338 45266 442894
rect 45822 442338 45854 442894
rect 45234 406894 45854 442338
rect 45234 406338 45266 406894
rect 45822 406338 45854 406894
rect 45234 370894 45854 406338
rect 45234 370338 45266 370894
rect 45822 370338 45854 370894
rect 45234 334894 45854 370338
rect 45234 334338 45266 334894
rect 45822 334338 45854 334894
rect 45234 298894 45854 334338
rect 45234 298338 45266 298894
rect 45822 298338 45854 298894
rect 45234 262894 45854 298338
rect 45234 262338 45266 262894
rect 45822 262338 45854 262894
rect 45234 226894 45854 262338
rect 45234 226338 45266 226894
rect 45822 226338 45854 226894
rect 45234 190894 45854 226338
rect 45234 190338 45266 190894
rect 45822 190338 45854 190894
rect 45234 154894 45854 190338
rect 45234 154338 45266 154894
rect 45822 154338 45854 154894
rect 45234 118894 45854 154338
rect 45234 118338 45266 118894
rect 45822 118338 45854 118894
rect 45234 82894 45854 118338
rect 45234 82338 45266 82894
rect 45822 82338 45854 82894
rect 45234 46894 45854 82338
rect 45234 46338 45266 46894
rect 45822 46338 45854 46894
rect 45234 10894 45854 46338
rect 45234 10338 45266 10894
rect 45822 10338 45854 10894
rect 45234 -4186 45854 10338
rect 45234 -4742 45266 -4186
rect 45822 -4742 45854 -4186
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711002 66986 711558
rect 67542 711002 67574 711558
rect 63234 709638 63854 709670
rect 63234 709082 63266 709638
rect 63822 709082 63854 709638
rect 59514 707718 60134 707750
rect 59514 707162 59546 707718
rect 60102 707162 60134 707718
rect 48954 698058 48986 698614
rect 49542 698058 49574 698614
rect 48954 662614 49574 698058
rect 48954 662058 48986 662614
rect 49542 662058 49574 662614
rect 48954 626614 49574 662058
rect 48954 626058 48986 626614
rect 49542 626058 49574 626614
rect 48954 590614 49574 626058
rect 48954 590058 48986 590614
rect 49542 590058 49574 590614
rect 48954 554614 49574 590058
rect 48954 554058 48986 554614
rect 49542 554058 49574 554614
rect 48954 518614 49574 554058
rect 48954 518058 48986 518614
rect 49542 518058 49574 518614
rect 48954 482614 49574 518058
rect 48954 482058 48986 482614
rect 49542 482058 49574 482614
rect 48954 446614 49574 482058
rect 48954 446058 48986 446614
rect 49542 446058 49574 446614
rect 48954 410614 49574 446058
rect 48954 410058 48986 410614
rect 49542 410058 49574 410614
rect 48954 374614 49574 410058
rect 48954 374058 48986 374614
rect 49542 374058 49574 374614
rect 48954 338614 49574 374058
rect 48954 338058 48986 338614
rect 49542 338058 49574 338614
rect 48954 302614 49574 338058
rect 48954 302058 48986 302614
rect 49542 302058 49574 302614
rect 48954 266614 49574 302058
rect 48954 266058 48986 266614
rect 49542 266058 49574 266614
rect 48954 230614 49574 266058
rect 48954 230058 48986 230614
rect 49542 230058 49574 230614
rect 48954 194614 49574 230058
rect 48954 194058 48986 194614
rect 49542 194058 49574 194614
rect 48954 158614 49574 194058
rect 48954 158058 48986 158614
rect 49542 158058 49574 158614
rect 48954 122614 49574 158058
rect 48954 122058 48986 122614
rect 49542 122058 49574 122614
rect 48954 86614 49574 122058
rect 48954 86058 48986 86614
rect 49542 86058 49574 86614
rect 48954 50614 49574 86058
rect 48954 50058 48986 50614
rect 49542 50058 49574 50614
rect 48954 14614 49574 50058
rect 48954 14058 48986 14614
rect 49542 14058 49574 14614
rect 30954 -7622 30986 -7066
rect 31542 -7622 31574 -7066
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705242 55826 705798
rect 56382 705242 56414 705798
rect 55794 669454 56414 705242
rect 55794 668898 55826 669454
rect 56382 668898 56414 669454
rect 55794 633454 56414 668898
rect 55794 632898 55826 633454
rect 56382 632898 56414 633454
rect 55794 597454 56414 632898
rect 55794 596898 55826 597454
rect 56382 596898 56414 597454
rect 55794 561454 56414 596898
rect 55794 560898 55826 561454
rect 56382 560898 56414 561454
rect 55794 525454 56414 560898
rect 55794 524898 55826 525454
rect 56382 524898 56414 525454
rect 55794 489454 56414 524898
rect 55794 488898 55826 489454
rect 56382 488898 56414 489454
rect 55794 453454 56414 488898
rect 55794 452898 55826 453454
rect 56382 452898 56414 453454
rect 55794 417454 56414 452898
rect 55794 416898 55826 417454
rect 56382 416898 56414 417454
rect 55794 381454 56414 416898
rect 55794 380898 55826 381454
rect 56382 380898 56414 381454
rect 55794 345454 56414 380898
rect 55794 344898 55826 345454
rect 56382 344898 56414 345454
rect 55794 309454 56414 344898
rect 55794 308898 55826 309454
rect 56382 308898 56414 309454
rect 55794 273454 56414 308898
rect 55794 272898 55826 273454
rect 56382 272898 56414 273454
rect 55794 237454 56414 272898
rect 55794 236898 55826 237454
rect 56382 236898 56414 237454
rect 55794 201454 56414 236898
rect 55794 200898 55826 201454
rect 56382 200898 56414 201454
rect 55794 165454 56414 200898
rect 55794 164898 55826 165454
rect 56382 164898 56414 165454
rect 55794 129454 56414 164898
rect 55794 128898 55826 129454
rect 56382 128898 56414 129454
rect 55794 93454 56414 128898
rect 55794 92898 55826 93454
rect 56382 92898 56414 93454
rect 55794 57454 56414 92898
rect 55794 56898 55826 57454
rect 56382 56898 56414 57454
rect 55794 21454 56414 56898
rect 55794 20898 55826 21454
rect 56382 20898 56414 21454
rect 55794 -1306 56414 20898
rect 55794 -1862 55826 -1306
rect 56382 -1862 56414 -1306
rect 55794 -1894 56414 -1862
rect 59514 673174 60134 707162
rect 59514 672618 59546 673174
rect 60102 672618 60134 673174
rect 59514 637174 60134 672618
rect 59514 636618 59546 637174
rect 60102 636618 60134 637174
rect 59514 601174 60134 636618
rect 59514 600618 59546 601174
rect 60102 600618 60134 601174
rect 59514 565174 60134 600618
rect 59514 564618 59546 565174
rect 60102 564618 60134 565174
rect 59514 529174 60134 564618
rect 59514 528618 59546 529174
rect 60102 528618 60134 529174
rect 59514 493174 60134 528618
rect 59514 492618 59546 493174
rect 60102 492618 60134 493174
rect 59514 457174 60134 492618
rect 59514 456618 59546 457174
rect 60102 456618 60134 457174
rect 59514 421174 60134 456618
rect 59514 420618 59546 421174
rect 60102 420618 60134 421174
rect 59514 385174 60134 420618
rect 59514 384618 59546 385174
rect 60102 384618 60134 385174
rect 59514 349174 60134 384618
rect 59514 348618 59546 349174
rect 60102 348618 60134 349174
rect 59514 313174 60134 348618
rect 59514 312618 59546 313174
rect 60102 312618 60134 313174
rect 59514 277174 60134 312618
rect 59514 276618 59546 277174
rect 60102 276618 60134 277174
rect 59514 241174 60134 276618
rect 59514 240618 59546 241174
rect 60102 240618 60134 241174
rect 59514 205174 60134 240618
rect 59514 204618 59546 205174
rect 60102 204618 60134 205174
rect 59514 169174 60134 204618
rect 59514 168618 59546 169174
rect 60102 168618 60134 169174
rect 59514 133174 60134 168618
rect 59514 132618 59546 133174
rect 60102 132618 60134 133174
rect 59514 97174 60134 132618
rect 59514 96618 59546 97174
rect 60102 96618 60134 97174
rect 59514 61174 60134 96618
rect 59514 60618 59546 61174
rect 60102 60618 60134 61174
rect 59514 25174 60134 60618
rect 59514 24618 59546 25174
rect 60102 24618 60134 25174
rect 59514 -3226 60134 24618
rect 59514 -3782 59546 -3226
rect 60102 -3782 60134 -3226
rect 59514 -3814 60134 -3782
rect 63234 676894 63854 709082
rect 63234 676338 63266 676894
rect 63822 676338 63854 676894
rect 63234 640894 63854 676338
rect 63234 640338 63266 640894
rect 63822 640338 63854 640894
rect 63234 604894 63854 640338
rect 63234 604338 63266 604894
rect 63822 604338 63854 604894
rect 63234 568894 63854 604338
rect 63234 568338 63266 568894
rect 63822 568338 63854 568894
rect 63234 532894 63854 568338
rect 63234 532338 63266 532894
rect 63822 532338 63854 532894
rect 63234 496894 63854 532338
rect 63234 496338 63266 496894
rect 63822 496338 63854 496894
rect 63234 460894 63854 496338
rect 63234 460338 63266 460894
rect 63822 460338 63854 460894
rect 63234 424894 63854 460338
rect 63234 424338 63266 424894
rect 63822 424338 63854 424894
rect 63234 388894 63854 424338
rect 63234 388338 63266 388894
rect 63822 388338 63854 388894
rect 63234 352894 63854 388338
rect 63234 352338 63266 352894
rect 63822 352338 63854 352894
rect 63234 316894 63854 352338
rect 63234 316338 63266 316894
rect 63822 316338 63854 316894
rect 63234 280894 63854 316338
rect 63234 280338 63266 280894
rect 63822 280338 63854 280894
rect 63234 244894 63854 280338
rect 63234 244338 63266 244894
rect 63822 244338 63854 244894
rect 63234 208894 63854 244338
rect 63234 208338 63266 208894
rect 63822 208338 63854 208894
rect 63234 172894 63854 208338
rect 63234 172338 63266 172894
rect 63822 172338 63854 172894
rect 63234 136894 63854 172338
rect 63234 136338 63266 136894
rect 63822 136338 63854 136894
rect 63234 100894 63854 136338
rect 63234 100338 63266 100894
rect 63822 100338 63854 100894
rect 63234 64894 63854 100338
rect 63234 64338 63266 64894
rect 63822 64338 63854 64894
rect 63234 28894 63854 64338
rect 63234 28338 63266 28894
rect 63822 28338 63854 28894
rect 63234 -5146 63854 28338
rect 63234 -5702 63266 -5146
rect 63822 -5702 63854 -5146
rect 63234 -5734 63854 -5702
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710042 84986 710598
rect 85542 710042 85574 710598
rect 81234 708678 81854 709670
rect 81234 708122 81266 708678
rect 81822 708122 81854 708678
rect 77514 706758 78134 707750
rect 77514 706202 77546 706758
rect 78102 706202 78134 706758
rect 66954 680058 66986 680614
rect 67542 680058 67574 680614
rect 66954 644614 67574 680058
rect 66954 644058 66986 644614
rect 67542 644058 67574 644614
rect 66954 608614 67574 644058
rect 66954 608058 66986 608614
rect 67542 608058 67574 608614
rect 66954 572614 67574 608058
rect 66954 572058 66986 572614
rect 67542 572058 67574 572614
rect 66954 536614 67574 572058
rect 66954 536058 66986 536614
rect 67542 536058 67574 536614
rect 66954 500614 67574 536058
rect 66954 500058 66986 500614
rect 67542 500058 67574 500614
rect 66954 464614 67574 500058
rect 66954 464058 66986 464614
rect 67542 464058 67574 464614
rect 66954 428614 67574 464058
rect 66954 428058 66986 428614
rect 67542 428058 67574 428614
rect 66954 392614 67574 428058
rect 66954 392058 66986 392614
rect 67542 392058 67574 392614
rect 66954 356614 67574 392058
rect 66954 356058 66986 356614
rect 67542 356058 67574 356614
rect 66954 320614 67574 356058
rect 66954 320058 66986 320614
rect 67542 320058 67574 320614
rect 66954 284614 67574 320058
rect 66954 284058 66986 284614
rect 67542 284058 67574 284614
rect 66954 248614 67574 284058
rect 66954 248058 66986 248614
rect 67542 248058 67574 248614
rect 66954 212614 67574 248058
rect 66954 212058 66986 212614
rect 67542 212058 67574 212614
rect 66954 176614 67574 212058
rect 66954 176058 66986 176614
rect 67542 176058 67574 176614
rect 66954 140614 67574 176058
rect 66954 140058 66986 140614
rect 67542 140058 67574 140614
rect 66954 104614 67574 140058
rect 66954 104058 66986 104614
rect 67542 104058 67574 104614
rect 66954 68614 67574 104058
rect 66954 68058 66986 68614
rect 67542 68058 67574 68614
rect 66954 32614 67574 68058
rect 66954 32058 66986 32614
rect 67542 32058 67574 32614
rect 48954 -6662 48986 -6106
rect 49542 -6662 49574 -6106
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 704838 74414 705830
rect 73794 704282 73826 704838
rect 74382 704282 74414 704838
rect 73794 687454 74414 704282
rect 73794 686898 73826 687454
rect 74382 686898 74414 687454
rect 73794 651454 74414 686898
rect 73794 650898 73826 651454
rect 74382 650898 74414 651454
rect 73794 615454 74414 650898
rect 73794 614898 73826 615454
rect 74382 614898 74414 615454
rect 73794 579454 74414 614898
rect 73794 578898 73826 579454
rect 74382 578898 74414 579454
rect 73794 543454 74414 578898
rect 73794 542898 73826 543454
rect 74382 542898 74414 543454
rect 73794 507454 74414 542898
rect 73794 506898 73826 507454
rect 74382 506898 74414 507454
rect 73794 471454 74414 506898
rect 73794 470898 73826 471454
rect 74382 470898 74414 471454
rect 73794 435454 74414 470898
rect 73794 434898 73826 435454
rect 74382 434898 74414 435454
rect 73794 399454 74414 434898
rect 73794 398898 73826 399454
rect 74382 398898 74414 399454
rect 73794 363454 74414 398898
rect 73794 362898 73826 363454
rect 74382 362898 74414 363454
rect 73794 327454 74414 362898
rect 73794 326898 73826 327454
rect 74382 326898 74414 327454
rect 73794 291454 74414 326898
rect 73794 290898 73826 291454
rect 74382 290898 74414 291454
rect 73794 255454 74414 290898
rect 73794 254898 73826 255454
rect 74382 254898 74414 255454
rect 73794 219454 74414 254898
rect 73794 218898 73826 219454
rect 74382 218898 74414 219454
rect 73794 183454 74414 218898
rect 73794 182898 73826 183454
rect 74382 182898 74414 183454
rect 73794 147454 74414 182898
rect 73794 146898 73826 147454
rect 74382 146898 74414 147454
rect 73794 111454 74414 146898
rect 73794 110898 73826 111454
rect 74382 110898 74414 111454
rect 73794 75454 74414 110898
rect 73794 74898 73826 75454
rect 74382 74898 74414 75454
rect 73794 39454 74414 74898
rect 73794 38898 73826 39454
rect 74382 38898 74414 39454
rect 73794 3454 74414 38898
rect 73794 2898 73826 3454
rect 74382 2898 74414 3454
rect 73794 -346 74414 2898
rect 73794 -902 73826 -346
rect 74382 -902 74414 -346
rect 73794 -1894 74414 -902
rect 77514 691174 78134 706202
rect 77514 690618 77546 691174
rect 78102 690618 78134 691174
rect 77514 655174 78134 690618
rect 77514 654618 77546 655174
rect 78102 654618 78134 655174
rect 77514 619174 78134 654618
rect 77514 618618 77546 619174
rect 78102 618618 78134 619174
rect 77514 583174 78134 618618
rect 77514 582618 77546 583174
rect 78102 582618 78134 583174
rect 77514 547174 78134 582618
rect 77514 546618 77546 547174
rect 78102 546618 78134 547174
rect 77514 511174 78134 546618
rect 77514 510618 77546 511174
rect 78102 510618 78134 511174
rect 77514 475174 78134 510618
rect 77514 474618 77546 475174
rect 78102 474618 78134 475174
rect 77514 439174 78134 474618
rect 77514 438618 77546 439174
rect 78102 438618 78134 439174
rect 77514 403174 78134 438618
rect 77514 402618 77546 403174
rect 78102 402618 78134 403174
rect 77514 367174 78134 402618
rect 77514 366618 77546 367174
rect 78102 366618 78134 367174
rect 77514 331174 78134 366618
rect 77514 330618 77546 331174
rect 78102 330618 78134 331174
rect 77514 295174 78134 330618
rect 77514 294618 77546 295174
rect 78102 294618 78134 295174
rect 77514 259174 78134 294618
rect 77514 258618 77546 259174
rect 78102 258618 78134 259174
rect 77514 223174 78134 258618
rect 77514 222618 77546 223174
rect 78102 222618 78134 223174
rect 77514 187174 78134 222618
rect 77514 186618 77546 187174
rect 78102 186618 78134 187174
rect 77514 151174 78134 186618
rect 77514 150618 77546 151174
rect 78102 150618 78134 151174
rect 77514 115174 78134 150618
rect 77514 114618 77546 115174
rect 78102 114618 78134 115174
rect 77514 79174 78134 114618
rect 77514 78618 77546 79174
rect 78102 78618 78134 79174
rect 77514 43174 78134 78618
rect 77514 42618 77546 43174
rect 78102 42618 78134 43174
rect 77514 7174 78134 42618
rect 77514 6618 77546 7174
rect 78102 6618 78134 7174
rect 77514 -2266 78134 6618
rect 77514 -2822 77546 -2266
rect 78102 -2822 78134 -2266
rect 77514 -3814 78134 -2822
rect 81234 694894 81854 708122
rect 81234 694338 81266 694894
rect 81822 694338 81854 694894
rect 81234 658894 81854 694338
rect 81234 658338 81266 658894
rect 81822 658338 81854 658894
rect 81234 622894 81854 658338
rect 81234 622338 81266 622894
rect 81822 622338 81854 622894
rect 81234 586894 81854 622338
rect 81234 586338 81266 586894
rect 81822 586338 81854 586894
rect 81234 550894 81854 586338
rect 81234 550338 81266 550894
rect 81822 550338 81854 550894
rect 81234 514894 81854 550338
rect 81234 514338 81266 514894
rect 81822 514338 81854 514894
rect 81234 478894 81854 514338
rect 81234 478338 81266 478894
rect 81822 478338 81854 478894
rect 81234 442894 81854 478338
rect 81234 442338 81266 442894
rect 81822 442338 81854 442894
rect 81234 406894 81854 442338
rect 81234 406338 81266 406894
rect 81822 406338 81854 406894
rect 81234 370894 81854 406338
rect 81234 370338 81266 370894
rect 81822 370338 81854 370894
rect 81234 334894 81854 370338
rect 81234 334338 81266 334894
rect 81822 334338 81854 334894
rect 81234 298894 81854 334338
rect 81234 298338 81266 298894
rect 81822 298338 81854 298894
rect 81234 262894 81854 298338
rect 81234 262338 81266 262894
rect 81822 262338 81854 262894
rect 81234 226894 81854 262338
rect 81234 226338 81266 226894
rect 81822 226338 81854 226894
rect 81234 190894 81854 226338
rect 81234 190338 81266 190894
rect 81822 190338 81854 190894
rect 81234 154894 81854 190338
rect 81234 154338 81266 154894
rect 81822 154338 81854 154894
rect 81234 118894 81854 154338
rect 81234 118338 81266 118894
rect 81822 118338 81854 118894
rect 81234 82894 81854 118338
rect 81234 82338 81266 82894
rect 81822 82338 81854 82894
rect 81234 46894 81854 82338
rect 81234 46338 81266 46894
rect 81822 46338 81854 46894
rect 81234 10894 81854 46338
rect 81234 10338 81266 10894
rect 81822 10338 81854 10894
rect 81234 -4186 81854 10338
rect 81234 -4742 81266 -4186
rect 81822 -4742 81854 -4186
rect 81234 -5734 81854 -4742
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711002 102986 711558
rect 103542 711002 103574 711558
rect 99234 709638 99854 709670
rect 99234 709082 99266 709638
rect 99822 709082 99854 709638
rect 95514 707718 96134 707750
rect 95514 707162 95546 707718
rect 96102 707162 96134 707718
rect 84954 698058 84986 698614
rect 85542 698058 85574 698614
rect 84954 662614 85574 698058
rect 84954 662058 84986 662614
rect 85542 662058 85574 662614
rect 84954 626614 85574 662058
rect 84954 626058 84986 626614
rect 85542 626058 85574 626614
rect 84954 590614 85574 626058
rect 84954 590058 84986 590614
rect 85542 590058 85574 590614
rect 84954 554614 85574 590058
rect 84954 554058 84986 554614
rect 85542 554058 85574 554614
rect 84954 518614 85574 554058
rect 84954 518058 84986 518614
rect 85542 518058 85574 518614
rect 84954 482614 85574 518058
rect 84954 482058 84986 482614
rect 85542 482058 85574 482614
rect 84954 446614 85574 482058
rect 84954 446058 84986 446614
rect 85542 446058 85574 446614
rect 84954 410614 85574 446058
rect 84954 410058 84986 410614
rect 85542 410058 85574 410614
rect 84954 374614 85574 410058
rect 84954 374058 84986 374614
rect 85542 374058 85574 374614
rect 84954 338614 85574 374058
rect 84954 338058 84986 338614
rect 85542 338058 85574 338614
rect 84954 302614 85574 338058
rect 84954 302058 84986 302614
rect 85542 302058 85574 302614
rect 84954 266614 85574 302058
rect 84954 266058 84986 266614
rect 85542 266058 85574 266614
rect 84954 230614 85574 266058
rect 84954 230058 84986 230614
rect 85542 230058 85574 230614
rect 84954 194614 85574 230058
rect 84954 194058 84986 194614
rect 85542 194058 85574 194614
rect 84954 158614 85574 194058
rect 84954 158058 84986 158614
rect 85542 158058 85574 158614
rect 84954 122614 85574 158058
rect 84954 122058 84986 122614
rect 85542 122058 85574 122614
rect 84954 86614 85574 122058
rect 84954 86058 84986 86614
rect 85542 86058 85574 86614
rect 84954 50614 85574 86058
rect 84954 50058 84986 50614
rect 85542 50058 85574 50614
rect 84954 14614 85574 50058
rect 84954 14058 84986 14614
rect 85542 14058 85574 14614
rect 66954 -7622 66986 -7066
rect 67542 -7622 67574 -7066
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 705798 92414 705830
rect 91794 705242 91826 705798
rect 92382 705242 92414 705798
rect 91794 669454 92414 705242
rect 91794 668898 91826 669454
rect 92382 668898 92414 669454
rect 91794 633454 92414 668898
rect 91794 632898 91826 633454
rect 92382 632898 92414 633454
rect 91794 597454 92414 632898
rect 91794 596898 91826 597454
rect 92382 596898 92414 597454
rect 91794 561454 92414 596898
rect 91794 560898 91826 561454
rect 92382 560898 92414 561454
rect 91794 525454 92414 560898
rect 91794 524898 91826 525454
rect 92382 524898 92414 525454
rect 91794 489454 92414 524898
rect 91794 488898 91826 489454
rect 92382 488898 92414 489454
rect 91794 453454 92414 488898
rect 91794 452898 91826 453454
rect 92382 452898 92414 453454
rect 91794 417454 92414 452898
rect 91794 416898 91826 417454
rect 92382 416898 92414 417454
rect 91794 381454 92414 416898
rect 91794 380898 91826 381454
rect 92382 380898 92414 381454
rect 91794 345454 92414 380898
rect 91794 344898 91826 345454
rect 92382 344898 92414 345454
rect 91794 309454 92414 344898
rect 91794 308898 91826 309454
rect 92382 308898 92414 309454
rect 91794 273454 92414 308898
rect 91794 272898 91826 273454
rect 92382 272898 92414 273454
rect 91794 237454 92414 272898
rect 91794 236898 91826 237454
rect 92382 236898 92414 237454
rect 91794 201454 92414 236898
rect 91794 200898 91826 201454
rect 92382 200898 92414 201454
rect 91794 165454 92414 200898
rect 91794 164898 91826 165454
rect 92382 164898 92414 165454
rect 91794 129454 92414 164898
rect 91794 128898 91826 129454
rect 92382 128898 92414 129454
rect 91794 93454 92414 128898
rect 91794 92898 91826 93454
rect 92382 92898 92414 93454
rect 91794 57454 92414 92898
rect 91794 56898 91826 57454
rect 92382 56898 92414 57454
rect 91794 21454 92414 56898
rect 91794 20898 91826 21454
rect 92382 20898 92414 21454
rect 91794 -1306 92414 20898
rect 91794 -1862 91826 -1306
rect 92382 -1862 92414 -1306
rect 91794 -1894 92414 -1862
rect 95514 673174 96134 707162
rect 95514 672618 95546 673174
rect 96102 672618 96134 673174
rect 95514 637174 96134 672618
rect 95514 636618 95546 637174
rect 96102 636618 96134 637174
rect 95514 601174 96134 636618
rect 95514 600618 95546 601174
rect 96102 600618 96134 601174
rect 95514 565174 96134 600618
rect 95514 564618 95546 565174
rect 96102 564618 96134 565174
rect 95514 529174 96134 564618
rect 95514 528618 95546 529174
rect 96102 528618 96134 529174
rect 95514 493174 96134 528618
rect 95514 492618 95546 493174
rect 96102 492618 96134 493174
rect 95514 457174 96134 492618
rect 95514 456618 95546 457174
rect 96102 456618 96134 457174
rect 95514 421174 96134 456618
rect 95514 420618 95546 421174
rect 96102 420618 96134 421174
rect 95514 385174 96134 420618
rect 95514 384618 95546 385174
rect 96102 384618 96134 385174
rect 95514 349174 96134 384618
rect 95514 348618 95546 349174
rect 96102 348618 96134 349174
rect 95514 313174 96134 348618
rect 95514 312618 95546 313174
rect 96102 312618 96134 313174
rect 95514 277174 96134 312618
rect 95514 276618 95546 277174
rect 96102 276618 96134 277174
rect 95514 241174 96134 276618
rect 95514 240618 95546 241174
rect 96102 240618 96134 241174
rect 95514 205174 96134 240618
rect 95514 204618 95546 205174
rect 96102 204618 96134 205174
rect 95514 169174 96134 204618
rect 95514 168618 95546 169174
rect 96102 168618 96134 169174
rect 95514 133174 96134 168618
rect 95514 132618 95546 133174
rect 96102 132618 96134 133174
rect 95514 97174 96134 132618
rect 95514 96618 95546 97174
rect 96102 96618 96134 97174
rect 95514 61174 96134 96618
rect 95514 60618 95546 61174
rect 96102 60618 96134 61174
rect 95514 25174 96134 60618
rect 95514 24618 95546 25174
rect 96102 24618 96134 25174
rect 95514 -3226 96134 24618
rect 95514 -3782 95546 -3226
rect 96102 -3782 96134 -3226
rect 95514 -3814 96134 -3782
rect 99234 676894 99854 709082
rect 99234 676338 99266 676894
rect 99822 676338 99854 676894
rect 99234 640894 99854 676338
rect 99234 640338 99266 640894
rect 99822 640338 99854 640894
rect 99234 604894 99854 640338
rect 99234 604338 99266 604894
rect 99822 604338 99854 604894
rect 99234 568894 99854 604338
rect 99234 568338 99266 568894
rect 99822 568338 99854 568894
rect 99234 532894 99854 568338
rect 99234 532338 99266 532894
rect 99822 532338 99854 532894
rect 99234 496894 99854 532338
rect 99234 496338 99266 496894
rect 99822 496338 99854 496894
rect 99234 460894 99854 496338
rect 99234 460338 99266 460894
rect 99822 460338 99854 460894
rect 99234 424894 99854 460338
rect 99234 424338 99266 424894
rect 99822 424338 99854 424894
rect 99234 388894 99854 424338
rect 99234 388338 99266 388894
rect 99822 388338 99854 388894
rect 99234 352894 99854 388338
rect 99234 352338 99266 352894
rect 99822 352338 99854 352894
rect 99234 316894 99854 352338
rect 99234 316338 99266 316894
rect 99822 316338 99854 316894
rect 99234 280894 99854 316338
rect 99234 280338 99266 280894
rect 99822 280338 99854 280894
rect 99234 244894 99854 280338
rect 99234 244338 99266 244894
rect 99822 244338 99854 244894
rect 99234 208894 99854 244338
rect 99234 208338 99266 208894
rect 99822 208338 99854 208894
rect 99234 172894 99854 208338
rect 99234 172338 99266 172894
rect 99822 172338 99854 172894
rect 99234 136894 99854 172338
rect 99234 136338 99266 136894
rect 99822 136338 99854 136894
rect 99234 100894 99854 136338
rect 99234 100338 99266 100894
rect 99822 100338 99854 100894
rect 99234 64894 99854 100338
rect 99234 64338 99266 64894
rect 99822 64338 99854 64894
rect 99234 28894 99854 64338
rect 99234 28338 99266 28894
rect 99822 28338 99854 28894
rect 99234 -5146 99854 28338
rect 99234 -5702 99266 -5146
rect 99822 -5702 99854 -5146
rect 99234 -5734 99854 -5702
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710042 120986 710598
rect 121542 710042 121574 710598
rect 117234 708678 117854 709670
rect 117234 708122 117266 708678
rect 117822 708122 117854 708678
rect 113514 706758 114134 707750
rect 113514 706202 113546 706758
rect 114102 706202 114134 706758
rect 102954 680058 102986 680614
rect 103542 680058 103574 680614
rect 102954 644614 103574 680058
rect 102954 644058 102986 644614
rect 103542 644058 103574 644614
rect 102954 608614 103574 644058
rect 102954 608058 102986 608614
rect 103542 608058 103574 608614
rect 102954 572614 103574 608058
rect 102954 572058 102986 572614
rect 103542 572058 103574 572614
rect 102954 536614 103574 572058
rect 102954 536058 102986 536614
rect 103542 536058 103574 536614
rect 102954 500614 103574 536058
rect 102954 500058 102986 500614
rect 103542 500058 103574 500614
rect 102954 464614 103574 500058
rect 102954 464058 102986 464614
rect 103542 464058 103574 464614
rect 102954 428614 103574 464058
rect 102954 428058 102986 428614
rect 103542 428058 103574 428614
rect 102954 392614 103574 428058
rect 102954 392058 102986 392614
rect 103542 392058 103574 392614
rect 102954 356614 103574 392058
rect 102954 356058 102986 356614
rect 103542 356058 103574 356614
rect 102954 320614 103574 356058
rect 102954 320058 102986 320614
rect 103542 320058 103574 320614
rect 102954 284614 103574 320058
rect 102954 284058 102986 284614
rect 103542 284058 103574 284614
rect 102954 248614 103574 284058
rect 102954 248058 102986 248614
rect 103542 248058 103574 248614
rect 102954 212614 103574 248058
rect 102954 212058 102986 212614
rect 103542 212058 103574 212614
rect 102954 176614 103574 212058
rect 102954 176058 102986 176614
rect 103542 176058 103574 176614
rect 102954 140614 103574 176058
rect 102954 140058 102986 140614
rect 103542 140058 103574 140614
rect 102954 104614 103574 140058
rect 102954 104058 102986 104614
rect 103542 104058 103574 104614
rect 102954 68614 103574 104058
rect 102954 68058 102986 68614
rect 103542 68058 103574 68614
rect 102954 32614 103574 68058
rect 102954 32058 102986 32614
rect 103542 32058 103574 32614
rect 84954 -6662 84986 -6106
rect 85542 -6662 85574 -6106
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 704838 110414 705830
rect 109794 704282 109826 704838
rect 110382 704282 110414 704838
rect 109794 687454 110414 704282
rect 109794 686898 109826 687454
rect 110382 686898 110414 687454
rect 109794 651454 110414 686898
rect 109794 650898 109826 651454
rect 110382 650898 110414 651454
rect 109794 615454 110414 650898
rect 109794 614898 109826 615454
rect 110382 614898 110414 615454
rect 109794 579454 110414 614898
rect 109794 578898 109826 579454
rect 110382 578898 110414 579454
rect 109794 543454 110414 578898
rect 109794 542898 109826 543454
rect 110382 542898 110414 543454
rect 109794 507454 110414 542898
rect 109794 506898 109826 507454
rect 110382 506898 110414 507454
rect 109794 471454 110414 506898
rect 109794 470898 109826 471454
rect 110382 470898 110414 471454
rect 109794 435454 110414 470898
rect 109794 434898 109826 435454
rect 110382 434898 110414 435454
rect 109794 399454 110414 434898
rect 109794 398898 109826 399454
rect 110382 398898 110414 399454
rect 109794 363454 110414 398898
rect 109794 362898 109826 363454
rect 110382 362898 110414 363454
rect 109794 327454 110414 362898
rect 109794 326898 109826 327454
rect 110382 326898 110414 327454
rect 109794 291454 110414 326898
rect 109794 290898 109826 291454
rect 110382 290898 110414 291454
rect 109794 255454 110414 290898
rect 109794 254898 109826 255454
rect 110382 254898 110414 255454
rect 109794 219454 110414 254898
rect 109794 218898 109826 219454
rect 110382 218898 110414 219454
rect 109794 183454 110414 218898
rect 109794 182898 109826 183454
rect 110382 182898 110414 183454
rect 109794 147454 110414 182898
rect 109794 146898 109826 147454
rect 110382 146898 110414 147454
rect 109794 111454 110414 146898
rect 109794 110898 109826 111454
rect 110382 110898 110414 111454
rect 109794 75454 110414 110898
rect 109794 74898 109826 75454
rect 110382 74898 110414 75454
rect 109794 39454 110414 74898
rect 109794 38898 109826 39454
rect 110382 38898 110414 39454
rect 109794 3454 110414 38898
rect 109794 2898 109826 3454
rect 110382 2898 110414 3454
rect 109794 -346 110414 2898
rect 109794 -902 109826 -346
rect 110382 -902 110414 -346
rect 109794 -1894 110414 -902
rect 113514 691174 114134 706202
rect 113514 690618 113546 691174
rect 114102 690618 114134 691174
rect 113514 655174 114134 690618
rect 113514 654618 113546 655174
rect 114102 654618 114134 655174
rect 113514 619174 114134 654618
rect 113514 618618 113546 619174
rect 114102 618618 114134 619174
rect 113514 583174 114134 618618
rect 113514 582618 113546 583174
rect 114102 582618 114134 583174
rect 113514 547174 114134 582618
rect 113514 546618 113546 547174
rect 114102 546618 114134 547174
rect 113514 511174 114134 546618
rect 113514 510618 113546 511174
rect 114102 510618 114134 511174
rect 113514 475174 114134 510618
rect 113514 474618 113546 475174
rect 114102 474618 114134 475174
rect 113514 439174 114134 474618
rect 113514 438618 113546 439174
rect 114102 438618 114134 439174
rect 113514 403174 114134 438618
rect 113514 402618 113546 403174
rect 114102 402618 114134 403174
rect 113514 367174 114134 402618
rect 113514 366618 113546 367174
rect 114102 366618 114134 367174
rect 113514 331174 114134 366618
rect 113514 330618 113546 331174
rect 114102 330618 114134 331174
rect 113514 295174 114134 330618
rect 113514 294618 113546 295174
rect 114102 294618 114134 295174
rect 113514 259174 114134 294618
rect 113514 258618 113546 259174
rect 114102 258618 114134 259174
rect 113514 223174 114134 258618
rect 113514 222618 113546 223174
rect 114102 222618 114134 223174
rect 113514 187174 114134 222618
rect 113514 186618 113546 187174
rect 114102 186618 114134 187174
rect 113514 151174 114134 186618
rect 113514 150618 113546 151174
rect 114102 150618 114134 151174
rect 113514 115174 114134 150618
rect 113514 114618 113546 115174
rect 114102 114618 114134 115174
rect 113514 79174 114134 114618
rect 113514 78618 113546 79174
rect 114102 78618 114134 79174
rect 113514 43174 114134 78618
rect 113514 42618 113546 43174
rect 114102 42618 114134 43174
rect 113514 7174 114134 42618
rect 113514 6618 113546 7174
rect 114102 6618 114134 7174
rect 113514 -2266 114134 6618
rect 113514 -2822 113546 -2266
rect 114102 -2822 114134 -2266
rect 113514 -3814 114134 -2822
rect 117234 694894 117854 708122
rect 117234 694338 117266 694894
rect 117822 694338 117854 694894
rect 117234 658894 117854 694338
rect 117234 658338 117266 658894
rect 117822 658338 117854 658894
rect 117234 622894 117854 658338
rect 117234 622338 117266 622894
rect 117822 622338 117854 622894
rect 117234 586894 117854 622338
rect 117234 586338 117266 586894
rect 117822 586338 117854 586894
rect 117234 550894 117854 586338
rect 117234 550338 117266 550894
rect 117822 550338 117854 550894
rect 117234 514894 117854 550338
rect 117234 514338 117266 514894
rect 117822 514338 117854 514894
rect 117234 478894 117854 514338
rect 117234 478338 117266 478894
rect 117822 478338 117854 478894
rect 117234 442894 117854 478338
rect 117234 442338 117266 442894
rect 117822 442338 117854 442894
rect 117234 406894 117854 442338
rect 117234 406338 117266 406894
rect 117822 406338 117854 406894
rect 117234 370894 117854 406338
rect 117234 370338 117266 370894
rect 117822 370338 117854 370894
rect 117234 334894 117854 370338
rect 117234 334338 117266 334894
rect 117822 334338 117854 334894
rect 117234 298894 117854 334338
rect 117234 298338 117266 298894
rect 117822 298338 117854 298894
rect 117234 262894 117854 298338
rect 117234 262338 117266 262894
rect 117822 262338 117854 262894
rect 117234 226894 117854 262338
rect 117234 226338 117266 226894
rect 117822 226338 117854 226894
rect 117234 190894 117854 226338
rect 117234 190338 117266 190894
rect 117822 190338 117854 190894
rect 117234 154894 117854 190338
rect 117234 154338 117266 154894
rect 117822 154338 117854 154894
rect 117234 118894 117854 154338
rect 117234 118338 117266 118894
rect 117822 118338 117854 118894
rect 117234 82894 117854 118338
rect 117234 82338 117266 82894
rect 117822 82338 117854 82894
rect 117234 46894 117854 82338
rect 117234 46338 117266 46894
rect 117822 46338 117854 46894
rect 117234 10894 117854 46338
rect 117234 10338 117266 10894
rect 117822 10338 117854 10894
rect 117234 -4186 117854 10338
rect 117234 -4742 117266 -4186
rect 117822 -4742 117854 -4186
rect 117234 -5734 117854 -4742
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711002 138986 711558
rect 139542 711002 139574 711558
rect 135234 709638 135854 709670
rect 135234 709082 135266 709638
rect 135822 709082 135854 709638
rect 131514 707718 132134 707750
rect 131514 707162 131546 707718
rect 132102 707162 132134 707718
rect 120954 698058 120986 698614
rect 121542 698058 121574 698614
rect 120954 662614 121574 698058
rect 120954 662058 120986 662614
rect 121542 662058 121574 662614
rect 120954 626614 121574 662058
rect 120954 626058 120986 626614
rect 121542 626058 121574 626614
rect 120954 590614 121574 626058
rect 120954 590058 120986 590614
rect 121542 590058 121574 590614
rect 120954 554614 121574 590058
rect 120954 554058 120986 554614
rect 121542 554058 121574 554614
rect 120954 518614 121574 554058
rect 120954 518058 120986 518614
rect 121542 518058 121574 518614
rect 120954 482614 121574 518058
rect 120954 482058 120986 482614
rect 121542 482058 121574 482614
rect 120954 446614 121574 482058
rect 120954 446058 120986 446614
rect 121542 446058 121574 446614
rect 120954 410614 121574 446058
rect 120954 410058 120986 410614
rect 121542 410058 121574 410614
rect 120954 374614 121574 410058
rect 120954 374058 120986 374614
rect 121542 374058 121574 374614
rect 120954 338614 121574 374058
rect 120954 338058 120986 338614
rect 121542 338058 121574 338614
rect 120954 302614 121574 338058
rect 120954 302058 120986 302614
rect 121542 302058 121574 302614
rect 120954 266614 121574 302058
rect 120954 266058 120986 266614
rect 121542 266058 121574 266614
rect 120954 230614 121574 266058
rect 120954 230058 120986 230614
rect 121542 230058 121574 230614
rect 120954 194614 121574 230058
rect 120954 194058 120986 194614
rect 121542 194058 121574 194614
rect 120954 158614 121574 194058
rect 120954 158058 120986 158614
rect 121542 158058 121574 158614
rect 120954 122614 121574 158058
rect 120954 122058 120986 122614
rect 121542 122058 121574 122614
rect 120954 86614 121574 122058
rect 120954 86058 120986 86614
rect 121542 86058 121574 86614
rect 120954 50614 121574 86058
rect 120954 50058 120986 50614
rect 121542 50058 121574 50614
rect 120954 14614 121574 50058
rect 120954 14058 120986 14614
rect 121542 14058 121574 14614
rect 102954 -7622 102986 -7066
rect 103542 -7622 103574 -7066
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 705798 128414 705830
rect 127794 705242 127826 705798
rect 128382 705242 128414 705798
rect 127794 669454 128414 705242
rect 127794 668898 127826 669454
rect 128382 668898 128414 669454
rect 127794 633454 128414 668898
rect 127794 632898 127826 633454
rect 128382 632898 128414 633454
rect 127794 597454 128414 632898
rect 127794 596898 127826 597454
rect 128382 596898 128414 597454
rect 127794 561454 128414 596898
rect 127794 560898 127826 561454
rect 128382 560898 128414 561454
rect 127794 525454 128414 560898
rect 127794 524898 127826 525454
rect 128382 524898 128414 525454
rect 127794 489454 128414 524898
rect 127794 488898 127826 489454
rect 128382 488898 128414 489454
rect 127794 453454 128414 488898
rect 127794 452898 127826 453454
rect 128382 452898 128414 453454
rect 127794 417454 128414 452898
rect 127794 416898 127826 417454
rect 128382 416898 128414 417454
rect 127794 381454 128414 416898
rect 127794 380898 127826 381454
rect 128382 380898 128414 381454
rect 127794 345454 128414 380898
rect 127794 344898 127826 345454
rect 128382 344898 128414 345454
rect 127794 309454 128414 344898
rect 127794 308898 127826 309454
rect 128382 308898 128414 309454
rect 127794 273454 128414 308898
rect 127794 272898 127826 273454
rect 128382 272898 128414 273454
rect 127794 237454 128414 272898
rect 127794 236898 127826 237454
rect 128382 236898 128414 237454
rect 127794 201454 128414 236898
rect 127794 200898 127826 201454
rect 128382 200898 128414 201454
rect 127794 165454 128414 200898
rect 127794 164898 127826 165454
rect 128382 164898 128414 165454
rect 127794 129454 128414 164898
rect 127794 128898 127826 129454
rect 128382 128898 128414 129454
rect 127794 93454 128414 128898
rect 127794 92898 127826 93454
rect 128382 92898 128414 93454
rect 127794 57454 128414 92898
rect 127794 56898 127826 57454
rect 128382 56898 128414 57454
rect 127794 21454 128414 56898
rect 127794 20898 127826 21454
rect 128382 20898 128414 21454
rect 127794 -1306 128414 20898
rect 127794 -1862 127826 -1306
rect 128382 -1862 128414 -1306
rect 127794 -1894 128414 -1862
rect 131514 673174 132134 707162
rect 131514 672618 131546 673174
rect 132102 672618 132134 673174
rect 131514 637174 132134 672618
rect 131514 636618 131546 637174
rect 132102 636618 132134 637174
rect 131514 601174 132134 636618
rect 131514 600618 131546 601174
rect 132102 600618 132134 601174
rect 131514 565174 132134 600618
rect 131514 564618 131546 565174
rect 132102 564618 132134 565174
rect 131514 529174 132134 564618
rect 131514 528618 131546 529174
rect 132102 528618 132134 529174
rect 131514 493174 132134 528618
rect 131514 492618 131546 493174
rect 132102 492618 132134 493174
rect 131514 457174 132134 492618
rect 131514 456618 131546 457174
rect 132102 456618 132134 457174
rect 131514 421174 132134 456618
rect 131514 420618 131546 421174
rect 132102 420618 132134 421174
rect 131514 385174 132134 420618
rect 131514 384618 131546 385174
rect 132102 384618 132134 385174
rect 131514 349174 132134 384618
rect 131514 348618 131546 349174
rect 132102 348618 132134 349174
rect 131514 313174 132134 348618
rect 131514 312618 131546 313174
rect 132102 312618 132134 313174
rect 131514 277174 132134 312618
rect 131514 276618 131546 277174
rect 132102 276618 132134 277174
rect 131514 241174 132134 276618
rect 131514 240618 131546 241174
rect 132102 240618 132134 241174
rect 131514 205174 132134 240618
rect 131514 204618 131546 205174
rect 132102 204618 132134 205174
rect 131514 169174 132134 204618
rect 131514 168618 131546 169174
rect 132102 168618 132134 169174
rect 131514 133174 132134 168618
rect 131514 132618 131546 133174
rect 132102 132618 132134 133174
rect 131514 97174 132134 132618
rect 131514 96618 131546 97174
rect 132102 96618 132134 97174
rect 131514 61174 132134 96618
rect 131514 60618 131546 61174
rect 132102 60618 132134 61174
rect 131514 25174 132134 60618
rect 131514 24618 131546 25174
rect 132102 24618 132134 25174
rect 131514 -3226 132134 24618
rect 131514 -3782 131546 -3226
rect 132102 -3782 132134 -3226
rect 131514 -3814 132134 -3782
rect 135234 676894 135854 709082
rect 135234 676338 135266 676894
rect 135822 676338 135854 676894
rect 135234 640894 135854 676338
rect 135234 640338 135266 640894
rect 135822 640338 135854 640894
rect 135234 604894 135854 640338
rect 135234 604338 135266 604894
rect 135822 604338 135854 604894
rect 135234 568894 135854 604338
rect 135234 568338 135266 568894
rect 135822 568338 135854 568894
rect 135234 532894 135854 568338
rect 135234 532338 135266 532894
rect 135822 532338 135854 532894
rect 135234 496894 135854 532338
rect 135234 496338 135266 496894
rect 135822 496338 135854 496894
rect 135234 460894 135854 496338
rect 135234 460338 135266 460894
rect 135822 460338 135854 460894
rect 135234 424894 135854 460338
rect 135234 424338 135266 424894
rect 135822 424338 135854 424894
rect 135234 388894 135854 424338
rect 135234 388338 135266 388894
rect 135822 388338 135854 388894
rect 135234 352894 135854 388338
rect 135234 352338 135266 352894
rect 135822 352338 135854 352894
rect 135234 316894 135854 352338
rect 135234 316338 135266 316894
rect 135822 316338 135854 316894
rect 135234 280894 135854 316338
rect 135234 280338 135266 280894
rect 135822 280338 135854 280894
rect 135234 244894 135854 280338
rect 135234 244338 135266 244894
rect 135822 244338 135854 244894
rect 135234 208894 135854 244338
rect 135234 208338 135266 208894
rect 135822 208338 135854 208894
rect 135234 172894 135854 208338
rect 135234 172338 135266 172894
rect 135822 172338 135854 172894
rect 135234 136894 135854 172338
rect 135234 136338 135266 136894
rect 135822 136338 135854 136894
rect 135234 100894 135854 136338
rect 135234 100338 135266 100894
rect 135822 100338 135854 100894
rect 135234 64894 135854 100338
rect 135234 64338 135266 64894
rect 135822 64338 135854 64894
rect 135234 28894 135854 64338
rect 135234 28338 135266 28894
rect 135822 28338 135854 28894
rect 135234 -5146 135854 28338
rect 135234 -5702 135266 -5146
rect 135822 -5702 135854 -5146
rect 135234 -5734 135854 -5702
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710042 156986 710598
rect 157542 710042 157574 710598
rect 153234 708678 153854 709670
rect 153234 708122 153266 708678
rect 153822 708122 153854 708678
rect 149514 706758 150134 707750
rect 149514 706202 149546 706758
rect 150102 706202 150134 706758
rect 138954 680058 138986 680614
rect 139542 680058 139574 680614
rect 138954 644614 139574 680058
rect 138954 644058 138986 644614
rect 139542 644058 139574 644614
rect 138954 608614 139574 644058
rect 138954 608058 138986 608614
rect 139542 608058 139574 608614
rect 138954 572614 139574 608058
rect 138954 572058 138986 572614
rect 139542 572058 139574 572614
rect 138954 536614 139574 572058
rect 138954 536058 138986 536614
rect 139542 536058 139574 536614
rect 138954 500614 139574 536058
rect 138954 500058 138986 500614
rect 139542 500058 139574 500614
rect 138954 464614 139574 500058
rect 138954 464058 138986 464614
rect 139542 464058 139574 464614
rect 138954 428614 139574 464058
rect 138954 428058 138986 428614
rect 139542 428058 139574 428614
rect 138954 392614 139574 428058
rect 138954 392058 138986 392614
rect 139542 392058 139574 392614
rect 138954 356614 139574 392058
rect 138954 356058 138986 356614
rect 139542 356058 139574 356614
rect 138954 320614 139574 356058
rect 138954 320058 138986 320614
rect 139542 320058 139574 320614
rect 138954 284614 139574 320058
rect 138954 284058 138986 284614
rect 139542 284058 139574 284614
rect 138954 248614 139574 284058
rect 138954 248058 138986 248614
rect 139542 248058 139574 248614
rect 138954 212614 139574 248058
rect 138954 212058 138986 212614
rect 139542 212058 139574 212614
rect 138954 176614 139574 212058
rect 138954 176058 138986 176614
rect 139542 176058 139574 176614
rect 138954 140614 139574 176058
rect 138954 140058 138986 140614
rect 139542 140058 139574 140614
rect 138954 104614 139574 140058
rect 138954 104058 138986 104614
rect 139542 104058 139574 104614
rect 138954 68614 139574 104058
rect 138954 68058 138986 68614
rect 139542 68058 139574 68614
rect 138954 32614 139574 68058
rect 138954 32058 138986 32614
rect 139542 32058 139574 32614
rect 120954 -6662 120986 -6106
rect 121542 -6662 121574 -6106
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 704838 146414 705830
rect 145794 704282 145826 704838
rect 146382 704282 146414 704838
rect 145794 687454 146414 704282
rect 145794 686898 145826 687454
rect 146382 686898 146414 687454
rect 145794 651454 146414 686898
rect 145794 650898 145826 651454
rect 146382 650898 146414 651454
rect 145794 615454 146414 650898
rect 145794 614898 145826 615454
rect 146382 614898 146414 615454
rect 145794 579454 146414 614898
rect 145794 578898 145826 579454
rect 146382 578898 146414 579454
rect 145794 543454 146414 578898
rect 145794 542898 145826 543454
rect 146382 542898 146414 543454
rect 145794 507454 146414 542898
rect 145794 506898 145826 507454
rect 146382 506898 146414 507454
rect 145794 471454 146414 506898
rect 145794 470898 145826 471454
rect 146382 470898 146414 471454
rect 145794 435454 146414 470898
rect 145794 434898 145826 435454
rect 146382 434898 146414 435454
rect 145794 399454 146414 434898
rect 145794 398898 145826 399454
rect 146382 398898 146414 399454
rect 145794 363454 146414 398898
rect 145794 362898 145826 363454
rect 146382 362898 146414 363454
rect 145794 327454 146414 362898
rect 145794 326898 145826 327454
rect 146382 326898 146414 327454
rect 145794 291454 146414 326898
rect 145794 290898 145826 291454
rect 146382 290898 146414 291454
rect 145794 255454 146414 290898
rect 145794 254898 145826 255454
rect 146382 254898 146414 255454
rect 145794 219454 146414 254898
rect 145794 218898 145826 219454
rect 146382 218898 146414 219454
rect 145794 183454 146414 218898
rect 145794 182898 145826 183454
rect 146382 182898 146414 183454
rect 145794 147454 146414 182898
rect 145794 146898 145826 147454
rect 146382 146898 146414 147454
rect 145794 111454 146414 146898
rect 145794 110898 145826 111454
rect 146382 110898 146414 111454
rect 145794 75454 146414 110898
rect 145794 74898 145826 75454
rect 146382 74898 146414 75454
rect 145794 39454 146414 74898
rect 145794 38898 145826 39454
rect 146382 38898 146414 39454
rect 145794 3454 146414 38898
rect 145794 2898 145826 3454
rect 146382 2898 146414 3454
rect 145794 -346 146414 2898
rect 145794 -902 145826 -346
rect 146382 -902 146414 -346
rect 145794 -1894 146414 -902
rect 149514 691174 150134 706202
rect 149514 690618 149546 691174
rect 150102 690618 150134 691174
rect 149514 655174 150134 690618
rect 149514 654618 149546 655174
rect 150102 654618 150134 655174
rect 149514 619174 150134 654618
rect 149514 618618 149546 619174
rect 150102 618618 150134 619174
rect 149514 583174 150134 618618
rect 149514 582618 149546 583174
rect 150102 582618 150134 583174
rect 149514 547174 150134 582618
rect 149514 546618 149546 547174
rect 150102 546618 150134 547174
rect 149514 511174 150134 546618
rect 149514 510618 149546 511174
rect 150102 510618 150134 511174
rect 149514 475174 150134 510618
rect 149514 474618 149546 475174
rect 150102 474618 150134 475174
rect 149514 439174 150134 474618
rect 149514 438618 149546 439174
rect 150102 438618 150134 439174
rect 149514 403174 150134 438618
rect 149514 402618 149546 403174
rect 150102 402618 150134 403174
rect 149514 367174 150134 402618
rect 149514 366618 149546 367174
rect 150102 366618 150134 367174
rect 149514 331174 150134 366618
rect 149514 330618 149546 331174
rect 150102 330618 150134 331174
rect 149514 295174 150134 330618
rect 149514 294618 149546 295174
rect 150102 294618 150134 295174
rect 149514 259174 150134 294618
rect 149514 258618 149546 259174
rect 150102 258618 150134 259174
rect 149514 223174 150134 258618
rect 149514 222618 149546 223174
rect 150102 222618 150134 223174
rect 149514 187174 150134 222618
rect 149514 186618 149546 187174
rect 150102 186618 150134 187174
rect 149514 151174 150134 186618
rect 149514 150618 149546 151174
rect 150102 150618 150134 151174
rect 149514 115174 150134 150618
rect 149514 114618 149546 115174
rect 150102 114618 150134 115174
rect 149514 79174 150134 114618
rect 149514 78618 149546 79174
rect 150102 78618 150134 79174
rect 149514 43174 150134 78618
rect 149514 42618 149546 43174
rect 150102 42618 150134 43174
rect 149514 7174 150134 42618
rect 149514 6618 149546 7174
rect 150102 6618 150134 7174
rect 149514 -2266 150134 6618
rect 149514 -2822 149546 -2266
rect 150102 -2822 150134 -2266
rect 149514 -3814 150134 -2822
rect 153234 694894 153854 708122
rect 153234 694338 153266 694894
rect 153822 694338 153854 694894
rect 153234 658894 153854 694338
rect 153234 658338 153266 658894
rect 153822 658338 153854 658894
rect 153234 622894 153854 658338
rect 153234 622338 153266 622894
rect 153822 622338 153854 622894
rect 153234 586894 153854 622338
rect 153234 586338 153266 586894
rect 153822 586338 153854 586894
rect 153234 550894 153854 586338
rect 153234 550338 153266 550894
rect 153822 550338 153854 550894
rect 153234 514894 153854 550338
rect 153234 514338 153266 514894
rect 153822 514338 153854 514894
rect 153234 478894 153854 514338
rect 153234 478338 153266 478894
rect 153822 478338 153854 478894
rect 153234 442894 153854 478338
rect 153234 442338 153266 442894
rect 153822 442338 153854 442894
rect 153234 406894 153854 442338
rect 153234 406338 153266 406894
rect 153822 406338 153854 406894
rect 153234 370894 153854 406338
rect 153234 370338 153266 370894
rect 153822 370338 153854 370894
rect 153234 334894 153854 370338
rect 153234 334338 153266 334894
rect 153822 334338 153854 334894
rect 153234 298894 153854 334338
rect 153234 298338 153266 298894
rect 153822 298338 153854 298894
rect 153234 262894 153854 298338
rect 153234 262338 153266 262894
rect 153822 262338 153854 262894
rect 153234 226894 153854 262338
rect 153234 226338 153266 226894
rect 153822 226338 153854 226894
rect 153234 190894 153854 226338
rect 153234 190338 153266 190894
rect 153822 190338 153854 190894
rect 153234 154894 153854 190338
rect 153234 154338 153266 154894
rect 153822 154338 153854 154894
rect 153234 118894 153854 154338
rect 153234 118338 153266 118894
rect 153822 118338 153854 118894
rect 153234 82894 153854 118338
rect 153234 82338 153266 82894
rect 153822 82338 153854 82894
rect 153234 46894 153854 82338
rect 153234 46338 153266 46894
rect 153822 46338 153854 46894
rect 153234 10894 153854 46338
rect 153234 10338 153266 10894
rect 153822 10338 153854 10894
rect 153234 -4186 153854 10338
rect 153234 -4742 153266 -4186
rect 153822 -4742 153854 -4186
rect 153234 -5734 153854 -4742
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711002 174986 711558
rect 175542 711002 175574 711558
rect 171234 709638 171854 709670
rect 171234 709082 171266 709638
rect 171822 709082 171854 709638
rect 167514 707718 168134 707750
rect 167514 707162 167546 707718
rect 168102 707162 168134 707718
rect 156954 698058 156986 698614
rect 157542 698058 157574 698614
rect 156954 662614 157574 698058
rect 156954 662058 156986 662614
rect 157542 662058 157574 662614
rect 156954 626614 157574 662058
rect 156954 626058 156986 626614
rect 157542 626058 157574 626614
rect 156954 590614 157574 626058
rect 156954 590058 156986 590614
rect 157542 590058 157574 590614
rect 156954 554614 157574 590058
rect 156954 554058 156986 554614
rect 157542 554058 157574 554614
rect 156954 518614 157574 554058
rect 156954 518058 156986 518614
rect 157542 518058 157574 518614
rect 156954 482614 157574 518058
rect 156954 482058 156986 482614
rect 157542 482058 157574 482614
rect 156954 446614 157574 482058
rect 156954 446058 156986 446614
rect 157542 446058 157574 446614
rect 156954 410614 157574 446058
rect 156954 410058 156986 410614
rect 157542 410058 157574 410614
rect 156954 374614 157574 410058
rect 156954 374058 156986 374614
rect 157542 374058 157574 374614
rect 156954 338614 157574 374058
rect 156954 338058 156986 338614
rect 157542 338058 157574 338614
rect 156954 302614 157574 338058
rect 156954 302058 156986 302614
rect 157542 302058 157574 302614
rect 156954 266614 157574 302058
rect 156954 266058 156986 266614
rect 157542 266058 157574 266614
rect 156954 230614 157574 266058
rect 156954 230058 156986 230614
rect 157542 230058 157574 230614
rect 156954 194614 157574 230058
rect 156954 194058 156986 194614
rect 157542 194058 157574 194614
rect 156954 158614 157574 194058
rect 156954 158058 156986 158614
rect 157542 158058 157574 158614
rect 156954 122614 157574 158058
rect 156954 122058 156986 122614
rect 157542 122058 157574 122614
rect 156954 86614 157574 122058
rect 156954 86058 156986 86614
rect 157542 86058 157574 86614
rect 156954 50614 157574 86058
rect 156954 50058 156986 50614
rect 157542 50058 157574 50614
rect 156954 14614 157574 50058
rect 156954 14058 156986 14614
rect 157542 14058 157574 14614
rect 138954 -7622 138986 -7066
rect 139542 -7622 139574 -7066
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 705798 164414 705830
rect 163794 705242 163826 705798
rect 164382 705242 164414 705798
rect 163794 669454 164414 705242
rect 163794 668898 163826 669454
rect 164382 668898 164414 669454
rect 163794 633454 164414 668898
rect 163794 632898 163826 633454
rect 164382 632898 164414 633454
rect 163794 597454 164414 632898
rect 163794 596898 163826 597454
rect 164382 596898 164414 597454
rect 163794 561454 164414 596898
rect 163794 560898 163826 561454
rect 164382 560898 164414 561454
rect 163794 525454 164414 560898
rect 163794 524898 163826 525454
rect 164382 524898 164414 525454
rect 163794 489454 164414 524898
rect 163794 488898 163826 489454
rect 164382 488898 164414 489454
rect 163794 453454 164414 488898
rect 163794 452898 163826 453454
rect 164382 452898 164414 453454
rect 163794 417454 164414 452898
rect 163794 416898 163826 417454
rect 164382 416898 164414 417454
rect 163794 381454 164414 416898
rect 163794 380898 163826 381454
rect 164382 380898 164414 381454
rect 163794 345454 164414 380898
rect 163794 344898 163826 345454
rect 164382 344898 164414 345454
rect 163794 309454 164414 344898
rect 163794 308898 163826 309454
rect 164382 308898 164414 309454
rect 163794 273454 164414 308898
rect 163794 272898 163826 273454
rect 164382 272898 164414 273454
rect 163794 237454 164414 272898
rect 163794 236898 163826 237454
rect 164382 236898 164414 237454
rect 163794 201454 164414 236898
rect 163794 200898 163826 201454
rect 164382 200898 164414 201454
rect 163794 165454 164414 200898
rect 163794 164898 163826 165454
rect 164382 164898 164414 165454
rect 163794 129454 164414 164898
rect 163794 128898 163826 129454
rect 164382 128898 164414 129454
rect 163794 93454 164414 128898
rect 163794 92898 163826 93454
rect 164382 92898 164414 93454
rect 163794 57454 164414 92898
rect 163794 56898 163826 57454
rect 164382 56898 164414 57454
rect 163794 21454 164414 56898
rect 163794 20898 163826 21454
rect 164382 20898 164414 21454
rect 163794 -1306 164414 20898
rect 163794 -1862 163826 -1306
rect 164382 -1862 164414 -1306
rect 163794 -1894 164414 -1862
rect 167514 673174 168134 707162
rect 167514 672618 167546 673174
rect 168102 672618 168134 673174
rect 167514 637174 168134 672618
rect 167514 636618 167546 637174
rect 168102 636618 168134 637174
rect 167514 601174 168134 636618
rect 167514 600618 167546 601174
rect 168102 600618 168134 601174
rect 167514 565174 168134 600618
rect 167514 564618 167546 565174
rect 168102 564618 168134 565174
rect 167514 529174 168134 564618
rect 167514 528618 167546 529174
rect 168102 528618 168134 529174
rect 167514 493174 168134 528618
rect 167514 492618 167546 493174
rect 168102 492618 168134 493174
rect 167514 457174 168134 492618
rect 167514 456618 167546 457174
rect 168102 456618 168134 457174
rect 167514 421174 168134 456618
rect 167514 420618 167546 421174
rect 168102 420618 168134 421174
rect 167514 385174 168134 420618
rect 167514 384618 167546 385174
rect 168102 384618 168134 385174
rect 167514 349174 168134 384618
rect 167514 348618 167546 349174
rect 168102 348618 168134 349174
rect 167514 313174 168134 348618
rect 167514 312618 167546 313174
rect 168102 312618 168134 313174
rect 167514 277174 168134 312618
rect 167514 276618 167546 277174
rect 168102 276618 168134 277174
rect 167514 241174 168134 276618
rect 167514 240618 167546 241174
rect 168102 240618 168134 241174
rect 167514 205174 168134 240618
rect 167514 204618 167546 205174
rect 168102 204618 168134 205174
rect 167514 169174 168134 204618
rect 167514 168618 167546 169174
rect 168102 168618 168134 169174
rect 167514 133174 168134 168618
rect 167514 132618 167546 133174
rect 168102 132618 168134 133174
rect 167514 97174 168134 132618
rect 167514 96618 167546 97174
rect 168102 96618 168134 97174
rect 167514 61174 168134 96618
rect 167514 60618 167546 61174
rect 168102 60618 168134 61174
rect 167514 25174 168134 60618
rect 167514 24618 167546 25174
rect 168102 24618 168134 25174
rect 167514 -3226 168134 24618
rect 167514 -3782 167546 -3226
rect 168102 -3782 168134 -3226
rect 167514 -3814 168134 -3782
rect 171234 676894 171854 709082
rect 171234 676338 171266 676894
rect 171822 676338 171854 676894
rect 171234 640894 171854 676338
rect 171234 640338 171266 640894
rect 171822 640338 171854 640894
rect 171234 604894 171854 640338
rect 171234 604338 171266 604894
rect 171822 604338 171854 604894
rect 171234 568894 171854 604338
rect 171234 568338 171266 568894
rect 171822 568338 171854 568894
rect 171234 532894 171854 568338
rect 171234 532338 171266 532894
rect 171822 532338 171854 532894
rect 171234 496894 171854 532338
rect 171234 496338 171266 496894
rect 171822 496338 171854 496894
rect 171234 460894 171854 496338
rect 171234 460338 171266 460894
rect 171822 460338 171854 460894
rect 171234 424894 171854 460338
rect 171234 424338 171266 424894
rect 171822 424338 171854 424894
rect 171234 388894 171854 424338
rect 171234 388338 171266 388894
rect 171822 388338 171854 388894
rect 171234 352894 171854 388338
rect 171234 352338 171266 352894
rect 171822 352338 171854 352894
rect 171234 316894 171854 352338
rect 171234 316338 171266 316894
rect 171822 316338 171854 316894
rect 171234 280894 171854 316338
rect 171234 280338 171266 280894
rect 171822 280338 171854 280894
rect 171234 244894 171854 280338
rect 171234 244338 171266 244894
rect 171822 244338 171854 244894
rect 171234 208894 171854 244338
rect 171234 208338 171266 208894
rect 171822 208338 171854 208894
rect 171234 172894 171854 208338
rect 171234 172338 171266 172894
rect 171822 172338 171854 172894
rect 171234 136894 171854 172338
rect 171234 136338 171266 136894
rect 171822 136338 171854 136894
rect 171234 100894 171854 136338
rect 171234 100338 171266 100894
rect 171822 100338 171854 100894
rect 171234 64894 171854 100338
rect 171234 64338 171266 64894
rect 171822 64338 171854 64894
rect 171234 28894 171854 64338
rect 171234 28338 171266 28894
rect 171822 28338 171854 28894
rect 171234 -5146 171854 28338
rect 171234 -5702 171266 -5146
rect 171822 -5702 171854 -5146
rect 171234 -5734 171854 -5702
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710042 192986 710598
rect 193542 710042 193574 710598
rect 189234 708678 189854 709670
rect 189234 708122 189266 708678
rect 189822 708122 189854 708678
rect 185514 706758 186134 707750
rect 185514 706202 185546 706758
rect 186102 706202 186134 706758
rect 174954 680058 174986 680614
rect 175542 680058 175574 680614
rect 174954 644614 175574 680058
rect 174954 644058 174986 644614
rect 175542 644058 175574 644614
rect 174954 608614 175574 644058
rect 174954 608058 174986 608614
rect 175542 608058 175574 608614
rect 174954 572614 175574 608058
rect 174954 572058 174986 572614
rect 175542 572058 175574 572614
rect 174954 536614 175574 572058
rect 174954 536058 174986 536614
rect 175542 536058 175574 536614
rect 174954 500614 175574 536058
rect 174954 500058 174986 500614
rect 175542 500058 175574 500614
rect 174954 464614 175574 500058
rect 174954 464058 174986 464614
rect 175542 464058 175574 464614
rect 174954 428614 175574 464058
rect 174954 428058 174986 428614
rect 175542 428058 175574 428614
rect 174954 392614 175574 428058
rect 174954 392058 174986 392614
rect 175542 392058 175574 392614
rect 174954 356614 175574 392058
rect 174954 356058 174986 356614
rect 175542 356058 175574 356614
rect 174954 320614 175574 356058
rect 174954 320058 174986 320614
rect 175542 320058 175574 320614
rect 174954 284614 175574 320058
rect 174954 284058 174986 284614
rect 175542 284058 175574 284614
rect 174954 248614 175574 284058
rect 174954 248058 174986 248614
rect 175542 248058 175574 248614
rect 174954 212614 175574 248058
rect 174954 212058 174986 212614
rect 175542 212058 175574 212614
rect 174954 176614 175574 212058
rect 174954 176058 174986 176614
rect 175542 176058 175574 176614
rect 174954 140614 175574 176058
rect 174954 140058 174986 140614
rect 175542 140058 175574 140614
rect 174954 104614 175574 140058
rect 174954 104058 174986 104614
rect 175542 104058 175574 104614
rect 174954 68614 175574 104058
rect 174954 68058 174986 68614
rect 175542 68058 175574 68614
rect 174954 32614 175574 68058
rect 174954 32058 174986 32614
rect 175542 32058 175574 32614
rect 156954 -6662 156986 -6106
rect 157542 -6662 157574 -6106
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 704838 182414 705830
rect 181794 704282 181826 704838
rect 182382 704282 182414 704838
rect 181794 687454 182414 704282
rect 181794 686898 181826 687454
rect 182382 686898 182414 687454
rect 181794 651454 182414 686898
rect 181794 650898 181826 651454
rect 182382 650898 182414 651454
rect 181794 615454 182414 650898
rect 181794 614898 181826 615454
rect 182382 614898 182414 615454
rect 181794 579454 182414 614898
rect 181794 578898 181826 579454
rect 182382 578898 182414 579454
rect 181794 543454 182414 578898
rect 181794 542898 181826 543454
rect 182382 542898 182414 543454
rect 181794 507454 182414 542898
rect 181794 506898 181826 507454
rect 182382 506898 182414 507454
rect 181794 471454 182414 506898
rect 181794 470898 181826 471454
rect 182382 470898 182414 471454
rect 181794 435454 182414 470898
rect 181794 434898 181826 435454
rect 182382 434898 182414 435454
rect 181794 399454 182414 434898
rect 181794 398898 181826 399454
rect 182382 398898 182414 399454
rect 181794 363454 182414 398898
rect 181794 362898 181826 363454
rect 182382 362898 182414 363454
rect 181794 327454 182414 362898
rect 181794 326898 181826 327454
rect 182382 326898 182414 327454
rect 181794 291454 182414 326898
rect 181794 290898 181826 291454
rect 182382 290898 182414 291454
rect 181794 255454 182414 290898
rect 181794 254898 181826 255454
rect 182382 254898 182414 255454
rect 181794 219454 182414 254898
rect 181794 218898 181826 219454
rect 182382 218898 182414 219454
rect 181794 183454 182414 218898
rect 181794 182898 181826 183454
rect 182382 182898 182414 183454
rect 181794 147454 182414 182898
rect 181794 146898 181826 147454
rect 182382 146898 182414 147454
rect 181794 111454 182414 146898
rect 181794 110898 181826 111454
rect 182382 110898 182414 111454
rect 181794 75454 182414 110898
rect 181794 74898 181826 75454
rect 182382 74898 182414 75454
rect 181794 39454 182414 74898
rect 181794 38898 181826 39454
rect 182382 38898 182414 39454
rect 181794 3454 182414 38898
rect 181794 2898 181826 3454
rect 182382 2898 182414 3454
rect 181794 -346 182414 2898
rect 181794 -902 181826 -346
rect 182382 -902 182414 -346
rect 181794 -1894 182414 -902
rect 185514 691174 186134 706202
rect 185514 690618 185546 691174
rect 186102 690618 186134 691174
rect 185514 655174 186134 690618
rect 185514 654618 185546 655174
rect 186102 654618 186134 655174
rect 185514 619174 186134 654618
rect 185514 618618 185546 619174
rect 186102 618618 186134 619174
rect 185514 583174 186134 618618
rect 185514 582618 185546 583174
rect 186102 582618 186134 583174
rect 185514 547174 186134 582618
rect 185514 546618 185546 547174
rect 186102 546618 186134 547174
rect 185514 511174 186134 546618
rect 185514 510618 185546 511174
rect 186102 510618 186134 511174
rect 185514 475174 186134 510618
rect 185514 474618 185546 475174
rect 186102 474618 186134 475174
rect 185514 439174 186134 474618
rect 185514 438618 185546 439174
rect 186102 438618 186134 439174
rect 185514 403174 186134 438618
rect 185514 402618 185546 403174
rect 186102 402618 186134 403174
rect 185514 367174 186134 402618
rect 185514 366618 185546 367174
rect 186102 366618 186134 367174
rect 185514 331174 186134 366618
rect 185514 330618 185546 331174
rect 186102 330618 186134 331174
rect 185514 295174 186134 330618
rect 185514 294618 185546 295174
rect 186102 294618 186134 295174
rect 185514 259174 186134 294618
rect 185514 258618 185546 259174
rect 186102 258618 186134 259174
rect 185514 223174 186134 258618
rect 185514 222618 185546 223174
rect 186102 222618 186134 223174
rect 185514 187174 186134 222618
rect 185514 186618 185546 187174
rect 186102 186618 186134 187174
rect 185514 151174 186134 186618
rect 185514 150618 185546 151174
rect 186102 150618 186134 151174
rect 185514 115174 186134 150618
rect 185514 114618 185546 115174
rect 186102 114618 186134 115174
rect 185514 79174 186134 114618
rect 185514 78618 185546 79174
rect 186102 78618 186134 79174
rect 185514 43174 186134 78618
rect 185514 42618 185546 43174
rect 186102 42618 186134 43174
rect 185514 7174 186134 42618
rect 185514 6618 185546 7174
rect 186102 6618 186134 7174
rect 185514 -2266 186134 6618
rect 185514 -2822 185546 -2266
rect 186102 -2822 186134 -2266
rect 185514 -3814 186134 -2822
rect 189234 694894 189854 708122
rect 189234 694338 189266 694894
rect 189822 694338 189854 694894
rect 189234 658894 189854 694338
rect 189234 658338 189266 658894
rect 189822 658338 189854 658894
rect 189234 622894 189854 658338
rect 189234 622338 189266 622894
rect 189822 622338 189854 622894
rect 189234 586894 189854 622338
rect 189234 586338 189266 586894
rect 189822 586338 189854 586894
rect 189234 550894 189854 586338
rect 189234 550338 189266 550894
rect 189822 550338 189854 550894
rect 189234 514894 189854 550338
rect 189234 514338 189266 514894
rect 189822 514338 189854 514894
rect 189234 478894 189854 514338
rect 189234 478338 189266 478894
rect 189822 478338 189854 478894
rect 189234 442894 189854 478338
rect 189234 442338 189266 442894
rect 189822 442338 189854 442894
rect 189234 406894 189854 442338
rect 189234 406338 189266 406894
rect 189822 406338 189854 406894
rect 189234 370894 189854 406338
rect 189234 370338 189266 370894
rect 189822 370338 189854 370894
rect 189234 334894 189854 370338
rect 189234 334338 189266 334894
rect 189822 334338 189854 334894
rect 189234 298894 189854 334338
rect 189234 298338 189266 298894
rect 189822 298338 189854 298894
rect 189234 262894 189854 298338
rect 189234 262338 189266 262894
rect 189822 262338 189854 262894
rect 189234 226894 189854 262338
rect 189234 226338 189266 226894
rect 189822 226338 189854 226894
rect 189234 190894 189854 226338
rect 189234 190338 189266 190894
rect 189822 190338 189854 190894
rect 189234 154894 189854 190338
rect 189234 154338 189266 154894
rect 189822 154338 189854 154894
rect 189234 118894 189854 154338
rect 189234 118338 189266 118894
rect 189822 118338 189854 118894
rect 189234 82894 189854 118338
rect 189234 82338 189266 82894
rect 189822 82338 189854 82894
rect 189234 46894 189854 82338
rect 189234 46338 189266 46894
rect 189822 46338 189854 46894
rect 189234 10894 189854 46338
rect 189234 10338 189266 10894
rect 189822 10338 189854 10894
rect 189234 -4186 189854 10338
rect 189234 -4742 189266 -4186
rect 189822 -4742 189854 -4186
rect 189234 -5734 189854 -4742
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711002 210986 711558
rect 211542 711002 211574 711558
rect 207234 709638 207854 709670
rect 207234 709082 207266 709638
rect 207822 709082 207854 709638
rect 203514 707718 204134 707750
rect 203514 707162 203546 707718
rect 204102 707162 204134 707718
rect 192954 698058 192986 698614
rect 193542 698058 193574 698614
rect 192954 662614 193574 698058
rect 192954 662058 192986 662614
rect 193542 662058 193574 662614
rect 192954 626614 193574 662058
rect 192954 626058 192986 626614
rect 193542 626058 193574 626614
rect 192954 590614 193574 626058
rect 192954 590058 192986 590614
rect 193542 590058 193574 590614
rect 192954 554614 193574 590058
rect 192954 554058 192986 554614
rect 193542 554058 193574 554614
rect 192954 518614 193574 554058
rect 192954 518058 192986 518614
rect 193542 518058 193574 518614
rect 192954 482614 193574 518058
rect 192954 482058 192986 482614
rect 193542 482058 193574 482614
rect 192954 446614 193574 482058
rect 192954 446058 192986 446614
rect 193542 446058 193574 446614
rect 192954 410614 193574 446058
rect 192954 410058 192986 410614
rect 193542 410058 193574 410614
rect 192954 374614 193574 410058
rect 192954 374058 192986 374614
rect 193542 374058 193574 374614
rect 192954 338614 193574 374058
rect 192954 338058 192986 338614
rect 193542 338058 193574 338614
rect 192954 302614 193574 338058
rect 192954 302058 192986 302614
rect 193542 302058 193574 302614
rect 192954 266614 193574 302058
rect 192954 266058 192986 266614
rect 193542 266058 193574 266614
rect 192954 230614 193574 266058
rect 192954 230058 192986 230614
rect 193542 230058 193574 230614
rect 192954 194614 193574 230058
rect 192954 194058 192986 194614
rect 193542 194058 193574 194614
rect 192954 158614 193574 194058
rect 192954 158058 192986 158614
rect 193542 158058 193574 158614
rect 192954 122614 193574 158058
rect 192954 122058 192986 122614
rect 193542 122058 193574 122614
rect 192954 86614 193574 122058
rect 192954 86058 192986 86614
rect 193542 86058 193574 86614
rect 192954 50614 193574 86058
rect 192954 50058 192986 50614
rect 193542 50058 193574 50614
rect 192954 14614 193574 50058
rect 192954 14058 192986 14614
rect 193542 14058 193574 14614
rect 174954 -7622 174986 -7066
rect 175542 -7622 175574 -7066
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 705798 200414 705830
rect 199794 705242 199826 705798
rect 200382 705242 200414 705798
rect 199794 669454 200414 705242
rect 199794 668898 199826 669454
rect 200382 668898 200414 669454
rect 199794 633454 200414 668898
rect 199794 632898 199826 633454
rect 200382 632898 200414 633454
rect 199794 597454 200414 632898
rect 199794 596898 199826 597454
rect 200382 596898 200414 597454
rect 199794 561454 200414 596898
rect 199794 560898 199826 561454
rect 200382 560898 200414 561454
rect 199794 525454 200414 560898
rect 199794 524898 199826 525454
rect 200382 524898 200414 525454
rect 199794 489454 200414 524898
rect 199794 488898 199826 489454
rect 200382 488898 200414 489454
rect 199794 453454 200414 488898
rect 199794 452898 199826 453454
rect 200382 452898 200414 453454
rect 199794 417454 200414 452898
rect 199794 416898 199826 417454
rect 200382 416898 200414 417454
rect 199794 381454 200414 416898
rect 199794 380898 199826 381454
rect 200382 380898 200414 381454
rect 199794 345454 200414 380898
rect 199794 344898 199826 345454
rect 200382 344898 200414 345454
rect 199794 309454 200414 344898
rect 199794 308898 199826 309454
rect 200382 308898 200414 309454
rect 199794 273454 200414 308898
rect 199794 272898 199826 273454
rect 200382 272898 200414 273454
rect 199794 237454 200414 272898
rect 199794 236898 199826 237454
rect 200382 236898 200414 237454
rect 199794 201454 200414 236898
rect 199794 200898 199826 201454
rect 200382 200898 200414 201454
rect 199794 165454 200414 200898
rect 199794 164898 199826 165454
rect 200382 164898 200414 165454
rect 199794 129454 200414 164898
rect 199794 128898 199826 129454
rect 200382 128898 200414 129454
rect 199794 93454 200414 128898
rect 199794 92898 199826 93454
rect 200382 92898 200414 93454
rect 199794 57454 200414 92898
rect 199794 56898 199826 57454
rect 200382 56898 200414 57454
rect 199794 21454 200414 56898
rect 199794 20898 199826 21454
rect 200382 20898 200414 21454
rect 199794 -1306 200414 20898
rect 199794 -1862 199826 -1306
rect 200382 -1862 200414 -1306
rect 199794 -1894 200414 -1862
rect 203514 673174 204134 707162
rect 203514 672618 203546 673174
rect 204102 672618 204134 673174
rect 203514 637174 204134 672618
rect 203514 636618 203546 637174
rect 204102 636618 204134 637174
rect 203514 601174 204134 636618
rect 203514 600618 203546 601174
rect 204102 600618 204134 601174
rect 203514 565174 204134 600618
rect 203514 564618 203546 565174
rect 204102 564618 204134 565174
rect 203514 529174 204134 564618
rect 203514 528618 203546 529174
rect 204102 528618 204134 529174
rect 203514 493174 204134 528618
rect 203514 492618 203546 493174
rect 204102 492618 204134 493174
rect 203514 457174 204134 492618
rect 203514 456618 203546 457174
rect 204102 456618 204134 457174
rect 203514 421174 204134 456618
rect 203514 420618 203546 421174
rect 204102 420618 204134 421174
rect 203514 385174 204134 420618
rect 203514 384618 203546 385174
rect 204102 384618 204134 385174
rect 203514 349174 204134 384618
rect 203514 348618 203546 349174
rect 204102 348618 204134 349174
rect 203514 313174 204134 348618
rect 203514 312618 203546 313174
rect 204102 312618 204134 313174
rect 203514 277174 204134 312618
rect 203514 276618 203546 277174
rect 204102 276618 204134 277174
rect 203514 241174 204134 276618
rect 203514 240618 203546 241174
rect 204102 240618 204134 241174
rect 203514 205174 204134 240618
rect 203514 204618 203546 205174
rect 204102 204618 204134 205174
rect 203514 169174 204134 204618
rect 203514 168618 203546 169174
rect 204102 168618 204134 169174
rect 203514 133174 204134 168618
rect 203514 132618 203546 133174
rect 204102 132618 204134 133174
rect 203514 97174 204134 132618
rect 203514 96618 203546 97174
rect 204102 96618 204134 97174
rect 203514 61174 204134 96618
rect 203514 60618 203546 61174
rect 204102 60618 204134 61174
rect 203514 25174 204134 60618
rect 203514 24618 203546 25174
rect 204102 24618 204134 25174
rect 203514 -3226 204134 24618
rect 203514 -3782 203546 -3226
rect 204102 -3782 204134 -3226
rect 203514 -3814 204134 -3782
rect 207234 676894 207854 709082
rect 207234 676338 207266 676894
rect 207822 676338 207854 676894
rect 207234 640894 207854 676338
rect 207234 640338 207266 640894
rect 207822 640338 207854 640894
rect 207234 604894 207854 640338
rect 207234 604338 207266 604894
rect 207822 604338 207854 604894
rect 207234 568894 207854 604338
rect 207234 568338 207266 568894
rect 207822 568338 207854 568894
rect 207234 532894 207854 568338
rect 207234 532338 207266 532894
rect 207822 532338 207854 532894
rect 207234 496894 207854 532338
rect 207234 496338 207266 496894
rect 207822 496338 207854 496894
rect 207234 460894 207854 496338
rect 207234 460338 207266 460894
rect 207822 460338 207854 460894
rect 207234 424894 207854 460338
rect 207234 424338 207266 424894
rect 207822 424338 207854 424894
rect 207234 388894 207854 424338
rect 207234 388338 207266 388894
rect 207822 388338 207854 388894
rect 207234 352894 207854 388338
rect 207234 352338 207266 352894
rect 207822 352338 207854 352894
rect 207234 316894 207854 352338
rect 207234 316338 207266 316894
rect 207822 316338 207854 316894
rect 207234 280894 207854 316338
rect 207234 280338 207266 280894
rect 207822 280338 207854 280894
rect 207234 244894 207854 280338
rect 207234 244338 207266 244894
rect 207822 244338 207854 244894
rect 207234 208894 207854 244338
rect 207234 208338 207266 208894
rect 207822 208338 207854 208894
rect 207234 172894 207854 208338
rect 207234 172338 207266 172894
rect 207822 172338 207854 172894
rect 207234 136894 207854 172338
rect 207234 136338 207266 136894
rect 207822 136338 207854 136894
rect 207234 100894 207854 136338
rect 207234 100338 207266 100894
rect 207822 100338 207854 100894
rect 207234 64894 207854 100338
rect 207234 64338 207266 64894
rect 207822 64338 207854 64894
rect 207234 28894 207854 64338
rect 207234 28338 207266 28894
rect 207822 28338 207854 28894
rect 207234 -5146 207854 28338
rect 207234 -5702 207266 -5146
rect 207822 -5702 207854 -5146
rect 207234 -5734 207854 -5702
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710042 228986 710598
rect 229542 710042 229574 710598
rect 225234 708678 225854 709670
rect 225234 708122 225266 708678
rect 225822 708122 225854 708678
rect 221514 706758 222134 707750
rect 221514 706202 221546 706758
rect 222102 706202 222134 706758
rect 210954 680058 210986 680614
rect 211542 680058 211574 680614
rect 210954 644614 211574 680058
rect 210954 644058 210986 644614
rect 211542 644058 211574 644614
rect 210954 608614 211574 644058
rect 210954 608058 210986 608614
rect 211542 608058 211574 608614
rect 210954 572614 211574 608058
rect 210954 572058 210986 572614
rect 211542 572058 211574 572614
rect 210954 536614 211574 572058
rect 210954 536058 210986 536614
rect 211542 536058 211574 536614
rect 210954 500614 211574 536058
rect 210954 500058 210986 500614
rect 211542 500058 211574 500614
rect 210954 464614 211574 500058
rect 210954 464058 210986 464614
rect 211542 464058 211574 464614
rect 210954 428614 211574 464058
rect 210954 428058 210986 428614
rect 211542 428058 211574 428614
rect 210954 392614 211574 428058
rect 210954 392058 210986 392614
rect 211542 392058 211574 392614
rect 210954 356614 211574 392058
rect 210954 356058 210986 356614
rect 211542 356058 211574 356614
rect 210954 320614 211574 356058
rect 210954 320058 210986 320614
rect 211542 320058 211574 320614
rect 210954 284614 211574 320058
rect 210954 284058 210986 284614
rect 211542 284058 211574 284614
rect 210954 248614 211574 284058
rect 210954 248058 210986 248614
rect 211542 248058 211574 248614
rect 210954 212614 211574 248058
rect 210954 212058 210986 212614
rect 211542 212058 211574 212614
rect 210954 176614 211574 212058
rect 210954 176058 210986 176614
rect 211542 176058 211574 176614
rect 210954 140614 211574 176058
rect 210954 140058 210986 140614
rect 211542 140058 211574 140614
rect 210954 104614 211574 140058
rect 210954 104058 210986 104614
rect 211542 104058 211574 104614
rect 210954 68614 211574 104058
rect 210954 68058 210986 68614
rect 211542 68058 211574 68614
rect 210954 32614 211574 68058
rect 210954 32058 210986 32614
rect 211542 32058 211574 32614
rect 192954 -6662 192986 -6106
rect 193542 -6662 193574 -6106
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 704838 218414 705830
rect 217794 704282 217826 704838
rect 218382 704282 218414 704838
rect 217794 687454 218414 704282
rect 217794 686898 217826 687454
rect 218382 686898 218414 687454
rect 217794 651454 218414 686898
rect 217794 650898 217826 651454
rect 218382 650898 218414 651454
rect 217794 615454 218414 650898
rect 217794 614898 217826 615454
rect 218382 614898 218414 615454
rect 217794 579454 218414 614898
rect 217794 578898 217826 579454
rect 218382 578898 218414 579454
rect 217794 543454 218414 578898
rect 217794 542898 217826 543454
rect 218382 542898 218414 543454
rect 217794 507454 218414 542898
rect 217794 506898 217826 507454
rect 218382 506898 218414 507454
rect 217794 471454 218414 506898
rect 217794 470898 217826 471454
rect 218382 470898 218414 471454
rect 217794 435454 218414 470898
rect 217794 434898 217826 435454
rect 218382 434898 218414 435454
rect 217794 399454 218414 434898
rect 217794 398898 217826 399454
rect 218382 398898 218414 399454
rect 217794 363454 218414 398898
rect 217794 362898 217826 363454
rect 218382 362898 218414 363454
rect 217794 327454 218414 362898
rect 217794 326898 217826 327454
rect 218382 326898 218414 327454
rect 217794 291454 218414 326898
rect 217794 290898 217826 291454
rect 218382 290898 218414 291454
rect 217794 255454 218414 290898
rect 217794 254898 217826 255454
rect 218382 254898 218414 255454
rect 217794 219454 218414 254898
rect 217794 218898 217826 219454
rect 218382 218898 218414 219454
rect 217794 183454 218414 218898
rect 217794 182898 217826 183454
rect 218382 182898 218414 183454
rect 217794 147454 218414 182898
rect 217794 146898 217826 147454
rect 218382 146898 218414 147454
rect 217794 111454 218414 146898
rect 217794 110898 217826 111454
rect 218382 110898 218414 111454
rect 217794 75454 218414 110898
rect 217794 74898 217826 75454
rect 218382 74898 218414 75454
rect 217794 39454 218414 74898
rect 217794 38898 217826 39454
rect 218382 38898 218414 39454
rect 217794 3454 218414 38898
rect 217794 2898 217826 3454
rect 218382 2898 218414 3454
rect 217794 -346 218414 2898
rect 217794 -902 217826 -346
rect 218382 -902 218414 -346
rect 217794 -1894 218414 -902
rect 221514 691174 222134 706202
rect 221514 690618 221546 691174
rect 222102 690618 222134 691174
rect 221514 655174 222134 690618
rect 221514 654618 221546 655174
rect 222102 654618 222134 655174
rect 221514 619174 222134 654618
rect 221514 618618 221546 619174
rect 222102 618618 222134 619174
rect 221514 583174 222134 618618
rect 221514 582618 221546 583174
rect 222102 582618 222134 583174
rect 221514 547174 222134 582618
rect 221514 546618 221546 547174
rect 222102 546618 222134 547174
rect 221514 511174 222134 546618
rect 221514 510618 221546 511174
rect 222102 510618 222134 511174
rect 221514 475174 222134 510618
rect 221514 474618 221546 475174
rect 222102 474618 222134 475174
rect 221514 439174 222134 474618
rect 221514 438618 221546 439174
rect 222102 438618 222134 439174
rect 221514 403174 222134 438618
rect 221514 402618 221546 403174
rect 222102 402618 222134 403174
rect 221514 367174 222134 402618
rect 221514 366618 221546 367174
rect 222102 366618 222134 367174
rect 221514 331174 222134 366618
rect 221514 330618 221546 331174
rect 222102 330618 222134 331174
rect 221514 295174 222134 330618
rect 221514 294618 221546 295174
rect 222102 294618 222134 295174
rect 221514 259174 222134 294618
rect 221514 258618 221546 259174
rect 222102 258618 222134 259174
rect 221514 223174 222134 258618
rect 221514 222618 221546 223174
rect 222102 222618 222134 223174
rect 221514 187174 222134 222618
rect 221514 186618 221546 187174
rect 222102 186618 222134 187174
rect 221514 151174 222134 186618
rect 221514 150618 221546 151174
rect 222102 150618 222134 151174
rect 221514 115174 222134 150618
rect 221514 114618 221546 115174
rect 222102 114618 222134 115174
rect 221514 79174 222134 114618
rect 221514 78618 221546 79174
rect 222102 78618 222134 79174
rect 221514 43174 222134 78618
rect 221514 42618 221546 43174
rect 222102 42618 222134 43174
rect 221514 7174 222134 42618
rect 221514 6618 221546 7174
rect 222102 6618 222134 7174
rect 221514 -2266 222134 6618
rect 221514 -2822 221546 -2266
rect 222102 -2822 222134 -2266
rect 221514 -3814 222134 -2822
rect 225234 694894 225854 708122
rect 225234 694338 225266 694894
rect 225822 694338 225854 694894
rect 225234 658894 225854 694338
rect 225234 658338 225266 658894
rect 225822 658338 225854 658894
rect 225234 622894 225854 658338
rect 225234 622338 225266 622894
rect 225822 622338 225854 622894
rect 225234 586894 225854 622338
rect 225234 586338 225266 586894
rect 225822 586338 225854 586894
rect 225234 550894 225854 586338
rect 225234 550338 225266 550894
rect 225822 550338 225854 550894
rect 225234 514894 225854 550338
rect 225234 514338 225266 514894
rect 225822 514338 225854 514894
rect 225234 478894 225854 514338
rect 225234 478338 225266 478894
rect 225822 478338 225854 478894
rect 225234 442894 225854 478338
rect 225234 442338 225266 442894
rect 225822 442338 225854 442894
rect 225234 406894 225854 442338
rect 225234 406338 225266 406894
rect 225822 406338 225854 406894
rect 225234 370894 225854 406338
rect 225234 370338 225266 370894
rect 225822 370338 225854 370894
rect 225234 334894 225854 370338
rect 225234 334338 225266 334894
rect 225822 334338 225854 334894
rect 225234 298894 225854 334338
rect 225234 298338 225266 298894
rect 225822 298338 225854 298894
rect 225234 262894 225854 298338
rect 225234 262338 225266 262894
rect 225822 262338 225854 262894
rect 225234 226894 225854 262338
rect 225234 226338 225266 226894
rect 225822 226338 225854 226894
rect 225234 190894 225854 226338
rect 225234 190338 225266 190894
rect 225822 190338 225854 190894
rect 225234 154894 225854 190338
rect 225234 154338 225266 154894
rect 225822 154338 225854 154894
rect 225234 118894 225854 154338
rect 225234 118338 225266 118894
rect 225822 118338 225854 118894
rect 225234 82894 225854 118338
rect 225234 82338 225266 82894
rect 225822 82338 225854 82894
rect 225234 46894 225854 82338
rect 225234 46338 225266 46894
rect 225822 46338 225854 46894
rect 225234 10894 225854 46338
rect 225234 10338 225266 10894
rect 225822 10338 225854 10894
rect 225234 -4186 225854 10338
rect 225234 -4742 225266 -4186
rect 225822 -4742 225854 -4186
rect 225234 -5734 225854 -4742
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711002 246986 711558
rect 247542 711002 247574 711558
rect 243234 709638 243854 709670
rect 243234 709082 243266 709638
rect 243822 709082 243854 709638
rect 239514 707718 240134 707750
rect 239514 707162 239546 707718
rect 240102 707162 240134 707718
rect 228954 698058 228986 698614
rect 229542 698058 229574 698614
rect 228954 662614 229574 698058
rect 228954 662058 228986 662614
rect 229542 662058 229574 662614
rect 228954 626614 229574 662058
rect 228954 626058 228986 626614
rect 229542 626058 229574 626614
rect 228954 590614 229574 626058
rect 228954 590058 228986 590614
rect 229542 590058 229574 590614
rect 228954 554614 229574 590058
rect 228954 554058 228986 554614
rect 229542 554058 229574 554614
rect 228954 518614 229574 554058
rect 228954 518058 228986 518614
rect 229542 518058 229574 518614
rect 228954 482614 229574 518058
rect 228954 482058 228986 482614
rect 229542 482058 229574 482614
rect 228954 446614 229574 482058
rect 235794 705798 236414 705830
rect 235794 705242 235826 705798
rect 236382 705242 236414 705798
rect 235794 669454 236414 705242
rect 235794 668898 235826 669454
rect 236382 668898 236414 669454
rect 235794 633454 236414 668898
rect 235794 632898 235826 633454
rect 236382 632898 236414 633454
rect 235794 597454 236414 632898
rect 235794 596898 235826 597454
rect 236382 596898 236414 597454
rect 235794 561454 236414 596898
rect 235794 560898 235826 561454
rect 236382 560898 236414 561454
rect 235794 525454 236414 560898
rect 235794 524898 235826 525454
rect 236382 524898 236414 525454
rect 235794 489454 236414 524898
rect 235794 488898 235826 489454
rect 236382 488898 236414 489454
rect 235794 460000 236414 488898
rect 239514 673174 240134 707162
rect 239514 672618 239546 673174
rect 240102 672618 240134 673174
rect 239514 637174 240134 672618
rect 239514 636618 239546 637174
rect 240102 636618 240134 637174
rect 239514 601174 240134 636618
rect 239514 600618 239546 601174
rect 240102 600618 240134 601174
rect 239514 565174 240134 600618
rect 239514 564618 239546 565174
rect 240102 564618 240134 565174
rect 239514 529174 240134 564618
rect 239514 528618 239546 529174
rect 240102 528618 240134 529174
rect 239514 493174 240134 528618
rect 239514 492618 239546 493174
rect 240102 492618 240134 493174
rect 239514 460000 240134 492618
rect 243234 676894 243854 709082
rect 243234 676338 243266 676894
rect 243822 676338 243854 676894
rect 243234 640894 243854 676338
rect 243234 640338 243266 640894
rect 243822 640338 243854 640894
rect 243234 604894 243854 640338
rect 243234 604338 243266 604894
rect 243822 604338 243854 604894
rect 243234 568894 243854 604338
rect 243234 568338 243266 568894
rect 243822 568338 243854 568894
rect 243234 532894 243854 568338
rect 243234 532338 243266 532894
rect 243822 532338 243854 532894
rect 243234 496894 243854 532338
rect 243234 496338 243266 496894
rect 243822 496338 243854 496894
rect 243234 460894 243854 496338
rect 243234 460338 243266 460894
rect 243822 460338 243854 460894
rect 243234 460000 243854 460338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710042 264986 710598
rect 265542 710042 265574 710598
rect 261234 708678 261854 709670
rect 261234 708122 261266 708678
rect 261822 708122 261854 708678
rect 257514 706758 258134 707750
rect 257514 706202 257546 706758
rect 258102 706202 258134 706758
rect 246954 680058 246986 680614
rect 247542 680058 247574 680614
rect 246954 644614 247574 680058
rect 246954 644058 246986 644614
rect 247542 644058 247574 644614
rect 246954 608614 247574 644058
rect 246954 608058 246986 608614
rect 247542 608058 247574 608614
rect 246954 572614 247574 608058
rect 246954 572058 246986 572614
rect 247542 572058 247574 572614
rect 246954 536614 247574 572058
rect 246954 536058 246986 536614
rect 247542 536058 247574 536614
rect 246954 500614 247574 536058
rect 246954 500058 246986 500614
rect 247542 500058 247574 500614
rect 246954 464614 247574 500058
rect 246954 464058 246986 464614
rect 247542 464058 247574 464614
rect 246954 460000 247574 464058
rect 253794 704838 254414 705830
rect 253794 704282 253826 704838
rect 254382 704282 254414 704838
rect 253794 687454 254414 704282
rect 253794 686898 253826 687454
rect 254382 686898 254414 687454
rect 253794 651454 254414 686898
rect 253794 650898 253826 651454
rect 254382 650898 254414 651454
rect 253794 615454 254414 650898
rect 253794 614898 253826 615454
rect 254382 614898 254414 615454
rect 253794 579454 254414 614898
rect 253794 578898 253826 579454
rect 254382 578898 254414 579454
rect 253794 543454 254414 578898
rect 253794 542898 253826 543454
rect 254382 542898 254414 543454
rect 253794 507454 254414 542898
rect 253794 506898 253826 507454
rect 254382 506898 254414 507454
rect 253794 471454 254414 506898
rect 253794 470898 253826 471454
rect 254382 470898 254414 471454
rect 253794 460000 254414 470898
rect 257514 691174 258134 706202
rect 257514 690618 257546 691174
rect 258102 690618 258134 691174
rect 257514 655174 258134 690618
rect 257514 654618 257546 655174
rect 258102 654618 258134 655174
rect 257514 619174 258134 654618
rect 257514 618618 257546 619174
rect 258102 618618 258134 619174
rect 257514 583174 258134 618618
rect 257514 582618 257546 583174
rect 258102 582618 258134 583174
rect 257514 547174 258134 582618
rect 257514 546618 257546 547174
rect 258102 546618 258134 547174
rect 257514 511174 258134 546618
rect 257514 510618 257546 511174
rect 258102 510618 258134 511174
rect 257514 475174 258134 510618
rect 257514 474618 257546 475174
rect 258102 474618 258134 475174
rect 257514 460000 258134 474618
rect 261234 694894 261854 708122
rect 261234 694338 261266 694894
rect 261822 694338 261854 694894
rect 261234 658894 261854 694338
rect 261234 658338 261266 658894
rect 261822 658338 261854 658894
rect 261234 622894 261854 658338
rect 261234 622338 261266 622894
rect 261822 622338 261854 622894
rect 261234 586894 261854 622338
rect 261234 586338 261266 586894
rect 261822 586338 261854 586894
rect 261234 550894 261854 586338
rect 261234 550338 261266 550894
rect 261822 550338 261854 550894
rect 261234 514894 261854 550338
rect 261234 514338 261266 514894
rect 261822 514338 261854 514894
rect 261234 478894 261854 514338
rect 261234 478338 261266 478894
rect 261822 478338 261854 478894
rect 261234 460000 261854 478338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711002 282986 711558
rect 283542 711002 283574 711558
rect 279234 709638 279854 709670
rect 279234 709082 279266 709638
rect 279822 709082 279854 709638
rect 275514 707718 276134 707750
rect 275514 707162 275546 707718
rect 276102 707162 276134 707718
rect 264954 698058 264986 698614
rect 265542 698058 265574 698614
rect 264954 662614 265574 698058
rect 264954 662058 264986 662614
rect 265542 662058 265574 662614
rect 264954 626614 265574 662058
rect 264954 626058 264986 626614
rect 265542 626058 265574 626614
rect 264954 590614 265574 626058
rect 264954 590058 264986 590614
rect 265542 590058 265574 590614
rect 264954 554614 265574 590058
rect 264954 554058 264986 554614
rect 265542 554058 265574 554614
rect 264954 518614 265574 554058
rect 264954 518058 264986 518614
rect 265542 518058 265574 518614
rect 264954 482614 265574 518058
rect 264954 482058 264986 482614
rect 265542 482058 265574 482614
rect 264954 460000 265574 482058
rect 271794 705798 272414 705830
rect 271794 705242 271826 705798
rect 272382 705242 272414 705798
rect 271794 669454 272414 705242
rect 271794 668898 271826 669454
rect 272382 668898 272414 669454
rect 271794 633454 272414 668898
rect 271794 632898 271826 633454
rect 272382 632898 272414 633454
rect 271794 597454 272414 632898
rect 271794 596898 271826 597454
rect 272382 596898 272414 597454
rect 271794 561454 272414 596898
rect 271794 560898 271826 561454
rect 272382 560898 272414 561454
rect 271794 525454 272414 560898
rect 271794 524898 271826 525454
rect 272382 524898 272414 525454
rect 271794 489454 272414 524898
rect 271794 488898 271826 489454
rect 272382 488898 272414 489454
rect 271794 460000 272414 488898
rect 275514 673174 276134 707162
rect 275514 672618 275546 673174
rect 276102 672618 276134 673174
rect 275514 637174 276134 672618
rect 275514 636618 275546 637174
rect 276102 636618 276134 637174
rect 275514 601174 276134 636618
rect 275514 600618 275546 601174
rect 276102 600618 276134 601174
rect 275514 565174 276134 600618
rect 275514 564618 275546 565174
rect 276102 564618 276134 565174
rect 275514 529174 276134 564618
rect 275514 528618 275546 529174
rect 276102 528618 276134 529174
rect 275514 493174 276134 528618
rect 275514 492618 275546 493174
rect 276102 492618 276134 493174
rect 275514 460000 276134 492618
rect 279234 676894 279854 709082
rect 279234 676338 279266 676894
rect 279822 676338 279854 676894
rect 279234 640894 279854 676338
rect 279234 640338 279266 640894
rect 279822 640338 279854 640894
rect 279234 604894 279854 640338
rect 279234 604338 279266 604894
rect 279822 604338 279854 604894
rect 279234 568894 279854 604338
rect 279234 568338 279266 568894
rect 279822 568338 279854 568894
rect 279234 532894 279854 568338
rect 279234 532338 279266 532894
rect 279822 532338 279854 532894
rect 279234 496894 279854 532338
rect 279234 496338 279266 496894
rect 279822 496338 279854 496894
rect 279234 460894 279854 496338
rect 279234 460338 279266 460894
rect 279822 460338 279854 460894
rect 279234 460000 279854 460338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710042 300986 710598
rect 301542 710042 301574 710598
rect 297234 708678 297854 709670
rect 297234 708122 297266 708678
rect 297822 708122 297854 708678
rect 293514 706758 294134 707750
rect 293514 706202 293546 706758
rect 294102 706202 294134 706758
rect 282954 680058 282986 680614
rect 283542 680058 283574 680614
rect 282954 644614 283574 680058
rect 282954 644058 282986 644614
rect 283542 644058 283574 644614
rect 282954 608614 283574 644058
rect 282954 608058 282986 608614
rect 283542 608058 283574 608614
rect 282954 572614 283574 608058
rect 282954 572058 282986 572614
rect 283542 572058 283574 572614
rect 282954 536614 283574 572058
rect 282954 536058 282986 536614
rect 283542 536058 283574 536614
rect 282954 500614 283574 536058
rect 282954 500058 282986 500614
rect 283542 500058 283574 500614
rect 282954 464614 283574 500058
rect 282954 464058 282986 464614
rect 283542 464058 283574 464614
rect 282954 460000 283574 464058
rect 289794 704838 290414 705830
rect 289794 704282 289826 704838
rect 290382 704282 290414 704838
rect 289794 687454 290414 704282
rect 289794 686898 289826 687454
rect 290382 686898 290414 687454
rect 289794 651454 290414 686898
rect 289794 650898 289826 651454
rect 290382 650898 290414 651454
rect 289794 615454 290414 650898
rect 289794 614898 289826 615454
rect 290382 614898 290414 615454
rect 289794 579454 290414 614898
rect 289794 578898 289826 579454
rect 290382 578898 290414 579454
rect 289794 543454 290414 578898
rect 289794 542898 289826 543454
rect 290382 542898 290414 543454
rect 289794 507454 290414 542898
rect 289794 506898 289826 507454
rect 290382 506898 290414 507454
rect 289794 471454 290414 506898
rect 289794 470898 289826 471454
rect 290382 470898 290414 471454
rect 289794 460000 290414 470898
rect 293514 691174 294134 706202
rect 293514 690618 293546 691174
rect 294102 690618 294134 691174
rect 293514 655174 294134 690618
rect 293514 654618 293546 655174
rect 294102 654618 294134 655174
rect 293514 619174 294134 654618
rect 293514 618618 293546 619174
rect 294102 618618 294134 619174
rect 293514 583174 294134 618618
rect 293514 582618 293546 583174
rect 294102 582618 294134 583174
rect 293514 547174 294134 582618
rect 293514 546618 293546 547174
rect 294102 546618 294134 547174
rect 293514 511174 294134 546618
rect 293514 510618 293546 511174
rect 294102 510618 294134 511174
rect 293514 475174 294134 510618
rect 293514 474618 293546 475174
rect 294102 474618 294134 475174
rect 293514 460000 294134 474618
rect 297234 694894 297854 708122
rect 297234 694338 297266 694894
rect 297822 694338 297854 694894
rect 297234 658894 297854 694338
rect 297234 658338 297266 658894
rect 297822 658338 297854 658894
rect 297234 622894 297854 658338
rect 297234 622338 297266 622894
rect 297822 622338 297854 622894
rect 297234 586894 297854 622338
rect 297234 586338 297266 586894
rect 297822 586338 297854 586894
rect 297234 550894 297854 586338
rect 297234 550338 297266 550894
rect 297822 550338 297854 550894
rect 297234 514894 297854 550338
rect 297234 514338 297266 514894
rect 297822 514338 297854 514894
rect 297234 478894 297854 514338
rect 297234 478338 297266 478894
rect 297822 478338 297854 478894
rect 297234 460000 297854 478338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711002 318986 711558
rect 319542 711002 319574 711558
rect 315234 709638 315854 709670
rect 315234 709082 315266 709638
rect 315822 709082 315854 709638
rect 311514 707718 312134 707750
rect 311514 707162 311546 707718
rect 312102 707162 312134 707718
rect 300954 698058 300986 698614
rect 301542 698058 301574 698614
rect 300954 662614 301574 698058
rect 300954 662058 300986 662614
rect 301542 662058 301574 662614
rect 300954 626614 301574 662058
rect 300954 626058 300986 626614
rect 301542 626058 301574 626614
rect 300954 590614 301574 626058
rect 300954 590058 300986 590614
rect 301542 590058 301574 590614
rect 300954 554614 301574 590058
rect 300954 554058 300986 554614
rect 301542 554058 301574 554614
rect 300954 518614 301574 554058
rect 300954 518058 300986 518614
rect 301542 518058 301574 518614
rect 300954 482614 301574 518058
rect 300954 482058 300986 482614
rect 301542 482058 301574 482614
rect 300954 460000 301574 482058
rect 307794 705798 308414 705830
rect 307794 705242 307826 705798
rect 308382 705242 308414 705798
rect 307794 669454 308414 705242
rect 307794 668898 307826 669454
rect 308382 668898 308414 669454
rect 307794 633454 308414 668898
rect 307794 632898 307826 633454
rect 308382 632898 308414 633454
rect 307794 597454 308414 632898
rect 307794 596898 307826 597454
rect 308382 596898 308414 597454
rect 307794 561454 308414 596898
rect 307794 560898 307826 561454
rect 308382 560898 308414 561454
rect 307794 525454 308414 560898
rect 307794 524898 307826 525454
rect 308382 524898 308414 525454
rect 307794 489454 308414 524898
rect 307794 488898 307826 489454
rect 308382 488898 308414 489454
rect 307794 460000 308414 488898
rect 311514 673174 312134 707162
rect 311514 672618 311546 673174
rect 312102 672618 312134 673174
rect 311514 637174 312134 672618
rect 311514 636618 311546 637174
rect 312102 636618 312134 637174
rect 311514 601174 312134 636618
rect 311514 600618 311546 601174
rect 312102 600618 312134 601174
rect 311514 565174 312134 600618
rect 311514 564618 311546 565174
rect 312102 564618 312134 565174
rect 311514 529174 312134 564618
rect 311514 528618 311546 529174
rect 312102 528618 312134 529174
rect 311514 493174 312134 528618
rect 311514 492618 311546 493174
rect 312102 492618 312134 493174
rect 311514 460000 312134 492618
rect 315234 676894 315854 709082
rect 315234 676338 315266 676894
rect 315822 676338 315854 676894
rect 315234 640894 315854 676338
rect 315234 640338 315266 640894
rect 315822 640338 315854 640894
rect 315234 604894 315854 640338
rect 315234 604338 315266 604894
rect 315822 604338 315854 604894
rect 315234 568894 315854 604338
rect 315234 568338 315266 568894
rect 315822 568338 315854 568894
rect 315234 532894 315854 568338
rect 315234 532338 315266 532894
rect 315822 532338 315854 532894
rect 315234 496894 315854 532338
rect 315234 496338 315266 496894
rect 315822 496338 315854 496894
rect 315234 460894 315854 496338
rect 315234 460338 315266 460894
rect 315822 460338 315854 460894
rect 315234 460000 315854 460338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710042 336986 710598
rect 337542 710042 337574 710598
rect 333234 708678 333854 709670
rect 333234 708122 333266 708678
rect 333822 708122 333854 708678
rect 329514 706758 330134 707750
rect 329514 706202 329546 706758
rect 330102 706202 330134 706758
rect 318954 680058 318986 680614
rect 319542 680058 319574 680614
rect 318954 644614 319574 680058
rect 318954 644058 318986 644614
rect 319542 644058 319574 644614
rect 318954 608614 319574 644058
rect 318954 608058 318986 608614
rect 319542 608058 319574 608614
rect 318954 572614 319574 608058
rect 318954 572058 318986 572614
rect 319542 572058 319574 572614
rect 318954 536614 319574 572058
rect 318954 536058 318986 536614
rect 319542 536058 319574 536614
rect 318954 500614 319574 536058
rect 318954 500058 318986 500614
rect 319542 500058 319574 500614
rect 318954 464614 319574 500058
rect 318954 464058 318986 464614
rect 319542 464058 319574 464614
rect 318954 460000 319574 464058
rect 325794 704838 326414 705830
rect 325794 704282 325826 704838
rect 326382 704282 326414 704838
rect 325794 687454 326414 704282
rect 325794 686898 325826 687454
rect 326382 686898 326414 687454
rect 325794 651454 326414 686898
rect 325794 650898 325826 651454
rect 326382 650898 326414 651454
rect 325794 615454 326414 650898
rect 325794 614898 325826 615454
rect 326382 614898 326414 615454
rect 325794 579454 326414 614898
rect 325794 578898 325826 579454
rect 326382 578898 326414 579454
rect 325794 543454 326414 578898
rect 325794 542898 325826 543454
rect 326382 542898 326414 543454
rect 325794 507454 326414 542898
rect 325794 506898 325826 507454
rect 326382 506898 326414 507454
rect 325794 471454 326414 506898
rect 325794 470898 325826 471454
rect 326382 470898 326414 471454
rect 325794 460000 326414 470898
rect 329514 691174 330134 706202
rect 329514 690618 329546 691174
rect 330102 690618 330134 691174
rect 329514 655174 330134 690618
rect 329514 654618 329546 655174
rect 330102 654618 330134 655174
rect 329514 619174 330134 654618
rect 329514 618618 329546 619174
rect 330102 618618 330134 619174
rect 329514 583174 330134 618618
rect 329514 582618 329546 583174
rect 330102 582618 330134 583174
rect 329514 547174 330134 582618
rect 329514 546618 329546 547174
rect 330102 546618 330134 547174
rect 329514 511174 330134 546618
rect 329514 510618 329546 511174
rect 330102 510618 330134 511174
rect 329514 475174 330134 510618
rect 329514 474618 329546 475174
rect 330102 474618 330134 475174
rect 329514 460000 330134 474618
rect 333234 694894 333854 708122
rect 333234 694338 333266 694894
rect 333822 694338 333854 694894
rect 333234 658894 333854 694338
rect 333234 658338 333266 658894
rect 333822 658338 333854 658894
rect 333234 622894 333854 658338
rect 333234 622338 333266 622894
rect 333822 622338 333854 622894
rect 333234 586894 333854 622338
rect 333234 586338 333266 586894
rect 333822 586338 333854 586894
rect 333234 550894 333854 586338
rect 333234 550338 333266 550894
rect 333822 550338 333854 550894
rect 333234 514894 333854 550338
rect 333234 514338 333266 514894
rect 333822 514338 333854 514894
rect 333234 478894 333854 514338
rect 333234 478338 333266 478894
rect 333822 478338 333854 478894
rect 333234 460000 333854 478338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711002 354986 711558
rect 355542 711002 355574 711558
rect 351234 709638 351854 709670
rect 351234 709082 351266 709638
rect 351822 709082 351854 709638
rect 347514 707718 348134 707750
rect 347514 707162 347546 707718
rect 348102 707162 348134 707718
rect 336954 698058 336986 698614
rect 337542 698058 337574 698614
rect 336954 662614 337574 698058
rect 336954 662058 336986 662614
rect 337542 662058 337574 662614
rect 336954 626614 337574 662058
rect 336954 626058 336986 626614
rect 337542 626058 337574 626614
rect 336954 590614 337574 626058
rect 336954 590058 336986 590614
rect 337542 590058 337574 590614
rect 336954 554614 337574 590058
rect 336954 554058 336986 554614
rect 337542 554058 337574 554614
rect 336954 518614 337574 554058
rect 336954 518058 336986 518614
rect 337542 518058 337574 518614
rect 336954 482614 337574 518058
rect 336954 482058 336986 482614
rect 337542 482058 337574 482614
rect 336954 460000 337574 482058
rect 343794 705798 344414 705830
rect 343794 705242 343826 705798
rect 344382 705242 344414 705798
rect 343794 669454 344414 705242
rect 343794 668898 343826 669454
rect 344382 668898 344414 669454
rect 343794 633454 344414 668898
rect 343794 632898 343826 633454
rect 344382 632898 344414 633454
rect 343794 597454 344414 632898
rect 343794 596898 343826 597454
rect 344382 596898 344414 597454
rect 343794 561454 344414 596898
rect 343794 560898 343826 561454
rect 344382 560898 344414 561454
rect 343794 525454 344414 560898
rect 343794 524898 343826 525454
rect 344382 524898 344414 525454
rect 343794 489454 344414 524898
rect 343794 488898 343826 489454
rect 344382 488898 344414 489454
rect 343794 460000 344414 488898
rect 347514 673174 348134 707162
rect 347514 672618 347546 673174
rect 348102 672618 348134 673174
rect 347514 637174 348134 672618
rect 347514 636618 347546 637174
rect 348102 636618 348134 637174
rect 347514 601174 348134 636618
rect 347514 600618 347546 601174
rect 348102 600618 348134 601174
rect 347514 565174 348134 600618
rect 347514 564618 347546 565174
rect 348102 564618 348134 565174
rect 347514 529174 348134 564618
rect 347514 528618 347546 529174
rect 348102 528618 348134 529174
rect 347514 493174 348134 528618
rect 347514 492618 347546 493174
rect 348102 492618 348134 493174
rect 347514 460000 348134 492618
rect 351234 676894 351854 709082
rect 351234 676338 351266 676894
rect 351822 676338 351854 676894
rect 351234 640894 351854 676338
rect 351234 640338 351266 640894
rect 351822 640338 351854 640894
rect 351234 604894 351854 640338
rect 351234 604338 351266 604894
rect 351822 604338 351854 604894
rect 351234 568894 351854 604338
rect 351234 568338 351266 568894
rect 351822 568338 351854 568894
rect 351234 532894 351854 568338
rect 351234 532338 351266 532894
rect 351822 532338 351854 532894
rect 351234 496894 351854 532338
rect 351234 496338 351266 496894
rect 351822 496338 351854 496894
rect 351234 460894 351854 496338
rect 351234 460338 351266 460894
rect 351822 460338 351854 460894
rect 351234 460000 351854 460338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710042 372986 710598
rect 373542 710042 373574 710598
rect 369234 708678 369854 709670
rect 369234 708122 369266 708678
rect 369822 708122 369854 708678
rect 365514 706758 366134 707750
rect 365514 706202 365546 706758
rect 366102 706202 366134 706758
rect 354954 680058 354986 680614
rect 355542 680058 355574 680614
rect 354954 644614 355574 680058
rect 354954 644058 354986 644614
rect 355542 644058 355574 644614
rect 354954 608614 355574 644058
rect 354954 608058 354986 608614
rect 355542 608058 355574 608614
rect 354954 572614 355574 608058
rect 354954 572058 354986 572614
rect 355542 572058 355574 572614
rect 354954 536614 355574 572058
rect 354954 536058 354986 536614
rect 355542 536058 355574 536614
rect 354954 500614 355574 536058
rect 354954 500058 354986 500614
rect 355542 500058 355574 500614
rect 354954 464614 355574 500058
rect 354954 464058 354986 464614
rect 355542 464058 355574 464614
rect 354954 460000 355574 464058
rect 361794 704838 362414 705830
rect 361794 704282 361826 704838
rect 362382 704282 362414 704838
rect 361794 687454 362414 704282
rect 361794 686898 361826 687454
rect 362382 686898 362414 687454
rect 361794 651454 362414 686898
rect 361794 650898 361826 651454
rect 362382 650898 362414 651454
rect 361794 615454 362414 650898
rect 361794 614898 361826 615454
rect 362382 614898 362414 615454
rect 361794 579454 362414 614898
rect 361794 578898 361826 579454
rect 362382 578898 362414 579454
rect 361794 543454 362414 578898
rect 361794 542898 361826 543454
rect 362382 542898 362414 543454
rect 361794 507454 362414 542898
rect 361794 506898 361826 507454
rect 362382 506898 362414 507454
rect 361794 471454 362414 506898
rect 361794 470898 361826 471454
rect 362382 470898 362414 471454
rect 361794 460000 362414 470898
rect 365514 691174 366134 706202
rect 365514 690618 365546 691174
rect 366102 690618 366134 691174
rect 365514 655174 366134 690618
rect 365514 654618 365546 655174
rect 366102 654618 366134 655174
rect 365514 619174 366134 654618
rect 365514 618618 365546 619174
rect 366102 618618 366134 619174
rect 365514 583174 366134 618618
rect 365514 582618 365546 583174
rect 366102 582618 366134 583174
rect 365514 547174 366134 582618
rect 365514 546618 365546 547174
rect 366102 546618 366134 547174
rect 365514 511174 366134 546618
rect 365514 510618 365546 511174
rect 366102 510618 366134 511174
rect 365514 475174 366134 510618
rect 365514 474618 365546 475174
rect 366102 474618 366134 475174
rect 365514 460000 366134 474618
rect 369234 694894 369854 708122
rect 369234 694338 369266 694894
rect 369822 694338 369854 694894
rect 369234 658894 369854 694338
rect 369234 658338 369266 658894
rect 369822 658338 369854 658894
rect 369234 622894 369854 658338
rect 369234 622338 369266 622894
rect 369822 622338 369854 622894
rect 369234 586894 369854 622338
rect 369234 586338 369266 586894
rect 369822 586338 369854 586894
rect 369234 550894 369854 586338
rect 369234 550338 369266 550894
rect 369822 550338 369854 550894
rect 369234 514894 369854 550338
rect 369234 514338 369266 514894
rect 369822 514338 369854 514894
rect 369234 478894 369854 514338
rect 369234 478338 369266 478894
rect 369822 478338 369854 478894
rect 369234 460000 369854 478338
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711002 390986 711558
rect 391542 711002 391574 711558
rect 387234 709638 387854 709670
rect 387234 709082 387266 709638
rect 387822 709082 387854 709638
rect 383514 707718 384134 707750
rect 383514 707162 383546 707718
rect 384102 707162 384134 707718
rect 372954 698058 372986 698614
rect 373542 698058 373574 698614
rect 372954 662614 373574 698058
rect 372954 662058 372986 662614
rect 373542 662058 373574 662614
rect 372954 626614 373574 662058
rect 372954 626058 372986 626614
rect 373542 626058 373574 626614
rect 372954 590614 373574 626058
rect 372954 590058 372986 590614
rect 373542 590058 373574 590614
rect 372954 554614 373574 590058
rect 372954 554058 372986 554614
rect 373542 554058 373574 554614
rect 372954 518614 373574 554058
rect 372954 518058 372986 518614
rect 373542 518058 373574 518614
rect 372954 482614 373574 518058
rect 372954 482058 372986 482614
rect 373542 482058 373574 482614
rect 372954 460000 373574 482058
rect 379794 705798 380414 705830
rect 379794 705242 379826 705798
rect 380382 705242 380414 705798
rect 379794 669454 380414 705242
rect 379794 668898 379826 669454
rect 380382 668898 380414 669454
rect 379794 633454 380414 668898
rect 379794 632898 379826 633454
rect 380382 632898 380414 633454
rect 379794 597454 380414 632898
rect 379794 596898 379826 597454
rect 380382 596898 380414 597454
rect 379794 561454 380414 596898
rect 379794 560898 379826 561454
rect 380382 560898 380414 561454
rect 379794 525454 380414 560898
rect 379794 524898 379826 525454
rect 380382 524898 380414 525454
rect 379794 489454 380414 524898
rect 379794 488898 379826 489454
rect 380382 488898 380414 489454
rect 379794 460000 380414 488898
rect 383514 673174 384134 707162
rect 383514 672618 383546 673174
rect 384102 672618 384134 673174
rect 383514 637174 384134 672618
rect 383514 636618 383546 637174
rect 384102 636618 384134 637174
rect 383514 601174 384134 636618
rect 383514 600618 383546 601174
rect 384102 600618 384134 601174
rect 383514 565174 384134 600618
rect 383514 564618 383546 565174
rect 384102 564618 384134 565174
rect 383514 529174 384134 564618
rect 383514 528618 383546 529174
rect 384102 528618 384134 529174
rect 383514 493174 384134 528618
rect 383514 492618 383546 493174
rect 384102 492618 384134 493174
rect 383514 460000 384134 492618
rect 387234 676894 387854 709082
rect 387234 676338 387266 676894
rect 387822 676338 387854 676894
rect 387234 640894 387854 676338
rect 387234 640338 387266 640894
rect 387822 640338 387854 640894
rect 387234 604894 387854 640338
rect 387234 604338 387266 604894
rect 387822 604338 387854 604894
rect 387234 568894 387854 604338
rect 387234 568338 387266 568894
rect 387822 568338 387854 568894
rect 387234 532894 387854 568338
rect 387234 532338 387266 532894
rect 387822 532338 387854 532894
rect 387234 496894 387854 532338
rect 387234 496338 387266 496894
rect 387822 496338 387854 496894
rect 387234 460894 387854 496338
rect 387234 460338 387266 460894
rect 387822 460338 387854 460894
rect 387234 460000 387854 460338
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710042 408986 710598
rect 409542 710042 409574 710598
rect 405234 708678 405854 709670
rect 405234 708122 405266 708678
rect 405822 708122 405854 708678
rect 401514 706758 402134 707750
rect 401514 706202 401546 706758
rect 402102 706202 402134 706758
rect 390954 680058 390986 680614
rect 391542 680058 391574 680614
rect 390954 644614 391574 680058
rect 390954 644058 390986 644614
rect 391542 644058 391574 644614
rect 390954 608614 391574 644058
rect 390954 608058 390986 608614
rect 391542 608058 391574 608614
rect 390954 572614 391574 608058
rect 390954 572058 390986 572614
rect 391542 572058 391574 572614
rect 390954 536614 391574 572058
rect 390954 536058 390986 536614
rect 391542 536058 391574 536614
rect 390954 500614 391574 536058
rect 390954 500058 390986 500614
rect 391542 500058 391574 500614
rect 390954 464614 391574 500058
rect 390954 464058 390986 464614
rect 391542 464058 391574 464614
rect 390954 460000 391574 464058
rect 397794 704838 398414 705830
rect 397794 704282 397826 704838
rect 398382 704282 398414 704838
rect 397794 687454 398414 704282
rect 397794 686898 397826 687454
rect 398382 686898 398414 687454
rect 397794 651454 398414 686898
rect 397794 650898 397826 651454
rect 398382 650898 398414 651454
rect 397794 615454 398414 650898
rect 397794 614898 397826 615454
rect 398382 614898 398414 615454
rect 397794 579454 398414 614898
rect 397794 578898 397826 579454
rect 398382 578898 398414 579454
rect 397794 543454 398414 578898
rect 397794 542898 397826 543454
rect 398382 542898 398414 543454
rect 397794 507454 398414 542898
rect 397794 506898 397826 507454
rect 398382 506898 398414 507454
rect 397794 471454 398414 506898
rect 397794 470898 397826 471454
rect 398382 470898 398414 471454
rect 397794 460000 398414 470898
rect 401514 691174 402134 706202
rect 401514 690618 401546 691174
rect 402102 690618 402134 691174
rect 401514 655174 402134 690618
rect 401514 654618 401546 655174
rect 402102 654618 402134 655174
rect 401514 619174 402134 654618
rect 401514 618618 401546 619174
rect 402102 618618 402134 619174
rect 401514 583174 402134 618618
rect 401514 582618 401546 583174
rect 402102 582618 402134 583174
rect 401514 547174 402134 582618
rect 401514 546618 401546 547174
rect 402102 546618 402134 547174
rect 401514 511174 402134 546618
rect 401514 510618 401546 511174
rect 402102 510618 402134 511174
rect 401514 475174 402134 510618
rect 401514 474618 401546 475174
rect 402102 474618 402134 475174
rect 401514 460000 402134 474618
rect 405234 694894 405854 708122
rect 405234 694338 405266 694894
rect 405822 694338 405854 694894
rect 405234 658894 405854 694338
rect 405234 658338 405266 658894
rect 405822 658338 405854 658894
rect 405234 622894 405854 658338
rect 405234 622338 405266 622894
rect 405822 622338 405854 622894
rect 405234 586894 405854 622338
rect 405234 586338 405266 586894
rect 405822 586338 405854 586894
rect 405234 550894 405854 586338
rect 405234 550338 405266 550894
rect 405822 550338 405854 550894
rect 405234 514894 405854 550338
rect 405234 514338 405266 514894
rect 405822 514338 405854 514894
rect 405234 478894 405854 514338
rect 405234 478338 405266 478894
rect 405822 478338 405854 478894
rect 405234 460000 405854 478338
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711002 426986 711558
rect 427542 711002 427574 711558
rect 423234 709638 423854 709670
rect 423234 709082 423266 709638
rect 423822 709082 423854 709638
rect 419514 707718 420134 707750
rect 419514 707162 419546 707718
rect 420102 707162 420134 707718
rect 408954 698058 408986 698614
rect 409542 698058 409574 698614
rect 408954 662614 409574 698058
rect 408954 662058 408986 662614
rect 409542 662058 409574 662614
rect 408954 626614 409574 662058
rect 408954 626058 408986 626614
rect 409542 626058 409574 626614
rect 408954 590614 409574 626058
rect 408954 590058 408986 590614
rect 409542 590058 409574 590614
rect 408954 554614 409574 590058
rect 408954 554058 408986 554614
rect 409542 554058 409574 554614
rect 408954 518614 409574 554058
rect 408954 518058 408986 518614
rect 409542 518058 409574 518614
rect 408954 482614 409574 518058
rect 408954 482058 408986 482614
rect 409542 482058 409574 482614
rect 408954 460000 409574 482058
rect 415794 705798 416414 705830
rect 415794 705242 415826 705798
rect 416382 705242 416414 705798
rect 415794 669454 416414 705242
rect 415794 668898 415826 669454
rect 416382 668898 416414 669454
rect 415794 633454 416414 668898
rect 415794 632898 415826 633454
rect 416382 632898 416414 633454
rect 415794 597454 416414 632898
rect 415794 596898 415826 597454
rect 416382 596898 416414 597454
rect 415794 561454 416414 596898
rect 415794 560898 415826 561454
rect 416382 560898 416414 561454
rect 415794 525454 416414 560898
rect 415794 524898 415826 525454
rect 416382 524898 416414 525454
rect 415794 489454 416414 524898
rect 415794 488898 415826 489454
rect 416382 488898 416414 489454
rect 415794 460000 416414 488898
rect 419514 673174 420134 707162
rect 419514 672618 419546 673174
rect 420102 672618 420134 673174
rect 419514 637174 420134 672618
rect 419514 636618 419546 637174
rect 420102 636618 420134 637174
rect 419514 601174 420134 636618
rect 419514 600618 419546 601174
rect 420102 600618 420134 601174
rect 419514 565174 420134 600618
rect 419514 564618 419546 565174
rect 420102 564618 420134 565174
rect 419514 529174 420134 564618
rect 419514 528618 419546 529174
rect 420102 528618 420134 529174
rect 419514 493174 420134 528618
rect 419514 492618 419546 493174
rect 420102 492618 420134 493174
rect 385355 457468 385421 457469
rect 385355 457404 385356 457468
rect 385420 457404 385421 457468
rect 385355 457403 385421 457404
rect 390139 457468 390205 457469
rect 390139 457404 390140 457468
rect 390204 457404 390205 457468
rect 390139 457403 390205 457404
rect 394923 457468 394989 457469
rect 394923 457404 394924 457468
rect 394988 457404 394989 457468
rect 394923 457403 394989 457404
rect 408723 457468 408789 457469
rect 408723 457404 408724 457468
rect 408788 457404 408789 457468
rect 408723 457403 408789 457404
rect 409827 457468 409893 457469
rect 409827 457404 409828 457468
rect 409892 457404 409893 457468
rect 409827 457403 409893 457404
rect 411299 457468 411365 457469
rect 411299 457404 411300 457468
rect 411364 457404 411365 457468
rect 411299 457403 411365 457404
rect 233739 456924 233805 456925
rect 233739 456860 233740 456924
rect 233804 456860 233805 456924
rect 233739 456859 233805 456860
rect 228954 446058 228986 446614
rect 229542 446058 229574 446614
rect 228954 410614 229574 446058
rect 228954 410058 228986 410614
rect 229542 410058 229574 410614
rect 228954 374614 229574 410058
rect 228954 374058 228986 374614
rect 229542 374058 229574 374614
rect 228954 338614 229574 374058
rect 228954 338058 228986 338614
rect 229542 338058 229574 338614
rect 228954 302614 229574 338058
rect 228954 302058 228986 302614
rect 229542 302058 229574 302614
rect 228954 266614 229574 302058
rect 228954 266058 228986 266614
rect 229542 266058 229574 266614
rect 228954 230614 229574 266058
rect 228954 230058 228986 230614
rect 229542 230058 229574 230614
rect 228954 194614 229574 230058
rect 228954 194058 228986 194614
rect 229542 194058 229574 194614
rect 228954 158614 229574 194058
rect 228954 158058 228986 158614
rect 229542 158058 229574 158614
rect 228954 122614 229574 158058
rect 228954 122058 228986 122614
rect 229542 122058 229574 122614
rect 228954 86614 229574 122058
rect 228954 86058 228986 86614
rect 229542 86058 229574 86614
rect 228954 50614 229574 86058
rect 228954 50058 228986 50614
rect 229542 50058 229574 50614
rect 228954 14614 229574 50058
rect 233742 44301 233802 456859
rect 385358 456381 385418 457403
rect 385355 456380 385421 456381
rect 385355 456316 385356 456380
rect 385420 456316 385421 456380
rect 385355 456315 385421 456316
rect 390142 456245 390202 457403
rect 390139 456244 390205 456245
rect 390139 456180 390140 456244
rect 390204 456180 390205 456244
rect 390139 456179 390205 456180
rect 394926 456109 394986 457403
rect 394923 456108 394989 456109
rect 394923 456044 394924 456108
rect 394988 456044 394989 456108
rect 394923 456043 394989 456044
rect 254568 453454 254888 453486
rect 254568 453218 254610 453454
rect 254846 453218 254888 453454
rect 254568 453134 254888 453218
rect 254568 452898 254610 453134
rect 254846 452898 254888 453134
rect 254568 452866 254888 452898
rect 285288 453454 285608 453486
rect 285288 453218 285330 453454
rect 285566 453218 285608 453454
rect 285288 453134 285608 453218
rect 285288 452898 285330 453134
rect 285566 452898 285608 453134
rect 285288 452866 285608 452898
rect 316008 453454 316328 453486
rect 316008 453218 316050 453454
rect 316286 453218 316328 453454
rect 316008 453134 316328 453218
rect 316008 452898 316050 453134
rect 316286 452898 316328 453134
rect 316008 452866 316328 452898
rect 346728 453454 347048 453486
rect 346728 453218 346770 453454
rect 347006 453218 347048 453454
rect 346728 453134 347048 453218
rect 346728 452898 346770 453134
rect 347006 452898 347048 453134
rect 346728 452866 347048 452898
rect 377448 453454 377768 453486
rect 377448 453218 377490 453454
rect 377726 453218 377768 453454
rect 377448 453134 377768 453218
rect 377448 452898 377490 453134
rect 377726 452898 377768 453134
rect 377448 452866 377768 452898
rect 408168 453454 408488 453486
rect 408168 453218 408210 453454
rect 408446 453218 408488 453454
rect 408168 453134 408488 453218
rect 408168 452898 408210 453134
rect 408446 452898 408488 453134
rect 408168 452866 408488 452898
rect 239208 435454 239528 435486
rect 239208 435218 239250 435454
rect 239486 435218 239528 435454
rect 239208 435134 239528 435218
rect 239208 434898 239250 435134
rect 239486 434898 239528 435134
rect 239208 434866 239528 434898
rect 269928 435454 270248 435486
rect 269928 435218 269970 435454
rect 270206 435218 270248 435454
rect 269928 435134 270248 435218
rect 269928 434898 269970 435134
rect 270206 434898 270248 435134
rect 269928 434866 270248 434898
rect 300648 435454 300968 435486
rect 300648 435218 300690 435454
rect 300926 435218 300968 435454
rect 300648 435134 300968 435218
rect 300648 434898 300690 435134
rect 300926 434898 300968 435134
rect 300648 434866 300968 434898
rect 331368 435454 331688 435486
rect 331368 435218 331410 435454
rect 331646 435218 331688 435454
rect 331368 435134 331688 435218
rect 331368 434898 331410 435134
rect 331646 434898 331688 435134
rect 331368 434866 331688 434898
rect 362088 435454 362408 435486
rect 362088 435218 362130 435454
rect 362366 435218 362408 435454
rect 362088 435134 362408 435218
rect 362088 434898 362130 435134
rect 362366 434898 362408 435134
rect 362088 434866 362408 434898
rect 392808 435454 393128 435486
rect 392808 435218 392850 435454
rect 393086 435218 393128 435454
rect 392808 435134 393128 435218
rect 392808 434898 392850 435134
rect 393086 434898 393128 435134
rect 392808 434866 393128 434898
rect 254568 417454 254888 417486
rect 254568 417218 254610 417454
rect 254846 417218 254888 417454
rect 254568 417134 254888 417218
rect 254568 416898 254610 417134
rect 254846 416898 254888 417134
rect 254568 416866 254888 416898
rect 285288 417454 285608 417486
rect 285288 417218 285330 417454
rect 285566 417218 285608 417454
rect 285288 417134 285608 417218
rect 285288 416898 285330 417134
rect 285566 416898 285608 417134
rect 285288 416866 285608 416898
rect 316008 417454 316328 417486
rect 316008 417218 316050 417454
rect 316286 417218 316328 417454
rect 316008 417134 316328 417218
rect 316008 416898 316050 417134
rect 316286 416898 316328 417134
rect 316008 416866 316328 416898
rect 346728 417454 347048 417486
rect 346728 417218 346770 417454
rect 347006 417218 347048 417454
rect 346728 417134 347048 417218
rect 346728 416898 346770 417134
rect 347006 416898 347048 417134
rect 346728 416866 347048 416898
rect 377448 417454 377768 417486
rect 377448 417218 377490 417454
rect 377726 417218 377768 417454
rect 377448 417134 377768 417218
rect 377448 416898 377490 417134
rect 377726 416898 377768 417134
rect 377448 416866 377768 416898
rect 408168 417454 408488 417486
rect 408168 417218 408210 417454
rect 408446 417218 408488 417454
rect 408168 417134 408488 417218
rect 408168 416898 408210 417134
rect 408446 416898 408488 417134
rect 408168 416866 408488 416898
rect 239208 399454 239528 399486
rect 239208 399218 239250 399454
rect 239486 399218 239528 399454
rect 239208 399134 239528 399218
rect 239208 398898 239250 399134
rect 239486 398898 239528 399134
rect 239208 398866 239528 398898
rect 269928 399454 270248 399486
rect 269928 399218 269970 399454
rect 270206 399218 270248 399454
rect 269928 399134 270248 399218
rect 269928 398898 269970 399134
rect 270206 398898 270248 399134
rect 269928 398866 270248 398898
rect 300648 399454 300968 399486
rect 300648 399218 300690 399454
rect 300926 399218 300968 399454
rect 300648 399134 300968 399218
rect 300648 398898 300690 399134
rect 300926 398898 300968 399134
rect 300648 398866 300968 398898
rect 331368 399454 331688 399486
rect 331368 399218 331410 399454
rect 331646 399218 331688 399454
rect 331368 399134 331688 399218
rect 331368 398898 331410 399134
rect 331646 398898 331688 399134
rect 331368 398866 331688 398898
rect 362088 399454 362408 399486
rect 362088 399218 362130 399454
rect 362366 399218 362408 399454
rect 362088 399134 362408 399218
rect 362088 398898 362130 399134
rect 362366 398898 362408 399134
rect 362088 398866 362408 398898
rect 392808 399454 393128 399486
rect 392808 399218 392850 399454
rect 393086 399218 393128 399454
rect 392808 399134 393128 399218
rect 392808 398898 392850 399134
rect 393086 398898 393128 399134
rect 392808 398866 393128 398898
rect 254568 381454 254888 381486
rect 254568 381218 254610 381454
rect 254846 381218 254888 381454
rect 254568 381134 254888 381218
rect 254568 380898 254610 381134
rect 254846 380898 254888 381134
rect 254568 380866 254888 380898
rect 285288 381454 285608 381486
rect 285288 381218 285330 381454
rect 285566 381218 285608 381454
rect 285288 381134 285608 381218
rect 285288 380898 285330 381134
rect 285566 380898 285608 381134
rect 285288 380866 285608 380898
rect 316008 381454 316328 381486
rect 316008 381218 316050 381454
rect 316286 381218 316328 381454
rect 316008 381134 316328 381218
rect 316008 380898 316050 381134
rect 316286 380898 316328 381134
rect 316008 380866 316328 380898
rect 346728 381454 347048 381486
rect 346728 381218 346770 381454
rect 347006 381218 347048 381454
rect 346728 381134 347048 381218
rect 346728 380898 346770 381134
rect 347006 380898 347048 381134
rect 346728 380866 347048 380898
rect 377448 381454 377768 381486
rect 377448 381218 377490 381454
rect 377726 381218 377768 381454
rect 377448 381134 377768 381218
rect 377448 380898 377490 381134
rect 377726 380898 377768 381134
rect 377448 380866 377768 380898
rect 408168 381454 408488 381486
rect 408168 381218 408210 381454
rect 408446 381218 408488 381454
rect 408168 381134 408488 381218
rect 408168 380898 408210 381134
rect 408446 380898 408488 381134
rect 408168 380866 408488 380898
rect 239208 363454 239528 363486
rect 239208 363218 239250 363454
rect 239486 363218 239528 363454
rect 239208 363134 239528 363218
rect 239208 362898 239250 363134
rect 239486 362898 239528 363134
rect 239208 362866 239528 362898
rect 269928 363454 270248 363486
rect 269928 363218 269970 363454
rect 270206 363218 270248 363454
rect 269928 363134 270248 363218
rect 269928 362898 269970 363134
rect 270206 362898 270248 363134
rect 269928 362866 270248 362898
rect 300648 363454 300968 363486
rect 300648 363218 300690 363454
rect 300926 363218 300968 363454
rect 300648 363134 300968 363218
rect 300648 362898 300690 363134
rect 300926 362898 300968 363134
rect 300648 362866 300968 362898
rect 331368 363454 331688 363486
rect 331368 363218 331410 363454
rect 331646 363218 331688 363454
rect 331368 363134 331688 363218
rect 331368 362898 331410 363134
rect 331646 362898 331688 363134
rect 331368 362866 331688 362898
rect 362088 363454 362408 363486
rect 362088 363218 362130 363454
rect 362366 363218 362408 363454
rect 362088 363134 362408 363218
rect 362088 362898 362130 363134
rect 362366 362898 362408 363134
rect 362088 362866 362408 362898
rect 392808 363454 393128 363486
rect 392808 363218 392850 363454
rect 393086 363218 393128 363454
rect 392808 363134 393128 363218
rect 392808 362898 392850 363134
rect 393086 362898 393128 363134
rect 392808 362866 393128 362898
rect 254568 345454 254888 345486
rect 254568 345218 254610 345454
rect 254846 345218 254888 345454
rect 254568 345134 254888 345218
rect 254568 344898 254610 345134
rect 254846 344898 254888 345134
rect 254568 344866 254888 344898
rect 285288 345454 285608 345486
rect 285288 345218 285330 345454
rect 285566 345218 285608 345454
rect 285288 345134 285608 345218
rect 285288 344898 285330 345134
rect 285566 344898 285608 345134
rect 285288 344866 285608 344898
rect 316008 345454 316328 345486
rect 316008 345218 316050 345454
rect 316286 345218 316328 345454
rect 316008 345134 316328 345218
rect 316008 344898 316050 345134
rect 316286 344898 316328 345134
rect 316008 344866 316328 344898
rect 346728 345454 347048 345486
rect 346728 345218 346770 345454
rect 347006 345218 347048 345454
rect 346728 345134 347048 345218
rect 346728 344898 346770 345134
rect 347006 344898 347048 345134
rect 346728 344866 347048 344898
rect 377448 345454 377768 345486
rect 377448 345218 377490 345454
rect 377726 345218 377768 345454
rect 377448 345134 377768 345218
rect 377448 344898 377490 345134
rect 377726 344898 377768 345134
rect 377448 344866 377768 344898
rect 408168 345454 408488 345486
rect 408168 345218 408210 345454
rect 408446 345218 408488 345454
rect 408168 345134 408488 345218
rect 408168 344898 408210 345134
rect 408446 344898 408488 345134
rect 408168 344866 408488 344898
rect 235794 309454 236414 336000
rect 235794 308898 235826 309454
rect 236382 308898 236414 309454
rect 235794 273454 236414 308898
rect 235794 272898 235826 273454
rect 236382 272898 236414 273454
rect 235794 237454 236414 272898
rect 235794 236898 235826 237454
rect 236382 236898 236414 237454
rect 235794 201454 236414 236898
rect 235794 200898 235826 201454
rect 236382 200898 236414 201454
rect 235794 165454 236414 200898
rect 235794 164898 235826 165454
rect 236382 164898 236414 165454
rect 235794 129454 236414 164898
rect 235794 128898 235826 129454
rect 236382 128898 236414 129454
rect 235794 93454 236414 128898
rect 235794 92898 235826 93454
rect 236382 92898 236414 93454
rect 235794 57454 236414 92898
rect 235794 56898 235826 57454
rect 236382 56898 236414 57454
rect 233739 44300 233805 44301
rect 233739 44236 233740 44300
rect 233804 44236 233805 44300
rect 233739 44235 233805 44236
rect 228954 14058 228986 14614
rect 229542 14058 229574 14614
rect 210954 -7622 210986 -7066
rect 211542 -7622 211574 -7066
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 21454 236414 56898
rect 235794 20898 235826 21454
rect 236382 20898 236414 21454
rect 235794 -1306 236414 20898
rect 235794 -1862 235826 -1306
rect 236382 -1862 236414 -1306
rect 235794 -1894 236414 -1862
rect 239514 313174 240134 336000
rect 239514 312618 239546 313174
rect 240102 312618 240134 313174
rect 239514 277174 240134 312618
rect 239514 276618 239546 277174
rect 240102 276618 240134 277174
rect 239514 241174 240134 276618
rect 239514 240618 239546 241174
rect 240102 240618 240134 241174
rect 239514 205174 240134 240618
rect 239514 204618 239546 205174
rect 240102 204618 240134 205174
rect 239514 169174 240134 204618
rect 239514 168618 239546 169174
rect 240102 168618 240134 169174
rect 239514 133174 240134 168618
rect 239514 132618 239546 133174
rect 240102 132618 240134 133174
rect 239514 97174 240134 132618
rect 239514 96618 239546 97174
rect 240102 96618 240134 97174
rect 239514 61174 240134 96618
rect 239514 60618 239546 61174
rect 240102 60618 240134 61174
rect 239514 25174 240134 60618
rect 239514 24618 239546 25174
rect 240102 24618 240134 25174
rect 239514 -3226 240134 24618
rect 239514 -3782 239546 -3226
rect 240102 -3782 240134 -3226
rect 239514 -3814 240134 -3782
rect 243234 316894 243854 336000
rect 243234 316338 243266 316894
rect 243822 316338 243854 316894
rect 243234 280894 243854 316338
rect 243234 280338 243266 280894
rect 243822 280338 243854 280894
rect 243234 244894 243854 280338
rect 243234 244338 243266 244894
rect 243822 244338 243854 244894
rect 243234 208894 243854 244338
rect 243234 208338 243266 208894
rect 243822 208338 243854 208894
rect 243234 172894 243854 208338
rect 243234 172338 243266 172894
rect 243822 172338 243854 172894
rect 243234 136894 243854 172338
rect 243234 136338 243266 136894
rect 243822 136338 243854 136894
rect 243234 100894 243854 136338
rect 243234 100338 243266 100894
rect 243822 100338 243854 100894
rect 243234 64894 243854 100338
rect 243234 64338 243266 64894
rect 243822 64338 243854 64894
rect 243234 28894 243854 64338
rect 243234 28338 243266 28894
rect 243822 28338 243854 28894
rect 243234 -5146 243854 28338
rect 243234 -5702 243266 -5146
rect 243822 -5702 243854 -5146
rect 243234 -5734 243854 -5702
rect 246954 320614 247574 336000
rect 246954 320058 246986 320614
rect 247542 320058 247574 320614
rect 246954 284614 247574 320058
rect 246954 284058 246986 284614
rect 247542 284058 247574 284614
rect 246954 248614 247574 284058
rect 246954 248058 246986 248614
rect 247542 248058 247574 248614
rect 246954 212614 247574 248058
rect 246954 212058 246986 212614
rect 247542 212058 247574 212614
rect 246954 176614 247574 212058
rect 246954 176058 246986 176614
rect 247542 176058 247574 176614
rect 246954 140614 247574 176058
rect 246954 140058 246986 140614
rect 247542 140058 247574 140614
rect 246954 104614 247574 140058
rect 246954 104058 246986 104614
rect 247542 104058 247574 104614
rect 246954 68614 247574 104058
rect 246954 68058 246986 68614
rect 247542 68058 247574 68614
rect 246954 32614 247574 68058
rect 246954 32058 246986 32614
rect 247542 32058 247574 32614
rect 228954 -6662 228986 -6106
rect 229542 -6662 229574 -6106
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 327454 254414 336000
rect 253794 326898 253826 327454
rect 254382 326898 254414 327454
rect 253794 291454 254414 326898
rect 253794 290898 253826 291454
rect 254382 290898 254414 291454
rect 253794 255454 254414 290898
rect 253794 254898 253826 255454
rect 254382 254898 254414 255454
rect 253794 219454 254414 254898
rect 253794 218898 253826 219454
rect 254382 218898 254414 219454
rect 253794 183454 254414 218898
rect 253794 182898 253826 183454
rect 254382 182898 254414 183454
rect 253794 147454 254414 182898
rect 253794 146898 253826 147454
rect 254382 146898 254414 147454
rect 253794 111454 254414 146898
rect 253794 110898 253826 111454
rect 254382 110898 254414 111454
rect 253794 75454 254414 110898
rect 253794 74898 253826 75454
rect 254382 74898 254414 75454
rect 253794 39454 254414 74898
rect 253794 38898 253826 39454
rect 254382 38898 254414 39454
rect 253794 3454 254414 38898
rect 253794 2898 253826 3454
rect 254382 2898 254414 3454
rect 253794 -346 254414 2898
rect 253794 -902 253826 -346
rect 254382 -902 254414 -346
rect 253794 -1894 254414 -902
rect 257514 331174 258134 336000
rect 257514 330618 257546 331174
rect 258102 330618 258134 331174
rect 257514 295174 258134 330618
rect 257514 294618 257546 295174
rect 258102 294618 258134 295174
rect 257514 259174 258134 294618
rect 257514 258618 257546 259174
rect 258102 258618 258134 259174
rect 257514 223174 258134 258618
rect 257514 222618 257546 223174
rect 258102 222618 258134 223174
rect 257514 187174 258134 222618
rect 257514 186618 257546 187174
rect 258102 186618 258134 187174
rect 257514 151174 258134 186618
rect 257514 150618 257546 151174
rect 258102 150618 258134 151174
rect 257514 115174 258134 150618
rect 257514 114618 257546 115174
rect 258102 114618 258134 115174
rect 257514 79174 258134 114618
rect 257514 78618 257546 79174
rect 258102 78618 258134 79174
rect 257514 43174 258134 78618
rect 257514 42618 257546 43174
rect 258102 42618 258134 43174
rect 257514 7174 258134 42618
rect 257514 6618 257546 7174
rect 258102 6618 258134 7174
rect 257514 -2266 258134 6618
rect 257514 -2822 257546 -2266
rect 258102 -2822 258134 -2266
rect 257514 -3814 258134 -2822
rect 261234 334894 261854 336000
rect 261234 334338 261266 334894
rect 261822 334338 261854 334894
rect 261234 298894 261854 334338
rect 261234 298338 261266 298894
rect 261822 298338 261854 298894
rect 261234 262894 261854 298338
rect 261234 262338 261266 262894
rect 261822 262338 261854 262894
rect 261234 226894 261854 262338
rect 261234 226338 261266 226894
rect 261822 226338 261854 226894
rect 261234 190894 261854 226338
rect 261234 190338 261266 190894
rect 261822 190338 261854 190894
rect 261234 154894 261854 190338
rect 261234 154338 261266 154894
rect 261822 154338 261854 154894
rect 261234 118894 261854 154338
rect 261234 118338 261266 118894
rect 261822 118338 261854 118894
rect 261234 82894 261854 118338
rect 261234 82338 261266 82894
rect 261822 82338 261854 82894
rect 261234 46894 261854 82338
rect 261234 46338 261266 46894
rect 261822 46338 261854 46894
rect 261234 10894 261854 46338
rect 261234 10338 261266 10894
rect 261822 10338 261854 10894
rect 261234 -4186 261854 10338
rect 261234 -4742 261266 -4186
rect 261822 -4742 261854 -4186
rect 261234 -5734 261854 -4742
rect 264954 302614 265574 336000
rect 264954 302058 264986 302614
rect 265542 302058 265574 302614
rect 264954 266614 265574 302058
rect 264954 266058 264986 266614
rect 265542 266058 265574 266614
rect 264954 230614 265574 266058
rect 264954 230058 264986 230614
rect 265542 230058 265574 230614
rect 264954 194614 265574 230058
rect 264954 194058 264986 194614
rect 265542 194058 265574 194614
rect 264954 158614 265574 194058
rect 264954 158058 264986 158614
rect 265542 158058 265574 158614
rect 264954 122614 265574 158058
rect 264954 122058 264986 122614
rect 265542 122058 265574 122614
rect 264954 86614 265574 122058
rect 264954 86058 264986 86614
rect 265542 86058 265574 86614
rect 264954 50614 265574 86058
rect 264954 50058 264986 50614
rect 265542 50058 265574 50614
rect 264954 14614 265574 50058
rect 264954 14058 264986 14614
rect 265542 14058 265574 14614
rect 246954 -7622 246986 -7066
rect 247542 -7622 247574 -7066
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 309454 272414 336000
rect 271794 308898 271826 309454
rect 272382 308898 272414 309454
rect 271794 273454 272414 308898
rect 271794 272898 271826 273454
rect 272382 272898 272414 273454
rect 271794 237454 272414 272898
rect 271794 236898 271826 237454
rect 272382 236898 272414 237454
rect 271794 201454 272414 236898
rect 271794 200898 271826 201454
rect 272382 200898 272414 201454
rect 271794 165454 272414 200898
rect 271794 164898 271826 165454
rect 272382 164898 272414 165454
rect 271794 129454 272414 164898
rect 271794 128898 271826 129454
rect 272382 128898 272414 129454
rect 271794 93454 272414 128898
rect 271794 92898 271826 93454
rect 272382 92898 272414 93454
rect 271794 57454 272414 92898
rect 271794 56898 271826 57454
rect 272382 56898 272414 57454
rect 271794 21454 272414 56898
rect 271794 20898 271826 21454
rect 272382 20898 272414 21454
rect 271794 -1306 272414 20898
rect 271794 -1862 271826 -1306
rect 272382 -1862 272414 -1306
rect 271794 -1894 272414 -1862
rect 275514 313174 276134 336000
rect 275514 312618 275546 313174
rect 276102 312618 276134 313174
rect 275514 277174 276134 312618
rect 275514 276618 275546 277174
rect 276102 276618 276134 277174
rect 275514 241174 276134 276618
rect 275514 240618 275546 241174
rect 276102 240618 276134 241174
rect 275514 205174 276134 240618
rect 275514 204618 275546 205174
rect 276102 204618 276134 205174
rect 275514 169174 276134 204618
rect 275514 168618 275546 169174
rect 276102 168618 276134 169174
rect 275514 133174 276134 168618
rect 275514 132618 275546 133174
rect 276102 132618 276134 133174
rect 275514 97174 276134 132618
rect 275514 96618 275546 97174
rect 276102 96618 276134 97174
rect 275514 61174 276134 96618
rect 275514 60618 275546 61174
rect 276102 60618 276134 61174
rect 275514 25174 276134 60618
rect 275514 24618 275546 25174
rect 276102 24618 276134 25174
rect 275514 -3226 276134 24618
rect 275514 -3782 275546 -3226
rect 276102 -3782 276134 -3226
rect 275514 -3814 276134 -3782
rect 279234 316894 279854 336000
rect 279234 316338 279266 316894
rect 279822 316338 279854 316894
rect 279234 280894 279854 316338
rect 279234 280338 279266 280894
rect 279822 280338 279854 280894
rect 279234 244894 279854 280338
rect 279234 244338 279266 244894
rect 279822 244338 279854 244894
rect 279234 208894 279854 244338
rect 279234 208338 279266 208894
rect 279822 208338 279854 208894
rect 279234 172894 279854 208338
rect 279234 172338 279266 172894
rect 279822 172338 279854 172894
rect 279234 136894 279854 172338
rect 279234 136338 279266 136894
rect 279822 136338 279854 136894
rect 279234 100894 279854 136338
rect 279234 100338 279266 100894
rect 279822 100338 279854 100894
rect 279234 64894 279854 100338
rect 279234 64338 279266 64894
rect 279822 64338 279854 64894
rect 279234 28894 279854 64338
rect 279234 28338 279266 28894
rect 279822 28338 279854 28894
rect 279234 -5146 279854 28338
rect 279234 -5702 279266 -5146
rect 279822 -5702 279854 -5146
rect 279234 -5734 279854 -5702
rect 282954 320614 283574 336000
rect 282954 320058 282986 320614
rect 283542 320058 283574 320614
rect 282954 284614 283574 320058
rect 282954 284058 282986 284614
rect 283542 284058 283574 284614
rect 282954 248614 283574 284058
rect 282954 248058 282986 248614
rect 283542 248058 283574 248614
rect 282954 212614 283574 248058
rect 282954 212058 282986 212614
rect 283542 212058 283574 212614
rect 282954 176614 283574 212058
rect 282954 176058 282986 176614
rect 283542 176058 283574 176614
rect 282954 140614 283574 176058
rect 282954 140058 282986 140614
rect 283542 140058 283574 140614
rect 282954 104614 283574 140058
rect 282954 104058 282986 104614
rect 283542 104058 283574 104614
rect 282954 68614 283574 104058
rect 282954 68058 282986 68614
rect 283542 68058 283574 68614
rect 282954 32614 283574 68058
rect 282954 32058 282986 32614
rect 283542 32058 283574 32614
rect 264954 -6662 264986 -6106
rect 265542 -6662 265574 -6106
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 327454 290414 336000
rect 289794 326898 289826 327454
rect 290382 326898 290414 327454
rect 289794 291454 290414 326898
rect 289794 290898 289826 291454
rect 290382 290898 290414 291454
rect 289794 255454 290414 290898
rect 289794 254898 289826 255454
rect 290382 254898 290414 255454
rect 289794 219454 290414 254898
rect 289794 218898 289826 219454
rect 290382 218898 290414 219454
rect 289794 183454 290414 218898
rect 289794 182898 289826 183454
rect 290382 182898 290414 183454
rect 289794 147454 290414 182898
rect 289794 146898 289826 147454
rect 290382 146898 290414 147454
rect 289794 111454 290414 146898
rect 289794 110898 289826 111454
rect 290382 110898 290414 111454
rect 289794 75454 290414 110898
rect 289794 74898 289826 75454
rect 290382 74898 290414 75454
rect 289794 39454 290414 74898
rect 289794 38898 289826 39454
rect 290382 38898 290414 39454
rect 289794 3454 290414 38898
rect 289794 2898 289826 3454
rect 290382 2898 290414 3454
rect 289794 -346 290414 2898
rect 289794 -902 289826 -346
rect 290382 -902 290414 -346
rect 289794 -1894 290414 -902
rect 293514 331174 294134 336000
rect 293514 330618 293546 331174
rect 294102 330618 294134 331174
rect 293514 295174 294134 330618
rect 293514 294618 293546 295174
rect 294102 294618 294134 295174
rect 293514 259174 294134 294618
rect 293514 258618 293546 259174
rect 294102 258618 294134 259174
rect 293514 223174 294134 258618
rect 293514 222618 293546 223174
rect 294102 222618 294134 223174
rect 293514 187174 294134 222618
rect 293514 186618 293546 187174
rect 294102 186618 294134 187174
rect 293514 151174 294134 186618
rect 293514 150618 293546 151174
rect 294102 150618 294134 151174
rect 293514 115174 294134 150618
rect 293514 114618 293546 115174
rect 294102 114618 294134 115174
rect 293514 79174 294134 114618
rect 293514 78618 293546 79174
rect 294102 78618 294134 79174
rect 293514 43174 294134 78618
rect 293514 42618 293546 43174
rect 294102 42618 294134 43174
rect 293514 7174 294134 42618
rect 293514 6618 293546 7174
rect 294102 6618 294134 7174
rect 293514 -2266 294134 6618
rect 293514 -2822 293546 -2266
rect 294102 -2822 294134 -2266
rect 293514 -3814 294134 -2822
rect 297234 334894 297854 336000
rect 297234 334338 297266 334894
rect 297822 334338 297854 334894
rect 297234 298894 297854 334338
rect 297234 298338 297266 298894
rect 297822 298338 297854 298894
rect 297234 262894 297854 298338
rect 297234 262338 297266 262894
rect 297822 262338 297854 262894
rect 297234 226894 297854 262338
rect 297234 226338 297266 226894
rect 297822 226338 297854 226894
rect 297234 190894 297854 226338
rect 297234 190338 297266 190894
rect 297822 190338 297854 190894
rect 297234 154894 297854 190338
rect 297234 154338 297266 154894
rect 297822 154338 297854 154894
rect 297234 118894 297854 154338
rect 297234 118338 297266 118894
rect 297822 118338 297854 118894
rect 297234 82894 297854 118338
rect 297234 82338 297266 82894
rect 297822 82338 297854 82894
rect 297234 46894 297854 82338
rect 297234 46338 297266 46894
rect 297822 46338 297854 46894
rect 297234 10894 297854 46338
rect 297234 10338 297266 10894
rect 297822 10338 297854 10894
rect 297234 -4186 297854 10338
rect 297234 -4742 297266 -4186
rect 297822 -4742 297854 -4186
rect 297234 -5734 297854 -4742
rect 300954 302614 301574 336000
rect 300954 302058 300986 302614
rect 301542 302058 301574 302614
rect 300954 266614 301574 302058
rect 300954 266058 300986 266614
rect 301542 266058 301574 266614
rect 300954 230614 301574 266058
rect 300954 230058 300986 230614
rect 301542 230058 301574 230614
rect 300954 194614 301574 230058
rect 300954 194058 300986 194614
rect 301542 194058 301574 194614
rect 300954 158614 301574 194058
rect 300954 158058 300986 158614
rect 301542 158058 301574 158614
rect 300954 122614 301574 158058
rect 300954 122058 300986 122614
rect 301542 122058 301574 122614
rect 300954 86614 301574 122058
rect 300954 86058 300986 86614
rect 301542 86058 301574 86614
rect 300954 50614 301574 86058
rect 300954 50058 300986 50614
rect 301542 50058 301574 50614
rect 300954 14614 301574 50058
rect 300954 14058 300986 14614
rect 301542 14058 301574 14614
rect 282954 -7622 282986 -7066
rect 283542 -7622 283574 -7066
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 309454 308414 336000
rect 307794 308898 307826 309454
rect 308382 308898 308414 309454
rect 307794 273454 308414 308898
rect 307794 272898 307826 273454
rect 308382 272898 308414 273454
rect 307794 237454 308414 272898
rect 307794 236898 307826 237454
rect 308382 236898 308414 237454
rect 307794 201454 308414 236898
rect 307794 200898 307826 201454
rect 308382 200898 308414 201454
rect 307794 165454 308414 200898
rect 307794 164898 307826 165454
rect 308382 164898 308414 165454
rect 307794 129454 308414 164898
rect 307794 128898 307826 129454
rect 308382 128898 308414 129454
rect 307794 93454 308414 128898
rect 307794 92898 307826 93454
rect 308382 92898 308414 93454
rect 307794 57454 308414 92898
rect 307794 56898 307826 57454
rect 308382 56898 308414 57454
rect 307794 21454 308414 56898
rect 307794 20898 307826 21454
rect 308382 20898 308414 21454
rect 307794 -1306 308414 20898
rect 307794 -1862 307826 -1306
rect 308382 -1862 308414 -1306
rect 307794 -1894 308414 -1862
rect 311514 313174 312134 336000
rect 311514 312618 311546 313174
rect 312102 312618 312134 313174
rect 311514 277174 312134 312618
rect 311514 276618 311546 277174
rect 312102 276618 312134 277174
rect 311514 241174 312134 276618
rect 311514 240618 311546 241174
rect 312102 240618 312134 241174
rect 311514 205174 312134 240618
rect 311514 204618 311546 205174
rect 312102 204618 312134 205174
rect 311514 169174 312134 204618
rect 311514 168618 311546 169174
rect 312102 168618 312134 169174
rect 311514 133174 312134 168618
rect 311514 132618 311546 133174
rect 312102 132618 312134 133174
rect 311514 97174 312134 132618
rect 311514 96618 311546 97174
rect 312102 96618 312134 97174
rect 311514 61174 312134 96618
rect 311514 60618 311546 61174
rect 312102 60618 312134 61174
rect 311514 25174 312134 60618
rect 311514 24618 311546 25174
rect 312102 24618 312134 25174
rect 311514 -3226 312134 24618
rect 311514 -3782 311546 -3226
rect 312102 -3782 312134 -3226
rect 311514 -3814 312134 -3782
rect 315234 316894 315854 336000
rect 315234 316338 315266 316894
rect 315822 316338 315854 316894
rect 315234 280894 315854 316338
rect 315234 280338 315266 280894
rect 315822 280338 315854 280894
rect 315234 244894 315854 280338
rect 315234 244338 315266 244894
rect 315822 244338 315854 244894
rect 315234 208894 315854 244338
rect 315234 208338 315266 208894
rect 315822 208338 315854 208894
rect 315234 172894 315854 208338
rect 315234 172338 315266 172894
rect 315822 172338 315854 172894
rect 315234 136894 315854 172338
rect 315234 136338 315266 136894
rect 315822 136338 315854 136894
rect 315234 100894 315854 136338
rect 315234 100338 315266 100894
rect 315822 100338 315854 100894
rect 315234 64894 315854 100338
rect 315234 64338 315266 64894
rect 315822 64338 315854 64894
rect 315234 28894 315854 64338
rect 315234 28338 315266 28894
rect 315822 28338 315854 28894
rect 315234 -5146 315854 28338
rect 315234 -5702 315266 -5146
rect 315822 -5702 315854 -5146
rect 315234 -5734 315854 -5702
rect 318954 320614 319574 336000
rect 318954 320058 318986 320614
rect 319542 320058 319574 320614
rect 318954 284614 319574 320058
rect 318954 284058 318986 284614
rect 319542 284058 319574 284614
rect 318954 248614 319574 284058
rect 318954 248058 318986 248614
rect 319542 248058 319574 248614
rect 318954 212614 319574 248058
rect 318954 212058 318986 212614
rect 319542 212058 319574 212614
rect 318954 176614 319574 212058
rect 318954 176058 318986 176614
rect 319542 176058 319574 176614
rect 318954 140614 319574 176058
rect 318954 140058 318986 140614
rect 319542 140058 319574 140614
rect 318954 104614 319574 140058
rect 318954 104058 318986 104614
rect 319542 104058 319574 104614
rect 318954 68614 319574 104058
rect 318954 68058 318986 68614
rect 319542 68058 319574 68614
rect 318954 32614 319574 68058
rect 318954 32058 318986 32614
rect 319542 32058 319574 32614
rect 300954 -6662 300986 -6106
rect 301542 -6662 301574 -6106
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 327454 326414 336000
rect 325794 326898 325826 327454
rect 326382 326898 326414 327454
rect 325794 291454 326414 326898
rect 325794 290898 325826 291454
rect 326382 290898 326414 291454
rect 325794 255454 326414 290898
rect 325794 254898 325826 255454
rect 326382 254898 326414 255454
rect 325794 219454 326414 254898
rect 325794 218898 325826 219454
rect 326382 218898 326414 219454
rect 325794 183454 326414 218898
rect 325794 182898 325826 183454
rect 326382 182898 326414 183454
rect 325794 147454 326414 182898
rect 325794 146898 325826 147454
rect 326382 146898 326414 147454
rect 325794 111454 326414 146898
rect 325794 110898 325826 111454
rect 326382 110898 326414 111454
rect 325794 75454 326414 110898
rect 325794 74898 325826 75454
rect 326382 74898 326414 75454
rect 325794 39454 326414 74898
rect 325794 38898 325826 39454
rect 326382 38898 326414 39454
rect 325794 3454 326414 38898
rect 325794 2898 325826 3454
rect 326382 2898 326414 3454
rect 325794 -346 326414 2898
rect 325794 -902 325826 -346
rect 326382 -902 326414 -346
rect 325794 -1894 326414 -902
rect 329514 331174 330134 336000
rect 329514 330618 329546 331174
rect 330102 330618 330134 331174
rect 329514 295174 330134 330618
rect 329514 294618 329546 295174
rect 330102 294618 330134 295174
rect 329514 259174 330134 294618
rect 329514 258618 329546 259174
rect 330102 258618 330134 259174
rect 329514 223174 330134 258618
rect 329514 222618 329546 223174
rect 330102 222618 330134 223174
rect 329514 187174 330134 222618
rect 329514 186618 329546 187174
rect 330102 186618 330134 187174
rect 329514 151174 330134 186618
rect 329514 150618 329546 151174
rect 330102 150618 330134 151174
rect 329514 115174 330134 150618
rect 329514 114618 329546 115174
rect 330102 114618 330134 115174
rect 329514 79174 330134 114618
rect 329514 78618 329546 79174
rect 330102 78618 330134 79174
rect 329514 43174 330134 78618
rect 329514 42618 329546 43174
rect 330102 42618 330134 43174
rect 329514 7174 330134 42618
rect 329514 6618 329546 7174
rect 330102 6618 330134 7174
rect 329514 -2266 330134 6618
rect 329514 -2822 329546 -2266
rect 330102 -2822 330134 -2266
rect 329514 -3814 330134 -2822
rect 333234 334894 333854 336000
rect 333234 334338 333266 334894
rect 333822 334338 333854 334894
rect 333234 298894 333854 334338
rect 333234 298338 333266 298894
rect 333822 298338 333854 298894
rect 333234 262894 333854 298338
rect 333234 262338 333266 262894
rect 333822 262338 333854 262894
rect 333234 226894 333854 262338
rect 333234 226338 333266 226894
rect 333822 226338 333854 226894
rect 333234 190894 333854 226338
rect 333234 190338 333266 190894
rect 333822 190338 333854 190894
rect 333234 154894 333854 190338
rect 333234 154338 333266 154894
rect 333822 154338 333854 154894
rect 333234 118894 333854 154338
rect 333234 118338 333266 118894
rect 333822 118338 333854 118894
rect 333234 82894 333854 118338
rect 333234 82338 333266 82894
rect 333822 82338 333854 82894
rect 333234 46894 333854 82338
rect 333234 46338 333266 46894
rect 333822 46338 333854 46894
rect 333234 10894 333854 46338
rect 333234 10338 333266 10894
rect 333822 10338 333854 10894
rect 333234 -4186 333854 10338
rect 333234 -4742 333266 -4186
rect 333822 -4742 333854 -4186
rect 333234 -5734 333854 -4742
rect 336954 302614 337574 336000
rect 336954 302058 336986 302614
rect 337542 302058 337574 302614
rect 336954 266614 337574 302058
rect 336954 266058 336986 266614
rect 337542 266058 337574 266614
rect 336954 230614 337574 266058
rect 336954 230058 336986 230614
rect 337542 230058 337574 230614
rect 336954 194614 337574 230058
rect 336954 194058 336986 194614
rect 337542 194058 337574 194614
rect 336954 158614 337574 194058
rect 336954 158058 336986 158614
rect 337542 158058 337574 158614
rect 336954 122614 337574 158058
rect 336954 122058 336986 122614
rect 337542 122058 337574 122614
rect 336954 86614 337574 122058
rect 336954 86058 336986 86614
rect 337542 86058 337574 86614
rect 336954 50614 337574 86058
rect 336954 50058 336986 50614
rect 337542 50058 337574 50614
rect 336954 14614 337574 50058
rect 336954 14058 336986 14614
rect 337542 14058 337574 14614
rect 318954 -7622 318986 -7066
rect 319542 -7622 319574 -7066
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 309454 344414 336000
rect 343794 308898 343826 309454
rect 344382 308898 344414 309454
rect 343794 273454 344414 308898
rect 343794 272898 343826 273454
rect 344382 272898 344414 273454
rect 343794 237454 344414 272898
rect 343794 236898 343826 237454
rect 344382 236898 344414 237454
rect 343794 201454 344414 236898
rect 343794 200898 343826 201454
rect 344382 200898 344414 201454
rect 343794 165454 344414 200898
rect 343794 164898 343826 165454
rect 344382 164898 344414 165454
rect 343794 129454 344414 164898
rect 343794 128898 343826 129454
rect 344382 128898 344414 129454
rect 343794 93454 344414 128898
rect 343794 92898 343826 93454
rect 344382 92898 344414 93454
rect 343794 57454 344414 92898
rect 343794 56898 343826 57454
rect 344382 56898 344414 57454
rect 343794 21454 344414 56898
rect 343794 20898 343826 21454
rect 344382 20898 344414 21454
rect 343794 -1306 344414 20898
rect 343794 -1862 343826 -1306
rect 344382 -1862 344414 -1306
rect 343794 -1894 344414 -1862
rect 347514 313174 348134 336000
rect 347514 312618 347546 313174
rect 348102 312618 348134 313174
rect 347514 277174 348134 312618
rect 347514 276618 347546 277174
rect 348102 276618 348134 277174
rect 347514 241174 348134 276618
rect 347514 240618 347546 241174
rect 348102 240618 348134 241174
rect 347514 205174 348134 240618
rect 347514 204618 347546 205174
rect 348102 204618 348134 205174
rect 347514 169174 348134 204618
rect 347514 168618 347546 169174
rect 348102 168618 348134 169174
rect 347514 133174 348134 168618
rect 347514 132618 347546 133174
rect 348102 132618 348134 133174
rect 347514 97174 348134 132618
rect 347514 96618 347546 97174
rect 348102 96618 348134 97174
rect 347514 61174 348134 96618
rect 347514 60618 347546 61174
rect 348102 60618 348134 61174
rect 347514 25174 348134 60618
rect 347514 24618 347546 25174
rect 348102 24618 348134 25174
rect 347514 -3226 348134 24618
rect 347514 -3782 347546 -3226
rect 348102 -3782 348134 -3226
rect 347514 -3814 348134 -3782
rect 351234 316894 351854 336000
rect 351234 316338 351266 316894
rect 351822 316338 351854 316894
rect 351234 280894 351854 316338
rect 351234 280338 351266 280894
rect 351822 280338 351854 280894
rect 351234 244894 351854 280338
rect 351234 244338 351266 244894
rect 351822 244338 351854 244894
rect 351234 208894 351854 244338
rect 351234 208338 351266 208894
rect 351822 208338 351854 208894
rect 351234 172894 351854 208338
rect 351234 172338 351266 172894
rect 351822 172338 351854 172894
rect 351234 136894 351854 172338
rect 351234 136338 351266 136894
rect 351822 136338 351854 136894
rect 351234 100894 351854 136338
rect 351234 100338 351266 100894
rect 351822 100338 351854 100894
rect 351234 64894 351854 100338
rect 351234 64338 351266 64894
rect 351822 64338 351854 64894
rect 351234 28894 351854 64338
rect 351234 28338 351266 28894
rect 351822 28338 351854 28894
rect 351234 -5146 351854 28338
rect 351234 -5702 351266 -5146
rect 351822 -5702 351854 -5146
rect 351234 -5734 351854 -5702
rect 354954 320614 355574 336000
rect 354954 320058 354986 320614
rect 355542 320058 355574 320614
rect 354954 284614 355574 320058
rect 354954 284058 354986 284614
rect 355542 284058 355574 284614
rect 354954 248614 355574 284058
rect 354954 248058 354986 248614
rect 355542 248058 355574 248614
rect 354954 212614 355574 248058
rect 354954 212058 354986 212614
rect 355542 212058 355574 212614
rect 354954 176614 355574 212058
rect 354954 176058 354986 176614
rect 355542 176058 355574 176614
rect 354954 140614 355574 176058
rect 354954 140058 354986 140614
rect 355542 140058 355574 140614
rect 354954 104614 355574 140058
rect 354954 104058 354986 104614
rect 355542 104058 355574 104614
rect 354954 68614 355574 104058
rect 354954 68058 354986 68614
rect 355542 68058 355574 68614
rect 354954 32614 355574 68058
rect 354954 32058 354986 32614
rect 355542 32058 355574 32614
rect 336954 -6662 336986 -6106
rect 337542 -6662 337574 -6106
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 327454 362414 336000
rect 361794 326898 361826 327454
rect 362382 326898 362414 327454
rect 361794 291454 362414 326898
rect 361794 290898 361826 291454
rect 362382 290898 362414 291454
rect 361794 255454 362414 290898
rect 361794 254898 361826 255454
rect 362382 254898 362414 255454
rect 361794 219454 362414 254898
rect 361794 218898 361826 219454
rect 362382 218898 362414 219454
rect 361794 183454 362414 218898
rect 361794 182898 361826 183454
rect 362382 182898 362414 183454
rect 361794 147454 362414 182898
rect 361794 146898 361826 147454
rect 362382 146898 362414 147454
rect 361794 111454 362414 146898
rect 361794 110898 361826 111454
rect 362382 110898 362414 111454
rect 361794 75454 362414 110898
rect 361794 74898 361826 75454
rect 362382 74898 362414 75454
rect 361794 39454 362414 74898
rect 361794 38898 361826 39454
rect 362382 38898 362414 39454
rect 361794 3454 362414 38898
rect 361794 2898 361826 3454
rect 362382 2898 362414 3454
rect 361794 -346 362414 2898
rect 361794 -902 361826 -346
rect 362382 -902 362414 -346
rect 361794 -1894 362414 -902
rect 365514 331174 366134 336000
rect 365514 330618 365546 331174
rect 366102 330618 366134 331174
rect 365514 295174 366134 330618
rect 365514 294618 365546 295174
rect 366102 294618 366134 295174
rect 365514 259174 366134 294618
rect 365514 258618 365546 259174
rect 366102 258618 366134 259174
rect 365514 223174 366134 258618
rect 365514 222618 365546 223174
rect 366102 222618 366134 223174
rect 365514 187174 366134 222618
rect 365514 186618 365546 187174
rect 366102 186618 366134 187174
rect 365514 151174 366134 186618
rect 365514 150618 365546 151174
rect 366102 150618 366134 151174
rect 365514 115174 366134 150618
rect 365514 114618 365546 115174
rect 366102 114618 366134 115174
rect 365514 79174 366134 114618
rect 365514 78618 365546 79174
rect 366102 78618 366134 79174
rect 365514 43174 366134 78618
rect 365514 42618 365546 43174
rect 366102 42618 366134 43174
rect 365514 7174 366134 42618
rect 365514 6618 365546 7174
rect 366102 6618 366134 7174
rect 365514 -2266 366134 6618
rect 365514 -2822 365546 -2266
rect 366102 -2822 366134 -2266
rect 365514 -3814 366134 -2822
rect 369234 334894 369854 336000
rect 369234 334338 369266 334894
rect 369822 334338 369854 334894
rect 369234 298894 369854 334338
rect 369234 298338 369266 298894
rect 369822 298338 369854 298894
rect 369234 262894 369854 298338
rect 369234 262338 369266 262894
rect 369822 262338 369854 262894
rect 369234 226894 369854 262338
rect 369234 226338 369266 226894
rect 369822 226338 369854 226894
rect 369234 190894 369854 226338
rect 369234 190338 369266 190894
rect 369822 190338 369854 190894
rect 369234 154894 369854 190338
rect 369234 154338 369266 154894
rect 369822 154338 369854 154894
rect 369234 118894 369854 154338
rect 369234 118338 369266 118894
rect 369822 118338 369854 118894
rect 369234 82894 369854 118338
rect 369234 82338 369266 82894
rect 369822 82338 369854 82894
rect 369234 46894 369854 82338
rect 369234 46338 369266 46894
rect 369822 46338 369854 46894
rect 369234 10894 369854 46338
rect 369234 10338 369266 10894
rect 369822 10338 369854 10894
rect 369234 -4186 369854 10338
rect 369234 -4742 369266 -4186
rect 369822 -4742 369854 -4186
rect 369234 -5734 369854 -4742
rect 372954 302614 373574 336000
rect 372954 302058 372986 302614
rect 373542 302058 373574 302614
rect 372954 266614 373574 302058
rect 372954 266058 372986 266614
rect 373542 266058 373574 266614
rect 372954 230614 373574 266058
rect 372954 230058 372986 230614
rect 373542 230058 373574 230614
rect 372954 194614 373574 230058
rect 372954 194058 372986 194614
rect 373542 194058 373574 194614
rect 372954 158614 373574 194058
rect 372954 158058 372986 158614
rect 373542 158058 373574 158614
rect 372954 122614 373574 158058
rect 372954 122058 372986 122614
rect 373542 122058 373574 122614
rect 372954 86614 373574 122058
rect 372954 86058 372986 86614
rect 373542 86058 373574 86614
rect 372954 50614 373574 86058
rect 372954 50058 372986 50614
rect 373542 50058 373574 50614
rect 372954 14614 373574 50058
rect 372954 14058 372986 14614
rect 373542 14058 373574 14614
rect 354954 -7622 354986 -7066
rect 355542 -7622 355574 -7066
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 309454 380414 336000
rect 379794 308898 379826 309454
rect 380382 308898 380414 309454
rect 379794 273454 380414 308898
rect 379794 272898 379826 273454
rect 380382 272898 380414 273454
rect 379794 237454 380414 272898
rect 379794 236898 379826 237454
rect 380382 236898 380414 237454
rect 379794 201454 380414 236898
rect 379794 200898 379826 201454
rect 380382 200898 380414 201454
rect 379794 165454 380414 200898
rect 379794 164898 379826 165454
rect 380382 164898 380414 165454
rect 379794 129454 380414 164898
rect 379794 128898 379826 129454
rect 380382 128898 380414 129454
rect 379794 93454 380414 128898
rect 379794 92898 379826 93454
rect 380382 92898 380414 93454
rect 379794 57454 380414 92898
rect 379794 56898 379826 57454
rect 380382 56898 380414 57454
rect 379794 21454 380414 56898
rect 379794 20898 379826 21454
rect 380382 20898 380414 21454
rect 379794 -1306 380414 20898
rect 379794 -1862 379826 -1306
rect 380382 -1862 380414 -1306
rect 379794 -1894 380414 -1862
rect 383514 313174 384134 336000
rect 383514 312618 383546 313174
rect 384102 312618 384134 313174
rect 383514 277174 384134 312618
rect 383514 276618 383546 277174
rect 384102 276618 384134 277174
rect 383514 241174 384134 276618
rect 383514 240618 383546 241174
rect 384102 240618 384134 241174
rect 383514 205174 384134 240618
rect 383514 204618 383546 205174
rect 384102 204618 384134 205174
rect 383514 169174 384134 204618
rect 383514 168618 383546 169174
rect 384102 168618 384134 169174
rect 383514 133174 384134 168618
rect 383514 132618 383546 133174
rect 384102 132618 384134 133174
rect 383514 97174 384134 132618
rect 383514 96618 383546 97174
rect 384102 96618 384134 97174
rect 383514 61174 384134 96618
rect 383514 60618 383546 61174
rect 384102 60618 384134 61174
rect 383514 25174 384134 60618
rect 383514 24618 383546 25174
rect 384102 24618 384134 25174
rect 383514 -3226 384134 24618
rect 383514 -3782 383546 -3226
rect 384102 -3782 384134 -3226
rect 383514 -3814 384134 -3782
rect 387234 316894 387854 336000
rect 387234 316338 387266 316894
rect 387822 316338 387854 316894
rect 387234 280894 387854 316338
rect 387234 280338 387266 280894
rect 387822 280338 387854 280894
rect 387234 244894 387854 280338
rect 387234 244338 387266 244894
rect 387822 244338 387854 244894
rect 387234 208894 387854 244338
rect 387234 208338 387266 208894
rect 387822 208338 387854 208894
rect 387234 172894 387854 208338
rect 387234 172338 387266 172894
rect 387822 172338 387854 172894
rect 387234 136894 387854 172338
rect 387234 136338 387266 136894
rect 387822 136338 387854 136894
rect 387234 100894 387854 136338
rect 387234 100338 387266 100894
rect 387822 100338 387854 100894
rect 387234 64894 387854 100338
rect 387234 64338 387266 64894
rect 387822 64338 387854 64894
rect 387234 28894 387854 64338
rect 387234 28338 387266 28894
rect 387822 28338 387854 28894
rect 387234 -5146 387854 28338
rect 387234 -5702 387266 -5146
rect 387822 -5702 387854 -5146
rect 387234 -5734 387854 -5702
rect 390954 320614 391574 336000
rect 390954 320058 390986 320614
rect 391542 320058 391574 320614
rect 390954 284614 391574 320058
rect 390954 284058 390986 284614
rect 391542 284058 391574 284614
rect 390954 248614 391574 284058
rect 390954 248058 390986 248614
rect 391542 248058 391574 248614
rect 390954 212614 391574 248058
rect 390954 212058 390986 212614
rect 391542 212058 391574 212614
rect 390954 176614 391574 212058
rect 390954 176058 390986 176614
rect 391542 176058 391574 176614
rect 390954 140614 391574 176058
rect 390954 140058 390986 140614
rect 391542 140058 391574 140614
rect 390954 104614 391574 140058
rect 390954 104058 390986 104614
rect 391542 104058 391574 104614
rect 390954 68614 391574 104058
rect 390954 68058 390986 68614
rect 391542 68058 391574 68614
rect 390954 32614 391574 68058
rect 390954 32058 390986 32614
rect 391542 32058 391574 32614
rect 372954 -6662 372986 -6106
rect 373542 -6662 373574 -6106
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 327454 398414 336000
rect 397794 326898 397826 327454
rect 398382 326898 398414 327454
rect 397794 291454 398414 326898
rect 397794 290898 397826 291454
rect 398382 290898 398414 291454
rect 397794 255454 398414 290898
rect 397794 254898 397826 255454
rect 398382 254898 398414 255454
rect 397794 219454 398414 254898
rect 397794 218898 397826 219454
rect 398382 218898 398414 219454
rect 397794 183454 398414 218898
rect 397794 182898 397826 183454
rect 398382 182898 398414 183454
rect 397794 147454 398414 182898
rect 397794 146898 397826 147454
rect 398382 146898 398414 147454
rect 397794 111454 398414 146898
rect 397794 110898 397826 111454
rect 398382 110898 398414 111454
rect 397794 75454 398414 110898
rect 397794 74898 397826 75454
rect 398382 74898 398414 75454
rect 397794 39454 398414 74898
rect 397794 38898 397826 39454
rect 398382 38898 398414 39454
rect 397794 3454 398414 38898
rect 397794 2898 397826 3454
rect 398382 2898 398414 3454
rect 397794 -346 398414 2898
rect 397794 -902 397826 -346
rect 398382 -902 398414 -346
rect 397794 -1894 398414 -902
rect 401514 331174 402134 336000
rect 401514 330618 401546 331174
rect 402102 330618 402134 331174
rect 401514 295174 402134 330618
rect 401514 294618 401546 295174
rect 402102 294618 402134 295174
rect 401514 259174 402134 294618
rect 401514 258618 401546 259174
rect 402102 258618 402134 259174
rect 401514 223174 402134 258618
rect 401514 222618 401546 223174
rect 402102 222618 402134 223174
rect 401514 187174 402134 222618
rect 401514 186618 401546 187174
rect 402102 186618 402134 187174
rect 401514 151174 402134 186618
rect 401514 150618 401546 151174
rect 402102 150618 402134 151174
rect 401514 115174 402134 150618
rect 401514 114618 401546 115174
rect 402102 114618 402134 115174
rect 401514 79174 402134 114618
rect 401514 78618 401546 79174
rect 402102 78618 402134 79174
rect 401514 43174 402134 78618
rect 401514 42618 401546 43174
rect 402102 42618 402134 43174
rect 401514 7174 402134 42618
rect 401514 6618 401546 7174
rect 402102 6618 402134 7174
rect 401514 -2266 402134 6618
rect 401514 -2822 401546 -2266
rect 402102 -2822 402134 -2266
rect 401514 -3814 402134 -2822
rect 405234 334894 405854 336000
rect 405234 334338 405266 334894
rect 405822 334338 405854 334894
rect 405234 298894 405854 334338
rect 405234 298338 405266 298894
rect 405822 298338 405854 298894
rect 405234 262894 405854 298338
rect 405234 262338 405266 262894
rect 405822 262338 405854 262894
rect 405234 226894 405854 262338
rect 405234 226338 405266 226894
rect 405822 226338 405854 226894
rect 405234 190894 405854 226338
rect 405234 190338 405266 190894
rect 405822 190338 405854 190894
rect 405234 154894 405854 190338
rect 405234 154338 405266 154894
rect 405822 154338 405854 154894
rect 405234 118894 405854 154338
rect 405234 118338 405266 118894
rect 405822 118338 405854 118894
rect 405234 82894 405854 118338
rect 405234 82338 405266 82894
rect 405822 82338 405854 82894
rect 405234 46894 405854 82338
rect 408726 58037 408786 457403
rect 408954 302614 409574 336000
rect 408954 302058 408986 302614
rect 409542 302058 409574 302614
rect 408954 266614 409574 302058
rect 408954 266058 408986 266614
rect 409542 266058 409574 266614
rect 408954 230614 409574 266058
rect 408954 230058 408986 230614
rect 409542 230058 409574 230614
rect 408954 194614 409574 230058
rect 408954 194058 408986 194614
rect 409542 194058 409574 194614
rect 408954 158614 409574 194058
rect 408954 158058 408986 158614
rect 409542 158058 409574 158614
rect 408954 122614 409574 158058
rect 408954 122058 408986 122614
rect 409542 122058 409574 122614
rect 408954 86614 409574 122058
rect 408954 86058 408986 86614
rect 409542 86058 409574 86614
rect 408723 58036 408789 58037
rect 408723 57972 408724 58036
rect 408788 57972 408789 58036
rect 408723 57971 408789 57972
rect 405234 46338 405266 46894
rect 405822 46338 405854 46894
rect 405234 10894 405854 46338
rect 405234 10338 405266 10894
rect 405822 10338 405854 10894
rect 405234 -4186 405854 10338
rect 405234 -4742 405266 -4186
rect 405822 -4742 405854 -4186
rect 405234 -5734 405854 -4742
rect 408954 50614 409574 86058
rect 408954 50058 408986 50614
rect 409542 50058 409574 50614
rect 408954 14614 409574 50058
rect 409830 31789 409890 457403
rect 409827 31788 409893 31789
rect 409827 31724 409828 31788
rect 409892 31724 409893 31788
rect 409827 31723 409893 31724
rect 411302 19957 411362 457403
rect 419514 457174 420134 492618
rect 419514 456618 419546 457174
rect 420102 456618 420134 457174
rect 419514 421174 420134 456618
rect 419514 420618 419546 421174
rect 420102 420618 420134 421174
rect 419514 385174 420134 420618
rect 419514 384618 419546 385174
rect 420102 384618 420134 385174
rect 419514 349174 420134 384618
rect 419514 348618 419546 349174
rect 420102 348618 420134 349174
rect 415794 309454 416414 336000
rect 415794 308898 415826 309454
rect 416382 308898 416414 309454
rect 415794 273454 416414 308898
rect 415794 272898 415826 273454
rect 416382 272898 416414 273454
rect 415794 237454 416414 272898
rect 415794 236898 415826 237454
rect 416382 236898 416414 237454
rect 415794 201454 416414 236898
rect 415794 200898 415826 201454
rect 416382 200898 416414 201454
rect 415794 165454 416414 200898
rect 415794 164898 415826 165454
rect 416382 164898 416414 165454
rect 415794 129454 416414 164898
rect 415794 128898 415826 129454
rect 416382 128898 416414 129454
rect 415794 93454 416414 128898
rect 415794 92898 415826 93454
rect 416382 92898 416414 93454
rect 415794 57454 416414 92898
rect 415794 56898 415826 57454
rect 416382 56898 416414 57454
rect 415794 21454 416414 56898
rect 415794 20898 415826 21454
rect 416382 20898 416414 21454
rect 411299 19956 411365 19957
rect 411299 19892 411300 19956
rect 411364 19892 411365 19956
rect 411299 19891 411365 19892
rect 408954 14058 408986 14614
rect 409542 14058 409574 14614
rect 390954 -7622 390986 -7066
rect 391542 -7622 391574 -7066
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 -1306 416414 20898
rect 415794 -1862 415826 -1306
rect 416382 -1862 416414 -1306
rect 415794 -1894 416414 -1862
rect 419514 313174 420134 348618
rect 419514 312618 419546 313174
rect 420102 312618 420134 313174
rect 419514 277174 420134 312618
rect 419514 276618 419546 277174
rect 420102 276618 420134 277174
rect 419514 241174 420134 276618
rect 419514 240618 419546 241174
rect 420102 240618 420134 241174
rect 419514 205174 420134 240618
rect 419514 204618 419546 205174
rect 420102 204618 420134 205174
rect 419514 169174 420134 204618
rect 419514 168618 419546 169174
rect 420102 168618 420134 169174
rect 419514 133174 420134 168618
rect 419514 132618 419546 133174
rect 420102 132618 420134 133174
rect 419514 97174 420134 132618
rect 419514 96618 419546 97174
rect 420102 96618 420134 97174
rect 419514 61174 420134 96618
rect 419514 60618 419546 61174
rect 420102 60618 420134 61174
rect 419514 25174 420134 60618
rect 419514 24618 419546 25174
rect 420102 24618 420134 25174
rect 419514 -3226 420134 24618
rect 419514 -3782 419546 -3226
rect 420102 -3782 420134 -3226
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676338 423266 676894
rect 423822 676338 423854 676894
rect 423234 640894 423854 676338
rect 423234 640338 423266 640894
rect 423822 640338 423854 640894
rect 423234 604894 423854 640338
rect 423234 604338 423266 604894
rect 423822 604338 423854 604894
rect 423234 568894 423854 604338
rect 423234 568338 423266 568894
rect 423822 568338 423854 568894
rect 423234 532894 423854 568338
rect 423234 532338 423266 532894
rect 423822 532338 423854 532894
rect 423234 496894 423854 532338
rect 423234 496338 423266 496894
rect 423822 496338 423854 496894
rect 423234 460894 423854 496338
rect 423234 460338 423266 460894
rect 423822 460338 423854 460894
rect 423234 424894 423854 460338
rect 423234 424338 423266 424894
rect 423822 424338 423854 424894
rect 423234 388894 423854 424338
rect 423234 388338 423266 388894
rect 423822 388338 423854 388894
rect 423234 352894 423854 388338
rect 423234 352338 423266 352894
rect 423822 352338 423854 352894
rect 423234 316894 423854 352338
rect 423234 316338 423266 316894
rect 423822 316338 423854 316894
rect 423234 280894 423854 316338
rect 423234 280338 423266 280894
rect 423822 280338 423854 280894
rect 423234 244894 423854 280338
rect 423234 244338 423266 244894
rect 423822 244338 423854 244894
rect 423234 208894 423854 244338
rect 423234 208338 423266 208894
rect 423822 208338 423854 208894
rect 423234 172894 423854 208338
rect 423234 172338 423266 172894
rect 423822 172338 423854 172894
rect 423234 136894 423854 172338
rect 423234 136338 423266 136894
rect 423822 136338 423854 136894
rect 423234 100894 423854 136338
rect 423234 100338 423266 100894
rect 423822 100338 423854 100894
rect 423234 64894 423854 100338
rect 423234 64338 423266 64894
rect 423822 64338 423854 64894
rect 423234 28894 423854 64338
rect 423234 28338 423266 28894
rect 423822 28338 423854 28894
rect 423234 -5146 423854 28338
rect 423234 -5702 423266 -5146
rect 423822 -5702 423854 -5146
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710042 444986 710598
rect 445542 710042 445574 710598
rect 441234 708678 441854 709670
rect 441234 708122 441266 708678
rect 441822 708122 441854 708678
rect 437514 706758 438134 707750
rect 437514 706202 437546 706758
rect 438102 706202 438134 706758
rect 426954 680058 426986 680614
rect 427542 680058 427574 680614
rect 426954 644614 427574 680058
rect 426954 644058 426986 644614
rect 427542 644058 427574 644614
rect 426954 608614 427574 644058
rect 426954 608058 426986 608614
rect 427542 608058 427574 608614
rect 426954 572614 427574 608058
rect 426954 572058 426986 572614
rect 427542 572058 427574 572614
rect 426954 536614 427574 572058
rect 426954 536058 426986 536614
rect 427542 536058 427574 536614
rect 426954 500614 427574 536058
rect 426954 500058 426986 500614
rect 427542 500058 427574 500614
rect 426954 464614 427574 500058
rect 426954 464058 426986 464614
rect 427542 464058 427574 464614
rect 426954 428614 427574 464058
rect 426954 428058 426986 428614
rect 427542 428058 427574 428614
rect 426954 392614 427574 428058
rect 426954 392058 426986 392614
rect 427542 392058 427574 392614
rect 426954 356614 427574 392058
rect 426954 356058 426986 356614
rect 427542 356058 427574 356614
rect 426954 320614 427574 356058
rect 426954 320058 426986 320614
rect 427542 320058 427574 320614
rect 426954 284614 427574 320058
rect 426954 284058 426986 284614
rect 427542 284058 427574 284614
rect 426954 248614 427574 284058
rect 426954 248058 426986 248614
rect 427542 248058 427574 248614
rect 426954 212614 427574 248058
rect 426954 212058 426986 212614
rect 427542 212058 427574 212614
rect 426954 176614 427574 212058
rect 426954 176058 426986 176614
rect 427542 176058 427574 176614
rect 426954 140614 427574 176058
rect 426954 140058 426986 140614
rect 427542 140058 427574 140614
rect 426954 104614 427574 140058
rect 426954 104058 426986 104614
rect 427542 104058 427574 104614
rect 426954 68614 427574 104058
rect 426954 68058 426986 68614
rect 427542 68058 427574 68614
rect 426954 32614 427574 68058
rect 426954 32058 426986 32614
rect 427542 32058 427574 32614
rect 408954 -6662 408986 -6106
rect 409542 -6662 409574 -6106
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704282 433826 704838
rect 434382 704282 434414 704838
rect 433794 687454 434414 704282
rect 433794 686898 433826 687454
rect 434382 686898 434414 687454
rect 433794 651454 434414 686898
rect 433794 650898 433826 651454
rect 434382 650898 434414 651454
rect 433794 615454 434414 650898
rect 433794 614898 433826 615454
rect 434382 614898 434414 615454
rect 433794 579454 434414 614898
rect 433794 578898 433826 579454
rect 434382 578898 434414 579454
rect 433794 543454 434414 578898
rect 433794 542898 433826 543454
rect 434382 542898 434414 543454
rect 433794 507454 434414 542898
rect 433794 506898 433826 507454
rect 434382 506898 434414 507454
rect 433794 471454 434414 506898
rect 433794 470898 433826 471454
rect 434382 470898 434414 471454
rect 433794 435454 434414 470898
rect 433794 434898 433826 435454
rect 434382 434898 434414 435454
rect 433794 399454 434414 434898
rect 433794 398898 433826 399454
rect 434382 398898 434414 399454
rect 433794 363454 434414 398898
rect 433794 362898 433826 363454
rect 434382 362898 434414 363454
rect 433794 327454 434414 362898
rect 433794 326898 433826 327454
rect 434382 326898 434414 327454
rect 433794 291454 434414 326898
rect 433794 290898 433826 291454
rect 434382 290898 434414 291454
rect 433794 255454 434414 290898
rect 433794 254898 433826 255454
rect 434382 254898 434414 255454
rect 433794 219454 434414 254898
rect 433794 218898 433826 219454
rect 434382 218898 434414 219454
rect 433794 183454 434414 218898
rect 433794 182898 433826 183454
rect 434382 182898 434414 183454
rect 433794 147454 434414 182898
rect 433794 146898 433826 147454
rect 434382 146898 434414 147454
rect 433794 111454 434414 146898
rect 433794 110898 433826 111454
rect 434382 110898 434414 111454
rect 433794 75454 434414 110898
rect 433794 74898 433826 75454
rect 434382 74898 434414 75454
rect 433794 39454 434414 74898
rect 433794 38898 433826 39454
rect 434382 38898 434414 39454
rect 433794 3454 434414 38898
rect 433794 2898 433826 3454
rect 434382 2898 434414 3454
rect 433794 -346 434414 2898
rect 433794 -902 433826 -346
rect 434382 -902 434414 -346
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690618 437546 691174
rect 438102 690618 438134 691174
rect 437514 655174 438134 690618
rect 437514 654618 437546 655174
rect 438102 654618 438134 655174
rect 437514 619174 438134 654618
rect 437514 618618 437546 619174
rect 438102 618618 438134 619174
rect 437514 583174 438134 618618
rect 437514 582618 437546 583174
rect 438102 582618 438134 583174
rect 437514 547174 438134 582618
rect 437514 546618 437546 547174
rect 438102 546618 438134 547174
rect 437514 511174 438134 546618
rect 437514 510618 437546 511174
rect 438102 510618 438134 511174
rect 437514 475174 438134 510618
rect 437514 474618 437546 475174
rect 438102 474618 438134 475174
rect 437514 439174 438134 474618
rect 437514 438618 437546 439174
rect 438102 438618 438134 439174
rect 437514 403174 438134 438618
rect 437514 402618 437546 403174
rect 438102 402618 438134 403174
rect 437514 367174 438134 402618
rect 437514 366618 437546 367174
rect 438102 366618 438134 367174
rect 437514 331174 438134 366618
rect 437514 330618 437546 331174
rect 438102 330618 438134 331174
rect 437514 295174 438134 330618
rect 437514 294618 437546 295174
rect 438102 294618 438134 295174
rect 437514 259174 438134 294618
rect 437514 258618 437546 259174
rect 438102 258618 438134 259174
rect 437514 223174 438134 258618
rect 437514 222618 437546 223174
rect 438102 222618 438134 223174
rect 437514 187174 438134 222618
rect 437514 186618 437546 187174
rect 438102 186618 438134 187174
rect 437514 151174 438134 186618
rect 437514 150618 437546 151174
rect 438102 150618 438134 151174
rect 437514 115174 438134 150618
rect 437514 114618 437546 115174
rect 438102 114618 438134 115174
rect 437514 79174 438134 114618
rect 437514 78618 437546 79174
rect 438102 78618 438134 79174
rect 437514 43174 438134 78618
rect 437514 42618 437546 43174
rect 438102 42618 438134 43174
rect 437514 7174 438134 42618
rect 437514 6618 437546 7174
rect 438102 6618 438134 7174
rect 437514 -2266 438134 6618
rect 437514 -2822 437546 -2266
rect 438102 -2822 438134 -2266
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694338 441266 694894
rect 441822 694338 441854 694894
rect 441234 658894 441854 694338
rect 441234 658338 441266 658894
rect 441822 658338 441854 658894
rect 441234 622894 441854 658338
rect 441234 622338 441266 622894
rect 441822 622338 441854 622894
rect 441234 586894 441854 622338
rect 441234 586338 441266 586894
rect 441822 586338 441854 586894
rect 441234 550894 441854 586338
rect 441234 550338 441266 550894
rect 441822 550338 441854 550894
rect 441234 514894 441854 550338
rect 441234 514338 441266 514894
rect 441822 514338 441854 514894
rect 441234 478894 441854 514338
rect 441234 478338 441266 478894
rect 441822 478338 441854 478894
rect 441234 442894 441854 478338
rect 441234 442338 441266 442894
rect 441822 442338 441854 442894
rect 441234 406894 441854 442338
rect 441234 406338 441266 406894
rect 441822 406338 441854 406894
rect 441234 370894 441854 406338
rect 441234 370338 441266 370894
rect 441822 370338 441854 370894
rect 441234 334894 441854 370338
rect 441234 334338 441266 334894
rect 441822 334338 441854 334894
rect 441234 298894 441854 334338
rect 441234 298338 441266 298894
rect 441822 298338 441854 298894
rect 441234 262894 441854 298338
rect 441234 262338 441266 262894
rect 441822 262338 441854 262894
rect 441234 226894 441854 262338
rect 441234 226338 441266 226894
rect 441822 226338 441854 226894
rect 441234 190894 441854 226338
rect 441234 190338 441266 190894
rect 441822 190338 441854 190894
rect 441234 154894 441854 190338
rect 441234 154338 441266 154894
rect 441822 154338 441854 154894
rect 441234 118894 441854 154338
rect 441234 118338 441266 118894
rect 441822 118338 441854 118894
rect 441234 82894 441854 118338
rect 441234 82338 441266 82894
rect 441822 82338 441854 82894
rect 441234 46894 441854 82338
rect 441234 46338 441266 46894
rect 441822 46338 441854 46894
rect 441234 10894 441854 46338
rect 441234 10338 441266 10894
rect 441822 10338 441854 10894
rect 441234 -4186 441854 10338
rect 441234 -4742 441266 -4186
rect 441822 -4742 441854 -4186
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711002 462986 711558
rect 463542 711002 463574 711558
rect 459234 709638 459854 709670
rect 459234 709082 459266 709638
rect 459822 709082 459854 709638
rect 455514 707718 456134 707750
rect 455514 707162 455546 707718
rect 456102 707162 456134 707718
rect 444954 698058 444986 698614
rect 445542 698058 445574 698614
rect 444954 662614 445574 698058
rect 444954 662058 444986 662614
rect 445542 662058 445574 662614
rect 444954 626614 445574 662058
rect 444954 626058 444986 626614
rect 445542 626058 445574 626614
rect 444954 590614 445574 626058
rect 444954 590058 444986 590614
rect 445542 590058 445574 590614
rect 444954 554614 445574 590058
rect 444954 554058 444986 554614
rect 445542 554058 445574 554614
rect 444954 518614 445574 554058
rect 444954 518058 444986 518614
rect 445542 518058 445574 518614
rect 444954 482614 445574 518058
rect 444954 482058 444986 482614
rect 445542 482058 445574 482614
rect 444954 446614 445574 482058
rect 444954 446058 444986 446614
rect 445542 446058 445574 446614
rect 444954 410614 445574 446058
rect 444954 410058 444986 410614
rect 445542 410058 445574 410614
rect 444954 374614 445574 410058
rect 444954 374058 444986 374614
rect 445542 374058 445574 374614
rect 444954 338614 445574 374058
rect 444954 338058 444986 338614
rect 445542 338058 445574 338614
rect 444954 302614 445574 338058
rect 444954 302058 444986 302614
rect 445542 302058 445574 302614
rect 444954 266614 445574 302058
rect 444954 266058 444986 266614
rect 445542 266058 445574 266614
rect 444954 230614 445574 266058
rect 444954 230058 444986 230614
rect 445542 230058 445574 230614
rect 444954 194614 445574 230058
rect 444954 194058 444986 194614
rect 445542 194058 445574 194614
rect 444954 158614 445574 194058
rect 444954 158058 444986 158614
rect 445542 158058 445574 158614
rect 444954 122614 445574 158058
rect 444954 122058 444986 122614
rect 445542 122058 445574 122614
rect 444954 86614 445574 122058
rect 444954 86058 444986 86614
rect 445542 86058 445574 86614
rect 444954 50614 445574 86058
rect 444954 50058 444986 50614
rect 445542 50058 445574 50614
rect 444954 14614 445574 50058
rect 444954 14058 444986 14614
rect 445542 14058 445574 14614
rect 426954 -7622 426986 -7066
rect 427542 -7622 427574 -7066
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705242 451826 705798
rect 452382 705242 452414 705798
rect 451794 669454 452414 705242
rect 451794 668898 451826 669454
rect 452382 668898 452414 669454
rect 451794 633454 452414 668898
rect 451794 632898 451826 633454
rect 452382 632898 452414 633454
rect 451794 597454 452414 632898
rect 451794 596898 451826 597454
rect 452382 596898 452414 597454
rect 451794 561454 452414 596898
rect 451794 560898 451826 561454
rect 452382 560898 452414 561454
rect 451794 525454 452414 560898
rect 451794 524898 451826 525454
rect 452382 524898 452414 525454
rect 451794 489454 452414 524898
rect 451794 488898 451826 489454
rect 452382 488898 452414 489454
rect 451794 453454 452414 488898
rect 451794 452898 451826 453454
rect 452382 452898 452414 453454
rect 451794 417454 452414 452898
rect 451794 416898 451826 417454
rect 452382 416898 452414 417454
rect 451794 381454 452414 416898
rect 451794 380898 451826 381454
rect 452382 380898 452414 381454
rect 451794 345454 452414 380898
rect 451794 344898 451826 345454
rect 452382 344898 452414 345454
rect 451794 309454 452414 344898
rect 451794 308898 451826 309454
rect 452382 308898 452414 309454
rect 451794 273454 452414 308898
rect 451794 272898 451826 273454
rect 452382 272898 452414 273454
rect 451794 237454 452414 272898
rect 451794 236898 451826 237454
rect 452382 236898 452414 237454
rect 451794 201454 452414 236898
rect 451794 200898 451826 201454
rect 452382 200898 452414 201454
rect 451794 165454 452414 200898
rect 451794 164898 451826 165454
rect 452382 164898 452414 165454
rect 451794 129454 452414 164898
rect 451794 128898 451826 129454
rect 452382 128898 452414 129454
rect 451794 93454 452414 128898
rect 451794 92898 451826 93454
rect 452382 92898 452414 93454
rect 451794 57454 452414 92898
rect 451794 56898 451826 57454
rect 452382 56898 452414 57454
rect 451794 21454 452414 56898
rect 451794 20898 451826 21454
rect 452382 20898 452414 21454
rect 451794 -1306 452414 20898
rect 451794 -1862 451826 -1306
rect 452382 -1862 452414 -1306
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672618 455546 673174
rect 456102 672618 456134 673174
rect 455514 637174 456134 672618
rect 455514 636618 455546 637174
rect 456102 636618 456134 637174
rect 455514 601174 456134 636618
rect 455514 600618 455546 601174
rect 456102 600618 456134 601174
rect 455514 565174 456134 600618
rect 455514 564618 455546 565174
rect 456102 564618 456134 565174
rect 455514 529174 456134 564618
rect 455514 528618 455546 529174
rect 456102 528618 456134 529174
rect 455514 493174 456134 528618
rect 455514 492618 455546 493174
rect 456102 492618 456134 493174
rect 455514 457174 456134 492618
rect 455514 456618 455546 457174
rect 456102 456618 456134 457174
rect 455514 421174 456134 456618
rect 455514 420618 455546 421174
rect 456102 420618 456134 421174
rect 455514 385174 456134 420618
rect 455514 384618 455546 385174
rect 456102 384618 456134 385174
rect 455514 349174 456134 384618
rect 455514 348618 455546 349174
rect 456102 348618 456134 349174
rect 455514 313174 456134 348618
rect 455514 312618 455546 313174
rect 456102 312618 456134 313174
rect 455514 277174 456134 312618
rect 455514 276618 455546 277174
rect 456102 276618 456134 277174
rect 455514 241174 456134 276618
rect 455514 240618 455546 241174
rect 456102 240618 456134 241174
rect 455514 205174 456134 240618
rect 455514 204618 455546 205174
rect 456102 204618 456134 205174
rect 455514 169174 456134 204618
rect 455514 168618 455546 169174
rect 456102 168618 456134 169174
rect 455514 133174 456134 168618
rect 455514 132618 455546 133174
rect 456102 132618 456134 133174
rect 455514 97174 456134 132618
rect 455514 96618 455546 97174
rect 456102 96618 456134 97174
rect 455514 61174 456134 96618
rect 455514 60618 455546 61174
rect 456102 60618 456134 61174
rect 455514 25174 456134 60618
rect 455514 24618 455546 25174
rect 456102 24618 456134 25174
rect 455514 -3226 456134 24618
rect 455514 -3782 455546 -3226
rect 456102 -3782 456134 -3226
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676338 459266 676894
rect 459822 676338 459854 676894
rect 459234 640894 459854 676338
rect 459234 640338 459266 640894
rect 459822 640338 459854 640894
rect 459234 604894 459854 640338
rect 459234 604338 459266 604894
rect 459822 604338 459854 604894
rect 459234 568894 459854 604338
rect 459234 568338 459266 568894
rect 459822 568338 459854 568894
rect 459234 532894 459854 568338
rect 459234 532338 459266 532894
rect 459822 532338 459854 532894
rect 459234 496894 459854 532338
rect 459234 496338 459266 496894
rect 459822 496338 459854 496894
rect 459234 460894 459854 496338
rect 459234 460338 459266 460894
rect 459822 460338 459854 460894
rect 459234 424894 459854 460338
rect 459234 424338 459266 424894
rect 459822 424338 459854 424894
rect 459234 388894 459854 424338
rect 459234 388338 459266 388894
rect 459822 388338 459854 388894
rect 459234 352894 459854 388338
rect 459234 352338 459266 352894
rect 459822 352338 459854 352894
rect 459234 316894 459854 352338
rect 459234 316338 459266 316894
rect 459822 316338 459854 316894
rect 459234 280894 459854 316338
rect 459234 280338 459266 280894
rect 459822 280338 459854 280894
rect 459234 244894 459854 280338
rect 459234 244338 459266 244894
rect 459822 244338 459854 244894
rect 459234 208894 459854 244338
rect 459234 208338 459266 208894
rect 459822 208338 459854 208894
rect 459234 172894 459854 208338
rect 459234 172338 459266 172894
rect 459822 172338 459854 172894
rect 459234 136894 459854 172338
rect 459234 136338 459266 136894
rect 459822 136338 459854 136894
rect 459234 100894 459854 136338
rect 459234 100338 459266 100894
rect 459822 100338 459854 100894
rect 459234 64894 459854 100338
rect 459234 64338 459266 64894
rect 459822 64338 459854 64894
rect 459234 28894 459854 64338
rect 459234 28338 459266 28894
rect 459822 28338 459854 28894
rect 459234 -5146 459854 28338
rect 459234 -5702 459266 -5146
rect 459822 -5702 459854 -5146
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710042 480986 710598
rect 481542 710042 481574 710598
rect 477234 708678 477854 709670
rect 477234 708122 477266 708678
rect 477822 708122 477854 708678
rect 473514 706758 474134 707750
rect 473514 706202 473546 706758
rect 474102 706202 474134 706758
rect 462954 680058 462986 680614
rect 463542 680058 463574 680614
rect 462954 644614 463574 680058
rect 462954 644058 462986 644614
rect 463542 644058 463574 644614
rect 462954 608614 463574 644058
rect 462954 608058 462986 608614
rect 463542 608058 463574 608614
rect 462954 572614 463574 608058
rect 462954 572058 462986 572614
rect 463542 572058 463574 572614
rect 462954 536614 463574 572058
rect 462954 536058 462986 536614
rect 463542 536058 463574 536614
rect 462954 500614 463574 536058
rect 462954 500058 462986 500614
rect 463542 500058 463574 500614
rect 462954 464614 463574 500058
rect 462954 464058 462986 464614
rect 463542 464058 463574 464614
rect 462954 428614 463574 464058
rect 462954 428058 462986 428614
rect 463542 428058 463574 428614
rect 462954 392614 463574 428058
rect 462954 392058 462986 392614
rect 463542 392058 463574 392614
rect 462954 356614 463574 392058
rect 462954 356058 462986 356614
rect 463542 356058 463574 356614
rect 462954 320614 463574 356058
rect 462954 320058 462986 320614
rect 463542 320058 463574 320614
rect 462954 284614 463574 320058
rect 462954 284058 462986 284614
rect 463542 284058 463574 284614
rect 462954 248614 463574 284058
rect 462954 248058 462986 248614
rect 463542 248058 463574 248614
rect 462954 212614 463574 248058
rect 462954 212058 462986 212614
rect 463542 212058 463574 212614
rect 462954 176614 463574 212058
rect 462954 176058 462986 176614
rect 463542 176058 463574 176614
rect 462954 140614 463574 176058
rect 462954 140058 462986 140614
rect 463542 140058 463574 140614
rect 462954 104614 463574 140058
rect 462954 104058 462986 104614
rect 463542 104058 463574 104614
rect 462954 68614 463574 104058
rect 462954 68058 462986 68614
rect 463542 68058 463574 68614
rect 462954 32614 463574 68058
rect 462954 32058 462986 32614
rect 463542 32058 463574 32614
rect 444954 -6662 444986 -6106
rect 445542 -6662 445574 -6106
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704282 469826 704838
rect 470382 704282 470414 704838
rect 469794 687454 470414 704282
rect 469794 686898 469826 687454
rect 470382 686898 470414 687454
rect 469794 651454 470414 686898
rect 469794 650898 469826 651454
rect 470382 650898 470414 651454
rect 469794 615454 470414 650898
rect 469794 614898 469826 615454
rect 470382 614898 470414 615454
rect 469794 579454 470414 614898
rect 469794 578898 469826 579454
rect 470382 578898 470414 579454
rect 469794 543454 470414 578898
rect 469794 542898 469826 543454
rect 470382 542898 470414 543454
rect 469794 507454 470414 542898
rect 469794 506898 469826 507454
rect 470382 506898 470414 507454
rect 469794 471454 470414 506898
rect 469794 470898 469826 471454
rect 470382 470898 470414 471454
rect 469794 435454 470414 470898
rect 469794 434898 469826 435454
rect 470382 434898 470414 435454
rect 469794 399454 470414 434898
rect 469794 398898 469826 399454
rect 470382 398898 470414 399454
rect 469794 363454 470414 398898
rect 469794 362898 469826 363454
rect 470382 362898 470414 363454
rect 469794 327454 470414 362898
rect 469794 326898 469826 327454
rect 470382 326898 470414 327454
rect 469794 291454 470414 326898
rect 469794 290898 469826 291454
rect 470382 290898 470414 291454
rect 469794 255454 470414 290898
rect 469794 254898 469826 255454
rect 470382 254898 470414 255454
rect 469794 219454 470414 254898
rect 469794 218898 469826 219454
rect 470382 218898 470414 219454
rect 469794 183454 470414 218898
rect 469794 182898 469826 183454
rect 470382 182898 470414 183454
rect 469794 147454 470414 182898
rect 469794 146898 469826 147454
rect 470382 146898 470414 147454
rect 469794 111454 470414 146898
rect 469794 110898 469826 111454
rect 470382 110898 470414 111454
rect 469794 75454 470414 110898
rect 469794 74898 469826 75454
rect 470382 74898 470414 75454
rect 469794 39454 470414 74898
rect 469794 38898 469826 39454
rect 470382 38898 470414 39454
rect 469794 3454 470414 38898
rect 469794 2898 469826 3454
rect 470382 2898 470414 3454
rect 469794 -346 470414 2898
rect 469794 -902 469826 -346
rect 470382 -902 470414 -346
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690618 473546 691174
rect 474102 690618 474134 691174
rect 473514 655174 474134 690618
rect 473514 654618 473546 655174
rect 474102 654618 474134 655174
rect 473514 619174 474134 654618
rect 473514 618618 473546 619174
rect 474102 618618 474134 619174
rect 473514 583174 474134 618618
rect 473514 582618 473546 583174
rect 474102 582618 474134 583174
rect 473514 547174 474134 582618
rect 473514 546618 473546 547174
rect 474102 546618 474134 547174
rect 473514 511174 474134 546618
rect 473514 510618 473546 511174
rect 474102 510618 474134 511174
rect 473514 475174 474134 510618
rect 473514 474618 473546 475174
rect 474102 474618 474134 475174
rect 473514 439174 474134 474618
rect 473514 438618 473546 439174
rect 474102 438618 474134 439174
rect 473514 403174 474134 438618
rect 473514 402618 473546 403174
rect 474102 402618 474134 403174
rect 473514 367174 474134 402618
rect 473514 366618 473546 367174
rect 474102 366618 474134 367174
rect 473514 331174 474134 366618
rect 473514 330618 473546 331174
rect 474102 330618 474134 331174
rect 473514 295174 474134 330618
rect 473514 294618 473546 295174
rect 474102 294618 474134 295174
rect 473514 259174 474134 294618
rect 473514 258618 473546 259174
rect 474102 258618 474134 259174
rect 473514 223174 474134 258618
rect 473514 222618 473546 223174
rect 474102 222618 474134 223174
rect 473514 187174 474134 222618
rect 473514 186618 473546 187174
rect 474102 186618 474134 187174
rect 473514 151174 474134 186618
rect 473514 150618 473546 151174
rect 474102 150618 474134 151174
rect 473514 115174 474134 150618
rect 473514 114618 473546 115174
rect 474102 114618 474134 115174
rect 473514 79174 474134 114618
rect 473514 78618 473546 79174
rect 474102 78618 474134 79174
rect 473514 43174 474134 78618
rect 473514 42618 473546 43174
rect 474102 42618 474134 43174
rect 473514 7174 474134 42618
rect 473514 6618 473546 7174
rect 474102 6618 474134 7174
rect 473514 -2266 474134 6618
rect 473514 -2822 473546 -2266
rect 474102 -2822 474134 -2266
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694338 477266 694894
rect 477822 694338 477854 694894
rect 477234 658894 477854 694338
rect 477234 658338 477266 658894
rect 477822 658338 477854 658894
rect 477234 622894 477854 658338
rect 477234 622338 477266 622894
rect 477822 622338 477854 622894
rect 477234 586894 477854 622338
rect 477234 586338 477266 586894
rect 477822 586338 477854 586894
rect 477234 550894 477854 586338
rect 477234 550338 477266 550894
rect 477822 550338 477854 550894
rect 477234 514894 477854 550338
rect 477234 514338 477266 514894
rect 477822 514338 477854 514894
rect 477234 478894 477854 514338
rect 477234 478338 477266 478894
rect 477822 478338 477854 478894
rect 477234 442894 477854 478338
rect 477234 442338 477266 442894
rect 477822 442338 477854 442894
rect 477234 406894 477854 442338
rect 477234 406338 477266 406894
rect 477822 406338 477854 406894
rect 477234 370894 477854 406338
rect 477234 370338 477266 370894
rect 477822 370338 477854 370894
rect 477234 334894 477854 370338
rect 477234 334338 477266 334894
rect 477822 334338 477854 334894
rect 477234 298894 477854 334338
rect 477234 298338 477266 298894
rect 477822 298338 477854 298894
rect 477234 262894 477854 298338
rect 477234 262338 477266 262894
rect 477822 262338 477854 262894
rect 477234 226894 477854 262338
rect 477234 226338 477266 226894
rect 477822 226338 477854 226894
rect 477234 190894 477854 226338
rect 477234 190338 477266 190894
rect 477822 190338 477854 190894
rect 477234 154894 477854 190338
rect 477234 154338 477266 154894
rect 477822 154338 477854 154894
rect 477234 118894 477854 154338
rect 477234 118338 477266 118894
rect 477822 118338 477854 118894
rect 477234 82894 477854 118338
rect 477234 82338 477266 82894
rect 477822 82338 477854 82894
rect 477234 46894 477854 82338
rect 477234 46338 477266 46894
rect 477822 46338 477854 46894
rect 477234 10894 477854 46338
rect 477234 10338 477266 10894
rect 477822 10338 477854 10894
rect 477234 -4186 477854 10338
rect 477234 -4742 477266 -4186
rect 477822 -4742 477854 -4186
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711002 498986 711558
rect 499542 711002 499574 711558
rect 495234 709638 495854 709670
rect 495234 709082 495266 709638
rect 495822 709082 495854 709638
rect 491514 707718 492134 707750
rect 491514 707162 491546 707718
rect 492102 707162 492134 707718
rect 480954 698058 480986 698614
rect 481542 698058 481574 698614
rect 480954 662614 481574 698058
rect 480954 662058 480986 662614
rect 481542 662058 481574 662614
rect 480954 626614 481574 662058
rect 480954 626058 480986 626614
rect 481542 626058 481574 626614
rect 480954 590614 481574 626058
rect 480954 590058 480986 590614
rect 481542 590058 481574 590614
rect 480954 554614 481574 590058
rect 480954 554058 480986 554614
rect 481542 554058 481574 554614
rect 480954 518614 481574 554058
rect 480954 518058 480986 518614
rect 481542 518058 481574 518614
rect 480954 482614 481574 518058
rect 480954 482058 480986 482614
rect 481542 482058 481574 482614
rect 480954 446614 481574 482058
rect 480954 446058 480986 446614
rect 481542 446058 481574 446614
rect 480954 410614 481574 446058
rect 480954 410058 480986 410614
rect 481542 410058 481574 410614
rect 480954 374614 481574 410058
rect 480954 374058 480986 374614
rect 481542 374058 481574 374614
rect 480954 338614 481574 374058
rect 480954 338058 480986 338614
rect 481542 338058 481574 338614
rect 480954 302614 481574 338058
rect 480954 302058 480986 302614
rect 481542 302058 481574 302614
rect 480954 266614 481574 302058
rect 480954 266058 480986 266614
rect 481542 266058 481574 266614
rect 480954 230614 481574 266058
rect 480954 230058 480986 230614
rect 481542 230058 481574 230614
rect 480954 194614 481574 230058
rect 480954 194058 480986 194614
rect 481542 194058 481574 194614
rect 480954 158614 481574 194058
rect 480954 158058 480986 158614
rect 481542 158058 481574 158614
rect 480954 122614 481574 158058
rect 480954 122058 480986 122614
rect 481542 122058 481574 122614
rect 480954 86614 481574 122058
rect 480954 86058 480986 86614
rect 481542 86058 481574 86614
rect 480954 50614 481574 86058
rect 480954 50058 480986 50614
rect 481542 50058 481574 50614
rect 480954 14614 481574 50058
rect 480954 14058 480986 14614
rect 481542 14058 481574 14614
rect 462954 -7622 462986 -7066
rect 463542 -7622 463574 -7066
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705242 487826 705798
rect 488382 705242 488414 705798
rect 487794 669454 488414 705242
rect 487794 668898 487826 669454
rect 488382 668898 488414 669454
rect 487794 633454 488414 668898
rect 487794 632898 487826 633454
rect 488382 632898 488414 633454
rect 487794 597454 488414 632898
rect 487794 596898 487826 597454
rect 488382 596898 488414 597454
rect 487794 561454 488414 596898
rect 487794 560898 487826 561454
rect 488382 560898 488414 561454
rect 487794 525454 488414 560898
rect 487794 524898 487826 525454
rect 488382 524898 488414 525454
rect 487794 489454 488414 524898
rect 487794 488898 487826 489454
rect 488382 488898 488414 489454
rect 487794 453454 488414 488898
rect 487794 452898 487826 453454
rect 488382 452898 488414 453454
rect 487794 417454 488414 452898
rect 487794 416898 487826 417454
rect 488382 416898 488414 417454
rect 487794 381454 488414 416898
rect 487794 380898 487826 381454
rect 488382 380898 488414 381454
rect 487794 345454 488414 380898
rect 487794 344898 487826 345454
rect 488382 344898 488414 345454
rect 487794 309454 488414 344898
rect 487794 308898 487826 309454
rect 488382 308898 488414 309454
rect 487794 273454 488414 308898
rect 487794 272898 487826 273454
rect 488382 272898 488414 273454
rect 487794 237454 488414 272898
rect 487794 236898 487826 237454
rect 488382 236898 488414 237454
rect 487794 201454 488414 236898
rect 487794 200898 487826 201454
rect 488382 200898 488414 201454
rect 487794 165454 488414 200898
rect 487794 164898 487826 165454
rect 488382 164898 488414 165454
rect 487794 129454 488414 164898
rect 487794 128898 487826 129454
rect 488382 128898 488414 129454
rect 487794 93454 488414 128898
rect 487794 92898 487826 93454
rect 488382 92898 488414 93454
rect 487794 57454 488414 92898
rect 487794 56898 487826 57454
rect 488382 56898 488414 57454
rect 487794 21454 488414 56898
rect 487794 20898 487826 21454
rect 488382 20898 488414 21454
rect 487794 -1306 488414 20898
rect 487794 -1862 487826 -1306
rect 488382 -1862 488414 -1306
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672618 491546 673174
rect 492102 672618 492134 673174
rect 491514 637174 492134 672618
rect 491514 636618 491546 637174
rect 492102 636618 492134 637174
rect 491514 601174 492134 636618
rect 491514 600618 491546 601174
rect 492102 600618 492134 601174
rect 491514 565174 492134 600618
rect 491514 564618 491546 565174
rect 492102 564618 492134 565174
rect 491514 529174 492134 564618
rect 491514 528618 491546 529174
rect 492102 528618 492134 529174
rect 491514 493174 492134 528618
rect 491514 492618 491546 493174
rect 492102 492618 492134 493174
rect 491514 457174 492134 492618
rect 491514 456618 491546 457174
rect 492102 456618 492134 457174
rect 491514 421174 492134 456618
rect 491514 420618 491546 421174
rect 492102 420618 492134 421174
rect 491514 385174 492134 420618
rect 491514 384618 491546 385174
rect 492102 384618 492134 385174
rect 491514 349174 492134 384618
rect 491514 348618 491546 349174
rect 492102 348618 492134 349174
rect 491514 313174 492134 348618
rect 491514 312618 491546 313174
rect 492102 312618 492134 313174
rect 491514 277174 492134 312618
rect 491514 276618 491546 277174
rect 492102 276618 492134 277174
rect 491514 241174 492134 276618
rect 491514 240618 491546 241174
rect 492102 240618 492134 241174
rect 491514 205174 492134 240618
rect 491514 204618 491546 205174
rect 492102 204618 492134 205174
rect 491514 169174 492134 204618
rect 491514 168618 491546 169174
rect 492102 168618 492134 169174
rect 491514 133174 492134 168618
rect 491514 132618 491546 133174
rect 492102 132618 492134 133174
rect 491514 97174 492134 132618
rect 491514 96618 491546 97174
rect 492102 96618 492134 97174
rect 491514 61174 492134 96618
rect 491514 60618 491546 61174
rect 492102 60618 492134 61174
rect 491514 25174 492134 60618
rect 491514 24618 491546 25174
rect 492102 24618 492134 25174
rect 491514 -3226 492134 24618
rect 491514 -3782 491546 -3226
rect 492102 -3782 492134 -3226
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676338 495266 676894
rect 495822 676338 495854 676894
rect 495234 640894 495854 676338
rect 495234 640338 495266 640894
rect 495822 640338 495854 640894
rect 495234 604894 495854 640338
rect 495234 604338 495266 604894
rect 495822 604338 495854 604894
rect 495234 568894 495854 604338
rect 495234 568338 495266 568894
rect 495822 568338 495854 568894
rect 495234 532894 495854 568338
rect 495234 532338 495266 532894
rect 495822 532338 495854 532894
rect 495234 496894 495854 532338
rect 495234 496338 495266 496894
rect 495822 496338 495854 496894
rect 495234 460894 495854 496338
rect 495234 460338 495266 460894
rect 495822 460338 495854 460894
rect 495234 424894 495854 460338
rect 495234 424338 495266 424894
rect 495822 424338 495854 424894
rect 495234 388894 495854 424338
rect 495234 388338 495266 388894
rect 495822 388338 495854 388894
rect 495234 352894 495854 388338
rect 495234 352338 495266 352894
rect 495822 352338 495854 352894
rect 495234 316894 495854 352338
rect 495234 316338 495266 316894
rect 495822 316338 495854 316894
rect 495234 280894 495854 316338
rect 495234 280338 495266 280894
rect 495822 280338 495854 280894
rect 495234 244894 495854 280338
rect 495234 244338 495266 244894
rect 495822 244338 495854 244894
rect 495234 208894 495854 244338
rect 495234 208338 495266 208894
rect 495822 208338 495854 208894
rect 495234 172894 495854 208338
rect 495234 172338 495266 172894
rect 495822 172338 495854 172894
rect 495234 136894 495854 172338
rect 495234 136338 495266 136894
rect 495822 136338 495854 136894
rect 495234 100894 495854 136338
rect 495234 100338 495266 100894
rect 495822 100338 495854 100894
rect 495234 64894 495854 100338
rect 495234 64338 495266 64894
rect 495822 64338 495854 64894
rect 495234 28894 495854 64338
rect 495234 28338 495266 28894
rect 495822 28338 495854 28894
rect 495234 -5146 495854 28338
rect 495234 -5702 495266 -5146
rect 495822 -5702 495854 -5146
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710042 516986 710598
rect 517542 710042 517574 710598
rect 513234 708678 513854 709670
rect 513234 708122 513266 708678
rect 513822 708122 513854 708678
rect 509514 706758 510134 707750
rect 509514 706202 509546 706758
rect 510102 706202 510134 706758
rect 498954 680058 498986 680614
rect 499542 680058 499574 680614
rect 498954 644614 499574 680058
rect 498954 644058 498986 644614
rect 499542 644058 499574 644614
rect 498954 608614 499574 644058
rect 498954 608058 498986 608614
rect 499542 608058 499574 608614
rect 498954 572614 499574 608058
rect 498954 572058 498986 572614
rect 499542 572058 499574 572614
rect 498954 536614 499574 572058
rect 498954 536058 498986 536614
rect 499542 536058 499574 536614
rect 498954 500614 499574 536058
rect 498954 500058 498986 500614
rect 499542 500058 499574 500614
rect 498954 464614 499574 500058
rect 498954 464058 498986 464614
rect 499542 464058 499574 464614
rect 498954 428614 499574 464058
rect 498954 428058 498986 428614
rect 499542 428058 499574 428614
rect 498954 392614 499574 428058
rect 498954 392058 498986 392614
rect 499542 392058 499574 392614
rect 498954 356614 499574 392058
rect 498954 356058 498986 356614
rect 499542 356058 499574 356614
rect 498954 320614 499574 356058
rect 498954 320058 498986 320614
rect 499542 320058 499574 320614
rect 498954 284614 499574 320058
rect 498954 284058 498986 284614
rect 499542 284058 499574 284614
rect 498954 248614 499574 284058
rect 498954 248058 498986 248614
rect 499542 248058 499574 248614
rect 498954 212614 499574 248058
rect 498954 212058 498986 212614
rect 499542 212058 499574 212614
rect 498954 176614 499574 212058
rect 498954 176058 498986 176614
rect 499542 176058 499574 176614
rect 498954 140614 499574 176058
rect 498954 140058 498986 140614
rect 499542 140058 499574 140614
rect 498954 104614 499574 140058
rect 498954 104058 498986 104614
rect 499542 104058 499574 104614
rect 498954 68614 499574 104058
rect 498954 68058 498986 68614
rect 499542 68058 499574 68614
rect 498954 32614 499574 68058
rect 498954 32058 498986 32614
rect 499542 32058 499574 32614
rect 480954 -6662 480986 -6106
rect 481542 -6662 481574 -6106
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704282 505826 704838
rect 506382 704282 506414 704838
rect 505794 687454 506414 704282
rect 505794 686898 505826 687454
rect 506382 686898 506414 687454
rect 505794 651454 506414 686898
rect 505794 650898 505826 651454
rect 506382 650898 506414 651454
rect 505794 615454 506414 650898
rect 505794 614898 505826 615454
rect 506382 614898 506414 615454
rect 505794 579454 506414 614898
rect 505794 578898 505826 579454
rect 506382 578898 506414 579454
rect 505794 543454 506414 578898
rect 505794 542898 505826 543454
rect 506382 542898 506414 543454
rect 505794 507454 506414 542898
rect 505794 506898 505826 507454
rect 506382 506898 506414 507454
rect 505794 471454 506414 506898
rect 505794 470898 505826 471454
rect 506382 470898 506414 471454
rect 505794 435454 506414 470898
rect 505794 434898 505826 435454
rect 506382 434898 506414 435454
rect 505794 399454 506414 434898
rect 505794 398898 505826 399454
rect 506382 398898 506414 399454
rect 505794 363454 506414 398898
rect 505794 362898 505826 363454
rect 506382 362898 506414 363454
rect 505794 327454 506414 362898
rect 505794 326898 505826 327454
rect 506382 326898 506414 327454
rect 505794 291454 506414 326898
rect 505794 290898 505826 291454
rect 506382 290898 506414 291454
rect 505794 255454 506414 290898
rect 505794 254898 505826 255454
rect 506382 254898 506414 255454
rect 505794 219454 506414 254898
rect 505794 218898 505826 219454
rect 506382 218898 506414 219454
rect 505794 183454 506414 218898
rect 505794 182898 505826 183454
rect 506382 182898 506414 183454
rect 505794 147454 506414 182898
rect 505794 146898 505826 147454
rect 506382 146898 506414 147454
rect 505794 111454 506414 146898
rect 505794 110898 505826 111454
rect 506382 110898 506414 111454
rect 505794 75454 506414 110898
rect 505794 74898 505826 75454
rect 506382 74898 506414 75454
rect 505794 39454 506414 74898
rect 505794 38898 505826 39454
rect 506382 38898 506414 39454
rect 505794 3454 506414 38898
rect 505794 2898 505826 3454
rect 506382 2898 506414 3454
rect 505794 -346 506414 2898
rect 505794 -902 505826 -346
rect 506382 -902 506414 -346
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690618 509546 691174
rect 510102 690618 510134 691174
rect 509514 655174 510134 690618
rect 509514 654618 509546 655174
rect 510102 654618 510134 655174
rect 509514 619174 510134 654618
rect 509514 618618 509546 619174
rect 510102 618618 510134 619174
rect 509514 583174 510134 618618
rect 509514 582618 509546 583174
rect 510102 582618 510134 583174
rect 509514 547174 510134 582618
rect 509514 546618 509546 547174
rect 510102 546618 510134 547174
rect 509514 511174 510134 546618
rect 509514 510618 509546 511174
rect 510102 510618 510134 511174
rect 509514 475174 510134 510618
rect 509514 474618 509546 475174
rect 510102 474618 510134 475174
rect 509514 439174 510134 474618
rect 509514 438618 509546 439174
rect 510102 438618 510134 439174
rect 509514 403174 510134 438618
rect 509514 402618 509546 403174
rect 510102 402618 510134 403174
rect 509514 367174 510134 402618
rect 509514 366618 509546 367174
rect 510102 366618 510134 367174
rect 509514 331174 510134 366618
rect 509514 330618 509546 331174
rect 510102 330618 510134 331174
rect 509514 295174 510134 330618
rect 509514 294618 509546 295174
rect 510102 294618 510134 295174
rect 509514 259174 510134 294618
rect 509514 258618 509546 259174
rect 510102 258618 510134 259174
rect 509514 223174 510134 258618
rect 509514 222618 509546 223174
rect 510102 222618 510134 223174
rect 509514 187174 510134 222618
rect 509514 186618 509546 187174
rect 510102 186618 510134 187174
rect 509514 151174 510134 186618
rect 509514 150618 509546 151174
rect 510102 150618 510134 151174
rect 509514 115174 510134 150618
rect 509514 114618 509546 115174
rect 510102 114618 510134 115174
rect 509514 79174 510134 114618
rect 509514 78618 509546 79174
rect 510102 78618 510134 79174
rect 509514 43174 510134 78618
rect 509514 42618 509546 43174
rect 510102 42618 510134 43174
rect 509514 7174 510134 42618
rect 509514 6618 509546 7174
rect 510102 6618 510134 7174
rect 509514 -2266 510134 6618
rect 509514 -2822 509546 -2266
rect 510102 -2822 510134 -2266
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694338 513266 694894
rect 513822 694338 513854 694894
rect 513234 658894 513854 694338
rect 513234 658338 513266 658894
rect 513822 658338 513854 658894
rect 513234 622894 513854 658338
rect 513234 622338 513266 622894
rect 513822 622338 513854 622894
rect 513234 586894 513854 622338
rect 513234 586338 513266 586894
rect 513822 586338 513854 586894
rect 513234 550894 513854 586338
rect 513234 550338 513266 550894
rect 513822 550338 513854 550894
rect 513234 514894 513854 550338
rect 513234 514338 513266 514894
rect 513822 514338 513854 514894
rect 513234 478894 513854 514338
rect 513234 478338 513266 478894
rect 513822 478338 513854 478894
rect 513234 442894 513854 478338
rect 513234 442338 513266 442894
rect 513822 442338 513854 442894
rect 513234 406894 513854 442338
rect 513234 406338 513266 406894
rect 513822 406338 513854 406894
rect 513234 370894 513854 406338
rect 513234 370338 513266 370894
rect 513822 370338 513854 370894
rect 513234 334894 513854 370338
rect 513234 334338 513266 334894
rect 513822 334338 513854 334894
rect 513234 298894 513854 334338
rect 513234 298338 513266 298894
rect 513822 298338 513854 298894
rect 513234 262894 513854 298338
rect 513234 262338 513266 262894
rect 513822 262338 513854 262894
rect 513234 226894 513854 262338
rect 513234 226338 513266 226894
rect 513822 226338 513854 226894
rect 513234 190894 513854 226338
rect 513234 190338 513266 190894
rect 513822 190338 513854 190894
rect 513234 154894 513854 190338
rect 513234 154338 513266 154894
rect 513822 154338 513854 154894
rect 513234 118894 513854 154338
rect 513234 118338 513266 118894
rect 513822 118338 513854 118894
rect 513234 82894 513854 118338
rect 513234 82338 513266 82894
rect 513822 82338 513854 82894
rect 513234 46894 513854 82338
rect 513234 46338 513266 46894
rect 513822 46338 513854 46894
rect 513234 10894 513854 46338
rect 513234 10338 513266 10894
rect 513822 10338 513854 10894
rect 513234 -4186 513854 10338
rect 513234 -4742 513266 -4186
rect 513822 -4742 513854 -4186
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711002 534986 711558
rect 535542 711002 535574 711558
rect 531234 709638 531854 709670
rect 531234 709082 531266 709638
rect 531822 709082 531854 709638
rect 527514 707718 528134 707750
rect 527514 707162 527546 707718
rect 528102 707162 528134 707718
rect 516954 698058 516986 698614
rect 517542 698058 517574 698614
rect 516954 662614 517574 698058
rect 516954 662058 516986 662614
rect 517542 662058 517574 662614
rect 516954 626614 517574 662058
rect 516954 626058 516986 626614
rect 517542 626058 517574 626614
rect 516954 590614 517574 626058
rect 516954 590058 516986 590614
rect 517542 590058 517574 590614
rect 516954 554614 517574 590058
rect 516954 554058 516986 554614
rect 517542 554058 517574 554614
rect 516954 518614 517574 554058
rect 516954 518058 516986 518614
rect 517542 518058 517574 518614
rect 516954 482614 517574 518058
rect 516954 482058 516986 482614
rect 517542 482058 517574 482614
rect 516954 446614 517574 482058
rect 516954 446058 516986 446614
rect 517542 446058 517574 446614
rect 516954 410614 517574 446058
rect 516954 410058 516986 410614
rect 517542 410058 517574 410614
rect 516954 374614 517574 410058
rect 516954 374058 516986 374614
rect 517542 374058 517574 374614
rect 516954 338614 517574 374058
rect 516954 338058 516986 338614
rect 517542 338058 517574 338614
rect 516954 302614 517574 338058
rect 516954 302058 516986 302614
rect 517542 302058 517574 302614
rect 516954 266614 517574 302058
rect 516954 266058 516986 266614
rect 517542 266058 517574 266614
rect 516954 230614 517574 266058
rect 516954 230058 516986 230614
rect 517542 230058 517574 230614
rect 516954 194614 517574 230058
rect 516954 194058 516986 194614
rect 517542 194058 517574 194614
rect 516954 158614 517574 194058
rect 516954 158058 516986 158614
rect 517542 158058 517574 158614
rect 516954 122614 517574 158058
rect 516954 122058 516986 122614
rect 517542 122058 517574 122614
rect 516954 86614 517574 122058
rect 516954 86058 516986 86614
rect 517542 86058 517574 86614
rect 516954 50614 517574 86058
rect 516954 50058 516986 50614
rect 517542 50058 517574 50614
rect 516954 14614 517574 50058
rect 516954 14058 516986 14614
rect 517542 14058 517574 14614
rect 498954 -7622 498986 -7066
rect 499542 -7622 499574 -7066
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705242 523826 705798
rect 524382 705242 524414 705798
rect 523794 669454 524414 705242
rect 523794 668898 523826 669454
rect 524382 668898 524414 669454
rect 523794 633454 524414 668898
rect 523794 632898 523826 633454
rect 524382 632898 524414 633454
rect 523794 597454 524414 632898
rect 523794 596898 523826 597454
rect 524382 596898 524414 597454
rect 523794 561454 524414 596898
rect 523794 560898 523826 561454
rect 524382 560898 524414 561454
rect 523794 525454 524414 560898
rect 523794 524898 523826 525454
rect 524382 524898 524414 525454
rect 523794 489454 524414 524898
rect 523794 488898 523826 489454
rect 524382 488898 524414 489454
rect 523794 453454 524414 488898
rect 523794 452898 523826 453454
rect 524382 452898 524414 453454
rect 523794 417454 524414 452898
rect 523794 416898 523826 417454
rect 524382 416898 524414 417454
rect 523794 381454 524414 416898
rect 523794 380898 523826 381454
rect 524382 380898 524414 381454
rect 523794 345454 524414 380898
rect 523794 344898 523826 345454
rect 524382 344898 524414 345454
rect 523794 309454 524414 344898
rect 523794 308898 523826 309454
rect 524382 308898 524414 309454
rect 523794 273454 524414 308898
rect 523794 272898 523826 273454
rect 524382 272898 524414 273454
rect 523794 237454 524414 272898
rect 523794 236898 523826 237454
rect 524382 236898 524414 237454
rect 523794 201454 524414 236898
rect 523794 200898 523826 201454
rect 524382 200898 524414 201454
rect 523794 165454 524414 200898
rect 523794 164898 523826 165454
rect 524382 164898 524414 165454
rect 523794 129454 524414 164898
rect 523794 128898 523826 129454
rect 524382 128898 524414 129454
rect 523794 93454 524414 128898
rect 523794 92898 523826 93454
rect 524382 92898 524414 93454
rect 523794 57454 524414 92898
rect 523794 56898 523826 57454
rect 524382 56898 524414 57454
rect 523794 21454 524414 56898
rect 523794 20898 523826 21454
rect 524382 20898 524414 21454
rect 523794 -1306 524414 20898
rect 523794 -1862 523826 -1306
rect 524382 -1862 524414 -1306
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672618 527546 673174
rect 528102 672618 528134 673174
rect 527514 637174 528134 672618
rect 527514 636618 527546 637174
rect 528102 636618 528134 637174
rect 527514 601174 528134 636618
rect 527514 600618 527546 601174
rect 528102 600618 528134 601174
rect 527514 565174 528134 600618
rect 527514 564618 527546 565174
rect 528102 564618 528134 565174
rect 527514 529174 528134 564618
rect 527514 528618 527546 529174
rect 528102 528618 528134 529174
rect 527514 493174 528134 528618
rect 527514 492618 527546 493174
rect 528102 492618 528134 493174
rect 527514 457174 528134 492618
rect 527514 456618 527546 457174
rect 528102 456618 528134 457174
rect 527514 421174 528134 456618
rect 527514 420618 527546 421174
rect 528102 420618 528134 421174
rect 527514 385174 528134 420618
rect 527514 384618 527546 385174
rect 528102 384618 528134 385174
rect 527514 349174 528134 384618
rect 527514 348618 527546 349174
rect 528102 348618 528134 349174
rect 527514 313174 528134 348618
rect 527514 312618 527546 313174
rect 528102 312618 528134 313174
rect 527514 277174 528134 312618
rect 527514 276618 527546 277174
rect 528102 276618 528134 277174
rect 527514 241174 528134 276618
rect 527514 240618 527546 241174
rect 528102 240618 528134 241174
rect 527514 205174 528134 240618
rect 527514 204618 527546 205174
rect 528102 204618 528134 205174
rect 527514 169174 528134 204618
rect 527514 168618 527546 169174
rect 528102 168618 528134 169174
rect 527514 133174 528134 168618
rect 527514 132618 527546 133174
rect 528102 132618 528134 133174
rect 527514 97174 528134 132618
rect 527514 96618 527546 97174
rect 528102 96618 528134 97174
rect 527514 61174 528134 96618
rect 527514 60618 527546 61174
rect 528102 60618 528134 61174
rect 527514 25174 528134 60618
rect 527514 24618 527546 25174
rect 528102 24618 528134 25174
rect 527514 -3226 528134 24618
rect 527514 -3782 527546 -3226
rect 528102 -3782 528134 -3226
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676338 531266 676894
rect 531822 676338 531854 676894
rect 531234 640894 531854 676338
rect 531234 640338 531266 640894
rect 531822 640338 531854 640894
rect 531234 604894 531854 640338
rect 531234 604338 531266 604894
rect 531822 604338 531854 604894
rect 531234 568894 531854 604338
rect 531234 568338 531266 568894
rect 531822 568338 531854 568894
rect 531234 532894 531854 568338
rect 531234 532338 531266 532894
rect 531822 532338 531854 532894
rect 531234 496894 531854 532338
rect 531234 496338 531266 496894
rect 531822 496338 531854 496894
rect 531234 460894 531854 496338
rect 531234 460338 531266 460894
rect 531822 460338 531854 460894
rect 531234 424894 531854 460338
rect 531234 424338 531266 424894
rect 531822 424338 531854 424894
rect 531234 388894 531854 424338
rect 531234 388338 531266 388894
rect 531822 388338 531854 388894
rect 531234 352894 531854 388338
rect 531234 352338 531266 352894
rect 531822 352338 531854 352894
rect 531234 316894 531854 352338
rect 531234 316338 531266 316894
rect 531822 316338 531854 316894
rect 531234 280894 531854 316338
rect 531234 280338 531266 280894
rect 531822 280338 531854 280894
rect 531234 244894 531854 280338
rect 531234 244338 531266 244894
rect 531822 244338 531854 244894
rect 531234 208894 531854 244338
rect 531234 208338 531266 208894
rect 531822 208338 531854 208894
rect 531234 172894 531854 208338
rect 531234 172338 531266 172894
rect 531822 172338 531854 172894
rect 531234 136894 531854 172338
rect 531234 136338 531266 136894
rect 531822 136338 531854 136894
rect 531234 100894 531854 136338
rect 531234 100338 531266 100894
rect 531822 100338 531854 100894
rect 531234 64894 531854 100338
rect 531234 64338 531266 64894
rect 531822 64338 531854 64894
rect 531234 28894 531854 64338
rect 531234 28338 531266 28894
rect 531822 28338 531854 28894
rect 531234 -5146 531854 28338
rect 531234 -5702 531266 -5146
rect 531822 -5702 531854 -5146
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710042 552986 710598
rect 553542 710042 553574 710598
rect 549234 708678 549854 709670
rect 549234 708122 549266 708678
rect 549822 708122 549854 708678
rect 545514 706758 546134 707750
rect 545514 706202 545546 706758
rect 546102 706202 546134 706758
rect 534954 680058 534986 680614
rect 535542 680058 535574 680614
rect 534954 644614 535574 680058
rect 534954 644058 534986 644614
rect 535542 644058 535574 644614
rect 534954 608614 535574 644058
rect 534954 608058 534986 608614
rect 535542 608058 535574 608614
rect 534954 572614 535574 608058
rect 534954 572058 534986 572614
rect 535542 572058 535574 572614
rect 534954 536614 535574 572058
rect 534954 536058 534986 536614
rect 535542 536058 535574 536614
rect 534954 500614 535574 536058
rect 534954 500058 534986 500614
rect 535542 500058 535574 500614
rect 534954 464614 535574 500058
rect 534954 464058 534986 464614
rect 535542 464058 535574 464614
rect 534954 428614 535574 464058
rect 534954 428058 534986 428614
rect 535542 428058 535574 428614
rect 534954 392614 535574 428058
rect 534954 392058 534986 392614
rect 535542 392058 535574 392614
rect 534954 356614 535574 392058
rect 534954 356058 534986 356614
rect 535542 356058 535574 356614
rect 534954 320614 535574 356058
rect 534954 320058 534986 320614
rect 535542 320058 535574 320614
rect 534954 284614 535574 320058
rect 534954 284058 534986 284614
rect 535542 284058 535574 284614
rect 534954 248614 535574 284058
rect 534954 248058 534986 248614
rect 535542 248058 535574 248614
rect 534954 212614 535574 248058
rect 534954 212058 534986 212614
rect 535542 212058 535574 212614
rect 534954 176614 535574 212058
rect 534954 176058 534986 176614
rect 535542 176058 535574 176614
rect 534954 140614 535574 176058
rect 534954 140058 534986 140614
rect 535542 140058 535574 140614
rect 534954 104614 535574 140058
rect 534954 104058 534986 104614
rect 535542 104058 535574 104614
rect 534954 68614 535574 104058
rect 534954 68058 534986 68614
rect 535542 68058 535574 68614
rect 534954 32614 535574 68058
rect 534954 32058 534986 32614
rect 535542 32058 535574 32614
rect 516954 -6662 516986 -6106
rect 517542 -6662 517574 -6106
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704282 541826 704838
rect 542382 704282 542414 704838
rect 541794 687454 542414 704282
rect 541794 686898 541826 687454
rect 542382 686898 542414 687454
rect 541794 651454 542414 686898
rect 541794 650898 541826 651454
rect 542382 650898 542414 651454
rect 541794 615454 542414 650898
rect 541794 614898 541826 615454
rect 542382 614898 542414 615454
rect 541794 579454 542414 614898
rect 541794 578898 541826 579454
rect 542382 578898 542414 579454
rect 541794 543454 542414 578898
rect 541794 542898 541826 543454
rect 542382 542898 542414 543454
rect 541794 507454 542414 542898
rect 541794 506898 541826 507454
rect 542382 506898 542414 507454
rect 541794 471454 542414 506898
rect 541794 470898 541826 471454
rect 542382 470898 542414 471454
rect 541794 435454 542414 470898
rect 541794 434898 541826 435454
rect 542382 434898 542414 435454
rect 541794 399454 542414 434898
rect 541794 398898 541826 399454
rect 542382 398898 542414 399454
rect 541794 363454 542414 398898
rect 541794 362898 541826 363454
rect 542382 362898 542414 363454
rect 541794 327454 542414 362898
rect 541794 326898 541826 327454
rect 542382 326898 542414 327454
rect 541794 291454 542414 326898
rect 541794 290898 541826 291454
rect 542382 290898 542414 291454
rect 541794 255454 542414 290898
rect 541794 254898 541826 255454
rect 542382 254898 542414 255454
rect 541794 219454 542414 254898
rect 541794 218898 541826 219454
rect 542382 218898 542414 219454
rect 541794 183454 542414 218898
rect 541794 182898 541826 183454
rect 542382 182898 542414 183454
rect 541794 147454 542414 182898
rect 541794 146898 541826 147454
rect 542382 146898 542414 147454
rect 541794 111454 542414 146898
rect 541794 110898 541826 111454
rect 542382 110898 542414 111454
rect 541794 75454 542414 110898
rect 541794 74898 541826 75454
rect 542382 74898 542414 75454
rect 541794 39454 542414 74898
rect 541794 38898 541826 39454
rect 542382 38898 542414 39454
rect 541794 3454 542414 38898
rect 541794 2898 541826 3454
rect 542382 2898 542414 3454
rect 541794 -346 542414 2898
rect 541794 -902 541826 -346
rect 542382 -902 542414 -346
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690618 545546 691174
rect 546102 690618 546134 691174
rect 545514 655174 546134 690618
rect 545514 654618 545546 655174
rect 546102 654618 546134 655174
rect 545514 619174 546134 654618
rect 545514 618618 545546 619174
rect 546102 618618 546134 619174
rect 545514 583174 546134 618618
rect 545514 582618 545546 583174
rect 546102 582618 546134 583174
rect 545514 547174 546134 582618
rect 545514 546618 545546 547174
rect 546102 546618 546134 547174
rect 545514 511174 546134 546618
rect 545514 510618 545546 511174
rect 546102 510618 546134 511174
rect 545514 475174 546134 510618
rect 545514 474618 545546 475174
rect 546102 474618 546134 475174
rect 545514 439174 546134 474618
rect 545514 438618 545546 439174
rect 546102 438618 546134 439174
rect 545514 403174 546134 438618
rect 545514 402618 545546 403174
rect 546102 402618 546134 403174
rect 545514 367174 546134 402618
rect 545514 366618 545546 367174
rect 546102 366618 546134 367174
rect 545514 331174 546134 366618
rect 545514 330618 545546 331174
rect 546102 330618 546134 331174
rect 545514 295174 546134 330618
rect 545514 294618 545546 295174
rect 546102 294618 546134 295174
rect 545514 259174 546134 294618
rect 545514 258618 545546 259174
rect 546102 258618 546134 259174
rect 545514 223174 546134 258618
rect 545514 222618 545546 223174
rect 546102 222618 546134 223174
rect 545514 187174 546134 222618
rect 545514 186618 545546 187174
rect 546102 186618 546134 187174
rect 545514 151174 546134 186618
rect 545514 150618 545546 151174
rect 546102 150618 546134 151174
rect 545514 115174 546134 150618
rect 545514 114618 545546 115174
rect 546102 114618 546134 115174
rect 545514 79174 546134 114618
rect 545514 78618 545546 79174
rect 546102 78618 546134 79174
rect 545514 43174 546134 78618
rect 545514 42618 545546 43174
rect 546102 42618 546134 43174
rect 545514 7174 546134 42618
rect 545514 6618 545546 7174
rect 546102 6618 546134 7174
rect 545514 -2266 546134 6618
rect 545514 -2822 545546 -2266
rect 546102 -2822 546134 -2266
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694338 549266 694894
rect 549822 694338 549854 694894
rect 549234 658894 549854 694338
rect 549234 658338 549266 658894
rect 549822 658338 549854 658894
rect 549234 622894 549854 658338
rect 549234 622338 549266 622894
rect 549822 622338 549854 622894
rect 549234 586894 549854 622338
rect 549234 586338 549266 586894
rect 549822 586338 549854 586894
rect 549234 550894 549854 586338
rect 549234 550338 549266 550894
rect 549822 550338 549854 550894
rect 549234 514894 549854 550338
rect 549234 514338 549266 514894
rect 549822 514338 549854 514894
rect 549234 478894 549854 514338
rect 549234 478338 549266 478894
rect 549822 478338 549854 478894
rect 549234 442894 549854 478338
rect 549234 442338 549266 442894
rect 549822 442338 549854 442894
rect 549234 406894 549854 442338
rect 549234 406338 549266 406894
rect 549822 406338 549854 406894
rect 549234 370894 549854 406338
rect 549234 370338 549266 370894
rect 549822 370338 549854 370894
rect 549234 334894 549854 370338
rect 549234 334338 549266 334894
rect 549822 334338 549854 334894
rect 549234 298894 549854 334338
rect 549234 298338 549266 298894
rect 549822 298338 549854 298894
rect 549234 262894 549854 298338
rect 549234 262338 549266 262894
rect 549822 262338 549854 262894
rect 549234 226894 549854 262338
rect 549234 226338 549266 226894
rect 549822 226338 549854 226894
rect 549234 190894 549854 226338
rect 549234 190338 549266 190894
rect 549822 190338 549854 190894
rect 549234 154894 549854 190338
rect 549234 154338 549266 154894
rect 549822 154338 549854 154894
rect 549234 118894 549854 154338
rect 549234 118338 549266 118894
rect 549822 118338 549854 118894
rect 549234 82894 549854 118338
rect 549234 82338 549266 82894
rect 549822 82338 549854 82894
rect 549234 46894 549854 82338
rect 549234 46338 549266 46894
rect 549822 46338 549854 46894
rect 549234 10894 549854 46338
rect 549234 10338 549266 10894
rect 549822 10338 549854 10894
rect 549234 -4186 549854 10338
rect 549234 -4742 549266 -4186
rect 549822 -4742 549854 -4186
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711002 570986 711558
rect 571542 711002 571574 711558
rect 567234 709638 567854 709670
rect 567234 709082 567266 709638
rect 567822 709082 567854 709638
rect 563514 707718 564134 707750
rect 563514 707162 563546 707718
rect 564102 707162 564134 707718
rect 552954 698058 552986 698614
rect 553542 698058 553574 698614
rect 552954 662614 553574 698058
rect 552954 662058 552986 662614
rect 553542 662058 553574 662614
rect 552954 626614 553574 662058
rect 552954 626058 552986 626614
rect 553542 626058 553574 626614
rect 552954 590614 553574 626058
rect 552954 590058 552986 590614
rect 553542 590058 553574 590614
rect 552954 554614 553574 590058
rect 552954 554058 552986 554614
rect 553542 554058 553574 554614
rect 552954 518614 553574 554058
rect 552954 518058 552986 518614
rect 553542 518058 553574 518614
rect 552954 482614 553574 518058
rect 552954 482058 552986 482614
rect 553542 482058 553574 482614
rect 552954 446614 553574 482058
rect 552954 446058 552986 446614
rect 553542 446058 553574 446614
rect 552954 410614 553574 446058
rect 552954 410058 552986 410614
rect 553542 410058 553574 410614
rect 552954 374614 553574 410058
rect 552954 374058 552986 374614
rect 553542 374058 553574 374614
rect 552954 338614 553574 374058
rect 552954 338058 552986 338614
rect 553542 338058 553574 338614
rect 552954 302614 553574 338058
rect 552954 302058 552986 302614
rect 553542 302058 553574 302614
rect 552954 266614 553574 302058
rect 552954 266058 552986 266614
rect 553542 266058 553574 266614
rect 552954 230614 553574 266058
rect 552954 230058 552986 230614
rect 553542 230058 553574 230614
rect 552954 194614 553574 230058
rect 552954 194058 552986 194614
rect 553542 194058 553574 194614
rect 552954 158614 553574 194058
rect 552954 158058 552986 158614
rect 553542 158058 553574 158614
rect 552954 122614 553574 158058
rect 552954 122058 552986 122614
rect 553542 122058 553574 122614
rect 552954 86614 553574 122058
rect 552954 86058 552986 86614
rect 553542 86058 553574 86614
rect 552954 50614 553574 86058
rect 552954 50058 552986 50614
rect 553542 50058 553574 50614
rect 552954 14614 553574 50058
rect 552954 14058 552986 14614
rect 553542 14058 553574 14614
rect 534954 -7622 534986 -7066
rect 535542 -7622 535574 -7066
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705242 559826 705798
rect 560382 705242 560414 705798
rect 559794 669454 560414 705242
rect 559794 668898 559826 669454
rect 560382 668898 560414 669454
rect 559794 633454 560414 668898
rect 559794 632898 559826 633454
rect 560382 632898 560414 633454
rect 559794 597454 560414 632898
rect 559794 596898 559826 597454
rect 560382 596898 560414 597454
rect 559794 561454 560414 596898
rect 559794 560898 559826 561454
rect 560382 560898 560414 561454
rect 559794 525454 560414 560898
rect 559794 524898 559826 525454
rect 560382 524898 560414 525454
rect 559794 489454 560414 524898
rect 559794 488898 559826 489454
rect 560382 488898 560414 489454
rect 559794 453454 560414 488898
rect 559794 452898 559826 453454
rect 560382 452898 560414 453454
rect 559794 417454 560414 452898
rect 559794 416898 559826 417454
rect 560382 416898 560414 417454
rect 559794 381454 560414 416898
rect 559794 380898 559826 381454
rect 560382 380898 560414 381454
rect 559794 345454 560414 380898
rect 559794 344898 559826 345454
rect 560382 344898 560414 345454
rect 559794 309454 560414 344898
rect 559794 308898 559826 309454
rect 560382 308898 560414 309454
rect 559794 273454 560414 308898
rect 559794 272898 559826 273454
rect 560382 272898 560414 273454
rect 559794 237454 560414 272898
rect 559794 236898 559826 237454
rect 560382 236898 560414 237454
rect 559794 201454 560414 236898
rect 559794 200898 559826 201454
rect 560382 200898 560414 201454
rect 559794 165454 560414 200898
rect 559794 164898 559826 165454
rect 560382 164898 560414 165454
rect 559794 129454 560414 164898
rect 559794 128898 559826 129454
rect 560382 128898 560414 129454
rect 559794 93454 560414 128898
rect 559794 92898 559826 93454
rect 560382 92898 560414 93454
rect 559794 57454 560414 92898
rect 559794 56898 559826 57454
rect 560382 56898 560414 57454
rect 559794 21454 560414 56898
rect 559794 20898 559826 21454
rect 560382 20898 560414 21454
rect 559794 -1306 560414 20898
rect 559794 -1862 559826 -1306
rect 560382 -1862 560414 -1306
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672618 563546 673174
rect 564102 672618 564134 673174
rect 563514 637174 564134 672618
rect 563514 636618 563546 637174
rect 564102 636618 564134 637174
rect 563514 601174 564134 636618
rect 563514 600618 563546 601174
rect 564102 600618 564134 601174
rect 563514 565174 564134 600618
rect 563514 564618 563546 565174
rect 564102 564618 564134 565174
rect 563514 529174 564134 564618
rect 563514 528618 563546 529174
rect 564102 528618 564134 529174
rect 563514 493174 564134 528618
rect 563514 492618 563546 493174
rect 564102 492618 564134 493174
rect 563514 457174 564134 492618
rect 563514 456618 563546 457174
rect 564102 456618 564134 457174
rect 563514 421174 564134 456618
rect 563514 420618 563546 421174
rect 564102 420618 564134 421174
rect 563514 385174 564134 420618
rect 563514 384618 563546 385174
rect 564102 384618 564134 385174
rect 563514 349174 564134 384618
rect 563514 348618 563546 349174
rect 564102 348618 564134 349174
rect 563514 313174 564134 348618
rect 563514 312618 563546 313174
rect 564102 312618 564134 313174
rect 563514 277174 564134 312618
rect 563514 276618 563546 277174
rect 564102 276618 564134 277174
rect 563514 241174 564134 276618
rect 563514 240618 563546 241174
rect 564102 240618 564134 241174
rect 563514 205174 564134 240618
rect 563514 204618 563546 205174
rect 564102 204618 564134 205174
rect 563514 169174 564134 204618
rect 563514 168618 563546 169174
rect 564102 168618 564134 169174
rect 563514 133174 564134 168618
rect 563514 132618 563546 133174
rect 564102 132618 564134 133174
rect 563514 97174 564134 132618
rect 563514 96618 563546 97174
rect 564102 96618 564134 97174
rect 563514 61174 564134 96618
rect 563514 60618 563546 61174
rect 564102 60618 564134 61174
rect 563514 25174 564134 60618
rect 563514 24618 563546 25174
rect 564102 24618 564134 25174
rect 563514 -3226 564134 24618
rect 563514 -3782 563546 -3226
rect 564102 -3782 564134 -3226
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676338 567266 676894
rect 567822 676338 567854 676894
rect 567234 640894 567854 676338
rect 567234 640338 567266 640894
rect 567822 640338 567854 640894
rect 567234 604894 567854 640338
rect 567234 604338 567266 604894
rect 567822 604338 567854 604894
rect 567234 568894 567854 604338
rect 567234 568338 567266 568894
rect 567822 568338 567854 568894
rect 567234 532894 567854 568338
rect 567234 532338 567266 532894
rect 567822 532338 567854 532894
rect 567234 496894 567854 532338
rect 567234 496338 567266 496894
rect 567822 496338 567854 496894
rect 567234 460894 567854 496338
rect 567234 460338 567266 460894
rect 567822 460338 567854 460894
rect 567234 424894 567854 460338
rect 567234 424338 567266 424894
rect 567822 424338 567854 424894
rect 567234 388894 567854 424338
rect 567234 388338 567266 388894
rect 567822 388338 567854 388894
rect 567234 352894 567854 388338
rect 567234 352338 567266 352894
rect 567822 352338 567854 352894
rect 567234 316894 567854 352338
rect 567234 316338 567266 316894
rect 567822 316338 567854 316894
rect 567234 280894 567854 316338
rect 567234 280338 567266 280894
rect 567822 280338 567854 280894
rect 567234 244894 567854 280338
rect 567234 244338 567266 244894
rect 567822 244338 567854 244894
rect 567234 208894 567854 244338
rect 567234 208338 567266 208894
rect 567822 208338 567854 208894
rect 567234 172894 567854 208338
rect 567234 172338 567266 172894
rect 567822 172338 567854 172894
rect 567234 136894 567854 172338
rect 567234 136338 567266 136894
rect 567822 136338 567854 136894
rect 567234 100894 567854 136338
rect 567234 100338 567266 100894
rect 567822 100338 567854 100894
rect 567234 64894 567854 100338
rect 567234 64338 567266 64894
rect 567822 64338 567854 64894
rect 567234 28894 567854 64338
rect 567234 28338 567266 28894
rect 567822 28338 567854 28894
rect 567234 -5146 567854 28338
rect 567234 -5702 567266 -5146
rect 567822 -5702 567854 -5146
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711002 592062 711558
rect 592618 711002 592650 711558
rect 591070 710598 591690 710630
rect 591070 710042 591102 710598
rect 591658 710042 591690 710598
rect 590110 709638 590730 709670
rect 590110 709082 590142 709638
rect 590698 709082 590730 709638
rect 589150 708678 589770 708710
rect 589150 708122 589182 708678
rect 589738 708122 589770 708678
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707162 588222 707718
rect 588778 707162 588810 707718
rect 581514 706202 581546 706758
rect 582102 706202 582134 706758
rect 570954 680058 570986 680614
rect 571542 680058 571574 680614
rect 570954 644614 571574 680058
rect 570954 644058 570986 644614
rect 571542 644058 571574 644614
rect 570954 608614 571574 644058
rect 570954 608058 570986 608614
rect 571542 608058 571574 608614
rect 570954 572614 571574 608058
rect 570954 572058 570986 572614
rect 571542 572058 571574 572614
rect 570954 536614 571574 572058
rect 570954 536058 570986 536614
rect 571542 536058 571574 536614
rect 570954 500614 571574 536058
rect 570954 500058 570986 500614
rect 571542 500058 571574 500614
rect 570954 464614 571574 500058
rect 570954 464058 570986 464614
rect 571542 464058 571574 464614
rect 570954 428614 571574 464058
rect 570954 428058 570986 428614
rect 571542 428058 571574 428614
rect 570954 392614 571574 428058
rect 570954 392058 570986 392614
rect 571542 392058 571574 392614
rect 570954 356614 571574 392058
rect 570954 356058 570986 356614
rect 571542 356058 571574 356614
rect 570954 320614 571574 356058
rect 570954 320058 570986 320614
rect 571542 320058 571574 320614
rect 570954 284614 571574 320058
rect 570954 284058 570986 284614
rect 571542 284058 571574 284614
rect 570954 248614 571574 284058
rect 570954 248058 570986 248614
rect 571542 248058 571574 248614
rect 570954 212614 571574 248058
rect 570954 212058 570986 212614
rect 571542 212058 571574 212614
rect 570954 176614 571574 212058
rect 570954 176058 570986 176614
rect 571542 176058 571574 176614
rect 570954 140614 571574 176058
rect 570954 140058 570986 140614
rect 571542 140058 571574 140614
rect 570954 104614 571574 140058
rect 570954 104058 570986 104614
rect 571542 104058 571574 104614
rect 570954 68614 571574 104058
rect 570954 68058 570986 68614
rect 571542 68058 571574 68614
rect 570954 32614 571574 68058
rect 570954 32058 570986 32614
rect 571542 32058 571574 32614
rect 552954 -6662 552986 -6106
rect 553542 -6662 553574 -6106
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704282 577826 704838
rect 578382 704282 578414 704838
rect 577794 687454 578414 704282
rect 577794 686898 577826 687454
rect 578382 686898 578414 687454
rect 577794 651454 578414 686898
rect 577794 650898 577826 651454
rect 578382 650898 578414 651454
rect 577794 615454 578414 650898
rect 577794 614898 577826 615454
rect 578382 614898 578414 615454
rect 577794 579454 578414 614898
rect 577794 578898 577826 579454
rect 578382 578898 578414 579454
rect 577794 543454 578414 578898
rect 577794 542898 577826 543454
rect 578382 542898 578414 543454
rect 577794 507454 578414 542898
rect 577794 506898 577826 507454
rect 578382 506898 578414 507454
rect 577794 471454 578414 506898
rect 577794 470898 577826 471454
rect 578382 470898 578414 471454
rect 577794 435454 578414 470898
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706202 587262 706758
rect 587818 706202 587850 706758
rect 586270 705798 586890 705830
rect 586270 705242 586302 705798
rect 586858 705242 586890 705798
rect 581514 690618 581546 691174
rect 582102 690618 582134 691174
rect 581514 655174 582134 690618
rect 581514 654618 581546 655174
rect 582102 654618 582134 655174
rect 581514 619174 582134 654618
rect 581514 618618 581546 619174
rect 582102 618618 582134 619174
rect 581514 583174 582134 618618
rect 581514 582618 581546 583174
rect 582102 582618 582134 583174
rect 581514 547174 582134 582618
rect 581514 546618 581546 547174
rect 582102 546618 582134 547174
rect 581514 511174 582134 546618
rect 581514 510618 581546 511174
rect 582102 510618 582134 511174
rect 581514 475174 582134 510618
rect 581514 474618 581546 475174
rect 582102 474618 582134 475174
rect 580395 458692 580461 458693
rect 580395 458628 580396 458692
rect 580460 458628 580461 458692
rect 580395 458627 580461 458628
rect 580211 458556 580277 458557
rect 580211 458492 580212 458556
rect 580276 458492 580277 458556
rect 580211 458491 580277 458492
rect 577794 434898 577826 435454
rect 578382 434898 578414 435454
rect 577794 399454 578414 434898
rect 577794 398898 577826 399454
rect 578382 398898 578414 399454
rect 577794 363454 578414 398898
rect 577794 362898 577826 363454
rect 578382 362898 578414 363454
rect 577794 327454 578414 362898
rect 577794 326898 577826 327454
rect 578382 326898 578414 327454
rect 577794 291454 578414 326898
rect 577794 290898 577826 291454
rect 578382 290898 578414 291454
rect 577794 255454 578414 290898
rect 577794 254898 577826 255454
rect 578382 254898 578414 255454
rect 577794 219454 578414 254898
rect 577794 218898 577826 219454
rect 578382 218898 578414 219454
rect 577794 183454 578414 218898
rect 577794 182898 577826 183454
rect 578382 182898 578414 183454
rect 577794 147454 578414 182898
rect 577794 146898 577826 147454
rect 578382 146898 578414 147454
rect 577794 111454 578414 146898
rect 577794 110898 577826 111454
rect 578382 110898 578414 111454
rect 577794 75454 578414 110898
rect 577794 74898 577826 75454
rect 578382 74898 578414 75454
rect 577794 39454 578414 74898
rect 580214 46341 580274 458491
rect 580398 86189 580458 458627
rect 581514 439174 582134 474618
rect 581514 438618 581546 439174
rect 582102 438618 582134 439174
rect 581514 403174 582134 438618
rect 581514 402618 581546 403174
rect 582102 402618 582134 403174
rect 581514 367174 582134 402618
rect 581514 366618 581546 367174
rect 582102 366618 582134 367174
rect 581514 331174 582134 366618
rect 581514 330618 581546 331174
rect 582102 330618 582134 331174
rect 581514 295174 582134 330618
rect 581514 294618 581546 295174
rect 582102 294618 582134 295174
rect 581514 259174 582134 294618
rect 581514 258618 581546 259174
rect 582102 258618 582134 259174
rect 581514 223174 582134 258618
rect 581514 222618 581546 223174
rect 582102 222618 582134 223174
rect 581514 187174 582134 222618
rect 581514 186618 581546 187174
rect 582102 186618 582134 187174
rect 581514 151174 582134 186618
rect 581514 150618 581546 151174
rect 582102 150618 582134 151174
rect 581514 115174 582134 150618
rect 581514 114618 581546 115174
rect 582102 114618 582134 115174
rect 580395 86188 580461 86189
rect 580395 86124 580396 86188
rect 580460 86124 580461 86188
rect 580395 86123 580461 86124
rect 581514 79174 582134 114618
rect 581514 78618 581546 79174
rect 582102 78618 582134 79174
rect 580211 46340 580277 46341
rect 580211 46276 580212 46340
rect 580276 46276 580277 46340
rect 580211 46275 580277 46276
rect 577794 38898 577826 39454
rect 578382 38898 578414 39454
rect 577794 3454 578414 38898
rect 577794 2898 577826 3454
rect 578382 2898 578414 3454
rect 577794 -346 578414 2898
rect 577794 -902 577826 -346
rect 578382 -902 578414 -346
rect 577794 -1894 578414 -902
rect 581514 43174 582134 78618
rect 581514 42618 581546 43174
rect 582102 42618 582134 43174
rect 581514 7174 582134 42618
rect 581514 6618 581546 7174
rect 582102 6618 582134 7174
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704282 585342 704838
rect 585898 704282 585930 704838
rect 585310 687454 585930 704282
rect 585310 686898 585342 687454
rect 585898 686898 585930 687454
rect 585310 651454 585930 686898
rect 585310 650898 585342 651454
rect 585898 650898 585930 651454
rect 585310 615454 585930 650898
rect 585310 614898 585342 615454
rect 585898 614898 585930 615454
rect 585310 579454 585930 614898
rect 585310 578898 585342 579454
rect 585898 578898 585930 579454
rect 585310 543454 585930 578898
rect 585310 542898 585342 543454
rect 585898 542898 585930 543454
rect 585310 507454 585930 542898
rect 585310 506898 585342 507454
rect 585898 506898 585930 507454
rect 585310 471454 585930 506898
rect 585310 470898 585342 471454
rect 585898 470898 585930 471454
rect 585310 435454 585930 470898
rect 585310 434898 585342 435454
rect 585898 434898 585930 435454
rect 585310 399454 585930 434898
rect 585310 398898 585342 399454
rect 585898 398898 585930 399454
rect 585310 363454 585930 398898
rect 585310 362898 585342 363454
rect 585898 362898 585930 363454
rect 585310 327454 585930 362898
rect 585310 326898 585342 327454
rect 585898 326898 585930 327454
rect 585310 291454 585930 326898
rect 585310 290898 585342 291454
rect 585898 290898 585930 291454
rect 585310 255454 585930 290898
rect 585310 254898 585342 255454
rect 585898 254898 585930 255454
rect 585310 219454 585930 254898
rect 585310 218898 585342 219454
rect 585898 218898 585930 219454
rect 585310 183454 585930 218898
rect 585310 182898 585342 183454
rect 585898 182898 585930 183454
rect 585310 147454 585930 182898
rect 585310 146898 585342 147454
rect 585898 146898 585930 147454
rect 585310 111454 585930 146898
rect 585310 110898 585342 111454
rect 585898 110898 585930 111454
rect 585310 75454 585930 110898
rect 585310 74898 585342 75454
rect 585898 74898 585930 75454
rect 585310 39454 585930 74898
rect 585310 38898 585342 39454
rect 585898 38898 585930 39454
rect 585310 3454 585930 38898
rect 585310 2898 585342 3454
rect 585898 2898 585930 3454
rect 585310 -346 585930 2898
rect 585310 -902 585342 -346
rect 585898 -902 585930 -346
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 668898 586302 669454
rect 586858 668898 586890 669454
rect 586270 633454 586890 668898
rect 586270 632898 586302 633454
rect 586858 632898 586890 633454
rect 586270 597454 586890 632898
rect 586270 596898 586302 597454
rect 586858 596898 586890 597454
rect 586270 561454 586890 596898
rect 586270 560898 586302 561454
rect 586858 560898 586890 561454
rect 586270 525454 586890 560898
rect 586270 524898 586302 525454
rect 586858 524898 586890 525454
rect 586270 489454 586890 524898
rect 586270 488898 586302 489454
rect 586858 488898 586890 489454
rect 586270 453454 586890 488898
rect 586270 452898 586302 453454
rect 586858 452898 586890 453454
rect 586270 417454 586890 452898
rect 586270 416898 586302 417454
rect 586858 416898 586890 417454
rect 586270 381454 586890 416898
rect 586270 380898 586302 381454
rect 586858 380898 586890 381454
rect 586270 345454 586890 380898
rect 586270 344898 586302 345454
rect 586858 344898 586890 345454
rect 586270 309454 586890 344898
rect 586270 308898 586302 309454
rect 586858 308898 586890 309454
rect 586270 273454 586890 308898
rect 586270 272898 586302 273454
rect 586858 272898 586890 273454
rect 586270 237454 586890 272898
rect 586270 236898 586302 237454
rect 586858 236898 586890 237454
rect 586270 201454 586890 236898
rect 586270 200898 586302 201454
rect 586858 200898 586890 201454
rect 586270 165454 586890 200898
rect 586270 164898 586302 165454
rect 586858 164898 586890 165454
rect 586270 129454 586890 164898
rect 586270 128898 586302 129454
rect 586858 128898 586890 129454
rect 586270 93454 586890 128898
rect 586270 92898 586302 93454
rect 586858 92898 586890 93454
rect 586270 57454 586890 92898
rect 586270 56898 586302 57454
rect 586858 56898 586890 57454
rect 586270 21454 586890 56898
rect 586270 20898 586302 21454
rect 586858 20898 586890 21454
rect 586270 -1306 586890 20898
rect 586270 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690618 587262 691174
rect 587818 690618 587850 691174
rect 587230 655174 587850 690618
rect 587230 654618 587262 655174
rect 587818 654618 587850 655174
rect 587230 619174 587850 654618
rect 587230 618618 587262 619174
rect 587818 618618 587850 619174
rect 587230 583174 587850 618618
rect 587230 582618 587262 583174
rect 587818 582618 587850 583174
rect 587230 547174 587850 582618
rect 587230 546618 587262 547174
rect 587818 546618 587850 547174
rect 587230 511174 587850 546618
rect 587230 510618 587262 511174
rect 587818 510618 587850 511174
rect 587230 475174 587850 510618
rect 587230 474618 587262 475174
rect 587818 474618 587850 475174
rect 587230 439174 587850 474618
rect 587230 438618 587262 439174
rect 587818 438618 587850 439174
rect 587230 403174 587850 438618
rect 587230 402618 587262 403174
rect 587818 402618 587850 403174
rect 587230 367174 587850 402618
rect 587230 366618 587262 367174
rect 587818 366618 587850 367174
rect 587230 331174 587850 366618
rect 587230 330618 587262 331174
rect 587818 330618 587850 331174
rect 587230 295174 587850 330618
rect 587230 294618 587262 295174
rect 587818 294618 587850 295174
rect 587230 259174 587850 294618
rect 587230 258618 587262 259174
rect 587818 258618 587850 259174
rect 587230 223174 587850 258618
rect 587230 222618 587262 223174
rect 587818 222618 587850 223174
rect 587230 187174 587850 222618
rect 587230 186618 587262 187174
rect 587818 186618 587850 187174
rect 587230 151174 587850 186618
rect 587230 150618 587262 151174
rect 587818 150618 587850 151174
rect 587230 115174 587850 150618
rect 587230 114618 587262 115174
rect 587818 114618 587850 115174
rect 587230 79174 587850 114618
rect 587230 78618 587262 79174
rect 587818 78618 587850 79174
rect 587230 43174 587850 78618
rect 587230 42618 587262 43174
rect 587818 42618 587850 43174
rect 587230 7174 587850 42618
rect 587230 6618 587262 7174
rect 587818 6618 587850 7174
rect 581514 -2822 581546 -2266
rect 582102 -2822 582134 -2266
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672618 588222 673174
rect 588778 672618 588810 673174
rect 588190 637174 588810 672618
rect 588190 636618 588222 637174
rect 588778 636618 588810 637174
rect 588190 601174 588810 636618
rect 588190 600618 588222 601174
rect 588778 600618 588810 601174
rect 588190 565174 588810 600618
rect 588190 564618 588222 565174
rect 588778 564618 588810 565174
rect 588190 529174 588810 564618
rect 588190 528618 588222 529174
rect 588778 528618 588810 529174
rect 588190 493174 588810 528618
rect 588190 492618 588222 493174
rect 588778 492618 588810 493174
rect 588190 457174 588810 492618
rect 588190 456618 588222 457174
rect 588778 456618 588810 457174
rect 588190 421174 588810 456618
rect 588190 420618 588222 421174
rect 588778 420618 588810 421174
rect 588190 385174 588810 420618
rect 588190 384618 588222 385174
rect 588778 384618 588810 385174
rect 588190 349174 588810 384618
rect 588190 348618 588222 349174
rect 588778 348618 588810 349174
rect 588190 313174 588810 348618
rect 588190 312618 588222 313174
rect 588778 312618 588810 313174
rect 588190 277174 588810 312618
rect 588190 276618 588222 277174
rect 588778 276618 588810 277174
rect 588190 241174 588810 276618
rect 588190 240618 588222 241174
rect 588778 240618 588810 241174
rect 588190 205174 588810 240618
rect 588190 204618 588222 205174
rect 588778 204618 588810 205174
rect 588190 169174 588810 204618
rect 588190 168618 588222 169174
rect 588778 168618 588810 169174
rect 588190 133174 588810 168618
rect 588190 132618 588222 133174
rect 588778 132618 588810 133174
rect 588190 97174 588810 132618
rect 588190 96618 588222 97174
rect 588778 96618 588810 97174
rect 588190 61174 588810 96618
rect 588190 60618 588222 61174
rect 588778 60618 588810 61174
rect 588190 25174 588810 60618
rect 588190 24618 588222 25174
rect 588778 24618 588810 25174
rect 588190 -3226 588810 24618
rect 588190 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694338 589182 694894
rect 589738 694338 589770 694894
rect 589150 658894 589770 694338
rect 589150 658338 589182 658894
rect 589738 658338 589770 658894
rect 589150 622894 589770 658338
rect 589150 622338 589182 622894
rect 589738 622338 589770 622894
rect 589150 586894 589770 622338
rect 589150 586338 589182 586894
rect 589738 586338 589770 586894
rect 589150 550894 589770 586338
rect 589150 550338 589182 550894
rect 589738 550338 589770 550894
rect 589150 514894 589770 550338
rect 589150 514338 589182 514894
rect 589738 514338 589770 514894
rect 589150 478894 589770 514338
rect 589150 478338 589182 478894
rect 589738 478338 589770 478894
rect 589150 442894 589770 478338
rect 589150 442338 589182 442894
rect 589738 442338 589770 442894
rect 589150 406894 589770 442338
rect 589150 406338 589182 406894
rect 589738 406338 589770 406894
rect 589150 370894 589770 406338
rect 589150 370338 589182 370894
rect 589738 370338 589770 370894
rect 589150 334894 589770 370338
rect 589150 334338 589182 334894
rect 589738 334338 589770 334894
rect 589150 298894 589770 334338
rect 589150 298338 589182 298894
rect 589738 298338 589770 298894
rect 589150 262894 589770 298338
rect 589150 262338 589182 262894
rect 589738 262338 589770 262894
rect 589150 226894 589770 262338
rect 589150 226338 589182 226894
rect 589738 226338 589770 226894
rect 589150 190894 589770 226338
rect 589150 190338 589182 190894
rect 589738 190338 589770 190894
rect 589150 154894 589770 190338
rect 589150 154338 589182 154894
rect 589738 154338 589770 154894
rect 589150 118894 589770 154338
rect 589150 118338 589182 118894
rect 589738 118338 589770 118894
rect 589150 82894 589770 118338
rect 589150 82338 589182 82894
rect 589738 82338 589770 82894
rect 589150 46894 589770 82338
rect 589150 46338 589182 46894
rect 589738 46338 589770 46894
rect 589150 10894 589770 46338
rect 589150 10338 589182 10894
rect 589738 10338 589770 10894
rect 589150 -4186 589770 10338
rect 589150 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676338 590142 676894
rect 590698 676338 590730 676894
rect 590110 640894 590730 676338
rect 590110 640338 590142 640894
rect 590698 640338 590730 640894
rect 590110 604894 590730 640338
rect 590110 604338 590142 604894
rect 590698 604338 590730 604894
rect 590110 568894 590730 604338
rect 590110 568338 590142 568894
rect 590698 568338 590730 568894
rect 590110 532894 590730 568338
rect 590110 532338 590142 532894
rect 590698 532338 590730 532894
rect 590110 496894 590730 532338
rect 590110 496338 590142 496894
rect 590698 496338 590730 496894
rect 590110 460894 590730 496338
rect 590110 460338 590142 460894
rect 590698 460338 590730 460894
rect 590110 424894 590730 460338
rect 590110 424338 590142 424894
rect 590698 424338 590730 424894
rect 590110 388894 590730 424338
rect 590110 388338 590142 388894
rect 590698 388338 590730 388894
rect 590110 352894 590730 388338
rect 590110 352338 590142 352894
rect 590698 352338 590730 352894
rect 590110 316894 590730 352338
rect 590110 316338 590142 316894
rect 590698 316338 590730 316894
rect 590110 280894 590730 316338
rect 590110 280338 590142 280894
rect 590698 280338 590730 280894
rect 590110 244894 590730 280338
rect 590110 244338 590142 244894
rect 590698 244338 590730 244894
rect 590110 208894 590730 244338
rect 590110 208338 590142 208894
rect 590698 208338 590730 208894
rect 590110 172894 590730 208338
rect 590110 172338 590142 172894
rect 590698 172338 590730 172894
rect 590110 136894 590730 172338
rect 590110 136338 590142 136894
rect 590698 136338 590730 136894
rect 590110 100894 590730 136338
rect 590110 100338 590142 100894
rect 590698 100338 590730 100894
rect 590110 64894 590730 100338
rect 590110 64338 590142 64894
rect 590698 64338 590730 64894
rect 590110 28894 590730 64338
rect 590110 28338 590142 28894
rect 590698 28338 590730 28894
rect 590110 -5146 590730 28338
rect 590110 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698058 591102 698614
rect 591658 698058 591690 698614
rect 591070 662614 591690 698058
rect 591070 662058 591102 662614
rect 591658 662058 591690 662614
rect 591070 626614 591690 662058
rect 591070 626058 591102 626614
rect 591658 626058 591690 626614
rect 591070 590614 591690 626058
rect 591070 590058 591102 590614
rect 591658 590058 591690 590614
rect 591070 554614 591690 590058
rect 591070 554058 591102 554614
rect 591658 554058 591690 554614
rect 591070 518614 591690 554058
rect 591070 518058 591102 518614
rect 591658 518058 591690 518614
rect 591070 482614 591690 518058
rect 591070 482058 591102 482614
rect 591658 482058 591690 482614
rect 591070 446614 591690 482058
rect 591070 446058 591102 446614
rect 591658 446058 591690 446614
rect 591070 410614 591690 446058
rect 591070 410058 591102 410614
rect 591658 410058 591690 410614
rect 591070 374614 591690 410058
rect 591070 374058 591102 374614
rect 591658 374058 591690 374614
rect 591070 338614 591690 374058
rect 591070 338058 591102 338614
rect 591658 338058 591690 338614
rect 591070 302614 591690 338058
rect 591070 302058 591102 302614
rect 591658 302058 591690 302614
rect 591070 266614 591690 302058
rect 591070 266058 591102 266614
rect 591658 266058 591690 266614
rect 591070 230614 591690 266058
rect 591070 230058 591102 230614
rect 591658 230058 591690 230614
rect 591070 194614 591690 230058
rect 591070 194058 591102 194614
rect 591658 194058 591690 194614
rect 591070 158614 591690 194058
rect 591070 158058 591102 158614
rect 591658 158058 591690 158614
rect 591070 122614 591690 158058
rect 591070 122058 591102 122614
rect 591658 122058 591690 122614
rect 591070 86614 591690 122058
rect 591070 86058 591102 86614
rect 591658 86058 591690 86614
rect 591070 50614 591690 86058
rect 591070 50058 591102 50614
rect 591658 50058 591690 50614
rect 591070 14614 591690 50058
rect 591070 14058 591102 14614
rect 591658 14058 591690 14614
rect 591070 -6106 591690 14058
rect 591070 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680058 592062 680614
rect 592618 680058 592650 680614
rect 592030 644614 592650 680058
rect 592030 644058 592062 644614
rect 592618 644058 592650 644614
rect 592030 608614 592650 644058
rect 592030 608058 592062 608614
rect 592618 608058 592650 608614
rect 592030 572614 592650 608058
rect 592030 572058 592062 572614
rect 592618 572058 592650 572614
rect 592030 536614 592650 572058
rect 592030 536058 592062 536614
rect 592618 536058 592650 536614
rect 592030 500614 592650 536058
rect 592030 500058 592062 500614
rect 592618 500058 592650 500614
rect 592030 464614 592650 500058
rect 592030 464058 592062 464614
rect 592618 464058 592650 464614
rect 592030 428614 592650 464058
rect 592030 428058 592062 428614
rect 592618 428058 592650 428614
rect 592030 392614 592650 428058
rect 592030 392058 592062 392614
rect 592618 392058 592650 392614
rect 592030 356614 592650 392058
rect 592030 356058 592062 356614
rect 592618 356058 592650 356614
rect 592030 320614 592650 356058
rect 592030 320058 592062 320614
rect 592618 320058 592650 320614
rect 592030 284614 592650 320058
rect 592030 284058 592062 284614
rect 592618 284058 592650 284614
rect 592030 248614 592650 284058
rect 592030 248058 592062 248614
rect 592618 248058 592650 248614
rect 592030 212614 592650 248058
rect 592030 212058 592062 212614
rect 592618 212058 592650 212614
rect 592030 176614 592650 212058
rect 592030 176058 592062 176614
rect 592618 176058 592650 176614
rect 592030 140614 592650 176058
rect 592030 140058 592062 140614
rect 592618 140058 592650 140614
rect 592030 104614 592650 140058
rect 592030 104058 592062 104614
rect 592618 104058 592650 104614
rect 592030 68614 592650 104058
rect 592030 68058 592062 68614
rect 592618 68058 592650 68614
rect 592030 32614 592650 68058
rect 592030 32058 592062 32614
rect 592618 32058 592650 32614
rect 570954 -7622 570986 -7066
rect 571542 -7622 571574 -7066
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711002 -8138 711558
rect -8694 680058 -8138 680614
rect -8694 644058 -8138 644614
rect -8694 608058 -8138 608614
rect -8694 572058 -8138 572614
rect -8694 536058 -8138 536614
rect -8694 500058 -8138 500614
rect -8694 464058 -8138 464614
rect -8694 428058 -8138 428614
rect -8694 392058 -8138 392614
rect -8694 356058 -8138 356614
rect -8694 320058 -8138 320614
rect -8694 284058 -8138 284614
rect -8694 248058 -8138 248614
rect -8694 212058 -8138 212614
rect -8694 176058 -8138 176614
rect -8694 140058 -8138 140614
rect -8694 104058 -8138 104614
rect -8694 68058 -8138 68614
rect -8694 32058 -8138 32614
rect -7734 710042 -7178 710598
rect 12986 710042 13542 710598
rect -7734 698058 -7178 698614
rect -7734 662058 -7178 662614
rect -7734 626058 -7178 626614
rect -7734 590058 -7178 590614
rect -7734 554058 -7178 554614
rect -7734 518058 -7178 518614
rect -7734 482058 -7178 482614
rect -7734 446058 -7178 446614
rect -7734 410058 -7178 410614
rect -7734 374058 -7178 374614
rect -7734 338058 -7178 338614
rect -7734 302058 -7178 302614
rect -7734 266058 -7178 266614
rect -7734 230058 -7178 230614
rect -7734 194058 -7178 194614
rect -7734 158058 -7178 158614
rect -7734 122058 -7178 122614
rect -7734 86058 -7178 86614
rect -7734 50058 -7178 50614
rect -7734 14058 -7178 14614
rect -6774 709082 -6218 709638
rect -6774 676338 -6218 676894
rect -6774 640338 -6218 640894
rect -6774 604338 -6218 604894
rect -6774 568338 -6218 568894
rect -6774 532338 -6218 532894
rect -6774 496338 -6218 496894
rect -6774 460338 -6218 460894
rect -6774 424338 -6218 424894
rect -6774 388338 -6218 388894
rect -6774 352338 -6218 352894
rect -6774 316338 -6218 316894
rect -6774 280338 -6218 280894
rect -6774 244338 -6218 244894
rect -6774 208338 -6218 208894
rect -6774 172338 -6218 172894
rect -6774 136338 -6218 136894
rect -6774 100338 -6218 100894
rect -6774 64338 -6218 64894
rect -6774 28338 -6218 28894
rect -5814 708122 -5258 708678
rect 9266 708122 9822 708678
rect -5814 694338 -5258 694894
rect -5814 658338 -5258 658894
rect -5814 622338 -5258 622894
rect -5814 586338 -5258 586894
rect -5814 550338 -5258 550894
rect -5814 514338 -5258 514894
rect -5814 478338 -5258 478894
rect -5814 442338 -5258 442894
rect -5814 406338 -5258 406894
rect -5814 370338 -5258 370894
rect -5814 334338 -5258 334894
rect -5814 298338 -5258 298894
rect -5814 262338 -5258 262894
rect -5814 226338 -5258 226894
rect -5814 190338 -5258 190894
rect -5814 154338 -5258 154894
rect -5814 118338 -5258 118894
rect -5814 82338 -5258 82894
rect -5814 46338 -5258 46894
rect -5814 10338 -5258 10894
rect -4854 707162 -4298 707718
rect -4854 672618 -4298 673174
rect -4854 636618 -4298 637174
rect -4854 600618 -4298 601174
rect -4854 564618 -4298 565174
rect -4854 528618 -4298 529174
rect -4854 492618 -4298 493174
rect -4854 456618 -4298 457174
rect -4854 420618 -4298 421174
rect -4854 384618 -4298 385174
rect -4854 348618 -4298 349174
rect -4854 312618 -4298 313174
rect -4854 276618 -4298 277174
rect -4854 240618 -4298 241174
rect -4854 204618 -4298 205174
rect -4854 168618 -4298 169174
rect -4854 132618 -4298 133174
rect -4854 96618 -4298 97174
rect -4854 60618 -4298 61174
rect -4854 24618 -4298 25174
rect -3894 706202 -3338 706758
rect 5546 706202 6102 706758
rect -3894 690618 -3338 691174
rect -3894 654618 -3338 655174
rect -3894 618618 -3338 619174
rect -3894 582618 -3338 583174
rect -3894 546618 -3338 547174
rect -3894 510618 -3338 511174
rect -3894 474618 -3338 475174
rect -3894 438618 -3338 439174
rect -3894 402618 -3338 403174
rect -3894 366618 -3338 367174
rect -3894 330618 -3338 331174
rect -3894 294618 -3338 295174
rect -3894 258618 -3338 259174
rect -3894 222618 -3338 223174
rect -3894 186618 -3338 187174
rect -3894 150618 -3338 151174
rect -3894 114618 -3338 115174
rect -3894 78618 -3338 79174
rect -3894 42618 -3338 43174
rect -3894 6618 -3338 7174
rect -2934 705242 -2378 705798
rect -2934 668898 -2378 669454
rect -2934 632898 -2378 633454
rect -2934 596898 -2378 597454
rect -2934 560898 -2378 561454
rect -2934 524898 -2378 525454
rect -2934 488898 -2378 489454
rect -2934 452898 -2378 453454
rect -2934 416898 -2378 417454
rect -2934 380898 -2378 381454
rect -2934 344898 -2378 345454
rect -2934 308898 -2378 309454
rect -2934 272898 -2378 273454
rect -2934 236898 -2378 237454
rect -2934 200898 -2378 201454
rect -2934 164898 -2378 165454
rect -2934 128898 -2378 129454
rect -2934 92898 -2378 93454
rect -2934 56898 -2378 57454
rect -2934 20898 -2378 21454
rect -1974 704282 -1418 704838
rect -1974 686898 -1418 687454
rect -1974 650898 -1418 651454
rect -1974 614898 -1418 615454
rect -1974 578898 -1418 579454
rect -1974 542898 -1418 543454
rect -1974 506898 -1418 507454
rect -1974 470898 -1418 471454
rect -1974 434898 -1418 435454
rect -1974 398898 -1418 399454
rect -1974 362898 -1418 363454
rect -1974 326898 -1418 327454
rect -1974 290898 -1418 291454
rect -1974 254898 -1418 255454
rect -1974 218898 -1418 219454
rect -1974 182898 -1418 183454
rect -1974 146898 -1418 147454
rect -1974 110898 -1418 111454
rect -1974 74898 -1418 75454
rect -1974 38898 -1418 39454
rect -1974 2898 -1418 3454
rect -1974 -902 -1418 -346
rect 1826 704282 2382 704838
rect 1826 686898 2382 687454
rect 1826 650898 2382 651454
rect 1826 614898 2382 615454
rect 1826 578898 2382 579454
rect 1826 542898 2382 543454
rect 1826 506898 2382 507454
rect 1826 470898 2382 471454
rect 5546 690618 6102 691174
rect 5546 654618 6102 655174
rect 5546 618618 6102 619174
rect 5546 582618 6102 583174
rect 5546 546618 6102 547174
rect 5546 510618 6102 511174
rect 5546 474618 6102 475174
rect 1826 434898 2382 435454
rect 1826 398898 2382 399454
rect 1826 362898 2382 363454
rect 1826 326898 2382 327454
rect 1826 290898 2382 291454
rect 1826 254898 2382 255454
rect 1826 218898 2382 219454
rect 1826 182898 2382 183454
rect 1826 146898 2382 147454
rect 1826 110898 2382 111454
rect 5546 438618 6102 439174
rect 5546 402618 6102 403174
rect 5546 366618 6102 367174
rect 5546 330618 6102 331174
rect 5546 294618 6102 295174
rect 5546 258618 6102 259174
rect 5546 222618 6102 223174
rect 5546 186618 6102 187174
rect 5546 150618 6102 151174
rect 5546 114618 6102 115174
rect 1826 74898 2382 75454
rect 1826 38898 2382 39454
rect 1826 2898 2382 3454
rect 1826 -902 2382 -346
rect -2934 -1862 -2378 -1306
rect 5546 78618 6102 79174
rect 5546 42618 6102 43174
rect 5546 6618 6102 7174
rect -3894 -2822 -3338 -2266
rect 5546 -2822 6102 -2266
rect -4854 -3782 -4298 -3226
rect 9266 694338 9822 694894
rect 9266 658338 9822 658894
rect 9266 622338 9822 622894
rect 9266 586338 9822 586894
rect 9266 550338 9822 550894
rect 9266 514338 9822 514894
rect 9266 478338 9822 478894
rect 9266 442338 9822 442894
rect 9266 406338 9822 406894
rect 9266 370338 9822 370894
rect 9266 334338 9822 334894
rect 9266 298338 9822 298894
rect 9266 262338 9822 262894
rect 9266 226338 9822 226894
rect 9266 190338 9822 190894
rect 9266 154338 9822 154894
rect 9266 118338 9822 118894
rect 9266 82338 9822 82894
rect 9266 46338 9822 46894
rect 9266 10338 9822 10894
rect -5814 -4742 -5258 -4186
rect 9266 -4742 9822 -4186
rect -6774 -5702 -6218 -5146
rect 30986 711002 31542 711558
rect 27266 709082 27822 709638
rect 23546 707162 24102 707718
rect 12986 698058 13542 698614
rect 12986 662058 13542 662614
rect 12986 626058 13542 626614
rect 12986 590058 13542 590614
rect 12986 554058 13542 554614
rect 12986 518058 13542 518614
rect 12986 482058 13542 482614
rect 12986 446058 13542 446614
rect 12986 410058 13542 410614
rect 12986 374058 13542 374614
rect 12986 338058 13542 338614
rect 12986 302058 13542 302614
rect 12986 266058 13542 266614
rect 12986 230058 13542 230614
rect 12986 194058 13542 194614
rect 12986 158058 13542 158614
rect 12986 122058 13542 122614
rect 12986 86058 13542 86614
rect 12986 50058 13542 50614
rect 12986 14058 13542 14614
rect -7734 -6662 -7178 -6106
rect 19826 705242 20382 705798
rect 19826 668898 20382 669454
rect 19826 632898 20382 633454
rect 19826 596898 20382 597454
rect 19826 560898 20382 561454
rect 19826 524898 20382 525454
rect 19826 488898 20382 489454
rect 19826 452898 20382 453454
rect 19826 416898 20382 417454
rect 19826 380898 20382 381454
rect 19826 344898 20382 345454
rect 19826 308898 20382 309454
rect 19826 272898 20382 273454
rect 19826 236898 20382 237454
rect 19826 200898 20382 201454
rect 19826 164898 20382 165454
rect 19826 128898 20382 129454
rect 19826 92898 20382 93454
rect 19826 56898 20382 57454
rect 19826 20898 20382 21454
rect 19826 -1862 20382 -1306
rect 23546 672618 24102 673174
rect 23546 636618 24102 637174
rect 23546 600618 24102 601174
rect 23546 564618 24102 565174
rect 23546 528618 24102 529174
rect 23546 492618 24102 493174
rect 23546 456618 24102 457174
rect 23546 420618 24102 421174
rect 23546 384618 24102 385174
rect 23546 348618 24102 349174
rect 23546 312618 24102 313174
rect 23546 276618 24102 277174
rect 23546 240618 24102 241174
rect 23546 204618 24102 205174
rect 23546 168618 24102 169174
rect 23546 132618 24102 133174
rect 23546 96618 24102 97174
rect 23546 60618 24102 61174
rect 23546 24618 24102 25174
rect 23546 -3782 24102 -3226
rect 27266 676338 27822 676894
rect 27266 640338 27822 640894
rect 27266 604338 27822 604894
rect 27266 568338 27822 568894
rect 27266 532338 27822 532894
rect 27266 496338 27822 496894
rect 27266 460338 27822 460894
rect 27266 424338 27822 424894
rect 27266 388338 27822 388894
rect 27266 352338 27822 352894
rect 27266 316338 27822 316894
rect 27266 280338 27822 280894
rect 27266 244338 27822 244894
rect 27266 208338 27822 208894
rect 27266 172338 27822 172894
rect 27266 136338 27822 136894
rect 27266 100338 27822 100894
rect 27266 64338 27822 64894
rect 27266 28338 27822 28894
rect 27266 -5702 27822 -5146
rect 48986 710042 49542 710598
rect 45266 708122 45822 708678
rect 41546 706202 42102 706758
rect 30986 680058 31542 680614
rect 30986 644058 31542 644614
rect 30986 608058 31542 608614
rect 30986 572058 31542 572614
rect 30986 536058 31542 536614
rect 30986 500058 31542 500614
rect 30986 464058 31542 464614
rect 30986 428058 31542 428614
rect 30986 392058 31542 392614
rect 30986 356058 31542 356614
rect 30986 320058 31542 320614
rect 30986 284058 31542 284614
rect 30986 248058 31542 248614
rect 30986 212058 31542 212614
rect 30986 176058 31542 176614
rect 30986 140058 31542 140614
rect 30986 104058 31542 104614
rect 30986 68058 31542 68614
rect 30986 32058 31542 32614
rect 12986 -6662 13542 -6106
rect -8694 -7622 -8138 -7066
rect 37826 704282 38382 704838
rect 37826 686898 38382 687454
rect 37826 650898 38382 651454
rect 37826 614898 38382 615454
rect 37826 578898 38382 579454
rect 37826 542898 38382 543454
rect 37826 506898 38382 507454
rect 37826 470898 38382 471454
rect 37826 434898 38382 435454
rect 37826 398898 38382 399454
rect 37826 362898 38382 363454
rect 37826 326898 38382 327454
rect 37826 290898 38382 291454
rect 37826 254898 38382 255454
rect 37826 218898 38382 219454
rect 37826 182898 38382 183454
rect 37826 146898 38382 147454
rect 37826 110898 38382 111454
rect 37826 74898 38382 75454
rect 37826 38898 38382 39454
rect 37826 2898 38382 3454
rect 37826 -902 38382 -346
rect 41546 690618 42102 691174
rect 41546 654618 42102 655174
rect 41546 618618 42102 619174
rect 41546 582618 42102 583174
rect 41546 546618 42102 547174
rect 41546 510618 42102 511174
rect 41546 474618 42102 475174
rect 41546 438618 42102 439174
rect 41546 402618 42102 403174
rect 41546 366618 42102 367174
rect 41546 330618 42102 331174
rect 41546 294618 42102 295174
rect 41546 258618 42102 259174
rect 41546 222618 42102 223174
rect 41546 186618 42102 187174
rect 41546 150618 42102 151174
rect 41546 114618 42102 115174
rect 41546 78618 42102 79174
rect 41546 42618 42102 43174
rect 41546 6618 42102 7174
rect 41546 -2822 42102 -2266
rect 45266 694338 45822 694894
rect 45266 658338 45822 658894
rect 45266 622338 45822 622894
rect 45266 586338 45822 586894
rect 45266 550338 45822 550894
rect 45266 514338 45822 514894
rect 45266 478338 45822 478894
rect 45266 442338 45822 442894
rect 45266 406338 45822 406894
rect 45266 370338 45822 370894
rect 45266 334338 45822 334894
rect 45266 298338 45822 298894
rect 45266 262338 45822 262894
rect 45266 226338 45822 226894
rect 45266 190338 45822 190894
rect 45266 154338 45822 154894
rect 45266 118338 45822 118894
rect 45266 82338 45822 82894
rect 45266 46338 45822 46894
rect 45266 10338 45822 10894
rect 45266 -4742 45822 -4186
rect 66986 711002 67542 711558
rect 63266 709082 63822 709638
rect 59546 707162 60102 707718
rect 48986 698058 49542 698614
rect 48986 662058 49542 662614
rect 48986 626058 49542 626614
rect 48986 590058 49542 590614
rect 48986 554058 49542 554614
rect 48986 518058 49542 518614
rect 48986 482058 49542 482614
rect 48986 446058 49542 446614
rect 48986 410058 49542 410614
rect 48986 374058 49542 374614
rect 48986 338058 49542 338614
rect 48986 302058 49542 302614
rect 48986 266058 49542 266614
rect 48986 230058 49542 230614
rect 48986 194058 49542 194614
rect 48986 158058 49542 158614
rect 48986 122058 49542 122614
rect 48986 86058 49542 86614
rect 48986 50058 49542 50614
rect 48986 14058 49542 14614
rect 30986 -7622 31542 -7066
rect 55826 705242 56382 705798
rect 55826 668898 56382 669454
rect 55826 632898 56382 633454
rect 55826 596898 56382 597454
rect 55826 560898 56382 561454
rect 55826 524898 56382 525454
rect 55826 488898 56382 489454
rect 55826 452898 56382 453454
rect 55826 416898 56382 417454
rect 55826 380898 56382 381454
rect 55826 344898 56382 345454
rect 55826 308898 56382 309454
rect 55826 272898 56382 273454
rect 55826 236898 56382 237454
rect 55826 200898 56382 201454
rect 55826 164898 56382 165454
rect 55826 128898 56382 129454
rect 55826 92898 56382 93454
rect 55826 56898 56382 57454
rect 55826 20898 56382 21454
rect 55826 -1862 56382 -1306
rect 59546 672618 60102 673174
rect 59546 636618 60102 637174
rect 59546 600618 60102 601174
rect 59546 564618 60102 565174
rect 59546 528618 60102 529174
rect 59546 492618 60102 493174
rect 59546 456618 60102 457174
rect 59546 420618 60102 421174
rect 59546 384618 60102 385174
rect 59546 348618 60102 349174
rect 59546 312618 60102 313174
rect 59546 276618 60102 277174
rect 59546 240618 60102 241174
rect 59546 204618 60102 205174
rect 59546 168618 60102 169174
rect 59546 132618 60102 133174
rect 59546 96618 60102 97174
rect 59546 60618 60102 61174
rect 59546 24618 60102 25174
rect 59546 -3782 60102 -3226
rect 63266 676338 63822 676894
rect 63266 640338 63822 640894
rect 63266 604338 63822 604894
rect 63266 568338 63822 568894
rect 63266 532338 63822 532894
rect 63266 496338 63822 496894
rect 63266 460338 63822 460894
rect 63266 424338 63822 424894
rect 63266 388338 63822 388894
rect 63266 352338 63822 352894
rect 63266 316338 63822 316894
rect 63266 280338 63822 280894
rect 63266 244338 63822 244894
rect 63266 208338 63822 208894
rect 63266 172338 63822 172894
rect 63266 136338 63822 136894
rect 63266 100338 63822 100894
rect 63266 64338 63822 64894
rect 63266 28338 63822 28894
rect 63266 -5702 63822 -5146
rect 84986 710042 85542 710598
rect 81266 708122 81822 708678
rect 77546 706202 78102 706758
rect 66986 680058 67542 680614
rect 66986 644058 67542 644614
rect 66986 608058 67542 608614
rect 66986 572058 67542 572614
rect 66986 536058 67542 536614
rect 66986 500058 67542 500614
rect 66986 464058 67542 464614
rect 66986 428058 67542 428614
rect 66986 392058 67542 392614
rect 66986 356058 67542 356614
rect 66986 320058 67542 320614
rect 66986 284058 67542 284614
rect 66986 248058 67542 248614
rect 66986 212058 67542 212614
rect 66986 176058 67542 176614
rect 66986 140058 67542 140614
rect 66986 104058 67542 104614
rect 66986 68058 67542 68614
rect 66986 32058 67542 32614
rect 48986 -6662 49542 -6106
rect 73826 704282 74382 704838
rect 73826 686898 74382 687454
rect 73826 650898 74382 651454
rect 73826 614898 74382 615454
rect 73826 578898 74382 579454
rect 73826 542898 74382 543454
rect 73826 506898 74382 507454
rect 73826 470898 74382 471454
rect 73826 434898 74382 435454
rect 73826 398898 74382 399454
rect 73826 362898 74382 363454
rect 73826 326898 74382 327454
rect 73826 290898 74382 291454
rect 73826 254898 74382 255454
rect 73826 218898 74382 219454
rect 73826 182898 74382 183454
rect 73826 146898 74382 147454
rect 73826 110898 74382 111454
rect 73826 74898 74382 75454
rect 73826 38898 74382 39454
rect 73826 2898 74382 3454
rect 73826 -902 74382 -346
rect 77546 690618 78102 691174
rect 77546 654618 78102 655174
rect 77546 618618 78102 619174
rect 77546 582618 78102 583174
rect 77546 546618 78102 547174
rect 77546 510618 78102 511174
rect 77546 474618 78102 475174
rect 77546 438618 78102 439174
rect 77546 402618 78102 403174
rect 77546 366618 78102 367174
rect 77546 330618 78102 331174
rect 77546 294618 78102 295174
rect 77546 258618 78102 259174
rect 77546 222618 78102 223174
rect 77546 186618 78102 187174
rect 77546 150618 78102 151174
rect 77546 114618 78102 115174
rect 77546 78618 78102 79174
rect 77546 42618 78102 43174
rect 77546 6618 78102 7174
rect 77546 -2822 78102 -2266
rect 81266 694338 81822 694894
rect 81266 658338 81822 658894
rect 81266 622338 81822 622894
rect 81266 586338 81822 586894
rect 81266 550338 81822 550894
rect 81266 514338 81822 514894
rect 81266 478338 81822 478894
rect 81266 442338 81822 442894
rect 81266 406338 81822 406894
rect 81266 370338 81822 370894
rect 81266 334338 81822 334894
rect 81266 298338 81822 298894
rect 81266 262338 81822 262894
rect 81266 226338 81822 226894
rect 81266 190338 81822 190894
rect 81266 154338 81822 154894
rect 81266 118338 81822 118894
rect 81266 82338 81822 82894
rect 81266 46338 81822 46894
rect 81266 10338 81822 10894
rect 81266 -4742 81822 -4186
rect 102986 711002 103542 711558
rect 99266 709082 99822 709638
rect 95546 707162 96102 707718
rect 84986 698058 85542 698614
rect 84986 662058 85542 662614
rect 84986 626058 85542 626614
rect 84986 590058 85542 590614
rect 84986 554058 85542 554614
rect 84986 518058 85542 518614
rect 84986 482058 85542 482614
rect 84986 446058 85542 446614
rect 84986 410058 85542 410614
rect 84986 374058 85542 374614
rect 84986 338058 85542 338614
rect 84986 302058 85542 302614
rect 84986 266058 85542 266614
rect 84986 230058 85542 230614
rect 84986 194058 85542 194614
rect 84986 158058 85542 158614
rect 84986 122058 85542 122614
rect 84986 86058 85542 86614
rect 84986 50058 85542 50614
rect 84986 14058 85542 14614
rect 66986 -7622 67542 -7066
rect 91826 705242 92382 705798
rect 91826 668898 92382 669454
rect 91826 632898 92382 633454
rect 91826 596898 92382 597454
rect 91826 560898 92382 561454
rect 91826 524898 92382 525454
rect 91826 488898 92382 489454
rect 91826 452898 92382 453454
rect 91826 416898 92382 417454
rect 91826 380898 92382 381454
rect 91826 344898 92382 345454
rect 91826 308898 92382 309454
rect 91826 272898 92382 273454
rect 91826 236898 92382 237454
rect 91826 200898 92382 201454
rect 91826 164898 92382 165454
rect 91826 128898 92382 129454
rect 91826 92898 92382 93454
rect 91826 56898 92382 57454
rect 91826 20898 92382 21454
rect 91826 -1862 92382 -1306
rect 95546 672618 96102 673174
rect 95546 636618 96102 637174
rect 95546 600618 96102 601174
rect 95546 564618 96102 565174
rect 95546 528618 96102 529174
rect 95546 492618 96102 493174
rect 95546 456618 96102 457174
rect 95546 420618 96102 421174
rect 95546 384618 96102 385174
rect 95546 348618 96102 349174
rect 95546 312618 96102 313174
rect 95546 276618 96102 277174
rect 95546 240618 96102 241174
rect 95546 204618 96102 205174
rect 95546 168618 96102 169174
rect 95546 132618 96102 133174
rect 95546 96618 96102 97174
rect 95546 60618 96102 61174
rect 95546 24618 96102 25174
rect 95546 -3782 96102 -3226
rect 99266 676338 99822 676894
rect 99266 640338 99822 640894
rect 99266 604338 99822 604894
rect 99266 568338 99822 568894
rect 99266 532338 99822 532894
rect 99266 496338 99822 496894
rect 99266 460338 99822 460894
rect 99266 424338 99822 424894
rect 99266 388338 99822 388894
rect 99266 352338 99822 352894
rect 99266 316338 99822 316894
rect 99266 280338 99822 280894
rect 99266 244338 99822 244894
rect 99266 208338 99822 208894
rect 99266 172338 99822 172894
rect 99266 136338 99822 136894
rect 99266 100338 99822 100894
rect 99266 64338 99822 64894
rect 99266 28338 99822 28894
rect 99266 -5702 99822 -5146
rect 120986 710042 121542 710598
rect 117266 708122 117822 708678
rect 113546 706202 114102 706758
rect 102986 680058 103542 680614
rect 102986 644058 103542 644614
rect 102986 608058 103542 608614
rect 102986 572058 103542 572614
rect 102986 536058 103542 536614
rect 102986 500058 103542 500614
rect 102986 464058 103542 464614
rect 102986 428058 103542 428614
rect 102986 392058 103542 392614
rect 102986 356058 103542 356614
rect 102986 320058 103542 320614
rect 102986 284058 103542 284614
rect 102986 248058 103542 248614
rect 102986 212058 103542 212614
rect 102986 176058 103542 176614
rect 102986 140058 103542 140614
rect 102986 104058 103542 104614
rect 102986 68058 103542 68614
rect 102986 32058 103542 32614
rect 84986 -6662 85542 -6106
rect 109826 704282 110382 704838
rect 109826 686898 110382 687454
rect 109826 650898 110382 651454
rect 109826 614898 110382 615454
rect 109826 578898 110382 579454
rect 109826 542898 110382 543454
rect 109826 506898 110382 507454
rect 109826 470898 110382 471454
rect 109826 434898 110382 435454
rect 109826 398898 110382 399454
rect 109826 362898 110382 363454
rect 109826 326898 110382 327454
rect 109826 290898 110382 291454
rect 109826 254898 110382 255454
rect 109826 218898 110382 219454
rect 109826 182898 110382 183454
rect 109826 146898 110382 147454
rect 109826 110898 110382 111454
rect 109826 74898 110382 75454
rect 109826 38898 110382 39454
rect 109826 2898 110382 3454
rect 109826 -902 110382 -346
rect 113546 690618 114102 691174
rect 113546 654618 114102 655174
rect 113546 618618 114102 619174
rect 113546 582618 114102 583174
rect 113546 546618 114102 547174
rect 113546 510618 114102 511174
rect 113546 474618 114102 475174
rect 113546 438618 114102 439174
rect 113546 402618 114102 403174
rect 113546 366618 114102 367174
rect 113546 330618 114102 331174
rect 113546 294618 114102 295174
rect 113546 258618 114102 259174
rect 113546 222618 114102 223174
rect 113546 186618 114102 187174
rect 113546 150618 114102 151174
rect 113546 114618 114102 115174
rect 113546 78618 114102 79174
rect 113546 42618 114102 43174
rect 113546 6618 114102 7174
rect 113546 -2822 114102 -2266
rect 117266 694338 117822 694894
rect 117266 658338 117822 658894
rect 117266 622338 117822 622894
rect 117266 586338 117822 586894
rect 117266 550338 117822 550894
rect 117266 514338 117822 514894
rect 117266 478338 117822 478894
rect 117266 442338 117822 442894
rect 117266 406338 117822 406894
rect 117266 370338 117822 370894
rect 117266 334338 117822 334894
rect 117266 298338 117822 298894
rect 117266 262338 117822 262894
rect 117266 226338 117822 226894
rect 117266 190338 117822 190894
rect 117266 154338 117822 154894
rect 117266 118338 117822 118894
rect 117266 82338 117822 82894
rect 117266 46338 117822 46894
rect 117266 10338 117822 10894
rect 117266 -4742 117822 -4186
rect 138986 711002 139542 711558
rect 135266 709082 135822 709638
rect 131546 707162 132102 707718
rect 120986 698058 121542 698614
rect 120986 662058 121542 662614
rect 120986 626058 121542 626614
rect 120986 590058 121542 590614
rect 120986 554058 121542 554614
rect 120986 518058 121542 518614
rect 120986 482058 121542 482614
rect 120986 446058 121542 446614
rect 120986 410058 121542 410614
rect 120986 374058 121542 374614
rect 120986 338058 121542 338614
rect 120986 302058 121542 302614
rect 120986 266058 121542 266614
rect 120986 230058 121542 230614
rect 120986 194058 121542 194614
rect 120986 158058 121542 158614
rect 120986 122058 121542 122614
rect 120986 86058 121542 86614
rect 120986 50058 121542 50614
rect 120986 14058 121542 14614
rect 102986 -7622 103542 -7066
rect 127826 705242 128382 705798
rect 127826 668898 128382 669454
rect 127826 632898 128382 633454
rect 127826 596898 128382 597454
rect 127826 560898 128382 561454
rect 127826 524898 128382 525454
rect 127826 488898 128382 489454
rect 127826 452898 128382 453454
rect 127826 416898 128382 417454
rect 127826 380898 128382 381454
rect 127826 344898 128382 345454
rect 127826 308898 128382 309454
rect 127826 272898 128382 273454
rect 127826 236898 128382 237454
rect 127826 200898 128382 201454
rect 127826 164898 128382 165454
rect 127826 128898 128382 129454
rect 127826 92898 128382 93454
rect 127826 56898 128382 57454
rect 127826 20898 128382 21454
rect 127826 -1862 128382 -1306
rect 131546 672618 132102 673174
rect 131546 636618 132102 637174
rect 131546 600618 132102 601174
rect 131546 564618 132102 565174
rect 131546 528618 132102 529174
rect 131546 492618 132102 493174
rect 131546 456618 132102 457174
rect 131546 420618 132102 421174
rect 131546 384618 132102 385174
rect 131546 348618 132102 349174
rect 131546 312618 132102 313174
rect 131546 276618 132102 277174
rect 131546 240618 132102 241174
rect 131546 204618 132102 205174
rect 131546 168618 132102 169174
rect 131546 132618 132102 133174
rect 131546 96618 132102 97174
rect 131546 60618 132102 61174
rect 131546 24618 132102 25174
rect 131546 -3782 132102 -3226
rect 135266 676338 135822 676894
rect 135266 640338 135822 640894
rect 135266 604338 135822 604894
rect 135266 568338 135822 568894
rect 135266 532338 135822 532894
rect 135266 496338 135822 496894
rect 135266 460338 135822 460894
rect 135266 424338 135822 424894
rect 135266 388338 135822 388894
rect 135266 352338 135822 352894
rect 135266 316338 135822 316894
rect 135266 280338 135822 280894
rect 135266 244338 135822 244894
rect 135266 208338 135822 208894
rect 135266 172338 135822 172894
rect 135266 136338 135822 136894
rect 135266 100338 135822 100894
rect 135266 64338 135822 64894
rect 135266 28338 135822 28894
rect 135266 -5702 135822 -5146
rect 156986 710042 157542 710598
rect 153266 708122 153822 708678
rect 149546 706202 150102 706758
rect 138986 680058 139542 680614
rect 138986 644058 139542 644614
rect 138986 608058 139542 608614
rect 138986 572058 139542 572614
rect 138986 536058 139542 536614
rect 138986 500058 139542 500614
rect 138986 464058 139542 464614
rect 138986 428058 139542 428614
rect 138986 392058 139542 392614
rect 138986 356058 139542 356614
rect 138986 320058 139542 320614
rect 138986 284058 139542 284614
rect 138986 248058 139542 248614
rect 138986 212058 139542 212614
rect 138986 176058 139542 176614
rect 138986 140058 139542 140614
rect 138986 104058 139542 104614
rect 138986 68058 139542 68614
rect 138986 32058 139542 32614
rect 120986 -6662 121542 -6106
rect 145826 704282 146382 704838
rect 145826 686898 146382 687454
rect 145826 650898 146382 651454
rect 145826 614898 146382 615454
rect 145826 578898 146382 579454
rect 145826 542898 146382 543454
rect 145826 506898 146382 507454
rect 145826 470898 146382 471454
rect 145826 434898 146382 435454
rect 145826 398898 146382 399454
rect 145826 362898 146382 363454
rect 145826 326898 146382 327454
rect 145826 290898 146382 291454
rect 145826 254898 146382 255454
rect 145826 218898 146382 219454
rect 145826 182898 146382 183454
rect 145826 146898 146382 147454
rect 145826 110898 146382 111454
rect 145826 74898 146382 75454
rect 145826 38898 146382 39454
rect 145826 2898 146382 3454
rect 145826 -902 146382 -346
rect 149546 690618 150102 691174
rect 149546 654618 150102 655174
rect 149546 618618 150102 619174
rect 149546 582618 150102 583174
rect 149546 546618 150102 547174
rect 149546 510618 150102 511174
rect 149546 474618 150102 475174
rect 149546 438618 150102 439174
rect 149546 402618 150102 403174
rect 149546 366618 150102 367174
rect 149546 330618 150102 331174
rect 149546 294618 150102 295174
rect 149546 258618 150102 259174
rect 149546 222618 150102 223174
rect 149546 186618 150102 187174
rect 149546 150618 150102 151174
rect 149546 114618 150102 115174
rect 149546 78618 150102 79174
rect 149546 42618 150102 43174
rect 149546 6618 150102 7174
rect 149546 -2822 150102 -2266
rect 153266 694338 153822 694894
rect 153266 658338 153822 658894
rect 153266 622338 153822 622894
rect 153266 586338 153822 586894
rect 153266 550338 153822 550894
rect 153266 514338 153822 514894
rect 153266 478338 153822 478894
rect 153266 442338 153822 442894
rect 153266 406338 153822 406894
rect 153266 370338 153822 370894
rect 153266 334338 153822 334894
rect 153266 298338 153822 298894
rect 153266 262338 153822 262894
rect 153266 226338 153822 226894
rect 153266 190338 153822 190894
rect 153266 154338 153822 154894
rect 153266 118338 153822 118894
rect 153266 82338 153822 82894
rect 153266 46338 153822 46894
rect 153266 10338 153822 10894
rect 153266 -4742 153822 -4186
rect 174986 711002 175542 711558
rect 171266 709082 171822 709638
rect 167546 707162 168102 707718
rect 156986 698058 157542 698614
rect 156986 662058 157542 662614
rect 156986 626058 157542 626614
rect 156986 590058 157542 590614
rect 156986 554058 157542 554614
rect 156986 518058 157542 518614
rect 156986 482058 157542 482614
rect 156986 446058 157542 446614
rect 156986 410058 157542 410614
rect 156986 374058 157542 374614
rect 156986 338058 157542 338614
rect 156986 302058 157542 302614
rect 156986 266058 157542 266614
rect 156986 230058 157542 230614
rect 156986 194058 157542 194614
rect 156986 158058 157542 158614
rect 156986 122058 157542 122614
rect 156986 86058 157542 86614
rect 156986 50058 157542 50614
rect 156986 14058 157542 14614
rect 138986 -7622 139542 -7066
rect 163826 705242 164382 705798
rect 163826 668898 164382 669454
rect 163826 632898 164382 633454
rect 163826 596898 164382 597454
rect 163826 560898 164382 561454
rect 163826 524898 164382 525454
rect 163826 488898 164382 489454
rect 163826 452898 164382 453454
rect 163826 416898 164382 417454
rect 163826 380898 164382 381454
rect 163826 344898 164382 345454
rect 163826 308898 164382 309454
rect 163826 272898 164382 273454
rect 163826 236898 164382 237454
rect 163826 200898 164382 201454
rect 163826 164898 164382 165454
rect 163826 128898 164382 129454
rect 163826 92898 164382 93454
rect 163826 56898 164382 57454
rect 163826 20898 164382 21454
rect 163826 -1862 164382 -1306
rect 167546 672618 168102 673174
rect 167546 636618 168102 637174
rect 167546 600618 168102 601174
rect 167546 564618 168102 565174
rect 167546 528618 168102 529174
rect 167546 492618 168102 493174
rect 167546 456618 168102 457174
rect 167546 420618 168102 421174
rect 167546 384618 168102 385174
rect 167546 348618 168102 349174
rect 167546 312618 168102 313174
rect 167546 276618 168102 277174
rect 167546 240618 168102 241174
rect 167546 204618 168102 205174
rect 167546 168618 168102 169174
rect 167546 132618 168102 133174
rect 167546 96618 168102 97174
rect 167546 60618 168102 61174
rect 167546 24618 168102 25174
rect 167546 -3782 168102 -3226
rect 171266 676338 171822 676894
rect 171266 640338 171822 640894
rect 171266 604338 171822 604894
rect 171266 568338 171822 568894
rect 171266 532338 171822 532894
rect 171266 496338 171822 496894
rect 171266 460338 171822 460894
rect 171266 424338 171822 424894
rect 171266 388338 171822 388894
rect 171266 352338 171822 352894
rect 171266 316338 171822 316894
rect 171266 280338 171822 280894
rect 171266 244338 171822 244894
rect 171266 208338 171822 208894
rect 171266 172338 171822 172894
rect 171266 136338 171822 136894
rect 171266 100338 171822 100894
rect 171266 64338 171822 64894
rect 171266 28338 171822 28894
rect 171266 -5702 171822 -5146
rect 192986 710042 193542 710598
rect 189266 708122 189822 708678
rect 185546 706202 186102 706758
rect 174986 680058 175542 680614
rect 174986 644058 175542 644614
rect 174986 608058 175542 608614
rect 174986 572058 175542 572614
rect 174986 536058 175542 536614
rect 174986 500058 175542 500614
rect 174986 464058 175542 464614
rect 174986 428058 175542 428614
rect 174986 392058 175542 392614
rect 174986 356058 175542 356614
rect 174986 320058 175542 320614
rect 174986 284058 175542 284614
rect 174986 248058 175542 248614
rect 174986 212058 175542 212614
rect 174986 176058 175542 176614
rect 174986 140058 175542 140614
rect 174986 104058 175542 104614
rect 174986 68058 175542 68614
rect 174986 32058 175542 32614
rect 156986 -6662 157542 -6106
rect 181826 704282 182382 704838
rect 181826 686898 182382 687454
rect 181826 650898 182382 651454
rect 181826 614898 182382 615454
rect 181826 578898 182382 579454
rect 181826 542898 182382 543454
rect 181826 506898 182382 507454
rect 181826 470898 182382 471454
rect 181826 434898 182382 435454
rect 181826 398898 182382 399454
rect 181826 362898 182382 363454
rect 181826 326898 182382 327454
rect 181826 290898 182382 291454
rect 181826 254898 182382 255454
rect 181826 218898 182382 219454
rect 181826 182898 182382 183454
rect 181826 146898 182382 147454
rect 181826 110898 182382 111454
rect 181826 74898 182382 75454
rect 181826 38898 182382 39454
rect 181826 2898 182382 3454
rect 181826 -902 182382 -346
rect 185546 690618 186102 691174
rect 185546 654618 186102 655174
rect 185546 618618 186102 619174
rect 185546 582618 186102 583174
rect 185546 546618 186102 547174
rect 185546 510618 186102 511174
rect 185546 474618 186102 475174
rect 185546 438618 186102 439174
rect 185546 402618 186102 403174
rect 185546 366618 186102 367174
rect 185546 330618 186102 331174
rect 185546 294618 186102 295174
rect 185546 258618 186102 259174
rect 185546 222618 186102 223174
rect 185546 186618 186102 187174
rect 185546 150618 186102 151174
rect 185546 114618 186102 115174
rect 185546 78618 186102 79174
rect 185546 42618 186102 43174
rect 185546 6618 186102 7174
rect 185546 -2822 186102 -2266
rect 189266 694338 189822 694894
rect 189266 658338 189822 658894
rect 189266 622338 189822 622894
rect 189266 586338 189822 586894
rect 189266 550338 189822 550894
rect 189266 514338 189822 514894
rect 189266 478338 189822 478894
rect 189266 442338 189822 442894
rect 189266 406338 189822 406894
rect 189266 370338 189822 370894
rect 189266 334338 189822 334894
rect 189266 298338 189822 298894
rect 189266 262338 189822 262894
rect 189266 226338 189822 226894
rect 189266 190338 189822 190894
rect 189266 154338 189822 154894
rect 189266 118338 189822 118894
rect 189266 82338 189822 82894
rect 189266 46338 189822 46894
rect 189266 10338 189822 10894
rect 189266 -4742 189822 -4186
rect 210986 711002 211542 711558
rect 207266 709082 207822 709638
rect 203546 707162 204102 707718
rect 192986 698058 193542 698614
rect 192986 662058 193542 662614
rect 192986 626058 193542 626614
rect 192986 590058 193542 590614
rect 192986 554058 193542 554614
rect 192986 518058 193542 518614
rect 192986 482058 193542 482614
rect 192986 446058 193542 446614
rect 192986 410058 193542 410614
rect 192986 374058 193542 374614
rect 192986 338058 193542 338614
rect 192986 302058 193542 302614
rect 192986 266058 193542 266614
rect 192986 230058 193542 230614
rect 192986 194058 193542 194614
rect 192986 158058 193542 158614
rect 192986 122058 193542 122614
rect 192986 86058 193542 86614
rect 192986 50058 193542 50614
rect 192986 14058 193542 14614
rect 174986 -7622 175542 -7066
rect 199826 705242 200382 705798
rect 199826 668898 200382 669454
rect 199826 632898 200382 633454
rect 199826 596898 200382 597454
rect 199826 560898 200382 561454
rect 199826 524898 200382 525454
rect 199826 488898 200382 489454
rect 199826 452898 200382 453454
rect 199826 416898 200382 417454
rect 199826 380898 200382 381454
rect 199826 344898 200382 345454
rect 199826 308898 200382 309454
rect 199826 272898 200382 273454
rect 199826 236898 200382 237454
rect 199826 200898 200382 201454
rect 199826 164898 200382 165454
rect 199826 128898 200382 129454
rect 199826 92898 200382 93454
rect 199826 56898 200382 57454
rect 199826 20898 200382 21454
rect 199826 -1862 200382 -1306
rect 203546 672618 204102 673174
rect 203546 636618 204102 637174
rect 203546 600618 204102 601174
rect 203546 564618 204102 565174
rect 203546 528618 204102 529174
rect 203546 492618 204102 493174
rect 203546 456618 204102 457174
rect 203546 420618 204102 421174
rect 203546 384618 204102 385174
rect 203546 348618 204102 349174
rect 203546 312618 204102 313174
rect 203546 276618 204102 277174
rect 203546 240618 204102 241174
rect 203546 204618 204102 205174
rect 203546 168618 204102 169174
rect 203546 132618 204102 133174
rect 203546 96618 204102 97174
rect 203546 60618 204102 61174
rect 203546 24618 204102 25174
rect 203546 -3782 204102 -3226
rect 207266 676338 207822 676894
rect 207266 640338 207822 640894
rect 207266 604338 207822 604894
rect 207266 568338 207822 568894
rect 207266 532338 207822 532894
rect 207266 496338 207822 496894
rect 207266 460338 207822 460894
rect 207266 424338 207822 424894
rect 207266 388338 207822 388894
rect 207266 352338 207822 352894
rect 207266 316338 207822 316894
rect 207266 280338 207822 280894
rect 207266 244338 207822 244894
rect 207266 208338 207822 208894
rect 207266 172338 207822 172894
rect 207266 136338 207822 136894
rect 207266 100338 207822 100894
rect 207266 64338 207822 64894
rect 207266 28338 207822 28894
rect 207266 -5702 207822 -5146
rect 228986 710042 229542 710598
rect 225266 708122 225822 708678
rect 221546 706202 222102 706758
rect 210986 680058 211542 680614
rect 210986 644058 211542 644614
rect 210986 608058 211542 608614
rect 210986 572058 211542 572614
rect 210986 536058 211542 536614
rect 210986 500058 211542 500614
rect 210986 464058 211542 464614
rect 210986 428058 211542 428614
rect 210986 392058 211542 392614
rect 210986 356058 211542 356614
rect 210986 320058 211542 320614
rect 210986 284058 211542 284614
rect 210986 248058 211542 248614
rect 210986 212058 211542 212614
rect 210986 176058 211542 176614
rect 210986 140058 211542 140614
rect 210986 104058 211542 104614
rect 210986 68058 211542 68614
rect 210986 32058 211542 32614
rect 192986 -6662 193542 -6106
rect 217826 704282 218382 704838
rect 217826 686898 218382 687454
rect 217826 650898 218382 651454
rect 217826 614898 218382 615454
rect 217826 578898 218382 579454
rect 217826 542898 218382 543454
rect 217826 506898 218382 507454
rect 217826 470898 218382 471454
rect 217826 434898 218382 435454
rect 217826 398898 218382 399454
rect 217826 362898 218382 363454
rect 217826 326898 218382 327454
rect 217826 290898 218382 291454
rect 217826 254898 218382 255454
rect 217826 218898 218382 219454
rect 217826 182898 218382 183454
rect 217826 146898 218382 147454
rect 217826 110898 218382 111454
rect 217826 74898 218382 75454
rect 217826 38898 218382 39454
rect 217826 2898 218382 3454
rect 217826 -902 218382 -346
rect 221546 690618 222102 691174
rect 221546 654618 222102 655174
rect 221546 618618 222102 619174
rect 221546 582618 222102 583174
rect 221546 546618 222102 547174
rect 221546 510618 222102 511174
rect 221546 474618 222102 475174
rect 221546 438618 222102 439174
rect 221546 402618 222102 403174
rect 221546 366618 222102 367174
rect 221546 330618 222102 331174
rect 221546 294618 222102 295174
rect 221546 258618 222102 259174
rect 221546 222618 222102 223174
rect 221546 186618 222102 187174
rect 221546 150618 222102 151174
rect 221546 114618 222102 115174
rect 221546 78618 222102 79174
rect 221546 42618 222102 43174
rect 221546 6618 222102 7174
rect 221546 -2822 222102 -2266
rect 225266 694338 225822 694894
rect 225266 658338 225822 658894
rect 225266 622338 225822 622894
rect 225266 586338 225822 586894
rect 225266 550338 225822 550894
rect 225266 514338 225822 514894
rect 225266 478338 225822 478894
rect 225266 442338 225822 442894
rect 225266 406338 225822 406894
rect 225266 370338 225822 370894
rect 225266 334338 225822 334894
rect 225266 298338 225822 298894
rect 225266 262338 225822 262894
rect 225266 226338 225822 226894
rect 225266 190338 225822 190894
rect 225266 154338 225822 154894
rect 225266 118338 225822 118894
rect 225266 82338 225822 82894
rect 225266 46338 225822 46894
rect 225266 10338 225822 10894
rect 225266 -4742 225822 -4186
rect 246986 711002 247542 711558
rect 243266 709082 243822 709638
rect 239546 707162 240102 707718
rect 228986 698058 229542 698614
rect 228986 662058 229542 662614
rect 228986 626058 229542 626614
rect 228986 590058 229542 590614
rect 228986 554058 229542 554614
rect 228986 518058 229542 518614
rect 228986 482058 229542 482614
rect 235826 705242 236382 705798
rect 235826 668898 236382 669454
rect 235826 632898 236382 633454
rect 235826 596898 236382 597454
rect 235826 560898 236382 561454
rect 235826 524898 236382 525454
rect 235826 488898 236382 489454
rect 239546 672618 240102 673174
rect 239546 636618 240102 637174
rect 239546 600618 240102 601174
rect 239546 564618 240102 565174
rect 239546 528618 240102 529174
rect 239546 492618 240102 493174
rect 243266 676338 243822 676894
rect 243266 640338 243822 640894
rect 243266 604338 243822 604894
rect 243266 568338 243822 568894
rect 243266 532338 243822 532894
rect 243266 496338 243822 496894
rect 243266 460338 243822 460894
rect 264986 710042 265542 710598
rect 261266 708122 261822 708678
rect 257546 706202 258102 706758
rect 246986 680058 247542 680614
rect 246986 644058 247542 644614
rect 246986 608058 247542 608614
rect 246986 572058 247542 572614
rect 246986 536058 247542 536614
rect 246986 500058 247542 500614
rect 246986 464058 247542 464614
rect 253826 704282 254382 704838
rect 253826 686898 254382 687454
rect 253826 650898 254382 651454
rect 253826 614898 254382 615454
rect 253826 578898 254382 579454
rect 253826 542898 254382 543454
rect 253826 506898 254382 507454
rect 253826 470898 254382 471454
rect 257546 690618 258102 691174
rect 257546 654618 258102 655174
rect 257546 618618 258102 619174
rect 257546 582618 258102 583174
rect 257546 546618 258102 547174
rect 257546 510618 258102 511174
rect 257546 474618 258102 475174
rect 261266 694338 261822 694894
rect 261266 658338 261822 658894
rect 261266 622338 261822 622894
rect 261266 586338 261822 586894
rect 261266 550338 261822 550894
rect 261266 514338 261822 514894
rect 261266 478338 261822 478894
rect 282986 711002 283542 711558
rect 279266 709082 279822 709638
rect 275546 707162 276102 707718
rect 264986 698058 265542 698614
rect 264986 662058 265542 662614
rect 264986 626058 265542 626614
rect 264986 590058 265542 590614
rect 264986 554058 265542 554614
rect 264986 518058 265542 518614
rect 264986 482058 265542 482614
rect 271826 705242 272382 705798
rect 271826 668898 272382 669454
rect 271826 632898 272382 633454
rect 271826 596898 272382 597454
rect 271826 560898 272382 561454
rect 271826 524898 272382 525454
rect 271826 488898 272382 489454
rect 275546 672618 276102 673174
rect 275546 636618 276102 637174
rect 275546 600618 276102 601174
rect 275546 564618 276102 565174
rect 275546 528618 276102 529174
rect 275546 492618 276102 493174
rect 279266 676338 279822 676894
rect 279266 640338 279822 640894
rect 279266 604338 279822 604894
rect 279266 568338 279822 568894
rect 279266 532338 279822 532894
rect 279266 496338 279822 496894
rect 279266 460338 279822 460894
rect 300986 710042 301542 710598
rect 297266 708122 297822 708678
rect 293546 706202 294102 706758
rect 282986 680058 283542 680614
rect 282986 644058 283542 644614
rect 282986 608058 283542 608614
rect 282986 572058 283542 572614
rect 282986 536058 283542 536614
rect 282986 500058 283542 500614
rect 282986 464058 283542 464614
rect 289826 704282 290382 704838
rect 289826 686898 290382 687454
rect 289826 650898 290382 651454
rect 289826 614898 290382 615454
rect 289826 578898 290382 579454
rect 289826 542898 290382 543454
rect 289826 506898 290382 507454
rect 289826 470898 290382 471454
rect 293546 690618 294102 691174
rect 293546 654618 294102 655174
rect 293546 618618 294102 619174
rect 293546 582618 294102 583174
rect 293546 546618 294102 547174
rect 293546 510618 294102 511174
rect 293546 474618 294102 475174
rect 297266 694338 297822 694894
rect 297266 658338 297822 658894
rect 297266 622338 297822 622894
rect 297266 586338 297822 586894
rect 297266 550338 297822 550894
rect 297266 514338 297822 514894
rect 297266 478338 297822 478894
rect 318986 711002 319542 711558
rect 315266 709082 315822 709638
rect 311546 707162 312102 707718
rect 300986 698058 301542 698614
rect 300986 662058 301542 662614
rect 300986 626058 301542 626614
rect 300986 590058 301542 590614
rect 300986 554058 301542 554614
rect 300986 518058 301542 518614
rect 300986 482058 301542 482614
rect 307826 705242 308382 705798
rect 307826 668898 308382 669454
rect 307826 632898 308382 633454
rect 307826 596898 308382 597454
rect 307826 560898 308382 561454
rect 307826 524898 308382 525454
rect 307826 488898 308382 489454
rect 311546 672618 312102 673174
rect 311546 636618 312102 637174
rect 311546 600618 312102 601174
rect 311546 564618 312102 565174
rect 311546 528618 312102 529174
rect 311546 492618 312102 493174
rect 315266 676338 315822 676894
rect 315266 640338 315822 640894
rect 315266 604338 315822 604894
rect 315266 568338 315822 568894
rect 315266 532338 315822 532894
rect 315266 496338 315822 496894
rect 315266 460338 315822 460894
rect 336986 710042 337542 710598
rect 333266 708122 333822 708678
rect 329546 706202 330102 706758
rect 318986 680058 319542 680614
rect 318986 644058 319542 644614
rect 318986 608058 319542 608614
rect 318986 572058 319542 572614
rect 318986 536058 319542 536614
rect 318986 500058 319542 500614
rect 318986 464058 319542 464614
rect 325826 704282 326382 704838
rect 325826 686898 326382 687454
rect 325826 650898 326382 651454
rect 325826 614898 326382 615454
rect 325826 578898 326382 579454
rect 325826 542898 326382 543454
rect 325826 506898 326382 507454
rect 325826 470898 326382 471454
rect 329546 690618 330102 691174
rect 329546 654618 330102 655174
rect 329546 618618 330102 619174
rect 329546 582618 330102 583174
rect 329546 546618 330102 547174
rect 329546 510618 330102 511174
rect 329546 474618 330102 475174
rect 333266 694338 333822 694894
rect 333266 658338 333822 658894
rect 333266 622338 333822 622894
rect 333266 586338 333822 586894
rect 333266 550338 333822 550894
rect 333266 514338 333822 514894
rect 333266 478338 333822 478894
rect 354986 711002 355542 711558
rect 351266 709082 351822 709638
rect 347546 707162 348102 707718
rect 336986 698058 337542 698614
rect 336986 662058 337542 662614
rect 336986 626058 337542 626614
rect 336986 590058 337542 590614
rect 336986 554058 337542 554614
rect 336986 518058 337542 518614
rect 336986 482058 337542 482614
rect 343826 705242 344382 705798
rect 343826 668898 344382 669454
rect 343826 632898 344382 633454
rect 343826 596898 344382 597454
rect 343826 560898 344382 561454
rect 343826 524898 344382 525454
rect 343826 488898 344382 489454
rect 347546 672618 348102 673174
rect 347546 636618 348102 637174
rect 347546 600618 348102 601174
rect 347546 564618 348102 565174
rect 347546 528618 348102 529174
rect 347546 492618 348102 493174
rect 351266 676338 351822 676894
rect 351266 640338 351822 640894
rect 351266 604338 351822 604894
rect 351266 568338 351822 568894
rect 351266 532338 351822 532894
rect 351266 496338 351822 496894
rect 351266 460338 351822 460894
rect 372986 710042 373542 710598
rect 369266 708122 369822 708678
rect 365546 706202 366102 706758
rect 354986 680058 355542 680614
rect 354986 644058 355542 644614
rect 354986 608058 355542 608614
rect 354986 572058 355542 572614
rect 354986 536058 355542 536614
rect 354986 500058 355542 500614
rect 354986 464058 355542 464614
rect 361826 704282 362382 704838
rect 361826 686898 362382 687454
rect 361826 650898 362382 651454
rect 361826 614898 362382 615454
rect 361826 578898 362382 579454
rect 361826 542898 362382 543454
rect 361826 506898 362382 507454
rect 361826 470898 362382 471454
rect 365546 690618 366102 691174
rect 365546 654618 366102 655174
rect 365546 618618 366102 619174
rect 365546 582618 366102 583174
rect 365546 546618 366102 547174
rect 365546 510618 366102 511174
rect 365546 474618 366102 475174
rect 369266 694338 369822 694894
rect 369266 658338 369822 658894
rect 369266 622338 369822 622894
rect 369266 586338 369822 586894
rect 369266 550338 369822 550894
rect 369266 514338 369822 514894
rect 369266 478338 369822 478894
rect 390986 711002 391542 711558
rect 387266 709082 387822 709638
rect 383546 707162 384102 707718
rect 372986 698058 373542 698614
rect 372986 662058 373542 662614
rect 372986 626058 373542 626614
rect 372986 590058 373542 590614
rect 372986 554058 373542 554614
rect 372986 518058 373542 518614
rect 372986 482058 373542 482614
rect 379826 705242 380382 705798
rect 379826 668898 380382 669454
rect 379826 632898 380382 633454
rect 379826 596898 380382 597454
rect 379826 560898 380382 561454
rect 379826 524898 380382 525454
rect 379826 488898 380382 489454
rect 383546 672618 384102 673174
rect 383546 636618 384102 637174
rect 383546 600618 384102 601174
rect 383546 564618 384102 565174
rect 383546 528618 384102 529174
rect 383546 492618 384102 493174
rect 387266 676338 387822 676894
rect 387266 640338 387822 640894
rect 387266 604338 387822 604894
rect 387266 568338 387822 568894
rect 387266 532338 387822 532894
rect 387266 496338 387822 496894
rect 387266 460338 387822 460894
rect 408986 710042 409542 710598
rect 405266 708122 405822 708678
rect 401546 706202 402102 706758
rect 390986 680058 391542 680614
rect 390986 644058 391542 644614
rect 390986 608058 391542 608614
rect 390986 572058 391542 572614
rect 390986 536058 391542 536614
rect 390986 500058 391542 500614
rect 390986 464058 391542 464614
rect 397826 704282 398382 704838
rect 397826 686898 398382 687454
rect 397826 650898 398382 651454
rect 397826 614898 398382 615454
rect 397826 578898 398382 579454
rect 397826 542898 398382 543454
rect 397826 506898 398382 507454
rect 397826 470898 398382 471454
rect 401546 690618 402102 691174
rect 401546 654618 402102 655174
rect 401546 618618 402102 619174
rect 401546 582618 402102 583174
rect 401546 546618 402102 547174
rect 401546 510618 402102 511174
rect 401546 474618 402102 475174
rect 405266 694338 405822 694894
rect 405266 658338 405822 658894
rect 405266 622338 405822 622894
rect 405266 586338 405822 586894
rect 405266 550338 405822 550894
rect 405266 514338 405822 514894
rect 405266 478338 405822 478894
rect 426986 711002 427542 711558
rect 423266 709082 423822 709638
rect 419546 707162 420102 707718
rect 408986 698058 409542 698614
rect 408986 662058 409542 662614
rect 408986 626058 409542 626614
rect 408986 590058 409542 590614
rect 408986 554058 409542 554614
rect 408986 518058 409542 518614
rect 408986 482058 409542 482614
rect 415826 705242 416382 705798
rect 415826 668898 416382 669454
rect 415826 632898 416382 633454
rect 415826 596898 416382 597454
rect 415826 560898 416382 561454
rect 415826 524898 416382 525454
rect 415826 488898 416382 489454
rect 419546 672618 420102 673174
rect 419546 636618 420102 637174
rect 419546 600618 420102 601174
rect 419546 564618 420102 565174
rect 419546 528618 420102 529174
rect 419546 492618 420102 493174
rect 228986 446058 229542 446614
rect 228986 410058 229542 410614
rect 228986 374058 229542 374614
rect 228986 338058 229542 338614
rect 228986 302058 229542 302614
rect 228986 266058 229542 266614
rect 228986 230058 229542 230614
rect 228986 194058 229542 194614
rect 228986 158058 229542 158614
rect 228986 122058 229542 122614
rect 228986 86058 229542 86614
rect 228986 50058 229542 50614
rect 254610 453218 254846 453454
rect 254610 452898 254846 453134
rect 285330 453218 285566 453454
rect 285330 452898 285566 453134
rect 316050 453218 316286 453454
rect 316050 452898 316286 453134
rect 346770 453218 347006 453454
rect 346770 452898 347006 453134
rect 377490 453218 377726 453454
rect 377490 452898 377726 453134
rect 408210 453218 408446 453454
rect 408210 452898 408446 453134
rect 239250 435218 239486 435454
rect 239250 434898 239486 435134
rect 269970 435218 270206 435454
rect 269970 434898 270206 435134
rect 300690 435218 300926 435454
rect 300690 434898 300926 435134
rect 331410 435218 331646 435454
rect 331410 434898 331646 435134
rect 362130 435218 362366 435454
rect 362130 434898 362366 435134
rect 392850 435218 393086 435454
rect 392850 434898 393086 435134
rect 254610 417218 254846 417454
rect 254610 416898 254846 417134
rect 285330 417218 285566 417454
rect 285330 416898 285566 417134
rect 316050 417218 316286 417454
rect 316050 416898 316286 417134
rect 346770 417218 347006 417454
rect 346770 416898 347006 417134
rect 377490 417218 377726 417454
rect 377490 416898 377726 417134
rect 408210 417218 408446 417454
rect 408210 416898 408446 417134
rect 239250 399218 239486 399454
rect 239250 398898 239486 399134
rect 269970 399218 270206 399454
rect 269970 398898 270206 399134
rect 300690 399218 300926 399454
rect 300690 398898 300926 399134
rect 331410 399218 331646 399454
rect 331410 398898 331646 399134
rect 362130 399218 362366 399454
rect 362130 398898 362366 399134
rect 392850 399218 393086 399454
rect 392850 398898 393086 399134
rect 254610 381218 254846 381454
rect 254610 380898 254846 381134
rect 285330 381218 285566 381454
rect 285330 380898 285566 381134
rect 316050 381218 316286 381454
rect 316050 380898 316286 381134
rect 346770 381218 347006 381454
rect 346770 380898 347006 381134
rect 377490 381218 377726 381454
rect 377490 380898 377726 381134
rect 408210 381218 408446 381454
rect 408210 380898 408446 381134
rect 239250 363218 239486 363454
rect 239250 362898 239486 363134
rect 269970 363218 270206 363454
rect 269970 362898 270206 363134
rect 300690 363218 300926 363454
rect 300690 362898 300926 363134
rect 331410 363218 331646 363454
rect 331410 362898 331646 363134
rect 362130 363218 362366 363454
rect 362130 362898 362366 363134
rect 392850 363218 393086 363454
rect 392850 362898 393086 363134
rect 254610 345218 254846 345454
rect 254610 344898 254846 345134
rect 285330 345218 285566 345454
rect 285330 344898 285566 345134
rect 316050 345218 316286 345454
rect 316050 344898 316286 345134
rect 346770 345218 347006 345454
rect 346770 344898 347006 345134
rect 377490 345218 377726 345454
rect 377490 344898 377726 345134
rect 408210 345218 408446 345454
rect 408210 344898 408446 345134
rect 235826 308898 236382 309454
rect 235826 272898 236382 273454
rect 235826 236898 236382 237454
rect 235826 200898 236382 201454
rect 235826 164898 236382 165454
rect 235826 128898 236382 129454
rect 235826 92898 236382 93454
rect 235826 56898 236382 57454
rect 228986 14058 229542 14614
rect 210986 -7622 211542 -7066
rect 235826 20898 236382 21454
rect 235826 -1862 236382 -1306
rect 239546 312618 240102 313174
rect 239546 276618 240102 277174
rect 239546 240618 240102 241174
rect 239546 204618 240102 205174
rect 239546 168618 240102 169174
rect 239546 132618 240102 133174
rect 239546 96618 240102 97174
rect 239546 60618 240102 61174
rect 239546 24618 240102 25174
rect 239546 -3782 240102 -3226
rect 243266 316338 243822 316894
rect 243266 280338 243822 280894
rect 243266 244338 243822 244894
rect 243266 208338 243822 208894
rect 243266 172338 243822 172894
rect 243266 136338 243822 136894
rect 243266 100338 243822 100894
rect 243266 64338 243822 64894
rect 243266 28338 243822 28894
rect 243266 -5702 243822 -5146
rect 246986 320058 247542 320614
rect 246986 284058 247542 284614
rect 246986 248058 247542 248614
rect 246986 212058 247542 212614
rect 246986 176058 247542 176614
rect 246986 140058 247542 140614
rect 246986 104058 247542 104614
rect 246986 68058 247542 68614
rect 246986 32058 247542 32614
rect 228986 -6662 229542 -6106
rect 253826 326898 254382 327454
rect 253826 290898 254382 291454
rect 253826 254898 254382 255454
rect 253826 218898 254382 219454
rect 253826 182898 254382 183454
rect 253826 146898 254382 147454
rect 253826 110898 254382 111454
rect 253826 74898 254382 75454
rect 253826 38898 254382 39454
rect 253826 2898 254382 3454
rect 253826 -902 254382 -346
rect 257546 330618 258102 331174
rect 257546 294618 258102 295174
rect 257546 258618 258102 259174
rect 257546 222618 258102 223174
rect 257546 186618 258102 187174
rect 257546 150618 258102 151174
rect 257546 114618 258102 115174
rect 257546 78618 258102 79174
rect 257546 42618 258102 43174
rect 257546 6618 258102 7174
rect 257546 -2822 258102 -2266
rect 261266 334338 261822 334894
rect 261266 298338 261822 298894
rect 261266 262338 261822 262894
rect 261266 226338 261822 226894
rect 261266 190338 261822 190894
rect 261266 154338 261822 154894
rect 261266 118338 261822 118894
rect 261266 82338 261822 82894
rect 261266 46338 261822 46894
rect 261266 10338 261822 10894
rect 261266 -4742 261822 -4186
rect 264986 302058 265542 302614
rect 264986 266058 265542 266614
rect 264986 230058 265542 230614
rect 264986 194058 265542 194614
rect 264986 158058 265542 158614
rect 264986 122058 265542 122614
rect 264986 86058 265542 86614
rect 264986 50058 265542 50614
rect 264986 14058 265542 14614
rect 246986 -7622 247542 -7066
rect 271826 308898 272382 309454
rect 271826 272898 272382 273454
rect 271826 236898 272382 237454
rect 271826 200898 272382 201454
rect 271826 164898 272382 165454
rect 271826 128898 272382 129454
rect 271826 92898 272382 93454
rect 271826 56898 272382 57454
rect 271826 20898 272382 21454
rect 271826 -1862 272382 -1306
rect 275546 312618 276102 313174
rect 275546 276618 276102 277174
rect 275546 240618 276102 241174
rect 275546 204618 276102 205174
rect 275546 168618 276102 169174
rect 275546 132618 276102 133174
rect 275546 96618 276102 97174
rect 275546 60618 276102 61174
rect 275546 24618 276102 25174
rect 275546 -3782 276102 -3226
rect 279266 316338 279822 316894
rect 279266 280338 279822 280894
rect 279266 244338 279822 244894
rect 279266 208338 279822 208894
rect 279266 172338 279822 172894
rect 279266 136338 279822 136894
rect 279266 100338 279822 100894
rect 279266 64338 279822 64894
rect 279266 28338 279822 28894
rect 279266 -5702 279822 -5146
rect 282986 320058 283542 320614
rect 282986 284058 283542 284614
rect 282986 248058 283542 248614
rect 282986 212058 283542 212614
rect 282986 176058 283542 176614
rect 282986 140058 283542 140614
rect 282986 104058 283542 104614
rect 282986 68058 283542 68614
rect 282986 32058 283542 32614
rect 264986 -6662 265542 -6106
rect 289826 326898 290382 327454
rect 289826 290898 290382 291454
rect 289826 254898 290382 255454
rect 289826 218898 290382 219454
rect 289826 182898 290382 183454
rect 289826 146898 290382 147454
rect 289826 110898 290382 111454
rect 289826 74898 290382 75454
rect 289826 38898 290382 39454
rect 289826 2898 290382 3454
rect 289826 -902 290382 -346
rect 293546 330618 294102 331174
rect 293546 294618 294102 295174
rect 293546 258618 294102 259174
rect 293546 222618 294102 223174
rect 293546 186618 294102 187174
rect 293546 150618 294102 151174
rect 293546 114618 294102 115174
rect 293546 78618 294102 79174
rect 293546 42618 294102 43174
rect 293546 6618 294102 7174
rect 293546 -2822 294102 -2266
rect 297266 334338 297822 334894
rect 297266 298338 297822 298894
rect 297266 262338 297822 262894
rect 297266 226338 297822 226894
rect 297266 190338 297822 190894
rect 297266 154338 297822 154894
rect 297266 118338 297822 118894
rect 297266 82338 297822 82894
rect 297266 46338 297822 46894
rect 297266 10338 297822 10894
rect 297266 -4742 297822 -4186
rect 300986 302058 301542 302614
rect 300986 266058 301542 266614
rect 300986 230058 301542 230614
rect 300986 194058 301542 194614
rect 300986 158058 301542 158614
rect 300986 122058 301542 122614
rect 300986 86058 301542 86614
rect 300986 50058 301542 50614
rect 300986 14058 301542 14614
rect 282986 -7622 283542 -7066
rect 307826 308898 308382 309454
rect 307826 272898 308382 273454
rect 307826 236898 308382 237454
rect 307826 200898 308382 201454
rect 307826 164898 308382 165454
rect 307826 128898 308382 129454
rect 307826 92898 308382 93454
rect 307826 56898 308382 57454
rect 307826 20898 308382 21454
rect 307826 -1862 308382 -1306
rect 311546 312618 312102 313174
rect 311546 276618 312102 277174
rect 311546 240618 312102 241174
rect 311546 204618 312102 205174
rect 311546 168618 312102 169174
rect 311546 132618 312102 133174
rect 311546 96618 312102 97174
rect 311546 60618 312102 61174
rect 311546 24618 312102 25174
rect 311546 -3782 312102 -3226
rect 315266 316338 315822 316894
rect 315266 280338 315822 280894
rect 315266 244338 315822 244894
rect 315266 208338 315822 208894
rect 315266 172338 315822 172894
rect 315266 136338 315822 136894
rect 315266 100338 315822 100894
rect 315266 64338 315822 64894
rect 315266 28338 315822 28894
rect 315266 -5702 315822 -5146
rect 318986 320058 319542 320614
rect 318986 284058 319542 284614
rect 318986 248058 319542 248614
rect 318986 212058 319542 212614
rect 318986 176058 319542 176614
rect 318986 140058 319542 140614
rect 318986 104058 319542 104614
rect 318986 68058 319542 68614
rect 318986 32058 319542 32614
rect 300986 -6662 301542 -6106
rect 325826 326898 326382 327454
rect 325826 290898 326382 291454
rect 325826 254898 326382 255454
rect 325826 218898 326382 219454
rect 325826 182898 326382 183454
rect 325826 146898 326382 147454
rect 325826 110898 326382 111454
rect 325826 74898 326382 75454
rect 325826 38898 326382 39454
rect 325826 2898 326382 3454
rect 325826 -902 326382 -346
rect 329546 330618 330102 331174
rect 329546 294618 330102 295174
rect 329546 258618 330102 259174
rect 329546 222618 330102 223174
rect 329546 186618 330102 187174
rect 329546 150618 330102 151174
rect 329546 114618 330102 115174
rect 329546 78618 330102 79174
rect 329546 42618 330102 43174
rect 329546 6618 330102 7174
rect 329546 -2822 330102 -2266
rect 333266 334338 333822 334894
rect 333266 298338 333822 298894
rect 333266 262338 333822 262894
rect 333266 226338 333822 226894
rect 333266 190338 333822 190894
rect 333266 154338 333822 154894
rect 333266 118338 333822 118894
rect 333266 82338 333822 82894
rect 333266 46338 333822 46894
rect 333266 10338 333822 10894
rect 333266 -4742 333822 -4186
rect 336986 302058 337542 302614
rect 336986 266058 337542 266614
rect 336986 230058 337542 230614
rect 336986 194058 337542 194614
rect 336986 158058 337542 158614
rect 336986 122058 337542 122614
rect 336986 86058 337542 86614
rect 336986 50058 337542 50614
rect 336986 14058 337542 14614
rect 318986 -7622 319542 -7066
rect 343826 308898 344382 309454
rect 343826 272898 344382 273454
rect 343826 236898 344382 237454
rect 343826 200898 344382 201454
rect 343826 164898 344382 165454
rect 343826 128898 344382 129454
rect 343826 92898 344382 93454
rect 343826 56898 344382 57454
rect 343826 20898 344382 21454
rect 343826 -1862 344382 -1306
rect 347546 312618 348102 313174
rect 347546 276618 348102 277174
rect 347546 240618 348102 241174
rect 347546 204618 348102 205174
rect 347546 168618 348102 169174
rect 347546 132618 348102 133174
rect 347546 96618 348102 97174
rect 347546 60618 348102 61174
rect 347546 24618 348102 25174
rect 347546 -3782 348102 -3226
rect 351266 316338 351822 316894
rect 351266 280338 351822 280894
rect 351266 244338 351822 244894
rect 351266 208338 351822 208894
rect 351266 172338 351822 172894
rect 351266 136338 351822 136894
rect 351266 100338 351822 100894
rect 351266 64338 351822 64894
rect 351266 28338 351822 28894
rect 351266 -5702 351822 -5146
rect 354986 320058 355542 320614
rect 354986 284058 355542 284614
rect 354986 248058 355542 248614
rect 354986 212058 355542 212614
rect 354986 176058 355542 176614
rect 354986 140058 355542 140614
rect 354986 104058 355542 104614
rect 354986 68058 355542 68614
rect 354986 32058 355542 32614
rect 336986 -6662 337542 -6106
rect 361826 326898 362382 327454
rect 361826 290898 362382 291454
rect 361826 254898 362382 255454
rect 361826 218898 362382 219454
rect 361826 182898 362382 183454
rect 361826 146898 362382 147454
rect 361826 110898 362382 111454
rect 361826 74898 362382 75454
rect 361826 38898 362382 39454
rect 361826 2898 362382 3454
rect 361826 -902 362382 -346
rect 365546 330618 366102 331174
rect 365546 294618 366102 295174
rect 365546 258618 366102 259174
rect 365546 222618 366102 223174
rect 365546 186618 366102 187174
rect 365546 150618 366102 151174
rect 365546 114618 366102 115174
rect 365546 78618 366102 79174
rect 365546 42618 366102 43174
rect 365546 6618 366102 7174
rect 365546 -2822 366102 -2266
rect 369266 334338 369822 334894
rect 369266 298338 369822 298894
rect 369266 262338 369822 262894
rect 369266 226338 369822 226894
rect 369266 190338 369822 190894
rect 369266 154338 369822 154894
rect 369266 118338 369822 118894
rect 369266 82338 369822 82894
rect 369266 46338 369822 46894
rect 369266 10338 369822 10894
rect 369266 -4742 369822 -4186
rect 372986 302058 373542 302614
rect 372986 266058 373542 266614
rect 372986 230058 373542 230614
rect 372986 194058 373542 194614
rect 372986 158058 373542 158614
rect 372986 122058 373542 122614
rect 372986 86058 373542 86614
rect 372986 50058 373542 50614
rect 372986 14058 373542 14614
rect 354986 -7622 355542 -7066
rect 379826 308898 380382 309454
rect 379826 272898 380382 273454
rect 379826 236898 380382 237454
rect 379826 200898 380382 201454
rect 379826 164898 380382 165454
rect 379826 128898 380382 129454
rect 379826 92898 380382 93454
rect 379826 56898 380382 57454
rect 379826 20898 380382 21454
rect 379826 -1862 380382 -1306
rect 383546 312618 384102 313174
rect 383546 276618 384102 277174
rect 383546 240618 384102 241174
rect 383546 204618 384102 205174
rect 383546 168618 384102 169174
rect 383546 132618 384102 133174
rect 383546 96618 384102 97174
rect 383546 60618 384102 61174
rect 383546 24618 384102 25174
rect 383546 -3782 384102 -3226
rect 387266 316338 387822 316894
rect 387266 280338 387822 280894
rect 387266 244338 387822 244894
rect 387266 208338 387822 208894
rect 387266 172338 387822 172894
rect 387266 136338 387822 136894
rect 387266 100338 387822 100894
rect 387266 64338 387822 64894
rect 387266 28338 387822 28894
rect 387266 -5702 387822 -5146
rect 390986 320058 391542 320614
rect 390986 284058 391542 284614
rect 390986 248058 391542 248614
rect 390986 212058 391542 212614
rect 390986 176058 391542 176614
rect 390986 140058 391542 140614
rect 390986 104058 391542 104614
rect 390986 68058 391542 68614
rect 390986 32058 391542 32614
rect 372986 -6662 373542 -6106
rect 397826 326898 398382 327454
rect 397826 290898 398382 291454
rect 397826 254898 398382 255454
rect 397826 218898 398382 219454
rect 397826 182898 398382 183454
rect 397826 146898 398382 147454
rect 397826 110898 398382 111454
rect 397826 74898 398382 75454
rect 397826 38898 398382 39454
rect 397826 2898 398382 3454
rect 397826 -902 398382 -346
rect 401546 330618 402102 331174
rect 401546 294618 402102 295174
rect 401546 258618 402102 259174
rect 401546 222618 402102 223174
rect 401546 186618 402102 187174
rect 401546 150618 402102 151174
rect 401546 114618 402102 115174
rect 401546 78618 402102 79174
rect 401546 42618 402102 43174
rect 401546 6618 402102 7174
rect 401546 -2822 402102 -2266
rect 405266 334338 405822 334894
rect 405266 298338 405822 298894
rect 405266 262338 405822 262894
rect 405266 226338 405822 226894
rect 405266 190338 405822 190894
rect 405266 154338 405822 154894
rect 405266 118338 405822 118894
rect 405266 82338 405822 82894
rect 408986 302058 409542 302614
rect 408986 266058 409542 266614
rect 408986 230058 409542 230614
rect 408986 194058 409542 194614
rect 408986 158058 409542 158614
rect 408986 122058 409542 122614
rect 408986 86058 409542 86614
rect 405266 46338 405822 46894
rect 405266 10338 405822 10894
rect 405266 -4742 405822 -4186
rect 408986 50058 409542 50614
rect 419546 456618 420102 457174
rect 419546 420618 420102 421174
rect 419546 384618 420102 385174
rect 419546 348618 420102 349174
rect 415826 308898 416382 309454
rect 415826 272898 416382 273454
rect 415826 236898 416382 237454
rect 415826 200898 416382 201454
rect 415826 164898 416382 165454
rect 415826 128898 416382 129454
rect 415826 92898 416382 93454
rect 415826 56898 416382 57454
rect 415826 20898 416382 21454
rect 408986 14058 409542 14614
rect 390986 -7622 391542 -7066
rect 415826 -1862 416382 -1306
rect 419546 312618 420102 313174
rect 419546 276618 420102 277174
rect 419546 240618 420102 241174
rect 419546 204618 420102 205174
rect 419546 168618 420102 169174
rect 419546 132618 420102 133174
rect 419546 96618 420102 97174
rect 419546 60618 420102 61174
rect 419546 24618 420102 25174
rect 419546 -3782 420102 -3226
rect 423266 676338 423822 676894
rect 423266 640338 423822 640894
rect 423266 604338 423822 604894
rect 423266 568338 423822 568894
rect 423266 532338 423822 532894
rect 423266 496338 423822 496894
rect 423266 460338 423822 460894
rect 423266 424338 423822 424894
rect 423266 388338 423822 388894
rect 423266 352338 423822 352894
rect 423266 316338 423822 316894
rect 423266 280338 423822 280894
rect 423266 244338 423822 244894
rect 423266 208338 423822 208894
rect 423266 172338 423822 172894
rect 423266 136338 423822 136894
rect 423266 100338 423822 100894
rect 423266 64338 423822 64894
rect 423266 28338 423822 28894
rect 423266 -5702 423822 -5146
rect 444986 710042 445542 710598
rect 441266 708122 441822 708678
rect 437546 706202 438102 706758
rect 426986 680058 427542 680614
rect 426986 644058 427542 644614
rect 426986 608058 427542 608614
rect 426986 572058 427542 572614
rect 426986 536058 427542 536614
rect 426986 500058 427542 500614
rect 426986 464058 427542 464614
rect 426986 428058 427542 428614
rect 426986 392058 427542 392614
rect 426986 356058 427542 356614
rect 426986 320058 427542 320614
rect 426986 284058 427542 284614
rect 426986 248058 427542 248614
rect 426986 212058 427542 212614
rect 426986 176058 427542 176614
rect 426986 140058 427542 140614
rect 426986 104058 427542 104614
rect 426986 68058 427542 68614
rect 426986 32058 427542 32614
rect 408986 -6662 409542 -6106
rect 433826 704282 434382 704838
rect 433826 686898 434382 687454
rect 433826 650898 434382 651454
rect 433826 614898 434382 615454
rect 433826 578898 434382 579454
rect 433826 542898 434382 543454
rect 433826 506898 434382 507454
rect 433826 470898 434382 471454
rect 433826 434898 434382 435454
rect 433826 398898 434382 399454
rect 433826 362898 434382 363454
rect 433826 326898 434382 327454
rect 433826 290898 434382 291454
rect 433826 254898 434382 255454
rect 433826 218898 434382 219454
rect 433826 182898 434382 183454
rect 433826 146898 434382 147454
rect 433826 110898 434382 111454
rect 433826 74898 434382 75454
rect 433826 38898 434382 39454
rect 433826 2898 434382 3454
rect 433826 -902 434382 -346
rect 437546 690618 438102 691174
rect 437546 654618 438102 655174
rect 437546 618618 438102 619174
rect 437546 582618 438102 583174
rect 437546 546618 438102 547174
rect 437546 510618 438102 511174
rect 437546 474618 438102 475174
rect 437546 438618 438102 439174
rect 437546 402618 438102 403174
rect 437546 366618 438102 367174
rect 437546 330618 438102 331174
rect 437546 294618 438102 295174
rect 437546 258618 438102 259174
rect 437546 222618 438102 223174
rect 437546 186618 438102 187174
rect 437546 150618 438102 151174
rect 437546 114618 438102 115174
rect 437546 78618 438102 79174
rect 437546 42618 438102 43174
rect 437546 6618 438102 7174
rect 437546 -2822 438102 -2266
rect 441266 694338 441822 694894
rect 441266 658338 441822 658894
rect 441266 622338 441822 622894
rect 441266 586338 441822 586894
rect 441266 550338 441822 550894
rect 441266 514338 441822 514894
rect 441266 478338 441822 478894
rect 441266 442338 441822 442894
rect 441266 406338 441822 406894
rect 441266 370338 441822 370894
rect 441266 334338 441822 334894
rect 441266 298338 441822 298894
rect 441266 262338 441822 262894
rect 441266 226338 441822 226894
rect 441266 190338 441822 190894
rect 441266 154338 441822 154894
rect 441266 118338 441822 118894
rect 441266 82338 441822 82894
rect 441266 46338 441822 46894
rect 441266 10338 441822 10894
rect 441266 -4742 441822 -4186
rect 462986 711002 463542 711558
rect 459266 709082 459822 709638
rect 455546 707162 456102 707718
rect 444986 698058 445542 698614
rect 444986 662058 445542 662614
rect 444986 626058 445542 626614
rect 444986 590058 445542 590614
rect 444986 554058 445542 554614
rect 444986 518058 445542 518614
rect 444986 482058 445542 482614
rect 444986 446058 445542 446614
rect 444986 410058 445542 410614
rect 444986 374058 445542 374614
rect 444986 338058 445542 338614
rect 444986 302058 445542 302614
rect 444986 266058 445542 266614
rect 444986 230058 445542 230614
rect 444986 194058 445542 194614
rect 444986 158058 445542 158614
rect 444986 122058 445542 122614
rect 444986 86058 445542 86614
rect 444986 50058 445542 50614
rect 444986 14058 445542 14614
rect 426986 -7622 427542 -7066
rect 451826 705242 452382 705798
rect 451826 668898 452382 669454
rect 451826 632898 452382 633454
rect 451826 596898 452382 597454
rect 451826 560898 452382 561454
rect 451826 524898 452382 525454
rect 451826 488898 452382 489454
rect 451826 452898 452382 453454
rect 451826 416898 452382 417454
rect 451826 380898 452382 381454
rect 451826 344898 452382 345454
rect 451826 308898 452382 309454
rect 451826 272898 452382 273454
rect 451826 236898 452382 237454
rect 451826 200898 452382 201454
rect 451826 164898 452382 165454
rect 451826 128898 452382 129454
rect 451826 92898 452382 93454
rect 451826 56898 452382 57454
rect 451826 20898 452382 21454
rect 451826 -1862 452382 -1306
rect 455546 672618 456102 673174
rect 455546 636618 456102 637174
rect 455546 600618 456102 601174
rect 455546 564618 456102 565174
rect 455546 528618 456102 529174
rect 455546 492618 456102 493174
rect 455546 456618 456102 457174
rect 455546 420618 456102 421174
rect 455546 384618 456102 385174
rect 455546 348618 456102 349174
rect 455546 312618 456102 313174
rect 455546 276618 456102 277174
rect 455546 240618 456102 241174
rect 455546 204618 456102 205174
rect 455546 168618 456102 169174
rect 455546 132618 456102 133174
rect 455546 96618 456102 97174
rect 455546 60618 456102 61174
rect 455546 24618 456102 25174
rect 455546 -3782 456102 -3226
rect 459266 676338 459822 676894
rect 459266 640338 459822 640894
rect 459266 604338 459822 604894
rect 459266 568338 459822 568894
rect 459266 532338 459822 532894
rect 459266 496338 459822 496894
rect 459266 460338 459822 460894
rect 459266 424338 459822 424894
rect 459266 388338 459822 388894
rect 459266 352338 459822 352894
rect 459266 316338 459822 316894
rect 459266 280338 459822 280894
rect 459266 244338 459822 244894
rect 459266 208338 459822 208894
rect 459266 172338 459822 172894
rect 459266 136338 459822 136894
rect 459266 100338 459822 100894
rect 459266 64338 459822 64894
rect 459266 28338 459822 28894
rect 459266 -5702 459822 -5146
rect 480986 710042 481542 710598
rect 477266 708122 477822 708678
rect 473546 706202 474102 706758
rect 462986 680058 463542 680614
rect 462986 644058 463542 644614
rect 462986 608058 463542 608614
rect 462986 572058 463542 572614
rect 462986 536058 463542 536614
rect 462986 500058 463542 500614
rect 462986 464058 463542 464614
rect 462986 428058 463542 428614
rect 462986 392058 463542 392614
rect 462986 356058 463542 356614
rect 462986 320058 463542 320614
rect 462986 284058 463542 284614
rect 462986 248058 463542 248614
rect 462986 212058 463542 212614
rect 462986 176058 463542 176614
rect 462986 140058 463542 140614
rect 462986 104058 463542 104614
rect 462986 68058 463542 68614
rect 462986 32058 463542 32614
rect 444986 -6662 445542 -6106
rect 469826 704282 470382 704838
rect 469826 686898 470382 687454
rect 469826 650898 470382 651454
rect 469826 614898 470382 615454
rect 469826 578898 470382 579454
rect 469826 542898 470382 543454
rect 469826 506898 470382 507454
rect 469826 470898 470382 471454
rect 469826 434898 470382 435454
rect 469826 398898 470382 399454
rect 469826 362898 470382 363454
rect 469826 326898 470382 327454
rect 469826 290898 470382 291454
rect 469826 254898 470382 255454
rect 469826 218898 470382 219454
rect 469826 182898 470382 183454
rect 469826 146898 470382 147454
rect 469826 110898 470382 111454
rect 469826 74898 470382 75454
rect 469826 38898 470382 39454
rect 469826 2898 470382 3454
rect 469826 -902 470382 -346
rect 473546 690618 474102 691174
rect 473546 654618 474102 655174
rect 473546 618618 474102 619174
rect 473546 582618 474102 583174
rect 473546 546618 474102 547174
rect 473546 510618 474102 511174
rect 473546 474618 474102 475174
rect 473546 438618 474102 439174
rect 473546 402618 474102 403174
rect 473546 366618 474102 367174
rect 473546 330618 474102 331174
rect 473546 294618 474102 295174
rect 473546 258618 474102 259174
rect 473546 222618 474102 223174
rect 473546 186618 474102 187174
rect 473546 150618 474102 151174
rect 473546 114618 474102 115174
rect 473546 78618 474102 79174
rect 473546 42618 474102 43174
rect 473546 6618 474102 7174
rect 473546 -2822 474102 -2266
rect 477266 694338 477822 694894
rect 477266 658338 477822 658894
rect 477266 622338 477822 622894
rect 477266 586338 477822 586894
rect 477266 550338 477822 550894
rect 477266 514338 477822 514894
rect 477266 478338 477822 478894
rect 477266 442338 477822 442894
rect 477266 406338 477822 406894
rect 477266 370338 477822 370894
rect 477266 334338 477822 334894
rect 477266 298338 477822 298894
rect 477266 262338 477822 262894
rect 477266 226338 477822 226894
rect 477266 190338 477822 190894
rect 477266 154338 477822 154894
rect 477266 118338 477822 118894
rect 477266 82338 477822 82894
rect 477266 46338 477822 46894
rect 477266 10338 477822 10894
rect 477266 -4742 477822 -4186
rect 498986 711002 499542 711558
rect 495266 709082 495822 709638
rect 491546 707162 492102 707718
rect 480986 698058 481542 698614
rect 480986 662058 481542 662614
rect 480986 626058 481542 626614
rect 480986 590058 481542 590614
rect 480986 554058 481542 554614
rect 480986 518058 481542 518614
rect 480986 482058 481542 482614
rect 480986 446058 481542 446614
rect 480986 410058 481542 410614
rect 480986 374058 481542 374614
rect 480986 338058 481542 338614
rect 480986 302058 481542 302614
rect 480986 266058 481542 266614
rect 480986 230058 481542 230614
rect 480986 194058 481542 194614
rect 480986 158058 481542 158614
rect 480986 122058 481542 122614
rect 480986 86058 481542 86614
rect 480986 50058 481542 50614
rect 480986 14058 481542 14614
rect 462986 -7622 463542 -7066
rect 487826 705242 488382 705798
rect 487826 668898 488382 669454
rect 487826 632898 488382 633454
rect 487826 596898 488382 597454
rect 487826 560898 488382 561454
rect 487826 524898 488382 525454
rect 487826 488898 488382 489454
rect 487826 452898 488382 453454
rect 487826 416898 488382 417454
rect 487826 380898 488382 381454
rect 487826 344898 488382 345454
rect 487826 308898 488382 309454
rect 487826 272898 488382 273454
rect 487826 236898 488382 237454
rect 487826 200898 488382 201454
rect 487826 164898 488382 165454
rect 487826 128898 488382 129454
rect 487826 92898 488382 93454
rect 487826 56898 488382 57454
rect 487826 20898 488382 21454
rect 487826 -1862 488382 -1306
rect 491546 672618 492102 673174
rect 491546 636618 492102 637174
rect 491546 600618 492102 601174
rect 491546 564618 492102 565174
rect 491546 528618 492102 529174
rect 491546 492618 492102 493174
rect 491546 456618 492102 457174
rect 491546 420618 492102 421174
rect 491546 384618 492102 385174
rect 491546 348618 492102 349174
rect 491546 312618 492102 313174
rect 491546 276618 492102 277174
rect 491546 240618 492102 241174
rect 491546 204618 492102 205174
rect 491546 168618 492102 169174
rect 491546 132618 492102 133174
rect 491546 96618 492102 97174
rect 491546 60618 492102 61174
rect 491546 24618 492102 25174
rect 491546 -3782 492102 -3226
rect 495266 676338 495822 676894
rect 495266 640338 495822 640894
rect 495266 604338 495822 604894
rect 495266 568338 495822 568894
rect 495266 532338 495822 532894
rect 495266 496338 495822 496894
rect 495266 460338 495822 460894
rect 495266 424338 495822 424894
rect 495266 388338 495822 388894
rect 495266 352338 495822 352894
rect 495266 316338 495822 316894
rect 495266 280338 495822 280894
rect 495266 244338 495822 244894
rect 495266 208338 495822 208894
rect 495266 172338 495822 172894
rect 495266 136338 495822 136894
rect 495266 100338 495822 100894
rect 495266 64338 495822 64894
rect 495266 28338 495822 28894
rect 495266 -5702 495822 -5146
rect 516986 710042 517542 710598
rect 513266 708122 513822 708678
rect 509546 706202 510102 706758
rect 498986 680058 499542 680614
rect 498986 644058 499542 644614
rect 498986 608058 499542 608614
rect 498986 572058 499542 572614
rect 498986 536058 499542 536614
rect 498986 500058 499542 500614
rect 498986 464058 499542 464614
rect 498986 428058 499542 428614
rect 498986 392058 499542 392614
rect 498986 356058 499542 356614
rect 498986 320058 499542 320614
rect 498986 284058 499542 284614
rect 498986 248058 499542 248614
rect 498986 212058 499542 212614
rect 498986 176058 499542 176614
rect 498986 140058 499542 140614
rect 498986 104058 499542 104614
rect 498986 68058 499542 68614
rect 498986 32058 499542 32614
rect 480986 -6662 481542 -6106
rect 505826 704282 506382 704838
rect 505826 686898 506382 687454
rect 505826 650898 506382 651454
rect 505826 614898 506382 615454
rect 505826 578898 506382 579454
rect 505826 542898 506382 543454
rect 505826 506898 506382 507454
rect 505826 470898 506382 471454
rect 505826 434898 506382 435454
rect 505826 398898 506382 399454
rect 505826 362898 506382 363454
rect 505826 326898 506382 327454
rect 505826 290898 506382 291454
rect 505826 254898 506382 255454
rect 505826 218898 506382 219454
rect 505826 182898 506382 183454
rect 505826 146898 506382 147454
rect 505826 110898 506382 111454
rect 505826 74898 506382 75454
rect 505826 38898 506382 39454
rect 505826 2898 506382 3454
rect 505826 -902 506382 -346
rect 509546 690618 510102 691174
rect 509546 654618 510102 655174
rect 509546 618618 510102 619174
rect 509546 582618 510102 583174
rect 509546 546618 510102 547174
rect 509546 510618 510102 511174
rect 509546 474618 510102 475174
rect 509546 438618 510102 439174
rect 509546 402618 510102 403174
rect 509546 366618 510102 367174
rect 509546 330618 510102 331174
rect 509546 294618 510102 295174
rect 509546 258618 510102 259174
rect 509546 222618 510102 223174
rect 509546 186618 510102 187174
rect 509546 150618 510102 151174
rect 509546 114618 510102 115174
rect 509546 78618 510102 79174
rect 509546 42618 510102 43174
rect 509546 6618 510102 7174
rect 509546 -2822 510102 -2266
rect 513266 694338 513822 694894
rect 513266 658338 513822 658894
rect 513266 622338 513822 622894
rect 513266 586338 513822 586894
rect 513266 550338 513822 550894
rect 513266 514338 513822 514894
rect 513266 478338 513822 478894
rect 513266 442338 513822 442894
rect 513266 406338 513822 406894
rect 513266 370338 513822 370894
rect 513266 334338 513822 334894
rect 513266 298338 513822 298894
rect 513266 262338 513822 262894
rect 513266 226338 513822 226894
rect 513266 190338 513822 190894
rect 513266 154338 513822 154894
rect 513266 118338 513822 118894
rect 513266 82338 513822 82894
rect 513266 46338 513822 46894
rect 513266 10338 513822 10894
rect 513266 -4742 513822 -4186
rect 534986 711002 535542 711558
rect 531266 709082 531822 709638
rect 527546 707162 528102 707718
rect 516986 698058 517542 698614
rect 516986 662058 517542 662614
rect 516986 626058 517542 626614
rect 516986 590058 517542 590614
rect 516986 554058 517542 554614
rect 516986 518058 517542 518614
rect 516986 482058 517542 482614
rect 516986 446058 517542 446614
rect 516986 410058 517542 410614
rect 516986 374058 517542 374614
rect 516986 338058 517542 338614
rect 516986 302058 517542 302614
rect 516986 266058 517542 266614
rect 516986 230058 517542 230614
rect 516986 194058 517542 194614
rect 516986 158058 517542 158614
rect 516986 122058 517542 122614
rect 516986 86058 517542 86614
rect 516986 50058 517542 50614
rect 516986 14058 517542 14614
rect 498986 -7622 499542 -7066
rect 523826 705242 524382 705798
rect 523826 668898 524382 669454
rect 523826 632898 524382 633454
rect 523826 596898 524382 597454
rect 523826 560898 524382 561454
rect 523826 524898 524382 525454
rect 523826 488898 524382 489454
rect 523826 452898 524382 453454
rect 523826 416898 524382 417454
rect 523826 380898 524382 381454
rect 523826 344898 524382 345454
rect 523826 308898 524382 309454
rect 523826 272898 524382 273454
rect 523826 236898 524382 237454
rect 523826 200898 524382 201454
rect 523826 164898 524382 165454
rect 523826 128898 524382 129454
rect 523826 92898 524382 93454
rect 523826 56898 524382 57454
rect 523826 20898 524382 21454
rect 523826 -1862 524382 -1306
rect 527546 672618 528102 673174
rect 527546 636618 528102 637174
rect 527546 600618 528102 601174
rect 527546 564618 528102 565174
rect 527546 528618 528102 529174
rect 527546 492618 528102 493174
rect 527546 456618 528102 457174
rect 527546 420618 528102 421174
rect 527546 384618 528102 385174
rect 527546 348618 528102 349174
rect 527546 312618 528102 313174
rect 527546 276618 528102 277174
rect 527546 240618 528102 241174
rect 527546 204618 528102 205174
rect 527546 168618 528102 169174
rect 527546 132618 528102 133174
rect 527546 96618 528102 97174
rect 527546 60618 528102 61174
rect 527546 24618 528102 25174
rect 527546 -3782 528102 -3226
rect 531266 676338 531822 676894
rect 531266 640338 531822 640894
rect 531266 604338 531822 604894
rect 531266 568338 531822 568894
rect 531266 532338 531822 532894
rect 531266 496338 531822 496894
rect 531266 460338 531822 460894
rect 531266 424338 531822 424894
rect 531266 388338 531822 388894
rect 531266 352338 531822 352894
rect 531266 316338 531822 316894
rect 531266 280338 531822 280894
rect 531266 244338 531822 244894
rect 531266 208338 531822 208894
rect 531266 172338 531822 172894
rect 531266 136338 531822 136894
rect 531266 100338 531822 100894
rect 531266 64338 531822 64894
rect 531266 28338 531822 28894
rect 531266 -5702 531822 -5146
rect 552986 710042 553542 710598
rect 549266 708122 549822 708678
rect 545546 706202 546102 706758
rect 534986 680058 535542 680614
rect 534986 644058 535542 644614
rect 534986 608058 535542 608614
rect 534986 572058 535542 572614
rect 534986 536058 535542 536614
rect 534986 500058 535542 500614
rect 534986 464058 535542 464614
rect 534986 428058 535542 428614
rect 534986 392058 535542 392614
rect 534986 356058 535542 356614
rect 534986 320058 535542 320614
rect 534986 284058 535542 284614
rect 534986 248058 535542 248614
rect 534986 212058 535542 212614
rect 534986 176058 535542 176614
rect 534986 140058 535542 140614
rect 534986 104058 535542 104614
rect 534986 68058 535542 68614
rect 534986 32058 535542 32614
rect 516986 -6662 517542 -6106
rect 541826 704282 542382 704838
rect 541826 686898 542382 687454
rect 541826 650898 542382 651454
rect 541826 614898 542382 615454
rect 541826 578898 542382 579454
rect 541826 542898 542382 543454
rect 541826 506898 542382 507454
rect 541826 470898 542382 471454
rect 541826 434898 542382 435454
rect 541826 398898 542382 399454
rect 541826 362898 542382 363454
rect 541826 326898 542382 327454
rect 541826 290898 542382 291454
rect 541826 254898 542382 255454
rect 541826 218898 542382 219454
rect 541826 182898 542382 183454
rect 541826 146898 542382 147454
rect 541826 110898 542382 111454
rect 541826 74898 542382 75454
rect 541826 38898 542382 39454
rect 541826 2898 542382 3454
rect 541826 -902 542382 -346
rect 545546 690618 546102 691174
rect 545546 654618 546102 655174
rect 545546 618618 546102 619174
rect 545546 582618 546102 583174
rect 545546 546618 546102 547174
rect 545546 510618 546102 511174
rect 545546 474618 546102 475174
rect 545546 438618 546102 439174
rect 545546 402618 546102 403174
rect 545546 366618 546102 367174
rect 545546 330618 546102 331174
rect 545546 294618 546102 295174
rect 545546 258618 546102 259174
rect 545546 222618 546102 223174
rect 545546 186618 546102 187174
rect 545546 150618 546102 151174
rect 545546 114618 546102 115174
rect 545546 78618 546102 79174
rect 545546 42618 546102 43174
rect 545546 6618 546102 7174
rect 545546 -2822 546102 -2266
rect 549266 694338 549822 694894
rect 549266 658338 549822 658894
rect 549266 622338 549822 622894
rect 549266 586338 549822 586894
rect 549266 550338 549822 550894
rect 549266 514338 549822 514894
rect 549266 478338 549822 478894
rect 549266 442338 549822 442894
rect 549266 406338 549822 406894
rect 549266 370338 549822 370894
rect 549266 334338 549822 334894
rect 549266 298338 549822 298894
rect 549266 262338 549822 262894
rect 549266 226338 549822 226894
rect 549266 190338 549822 190894
rect 549266 154338 549822 154894
rect 549266 118338 549822 118894
rect 549266 82338 549822 82894
rect 549266 46338 549822 46894
rect 549266 10338 549822 10894
rect 549266 -4742 549822 -4186
rect 570986 711002 571542 711558
rect 567266 709082 567822 709638
rect 563546 707162 564102 707718
rect 552986 698058 553542 698614
rect 552986 662058 553542 662614
rect 552986 626058 553542 626614
rect 552986 590058 553542 590614
rect 552986 554058 553542 554614
rect 552986 518058 553542 518614
rect 552986 482058 553542 482614
rect 552986 446058 553542 446614
rect 552986 410058 553542 410614
rect 552986 374058 553542 374614
rect 552986 338058 553542 338614
rect 552986 302058 553542 302614
rect 552986 266058 553542 266614
rect 552986 230058 553542 230614
rect 552986 194058 553542 194614
rect 552986 158058 553542 158614
rect 552986 122058 553542 122614
rect 552986 86058 553542 86614
rect 552986 50058 553542 50614
rect 552986 14058 553542 14614
rect 534986 -7622 535542 -7066
rect 559826 705242 560382 705798
rect 559826 668898 560382 669454
rect 559826 632898 560382 633454
rect 559826 596898 560382 597454
rect 559826 560898 560382 561454
rect 559826 524898 560382 525454
rect 559826 488898 560382 489454
rect 559826 452898 560382 453454
rect 559826 416898 560382 417454
rect 559826 380898 560382 381454
rect 559826 344898 560382 345454
rect 559826 308898 560382 309454
rect 559826 272898 560382 273454
rect 559826 236898 560382 237454
rect 559826 200898 560382 201454
rect 559826 164898 560382 165454
rect 559826 128898 560382 129454
rect 559826 92898 560382 93454
rect 559826 56898 560382 57454
rect 559826 20898 560382 21454
rect 559826 -1862 560382 -1306
rect 563546 672618 564102 673174
rect 563546 636618 564102 637174
rect 563546 600618 564102 601174
rect 563546 564618 564102 565174
rect 563546 528618 564102 529174
rect 563546 492618 564102 493174
rect 563546 456618 564102 457174
rect 563546 420618 564102 421174
rect 563546 384618 564102 385174
rect 563546 348618 564102 349174
rect 563546 312618 564102 313174
rect 563546 276618 564102 277174
rect 563546 240618 564102 241174
rect 563546 204618 564102 205174
rect 563546 168618 564102 169174
rect 563546 132618 564102 133174
rect 563546 96618 564102 97174
rect 563546 60618 564102 61174
rect 563546 24618 564102 25174
rect 563546 -3782 564102 -3226
rect 567266 676338 567822 676894
rect 567266 640338 567822 640894
rect 567266 604338 567822 604894
rect 567266 568338 567822 568894
rect 567266 532338 567822 532894
rect 567266 496338 567822 496894
rect 567266 460338 567822 460894
rect 567266 424338 567822 424894
rect 567266 388338 567822 388894
rect 567266 352338 567822 352894
rect 567266 316338 567822 316894
rect 567266 280338 567822 280894
rect 567266 244338 567822 244894
rect 567266 208338 567822 208894
rect 567266 172338 567822 172894
rect 567266 136338 567822 136894
rect 567266 100338 567822 100894
rect 567266 64338 567822 64894
rect 567266 28338 567822 28894
rect 567266 -5702 567822 -5146
rect 592062 711002 592618 711558
rect 591102 710042 591658 710598
rect 590142 709082 590698 709638
rect 589182 708122 589738 708678
rect 588222 707162 588778 707718
rect 581546 706202 582102 706758
rect 570986 680058 571542 680614
rect 570986 644058 571542 644614
rect 570986 608058 571542 608614
rect 570986 572058 571542 572614
rect 570986 536058 571542 536614
rect 570986 500058 571542 500614
rect 570986 464058 571542 464614
rect 570986 428058 571542 428614
rect 570986 392058 571542 392614
rect 570986 356058 571542 356614
rect 570986 320058 571542 320614
rect 570986 284058 571542 284614
rect 570986 248058 571542 248614
rect 570986 212058 571542 212614
rect 570986 176058 571542 176614
rect 570986 140058 571542 140614
rect 570986 104058 571542 104614
rect 570986 68058 571542 68614
rect 570986 32058 571542 32614
rect 552986 -6662 553542 -6106
rect 577826 704282 578382 704838
rect 577826 686898 578382 687454
rect 577826 650898 578382 651454
rect 577826 614898 578382 615454
rect 577826 578898 578382 579454
rect 577826 542898 578382 543454
rect 577826 506898 578382 507454
rect 577826 470898 578382 471454
rect 587262 706202 587818 706758
rect 586302 705242 586858 705798
rect 581546 690618 582102 691174
rect 581546 654618 582102 655174
rect 581546 618618 582102 619174
rect 581546 582618 582102 583174
rect 581546 546618 582102 547174
rect 581546 510618 582102 511174
rect 581546 474618 582102 475174
rect 577826 434898 578382 435454
rect 577826 398898 578382 399454
rect 577826 362898 578382 363454
rect 577826 326898 578382 327454
rect 577826 290898 578382 291454
rect 577826 254898 578382 255454
rect 577826 218898 578382 219454
rect 577826 182898 578382 183454
rect 577826 146898 578382 147454
rect 577826 110898 578382 111454
rect 577826 74898 578382 75454
rect 581546 438618 582102 439174
rect 581546 402618 582102 403174
rect 581546 366618 582102 367174
rect 581546 330618 582102 331174
rect 581546 294618 582102 295174
rect 581546 258618 582102 259174
rect 581546 222618 582102 223174
rect 581546 186618 582102 187174
rect 581546 150618 582102 151174
rect 581546 114618 582102 115174
rect 581546 78618 582102 79174
rect 577826 38898 578382 39454
rect 577826 2898 578382 3454
rect 577826 -902 578382 -346
rect 581546 42618 582102 43174
rect 581546 6618 582102 7174
rect 585342 704282 585898 704838
rect 585342 686898 585898 687454
rect 585342 650898 585898 651454
rect 585342 614898 585898 615454
rect 585342 578898 585898 579454
rect 585342 542898 585898 543454
rect 585342 506898 585898 507454
rect 585342 470898 585898 471454
rect 585342 434898 585898 435454
rect 585342 398898 585898 399454
rect 585342 362898 585898 363454
rect 585342 326898 585898 327454
rect 585342 290898 585898 291454
rect 585342 254898 585898 255454
rect 585342 218898 585898 219454
rect 585342 182898 585898 183454
rect 585342 146898 585898 147454
rect 585342 110898 585898 111454
rect 585342 74898 585898 75454
rect 585342 38898 585898 39454
rect 585342 2898 585898 3454
rect 585342 -902 585898 -346
rect 586302 668898 586858 669454
rect 586302 632898 586858 633454
rect 586302 596898 586858 597454
rect 586302 560898 586858 561454
rect 586302 524898 586858 525454
rect 586302 488898 586858 489454
rect 586302 452898 586858 453454
rect 586302 416898 586858 417454
rect 586302 380898 586858 381454
rect 586302 344898 586858 345454
rect 586302 308898 586858 309454
rect 586302 272898 586858 273454
rect 586302 236898 586858 237454
rect 586302 200898 586858 201454
rect 586302 164898 586858 165454
rect 586302 128898 586858 129454
rect 586302 92898 586858 93454
rect 586302 56898 586858 57454
rect 586302 20898 586858 21454
rect 586302 -1862 586858 -1306
rect 587262 690618 587818 691174
rect 587262 654618 587818 655174
rect 587262 618618 587818 619174
rect 587262 582618 587818 583174
rect 587262 546618 587818 547174
rect 587262 510618 587818 511174
rect 587262 474618 587818 475174
rect 587262 438618 587818 439174
rect 587262 402618 587818 403174
rect 587262 366618 587818 367174
rect 587262 330618 587818 331174
rect 587262 294618 587818 295174
rect 587262 258618 587818 259174
rect 587262 222618 587818 223174
rect 587262 186618 587818 187174
rect 587262 150618 587818 151174
rect 587262 114618 587818 115174
rect 587262 78618 587818 79174
rect 587262 42618 587818 43174
rect 587262 6618 587818 7174
rect 581546 -2822 582102 -2266
rect 587262 -2822 587818 -2266
rect 588222 672618 588778 673174
rect 588222 636618 588778 637174
rect 588222 600618 588778 601174
rect 588222 564618 588778 565174
rect 588222 528618 588778 529174
rect 588222 492618 588778 493174
rect 588222 456618 588778 457174
rect 588222 420618 588778 421174
rect 588222 384618 588778 385174
rect 588222 348618 588778 349174
rect 588222 312618 588778 313174
rect 588222 276618 588778 277174
rect 588222 240618 588778 241174
rect 588222 204618 588778 205174
rect 588222 168618 588778 169174
rect 588222 132618 588778 133174
rect 588222 96618 588778 97174
rect 588222 60618 588778 61174
rect 588222 24618 588778 25174
rect 588222 -3782 588778 -3226
rect 589182 694338 589738 694894
rect 589182 658338 589738 658894
rect 589182 622338 589738 622894
rect 589182 586338 589738 586894
rect 589182 550338 589738 550894
rect 589182 514338 589738 514894
rect 589182 478338 589738 478894
rect 589182 442338 589738 442894
rect 589182 406338 589738 406894
rect 589182 370338 589738 370894
rect 589182 334338 589738 334894
rect 589182 298338 589738 298894
rect 589182 262338 589738 262894
rect 589182 226338 589738 226894
rect 589182 190338 589738 190894
rect 589182 154338 589738 154894
rect 589182 118338 589738 118894
rect 589182 82338 589738 82894
rect 589182 46338 589738 46894
rect 589182 10338 589738 10894
rect 589182 -4742 589738 -4186
rect 590142 676338 590698 676894
rect 590142 640338 590698 640894
rect 590142 604338 590698 604894
rect 590142 568338 590698 568894
rect 590142 532338 590698 532894
rect 590142 496338 590698 496894
rect 590142 460338 590698 460894
rect 590142 424338 590698 424894
rect 590142 388338 590698 388894
rect 590142 352338 590698 352894
rect 590142 316338 590698 316894
rect 590142 280338 590698 280894
rect 590142 244338 590698 244894
rect 590142 208338 590698 208894
rect 590142 172338 590698 172894
rect 590142 136338 590698 136894
rect 590142 100338 590698 100894
rect 590142 64338 590698 64894
rect 590142 28338 590698 28894
rect 590142 -5702 590698 -5146
rect 591102 698058 591658 698614
rect 591102 662058 591658 662614
rect 591102 626058 591658 626614
rect 591102 590058 591658 590614
rect 591102 554058 591658 554614
rect 591102 518058 591658 518614
rect 591102 482058 591658 482614
rect 591102 446058 591658 446614
rect 591102 410058 591658 410614
rect 591102 374058 591658 374614
rect 591102 338058 591658 338614
rect 591102 302058 591658 302614
rect 591102 266058 591658 266614
rect 591102 230058 591658 230614
rect 591102 194058 591658 194614
rect 591102 158058 591658 158614
rect 591102 122058 591658 122614
rect 591102 86058 591658 86614
rect 591102 50058 591658 50614
rect 591102 14058 591658 14614
rect 591102 -6662 591658 -6106
rect 592062 680058 592618 680614
rect 592062 644058 592618 644614
rect 592062 608058 592618 608614
rect 592062 572058 592618 572614
rect 592062 536058 592618 536614
rect 592062 500058 592618 500614
rect 592062 464058 592618 464614
rect 592062 428058 592618 428614
rect 592062 392058 592618 392614
rect 592062 356058 592618 356614
rect 592062 320058 592618 320614
rect 592062 284058 592618 284614
rect 592062 248058 592618 248614
rect 592062 212058 592618 212614
rect 592062 176058 592618 176614
rect 592062 140058 592618 140614
rect 592062 104058 592618 104614
rect 592062 68058 592618 68614
rect 592062 32058 592618 32614
rect 570986 -7622 571542 -7066
rect 592062 -7622 592618 -7066
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711002 -8694 711558
rect -8138 711002 30986 711558
rect 31542 711002 66986 711558
rect 67542 711002 102986 711558
rect 103542 711002 138986 711558
rect 139542 711002 174986 711558
rect 175542 711002 210986 711558
rect 211542 711002 246986 711558
rect 247542 711002 282986 711558
rect 283542 711002 318986 711558
rect 319542 711002 354986 711558
rect 355542 711002 390986 711558
rect 391542 711002 426986 711558
rect 427542 711002 462986 711558
rect 463542 711002 498986 711558
rect 499542 711002 534986 711558
rect 535542 711002 570986 711558
rect 571542 711002 592062 711558
rect 592618 711002 592650 711558
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710042 -7734 710598
rect -7178 710042 12986 710598
rect 13542 710042 48986 710598
rect 49542 710042 84986 710598
rect 85542 710042 120986 710598
rect 121542 710042 156986 710598
rect 157542 710042 192986 710598
rect 193542 710042 228986 710598
rect 229542 710042 264986 710598
rect 265542 710042 300986 710598
rect 301542 710042 336986 710598
rect 337542 710042 372986 710598
rect 373542 710042 408986 710598
rect 409542 710042 444986 710598
rect 445542 710042 480986 710598
rect 481542 710042 516986 710598
rect 517542 710042 552986 710598
rect 553542 710042 591102 710598
rect 591658 710042 591690 710598
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709082 -6774 709638
rect -6218 709082 27266 709638
rect 27822 709082 63266 709638
rect 63822 709082 99266 709638
rect 99822 709082 135266 709638
rect 135822 709082 171266 709638
rect 171822 709082 207266 709638
rect 207822 709082 243266 709638
rect 243822 709082 279266 709638
rect 279822 709082 315266 709638
rect 315822 709082 351266 709638
rect 351822 709082 387266 709638
rect 387822 709082 423266 709638
rect 423822 709082 459266 709638
rect 459822 709082 495266 709638
rect 495822 709082 531266 709638
rect 531822 709082 567266 709638
rect 567822 709082 590142 709638
rect 590698 709082 590730 709638
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708122 -5814 708678
rect -5258 708122 9266 708678
rect 9822 708122 45266 708678
rect 45822 708122 81266 708678
rect 81822 708122 117266 708678
rect 117822 708122 153266 708678
rect 153822 708122 189266 708678
rect 189822 708122 225266 708678
rect 225822 708122 261266 708678
rect 261822 708122 297266 708678
rect 297822 708122 333266 708678
rect 333822 708122 369266 708678
rect 369822 708122 405266 708678
rect 405822 708122 441266 708678
rect 441822 708122 477266 708678
rect 477822 708122 513266 708678
rect 513822 708122 549266 708678
rect 549822 708122 589182 708678
rect 589738 708122 589770 708678
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707162 -4854 707718
rect -4298 707162 23546 707718
rect 24102 707162 59546 707718
rect 60102 707162 95546 707718
rect 96102 707162 131546 707718
rect 132102 707162 167546 707718
rect 168102 707162 203546 707718
rect 204102 707162 239546 707718
rect 240102 707162 275546 707718
rect 276102 707162 311546 707718
rect 312102 707162 347546 707718
rect 348102 707162 383546 707718
rect 384102 707162 419546 707718
rect 420102 707162 455546 707718
rect 456102 707162 491546 707718
rect 492102 707162 527546 707718
rect 528102 707162 563546 707718
rect 564102 707162 588222 707718
rect 588778 707162 588810 707718
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706202 -3894 706758
rect -3338 706202 5546 706758
rect 6102 706202 41546 706758
rect 42102 706202 77546 706758
rect 78102 706202 113546 706758
rect 114102 706202 149546 706758
rect 150102 706202 185546 706758
rect 186102 706202 221546 706758
rect 222102 706202 257546 706758
rect 258102 706202 293546 706758
rect 294102 706202 329546 706758
rect 330102 706202 365546 706758
rect 366102 706202 401546 706758
rect 402102 706202 437546 706758
rect 438102 706202 473546 706758
rect 474102 706202 509546 706758
rect 510102 706202 545546 706758
rect 546102 706202 581546 706758
rect 582102 706202 587262 706758
rect 587818 706202 587850 706758
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705242 -2934 705798
rect -2378 705242 19826 705798
rect 20382 705242 55826 705798
rect 56382 705242 91826 705798
rect 92382 705242 127826 705798
rect 128382 705242 163826 705798
rect 164382 705242 199826 705798
rect 200382 705242 235826 705798
rect 236382 705242 271826 705798
rect 272382 705242 307826 705798
rect 308382 705242 343826 705798
rect 344382 705242 379826 705798
rect 380382 705242 415826 705798
rect 416382 705242 451826 705798
rect 452382 705242 487826 705798
rect 488382 705242 523826 705798
rect 524382 705242 559826 705798
rect 560382 705242 586302 705798
rect 586858 705242 586890 705798
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704282 -1974 704838
rect -1418 704282 1826 704838
rect 2382 704282 37826 704838
rect 38382 704282 73826 704838
rect 74382 704282 109826 704838
rect 110382 704282 145826 704838
rect 146382 704282 181826 704838
rect 182382 704282 217826 704838
rect 218382 704282 253826 704838
rect 254382 704282 289826 704838
rect 290382 704282 325826 704838
rect 326382 704282 361826 704838
rect 362382 704282 397826 704838
rect 398382 704282 433826 704838
rect 434382 704282 469826 704838
rect 470382 704282 505826 704838
rect 506382 704282 541826 704838
rect 542382 704282 577826 704838
rect 578382 704282 585342 704838
rect 585898 704282 585930 704838
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698058 -7734 698614
rect -7178 698058 12986 698614
rect 13542 698058 48986 698614
rect 49542 698058 84986 698614
rect 85542 698058 120986 698614
rect 121542 698058 156986 698614
rect 157542 698058 192986 698614
rect 193542 698058 228986 698614
rect 229542 698058 264986 698614
rect 265542 698058 300986 698614
rect 301542 698058 336986 698614
rect 337542 698058 372986 698614
rect 373542 698058 408986 698614
rect 409542 698058 444986 698614
rect 445542 698058 480986 698614
rect 481542 698058 516986 698614
rect 517542 698058 552986 698614
rect 553542 698058 591102 698614
rect 591658 698058 592650 698614
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694338 -5814 694894
rect -5258 694338 9266 694894
rect 9822 694338 45266 694894
rect 45822 694338 81266 694894
rect 81822 694338 117266 694894
rect 117822 694338 153266 694894
rect 153822 694338 189266 694894
rect 189822 694338 225266 694894
rect 225822 694338 261266 694894
rect 261822 694338 297266 694894
rect 297822 694338 333266 694894
rect 333822 694338 369266 694894
rect 369822 694338 405266 694894
rect 405822 694338 441266 694894
rect 441822 694338 477266 694894
rect 477822 694338 513266 694894
rect 513822 694338 549266 694894
rect 549822 694338 589182 694894
rect 589738 694338 590730 694894
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690618 -3894 691174
rect -3338 690618 5546 691174
rect 6102 690618 41546 691174
rect 42102 690618 77546 691174
rect 78102 690618 113546 691174
rect 114102 690618 149546 691174
rect 150102 690618 185546 691174
rect 186102 690618 221546 691174
rect 222102 690618 257546 691174
rect 258102 690618 293546 691174
rect 294102 690618 329546 691174
rect 330102 690618 365546 691174
rect 366102 690618 401546 691174
rect 402102 690618 437546 691174
rect 438102 690618 473546 691174
rect 474102 690618 509546 691174
rect 510102 690618 545546 691174
rect 546102 690618 581546 691174
rect 582102 690618 587262 691174
rect 587818 690618 588810 691174
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 686898 -1974 687454
rect -1418 686898 1826 687454
rect 2382 686898 37826 687454
rect 38382 686898 73826 687454
rect 74382 686898 109826 687454
rect 110382 686898 145826 687454
rect 146382 686898 181826 687454
rect 182382 686898 217826 687454
rect 218382 686898 253826 687454
rect 254382 686898 289826 687454
rect 290382 686898 325826 687454
rect 326382 686898 361826 687454
rect 362382 686898 397826 687454
rect 398382 686898 433826 687454
rect 434382 686898 469826 687454
rect 470382 686898 505826 687454
rect 506382 686898 541826 687454
rect 542382 686898 577826 687454
rect 578382 686898 585342 687454
rect 585898 686898 586890 687454
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680058 -8694 680614
rect -8138 680058 30986 680614
rect 31542 680058 66986 680614
rect 67542 680058 102986 680614
rect 103542 680058 138986 680614
rect 139542 680058 174986 680614
rect 175542 680058 210986 680614
rect 211542 680058 246986 680614
rect 247542 680058 282986 680614
rect 283542 680058 318986 680614
rect 319542 680058 354986 680614
rect 355542 680058 390986 680614
rect 391542 680058 426986 680614
rect 427542 680058 462986 680614
rect 463542 680058 498986 680614
rect 499542 680058 534986 680614
rect 535542 680058 570986 680614
rect 571542 680058 592062 680614
rect 592618 680058 592650 680614
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676338 -6774 676894
rect -6218 676338 27266 676894
rect 27822 676338 63266 676894
rect 63822 676338 99266 676894
rect 99822 676338 135266 676894
rect 135822 676338 171266 676894
rect 171822 676338 207266 676894
rect 207822 676338 243266 676894
rect 243822 676338 279266 676894
rect 279822 676338 315266 676894
rect 315822 676338 351266 676894
rect 351822 676338 387266 676894
rect 387822 676338 423266 676894
rect 423822 676338 459266 676894
rect 459822 676338 495266 676894
rect 495822 676338 531266 676894
rect 531822 676338 567266 676894
rect 567822 676338 590142 676894
rect 590698 676338 590730 676894
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672618 -4854 673174
rect -4298 672618 23546 673174
rect 24102 672618 59546 673174
rect 60102 672618 95546 673174
rect 96102 672618 131546 673174
rect 132102 672618 167546 673174
rect 168102 672618 203546 673174
rect 204102 672618 239546 673174
rect 240102 672618 275546 673174
rect 276102 672618 311546 673174
rect 312102 672618 347546 673174
rect 348102 672618 383546 673174
rect 384102 672618 419546 673174
rect 420102 672618 455546 673174
rect 456102 672618 491546 673174
rect 492102 672618 527546 673174
rect 528102 672618 563546 673174
rect 564102 672618 588222 673174
rect 588778 672618 588810 673174
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 668898 -2934 669454
rect -2378 668898 19826 669454
rect 20382 668898 55826 669454
rect 56382 668898 91826 669454
rect 92382 668898 127826 669454
rect 128382 668898 163826 669454
rect 164382 668898 199826 669454
rect 200382 668898 235826 669454
rect 236382 668898 271826 669454
rect 272382 668898 307826 669454
rect 308382 668898 343826 669454
rect 344382 668898 379826 669454
rect 380382 668898 415826 669454
rect 416382 668898 451826 669454
rect 452382 668898 487826 669454
rect 488382 668898 523826 669454
rect 524382 668898 559826 669454
rect 560382 668898 586302 669454
rect 586858 668898 586890 669454
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662058 -7734 662614
rect -7178 662058 12986 662614
rect 13542 662058 48986 662614
rect 49542 662058 84986 662614
rect 85542 662058 120986 662614
rect 121542 662058 156986 662614
rect 157542 662058 192986 662614
rect 193542 662058 228986 662614
rect 229542 662058 264986 662614
rect 265542 662058 300986 662614
rect 301542 662058 336986 662614
rect 337542 662058 372986 662614
rect 373542 662058 408986 662614
rect 409542 662058 444986 662614
rect 445542 662058 480986 662614
rect 481542 662058 516986 662614
rect 517542 662058 552986 662614
rect 553542 662058 591102 662614
rect 591658 662058 592650 662614
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658338 -5814 658894
rect -5258 658338 9266 658894
rect 9822 658338 45266 658894
rect 45822 658338 81266 658894
rect 81822 658338 117266 658894
rect 117822 658338 153266 658894
rect 153822 658338 189266 658894
rect 189822 658338 225266 658894
rect 225822 658338 261266 658894
rect 261822 658338 297266 658894
rect 297822 658338 333266 658894
rect 333822 658338 369266 658894
rect 369822 658338 405266 658894
rect 405822 658338 441266 658894
rect 441822 658338 477266 658894
rect 477822 658338 513266 658894
rect 513822 658338 549266 658894
rect 549822 658338 589182 658894
rect 589738 658338 590730 658894
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654618 -3894 655174
rect -3338 654618 5546 655174
rect 6102 654618 41546 655174
rect 42102 654618 77546 655174
rect 78102 654618 113546 655174
rect 114102 654618 149546 655174
rect 150102 654618 185546 655174
rect 186102 654618 221546 655174
rect 222102 654618 257546 655174
rect 258102 654618 293546 655174
rect 294102 654618 329546 655174
rect 330102 654618 365546 655174
rect 366102 654618 401546 655174
rect 402102 654618 437546 655174
rect 438102 654618 473546 655174
rect 474102 654618 509546 655174
rect 510102 654618 545546 655174
rect 546102 654618 581546 655174
rect 582102 654618 587262 655174
rect 587818 654618 588810 655174
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 650898 -1974 651454
rect -1418 650898 1826 651454
rect 2382 650898 37826 651454
rect 38382 650898 73826 651454
rect 74382 650898 109826 651454
rect 110382 650898 145826 651454
rect 146382 650898 181826 651454
rect 182382 650898 217826 651454
rect 218382 650898 253826 651454
rect 254382 650898 289826 651454
rect 290382 650898 325826 651454
rect 326382 650898 361826 651454
rect 362382 650898 397826 651454
rect 398382 650898 433826 651454
rect 434382 650898 469826 651454
rect 470382 650898 505826 651454
rect 506382 650898 541826 651454
rect 542382 650898 577826 651454
rect 578382 650898 585342 651454
rect 585898 650898 586890 651454
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644058 -8694 644614
rect -8138 644058 30986 644614
rect 31542 644058 66986 644614
rect 67542 644058 102986 644614
rect 103542 644058 138986 644614
rect 139542 644058 174986 644614
rect 175542 644058 210986 644614
rect 211542 644058 246986 644614
rect 247542 644058 282986 644614
rect 283542 644058 318986 644614
rect 319542 644058 354986 644614
rect 355542 644058 390986 644614
rect 391542 644058 426986 644614
rect 427542 644058 462986 644614
rect 463542 644058 498986 644614
rect 499542 644058 534986 644614
rect 535542 644058 570986 644614
rect 571542 644058 592062 644614
rect 592618 644058 592650 644614
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640338 -6774 640894
rect -6218 640338 27266 640894
rect 27822 640338 63266 640894
rect 63822 640338 99266 640894
rect 99822 640338 135266 640894
rect 135822 640338 171266 640894
rect 171822 640338 207266 640894
rect 207822 640338 243266 640894
rect 243822 640338 279266 640894
rect 279822 640338 315266 640894
rect 315822 640338 351266 640894
rect 351822 640338 387266 640894
rect 387822 640338 423266 640894
rect 423822 640338 459266 640894
rect 459822 640338 495266 640894
rect 495822 640338 531266 640894
rect 531822 640338 567266 640894
rect 567822 640338 590142 640894
rect 590698 640338 590730 640894
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636618 -4854 637174
rect -4298 636618 23546 637174
rect 24102 636618 59546 637174
rect 60102 636618 95546 637174
rect 96102 636618 131546 637174
rect 132102 636618 167546 637174
rect 168102 636618 203546 637174
rect 204102 636618 239546 637174
rect 240102 636618 275546 637174
rect 276102 636618 311546 637174
rect 312102 636618 347546 637174
rect 348102 636618 383546 637174
rect 384102 636618 419546 637174
rect 420102 636618 455546 637174
rect 456102 636618 491546 637174
rect 492102 636618 527546 637174
rect 528102 636618 563546 637174
rect 564102 636618 588222 637174
rect 588778 636618 588810 637174
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 632898 -2934 633454
rect -2378 632898 19826 633454
rect 20382 632898 55826 633454
rect 56382 632898 91826 633454
rect 92382 632898 127826 633454
rect 128382 632898 163826 633454
rect 164382 632898 199826 633454
rect 200382 632898 235826 633454
rect 236382 632898 271826 633454
rect 272382 632898 307826 633454
rect 308382 632898 343826 633454
rect 344382 632898 379826 633454
rect 380382 632898 415826 633454
rect 416382 632898 451826 633454
rect 452382 632898 487826 633454
rect 488382 632898 523826 633454
rect 524382 632898 559826 633454
rect 560382 632898 586302 633454
rect 586858 632898 586890 633454
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626058 -7734 626614
rect -7178 626058 12986 626614
rect 13542 626058 48986 626614
rect 49542 626058 84986 626614
rect 85542 626058 120986 626614
rect 121542 626058 156986 626614
rect 157542 626058 192986 626614
rect 193542 626058 228986 626614
rect 229542 626058 264986 626614
rect 265542 626058 300986 626614
rect 301542 626058 336986 626614
rect 337542 626058 372986 626614
rect 373542 626058 408986 626614
rect 409542 626058 444986 626614
rect 445542 626058 480986 626614
rect 481542 626058 516986 626614
rect 517542 626058 552986 626614
rect 553542 626058 591102 626614
rect 591658 626058 592650 626614
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622338 -5814 622894
rect -5258 622338 9266 622894
rect 9822 622338 45266 622894
rect 45822 622338 81266 622894
rect 81822 622338 117266 622894
rect 117822 622338 153266 622894
rect 153822 622338 189266 622894
rect 189822 622338 225266 622894
rect 225822 622338 261266 622894
rect 261822 622338 297266 622894
rect 297822 622338 333266 622894
rect 333822 622338 369266 622894
rect 369822 622338 405266 622894
rect 405822 622338 441266 622894
rect 441822 622338 477266 622894
rect 477822 622338 513266 622894
rect 513822 622338 549266 622894
rect 549822 622338 589182 622894
rect 589738 622338 590730 622894
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618618 -3894 619174
rect -3338 618618 5546 619174
rect 6102 618618 41546 619174
rect 42102 618618 77546 619174
rect 78102 618618 113546 619174
rect 114102 618618 149546 619174
rect 150102 618618 185546 619174
rect 186102 618618 221546 619174
rect 222102 618618 257546 619174
rect 258102 618618 293546 619174
rect 294102 618618 329546 619174
rect 330102 618618 365546 619174
rect 366102 618618 401546 619174
rect 402102 618618 437546 619174
rect 438102 618618 473546 619174
rect 474102 618618 509546 619174
rect 510102 618618 545546 619174
rect 546102 618618 581546 619174
rect 582102 618618 587262 619174
rect 587818 618618 588810 619174
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 614898 -1974 615454
rect -1418 614898 1826 615454
rect 2382 614898 37826 615454
rect 38382 614898 73826 615454
rect 74382 614898 109826 615454
rect 110382 614898 145826 615454
rect 146382 614898 181826 615454
rect 182382 614898 217826 615454
rect 218382 614898 253826 615454
rect 254382 614898 289826 615454
rect 290382 614898 325826 615454
rect 326382 614898 361826 615454
rect 362382 614898 397826 615454
rect 398382 614898 433826 615454
rect 434382 614898 469826 615454
rect 470382 614898 505826 615454
rect 506382 614898 541826 615454
rect 542382 614898 577826 615454
rect 578382 614898 585342 615454
rect 585898 614898 586890 615454
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608058 -8694 608614
rect -8138 608058 30986 608614
rect 31542 608058 66986 608614
rect 67542 608058 102986 608614
rect 103542 608058 138986 608614
rect 139542 608058 174986 608614
rect 175542 608058 210986 608614
rect 211542 608058 246986 608614
rect 247542 608058 282986 608614
rect 283542 608058 318986 608614
rect 319542 608058 354986 608614
rect 355542 608058 390986 608614
rect 391542 608058 426986 608614
rect 427542 608058 462986 608614
rect 463542 608058 498986 608614
rect 499542 608058 534986 608614
rect 535542 608058 570986 608614
rect 571542 608058 592062 608614
rect 592618 608058 592650 608614
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604338 -6774 604894
rect -6218 604338 27266 604894
rect 27822 604338 63266 604894
rect 63822 604338 99266 604894
rect 99822 604338 135266 604894
rect 135822 604338 171266 604894
rect 171822 604338 207266 604894
rect 207822 604338 243266 604894
rect 243822 604338 279266 604894
rect 279822 604338 315266 604894
rect 315822 604338 351266 604894
rect 351822 604338 387266 604894
rect 387822 604338 423266 604894
rect 423822 604338 459266 604894
rect 459822 604338 495266 604894
rect 495822 604338 531266 604894
rect 531822 604338 567266 604894
rect 567822 604338 590142 604894
rect 590698 604338 590730 604894
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600618 -4854 601174
rect -4298 600618 23546 601174
rect 24102 600618 59546 601174
rect 60102 600618 95546 601174
rect 96102 600618 131546 601174
rect 132102 600618 167546 601174
rect 168102 600618 203546 601174
rect 204102 600618 239546 601174
rect 240102 600618 275546 601174
rect 276102 600618 311546 601174
rect 312102 600618 347546 601174
rect 348102 600618 383546 601174
rect 384102 600618 419546 601174
rect 420102 600618 455546 601174
rect 456102 600618 491546 601174
rect 492102 600618 527546 601174
rect 528102 600618 563546 601174
rect 564102 600618 588222 601174
rect 588778 600618 588810 601174
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 596898 -2934 597454
rect -2378 596898 19826 597454
rect 20382 596898 55826 597454
rect 56382 596898 91826 597454
rect 92382 596898 127826 597454
rect 128382 596898 163826 597454
rect 164382 596898 199826 597454
rect 200382 596898 235826 597454
rect 236382 596898 271826 597454
rect 272382 596898 307826 597454
rect 308382 596898 343826 597454
rect 344382 596898 379826 597454
rect 380382 596898 415826 597454
rect 416382 596898 451826 597454
rect 452382 596898 487826 597454
rect 488382 596898 523826 597454
rect 524382 596898 559826 597454
rect 560382 596898 586302 597454
rect 586858 596898 586890 597454
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590058 -7734 590614
rect -7178 590058 12986 590614
rect 13542 590058 48986 590614
rect 49542 590058 84986 590614
rect 85542 590058 120986 590614
rect 121542 590058 156986 590614
rect 157542 590058 192986 590614
rect 193542 590058 228986 590614
rect 229542 590058 264986 590614
rect 265542 590058 300986 590614
rect 301542 590058 336986 590614
rect 337542 590058 372986 590614
rect 373542 590058 408986 590614
rect 409542 590058 444986 590614
rect 445542 590058 480986 590614
rect 481542 590058 516986 590614
rect 517542 590058 552986 590614
rect 553542 590058 591102 590614
rect 591658 590058 592650 590614
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586338 -5814 586894
rect -5258 586338 9266 586894
rect 9822 586338 45266 586894
rect 45822 586338 81266 586894
rect 81822 586338 117266 586894
rect 117822 586338 153266 586894
rect 153822 586338 189266 586894
rect 189822 586338 225266 586894
rect 225822 586338 261266 586894
rect 261822 586338 297266 586894
rect 297822 586338 333266 586894
rect 333822 586338 369266 586894
rect 369822 586338 405266 586894
rect 405822 586338 441266 586894
rect 441822 586338 477266 586894
rect 477822 586338 513266 586894
rect 513822 586338 549266 586894
rect 549822 586338 589182 586894
rect 589738 586338 590730 586894
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582618 -3894 583174
rect -3338 582618 5546 583174
rect 6102 582618 41546 583174
rect 42102 582618 77546 583174
rect 78102 582618 113546 583174
rect 114102 582618 149546 583174
rect 150102 582618 185546 583174
rect 186102 582618 221546 583174
rect 222102 582618 257546 583174
rect 258102 582618 293546 583174
rect 294102 582618 329546 583174
rect 330102 582618 365546 583174
rect 366102 582618 401546 583174
rect 402102 582618 437546 583174
rect 438102 582618 473546 583174
rect 474102 582618 509546 583174
rect 510102 582618 545546 583174
rect 546102 582618 581546 583174
rect 582102 582618 587262 583174
rect 587818 582618 588810 583174
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 578898 -1974 579454
rect -1418 578898 1826 579454
rect 2382 578898 37826 579454
rect 38382 578898 73826 579454
rect 74382 578898 109826 579454
rect 110382 578898 145826 579454
rect 146382 578898 181826 579454
rect 182382 578898 217826 579454
rect 218382 578898 253826 579454
rect 254382 578898 289826 579454
rect 290382 578898 325826 579454
rect 326382 578898 361826 579454
rect 362382 578898 397826 579454
rect 398382 578898 433826 579454
rect 434382 578898 469826 579454
rect 470382 578898 505826 579454
rect 506382 578898 541826 579454
rect 542382 578898 577826 579454
rect 578382 578898 585342 579454
rect 585898 578898 586890 579454
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572058 -8694 572614
rect -8138 572058 30986 572614
rect 31542 572058 66986 572614
rect 67542 572058 102986 572614
rect 103542 572058 138986 572614
rect 139542 572058 174986 572614
rect 175542 572058 210986 572614
rect 211542 572058 246986 572614
rect 247542 572058 282986 572614
rect 283542 572058 318986 572614
rect 319542 572058 354986 572614
rect 355542 572058 390986 572614
rect 391542 572058 426986 572614
rect 427542 572058 462986 572614
rect 463542 572058 498986 572614
rect 499542 572058 534986 572614
rect 535542 572058 570986 572614
rect 571542 572058 592062 572614
rect 592618 572058 592650 572614
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568338 -6774 568894
rect -6218 568338 27266 568894
rect 27822 568338 63266 568894
rect 63822 568338 99266 568894
rect 99822 568338 135266 568894
rect 135822 568338 171266 568894
rect 171822 568338 207266 568894
rect 207822 568338 243266 568894
rect 243822 568338 279266 568894
rect 279822 568338 315266 568894
rect 315822 568338 351266 568894
rect 351822 568338 387266 568894
rect 387822 568338 423266 568894
rect 423822 568338 459266 568894
rect 459822 568338 495266 568894
rect 495822 568338 531266 568894
rect 531822 568338 567266 568894
rect 567822 568338 590142 568894
rect 590698 568338 590730 568894
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564618 -4854 565174
rect -4298 564618 23546 565174
rect 24102 564618 59546 565174
rect 60102 564618 95546 565174
rect 96102 564618 131546 565174
rect 132102 564618 167546 565174
rect 168102 564618 203546 565174
rect 204102 564618 239546 565174
rect 240102 564618 275546 565174
rect 276102 564618 311546 565174
rect 312102 564618 347546 565174
rect 348102 564618 383546 565174
rect 384102 564618 419546 565174
rect 420102 564618 455546 565174
rect 456102 564618 491546 565174
rect 492102 564618 527546 565174
rect 528102 564618 563546 565174
rect 564102 564618 588222 565174
rect 588778 564618 588810 565174
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 560898 -2934 561454
rect -2378 560898 19826 561454
rect 20382 560898 55826 561454
rect 56382 560898 91826 561454
rect 92382 560898 127826 561454
rect 128382 560898 163826 561454
rect 164382 560898 199826 561454
rect 200382 560898 235826 561454
rect 236382 560898 271826 561454
rect 272382 560898 307826 561454
rect 308382 560898 343826 561454
rect 344382 560898 379826 561454
rect 380382 560898 415826 561454
rect 416382 560898 451826 561454
rect 452382 560898 487826 561454
rect 488382 560898 523826 561454
rect 524382 560898 559826 561454
rect 560382 560898 586302 561454
rect 586858 560898 586890 561454
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554058 -7734 554614
rect -7178 554058 12986 554614
rect 13542 554058 48986 554614
rect 49542 554058 84986 554614
rect 85542 554058 120986 554614
rect 121542 554058 156986 554614
rect 157542 554058 192986 554614
rect 193542 554058 228986 554614
rect 229542 554058 264986 554614
rect 265542 554058 300986 554614
rect 301542 554058 336986 554614
rect 337542 554058 372986 554614
rect 373542 554058 408986 554614
rect 409542 554058 444986 554614
rect 445542 554058 480986 554614
rect 481542 554058 516986 554614
rect 517542 554058 552986 554614
rect 553542 554058 591102 554614
rect 591658 554058 592650 554614
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550338 -5814 550894
rect -5258 550338 9266 550894
rect 9822 550338 45266 550894
rect 45822 550338 81266 550894
rect 81822 550338 117266 550894
rect 117822 550338 153266 550894
rect 153822 550338 189266 550894
rect 189822 550338 225266 550894
rect 225822 550338 261266 550894
rect 261822 550338 297266 550894
rect 297822 550338 333266 550894
rect 333822 550338 369266 550894
rect 369822 550338 405266 550894
rect 405822 550338 441266 550894
rect 441822 550338 477266 550894
rect 477822 550338 513266 550894
rect 513822 550338 549266 550894
rect 549822 550338 589182 550894
rect 589738 550338 590730 550894
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546618 -3894 547174
rect -3338 546618 5546 547174
rect 6102 546618 41546 547174
rect 42102 546618 77546 547174
rect 78102 546618 113546 547174
rect 114102 546618 149546 547174
rect 150102 546618 185546 547174
rect 186102 546618 221546 547174
rect 222102 546618 257546 547174
rect 258102 546618 293546 547174
rect 294102 546618 329546 547174
rect 330102 546618 365546 547174
rect 366102 546618 401546 547174
rect 402102 546618 437546 547174
rect 438102 546618 473546 547174
rect 474102 546618 509546 547174
rect 510102 546618 545546 547174
rect 546102 546618 581546 547174
rect 582102 546618 587262 547174
rect 587818 546618 588810 547174
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 542898 -1974 543454
rect -1418 542898 1826 543454
rect 2382 542898 37826 543454
rect 38382 542898 73826 543454
rect 74382 542898 109826 543454
rect 110382 542898 145826 543454
rect 146382 542898 181826 543454
rect 182382 542898 217826 543454
rect 218382 542898 253826 543454
rect 254382 542898 289826 543454
rect 290382 542898 325826 543454
rect 326382 542898 361826 543454
rect 362382 542898 397826 543454
rect 398382 542898 433826 543454
rect 434382 542898 469826 543454
rect 470382 542898 505826 543454
rect 506382 542898 541826 543454
rect 542382 542898 577826 543454
rect 578382 542898 585342 543454
rect 585898 542898 586890 543454
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536058 -8694 536614
rect -8138 536058 30986 536614
rect 31542 536058 66986 536614
rect 67542 536058 102986 536614
rect 103542 536058 138986 536614
rect 139542 536058 174986 536614
rect 175542 536058 210986 536614
rect 211542 536058 246986 536614
rect 247542 536058 282986 536614
rect 283542 536058 318986 536614
rect 319542 536058 354986 536614
rect 355542 536058 390986 536614
rect 391542 536058 426986 536614
rect 427542 536058 462986 536614
rect 463542 536058 498986 536614
rect 499542 536058 534986 536614
rect 535542 536058 570986 536614
rect 571542 536058 592062 536614
rect 592618 536058 592650 536614
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532338 -6774 532894
rect -6218 532338 27266 532894
rect 27822 532338 63266 532894
rect 63822 532338 99266 532894
rect 99822 532338 135266 532894
rect 135822 532338 171266 532894
rect 171822 532338 207266 532894
rect 207822 532338 243266 532894
rect 243822 532338 279266 532894
rect 279822 532338 315266 532894
rect 315822 532338 351266 532894
rect 351822 532338 387266 532894
rect 387822 532338 423266 532894
rect 423822 532338 459266 532894
rect 459822 532338 495266 532894
rect 495822 532338 531266 532894
rect 531822 532338 567266 532894
rect 567822 532338 590142 532894
rect 590698 532338 590730 532894
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528618 -4854 529174
rect -4298 528618 23546 529174
rect 24102 528618 59546 529174
rect 60102 528618 95546 529174
rect 96102 528618 131546 529174
rect 132102 528618 167546 529174
rect 168102 528618 203546 529174
rect 204102 528618 239546 529174
rect 240102 528618 275546 529174
rect 276102 528618 311546 529174
rect 312102 528618 347546 529174
rect 348102 528618 383546 529174
rect 384102 528618 419546 529174
rect 420102 528618 455546 529174
rect 456102 528618 491546 529174
rect 492102 528618 527546 529174
rect 528102 528618 563546 529174
rect 564102 528618 588222 529174
rect 588778 528618 588810 529174
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 524898 -2934 525454
rect -2378 524898 19826 525454
rect 20382 524898 55826 525454
rect 56382 524898 91826 525454
rect 92382 524898 127826 525454
rect 128382 524898 163826 525454
rect 164382 524898 199826 525454
rect 200382 524898 235826 525454
rect 236382 524898 271826 525454
rect 272382 524898 307826 525454
rect 308382 524898 343826 525454
rect 344382 524898 379826 525454
rect 380382 524898 415826 525454
rect 416382 524898 451826 525454
rect 452382 524898 487826 525454
rect 488382 524898 523826 525454
rect 524382 524898 559826 525454
rect 560382 524898 586302 525454
rect 586858 524898 586890 525454
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518058 -7734 518614
rect -7178 518058 12986 518614
rect 13542 518058 48986 518614
rect 49542 518058 84986 518614
rect 85542 518058 120986 518614
rect 121542 518058 156986 518614
rect 157542 518058 192986 518614
rect 193542 518058 228986 518614
rect 229542 518058 264986 518614
rect 265542 518058 300986 518614
rect 301542 518058 336986 518614
rect 337542 518058 372986 518614
rect 373542 518058 408986 518614
rect 409542 518058 444986 518614
rect 445542 518058 480986 518614
rect 481542 518058 516986 518614
rect 517542 518058 552986 518614
rect 553542 518058 591102 518614
rect 591658 518058 592650 518614
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514338 -5814 514894
rect -5258 514338 9266 514894
rect 9822 514338 45266 514894
rect 45822 514338 81266 514894
rect 81822 514338 117266 514894
rect 117822 514338 153266 514894
rect 153822 514338 189266 514894
rect 189822 514338 225266 514894
rect 225822 514338 261266 514894
rect 261822 514338 297266 514894
rect 297822 514338 333266 514894
rect 333822 514338 369266 514894
rect 369822 514338 405266 514894
rect 405822 514338 441266 514894
rect 441822 514338 477266 514894
rect 477822 514338 513266 514894
rect 513822 514338 549266 514894
rect 549822 514338 589182 514894
rect 589738 514338 590730 514894
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510618 -3894 511174
rect -3338 510618 5546 511174
rect 6102 510618 41546 511174
rect 42102 510618 77546 511174
rect 78102 510618 113546 511174
rect 114102 510618 149546 511174
rect 150102 510618 185546 511174
rect 186102 510618 221546 511174
rect 222102 510618 257546 511174
rect 258102 510618 293546 511174
rect 294102 510618 329546 511174
rect 330102 510618 365546 511174
rect 366102 510618 401546 511174
rect 402102 510618 437546 511174
rect 438102 510618 473546 511174
rect 474102 510618 509546 511174
rect 510102 510618 545546 511174
rect 546102 510618 581546 511174
rect 582102 510618 587262 511174
rect 587818 510618 588810 511174
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 506898 -1974 507454
rect -1418 506898 1826 507454
rect 2382 506898 37826 507454
rect 38382 506898 73826 507454
rect 74382 506898 109826 507454
rect 110382 506898 145826 507454
rect 146382 506898 181826 507454
rect 182382 506898 217826 507454
rect 218382 506898 253826 507454
rect 254382 506898 289826 507454
rect 290382 506898 325826 507454
rect 326382 506898 361826 507454
rect 362382 506898 397826 507454
rect 398382 506898 433826 507454
rect 434382 506898 469826 507454
rect 470382 506898 505826 507454
rect 506382 506898 541826 507454
rect 542382 506898 577826 507454
rect 578382 506898 585342 507454
rect 585898 506898 586890 507454
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500058 -8694 500614
rect -8138 500058 30986 500614
rect 31542 500058 66986 500614
rect 67542 500058 102986 500614
rect 103542 500058 138986 500614
rect 139542 500058 174986 500614
rect 175542 500058 210986 500614
rect 211542 500058 246986 500614
rect 247542 500058 282986 500614
rect 283542 500058 318986 500614
rect 319542 500058 354986 500614
rect 355542 500058 390986 500614
rect 391542 500058 426986 500614
rect 427542 500058 462986 500614
rect 463542 500058 498986 500614
rect 499542 500058 534986 500614
rect 535542 500058 570986 500614
rect 571542 500058 592062 500614
rect 592618 500058 592650 500614
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496338 -6774 496894
rect -6218 496338 27266 496894
rect 27822 496338 63266 496894
rect 63822 496338 99266 496894
rect 99822 496338 135266 496894
rect 135822 496338 171266 496894
rect 171822 496338 207266 496894
rect 207822 496338 243266 496894
rect 243822 496338 279266 496894
rect 279822 496338 315266 496894
rect 315822 496338 351266 496894
rect 351822 496338 387266 496894
rect 387822 496338 423266 496894
rect 423822 496338 459266 496894
rect 459822 496338 495266 496894
rect 495822 496338 531266 496894
rect 531822 496338 567266 496894
rect 567822 496338 590142 496894
rect 590698 496338 590730 496894
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492618 -4854 493174
rect -4298 492618 23546 493174
rect 24102 492618 59546 493174
rect 60102 492618 95546 493174
rect 96102 492618 131546 493174
rect 132102 492618 167546 493174
rect 168102 492618 203546 493174
rect 204102 492618 239546 493174
rect 240102 492618 275546 493174
rect 276102 492618 311546 493174
rect 312102 492618 347546 493174
rect 348102 492618 383546 493174
rect 384102 492618 419546 493174
rect 420102 492618 455546 493174
rect 456102 492618 491546 493174
rect 492102 492618 527546 493174
rect 528102 492618 563546 493174
rect 564102 492618 588222 493174
rect 588778 492618 588810 493174
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 488898 -2934 489454
rect -2378 488898 19826 489454
rect 20382 488898 55826 489454
rect 56382 488898 91826 489454
rect 92382 488898 127826 489454
rect 128382 488898 163826 489454
rect 164382 488898 199826 489454
rect 200382 488898 235826 489454
rect 236382 488898 271826 489454
rect 272382 488898 307826 489454
rect 308382 488898 343826 489454
rect 344382 488898 379826 489454
rect 380382 488898 415826 489454
rect 416382 488898 451826 489454
rect 452382 488898 487826 489454
rect 488382 488898 523826 489454
rect 524382 488898 559826 489454
rect 560382 488898 586302 489454
rect 586858 488898 586890 489454
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482058 -7734 482614
rect -7178 482058 12986 482614
rect 13542 482058 48986 482614
rect 49542 482058 84986 482614
rect 85542 482058 120986 482614
rect 121542 482058 156986 482614
rect 157542 482058 192986 482614
rect 193542 482058 228986 482614
rect 229542 482058 264986 482614
rect 265542 482058 300986 482614
rect 301542 482058 336986 482614
rect 337542 482058 372986 482614
rect 373542 482058 408986 482614
rect 409542 482058 444986 482614
rect 445542 482058 480986 482614
rect 481542 482058 516986 482614
rect 517542 482058 552986 482614
rect 553542 482058 591102 482614
rect 591658 482058 592650 482614
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478338 -5814 478894
rect -5258 478338 9266 478894
rect 9822 478338 45266 478894
rect 45822 478338 81266 478894
rect 81822 478338 117266 478894
rect 117822 478338 153266 478894
rect 153822 478338 189266 478894
rect 189822 478338 225266 478894
rect 225822 478338 261266 478894
rect 261822 478338 297266 478894
rect 297822 478338 333266 478894
rect 333822 478338 369266 478894
rect 369822 478338 405266 478894
rect 405822 478338 441266 478894
rect 441822 478338 477266 478894
rect 477822 478338 513266 478894
rect 513822 478338 549266 478894
rect 549822 478338 589182 478894
rect 589738 478338 590730 478894
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474618 -3894 475174
rect -3338 474618 5546 475174
rect 6102 474618 41546 475174
rect 42102 474618 77546 475174
rect 78102 474618 113546 475174
rect 114102 474618 149546 475174
rect 150102 474618 185546 475174
rect 186102 474618 221546 475174
rect 222102 474618 257546 475174
rect 258102 474618 293546 475174
rect 294102 474618 329546 475174
rect 330102 474618 365546 475174
rect 366102 474618 401546 475174
rect 402102 474618 437546 475174
rect 438102 474618 473546 475174
rect 474102 474618 509546 475174
rect 510102 474618 545546 475174
rect 546102 474618 581546 475174
rect 582102 474618 587262 475174
rect 587818 474618 588810 475174
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 470898 -1974 471454
rect -1418 470898 1826 471454
rect 2382 470898 37826 471454
rect 38382 470898 73826 471454
rect 74382 470898 109826 471454
rect 110382 470898 145826 471454
rect 146382 470898 181826 471454
rect 182382 470898 217826 471454
rect 218382 470898 253826 471454
rect 254382 470898 289826 471454
rect 290382 470898 325826 471454
rect 326382 470898 361826 471454
rect 362382 470898 397826 471454
rect 398382 470898 433826 471454
rect 434382 470898 469826 471454
rect 470382 470898 505826 471454
rect 506382 470898 541826 471454
rect 542382 470898 577826 471454
rect 578382 470898 585342 471454
rect 585898 470898 586890 471454
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464058 -8694 464614
rect -8138 464058 30986 464614
rect 31542 464058 66986 464614
rect 67542 464058 102986 464614
rect 103542 464058 138986 464614
rect 139542 464058 174986 464614
rect 175542 464058 210986 464614
rect 211542 464058 246986 464614
rect 247542 464058 282986 464614
rect 283542 464058 318986 464614
rect 319542 464058 354986 464614
rect 355542 464058 390986 464614
rect 391542 464058 426986 464614
rect 427542 464058 462986 464614
rect 463542 464058 498986 464614
rect 499542 464058 534986 464614
rect 535542 464058 570986 464614
rect 571542 464058 592062 464614
rect 592618 464058 592650 464614
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460338 -6774 460894
rect -6218 460338 27266 460894
rect 27822 460338 63266 460894
rect 63822 460338 99266 460894
rect 99822 460338 135266 460894
rect 135822 460338 171266 460894
rect 171822 460338 207266 460894
rect 207822 460338 243266 460894
rect 243822 460338 279266 460894
rect 279822 460338 315266 460894
rect 315822 460338 351266 460894
rect 351822 460338 387266 460894
rect 387822 460338 423266 460894
rect 423822 460338 459266 460894
rect 459822 460338 495266 460894
rect 495822 460338 531266 460894
rect 531822 460338 567266 460894
rect 567822 460338 590142 460894
rect 590698 460338 590730 460894
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456618 -4854 457174
rect -4298 456618 23546 457174
rect 24102 456618 59546 457174
rect 60102 456618 95546 457174
rect 96102 456618 131546 457174
rect 132102 456618 167546 457174
rect 168102 456618 203546 457174
rect 204102 456618 419546 457174
rect 420102 456618 455546 457174
rect 456102 456618 491546 457174
rect 492102 456618 527546 457174
rect 528102 456618 563546 457174
rect 564102 456618 588222 457174
rect 588778 456618 588810 457174
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 452898 -2934 453454
rect -2378 452898 19826 453454
rect 20382 452898 55826 453454
rect 56382 452898 91826 453454
rect 92382 452898 127826 453454
rect 128382 452898 163826 453454
rect 164382 452898 199826 453454
rect 200382 453218 254610 453454
rect 254846 453218 285330 453454
rect 285566 453218 316050 453454
rect 316286 453218 346770 453454
rect 347006 453218 377490 453454
rect 377726 453218 408210 453454
rect 408446 453218 451826 453454
rect 200382 453134 451826 453218
rect 200382 452898 254610 453134
rect 254846 452898 285330 453134
rect 285566 452898 316050 453134
rect 316286 452898 346770 453134
rect 347006 452898 377490 453134
rect 377726 452898 408210 453134
rect 408446 452898 451826 453134
rect 452382 452898 487826 453454
rect 488382 452898 523826 453454
rect 524382 452898 559826 453454
rect 560382 452898 586302 453454
rect 586858 452898 586890 453454
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446058 -7734 446614
rect -7178 446058 12986 446614
rect 13542 446058 48986 446614
rect 49542 446058 84986 446614
rect 85542 446058 120986 446614
rect 121542 446058 156986 446614
rect 157542 446058 192986 446614
rect 193542 446058 228986 446614
rect 229542 446058 444986 446614
rect 445542 446058 480986 446614
rect 481542 446058 516986 446614
rect 517542 446058 552986 446614
rect 553542 446058 591102 446614
rect 591658 446058 592650 446614
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442338 -5814 442894
rect -5258 442338 9266 442894
rect 9822 442338 45266 442894
rect 45822 442338 81266 442894
rect 81822 442338 117266 442894
rect 117822 442338 153266 442894
rect 153822 442338 189266 442894
rect 189822 442338 225266 442894
rect 225822 442338 441266 442894
rect 441822 442338 477266 442894
rect 477822 442338 513266 442894
rect 513822 442338 549266 442894
rect 549822 442338 589182 442894
rect 589738 442338 590730 442894
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438618 -3894 439174
rect -3338 438618 5546 439174
rect 6102 438618 41546 439174
rect 42102 438618 77546 439174
rect 78102 438618 113546 439174
rect 114102 438618 149546 439174
rect 150102 438618 185546 439174
rect 186102 438618 221546 439174
rect 222102 438618 437546 439174
rect 438102 438618 473546 439174
rect 474102 438618 509546 439174
rect 510102 438618 545546 439174
rect 546102 438618 581546 439174
rect 582102 438618 587262 439174
rect 587818 438618 588810 439174
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 434898 -1974 435454
rect -1418 434898 1826 435454
rect 2382 434898 37826 435454
rect 38382 434898 73826 435454
rect 74382 434898 109826 435454
rect 110382 434898 145826 435454
rect 146382 434898 181826 435454
rect 182382 434898 217826 435454
rect 218382 435218 239250 435454
rect 239486 435218 269970 435454
rect 270206 435218 300690 435454
rect 300926 435218 331410 435454
rect 331646 435218 362130 435454
rect 362366 435218 392850 435454
rect 393086 435218 433826 435454
rect 218382 435134 433826 435218
rect 218382 434898 239250 435134
rect 239486 434898 269970 435134
rect 270206 434898 300690 435134
rect 300926 434898 331410 435134
rect 331646 434898 362130 435134
rect 362366 434898 392850 435134
rect 393086 434898 433826 435134
rect 434382 434898 469826 435454
rect 470382 434898 505826 435454
rect 506382 434898 541826 435454
rect 542382 434898 577826 435454
rect 578382 434898 585342 435454
rect 585898 434898 586890 435454
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428058 -8694 428614
rect -8138 428058 30986 428614
rect 31542 428058 66986 428614
rect 67542 428058 102986 428614
rect 103542 428058 138986 428614
rect 139542 428058 174986 428614
rect 175542 428058 210986 428614
rect 211542 428058 426986 428614
rect 427542 428058 462986 428614
rect 463542 428058 498986 428614
rect 499542 428058 534986 428614
rect 535542 428058 570986 428614
rect 571542 428058 592062 428614
rect 592618 428058 592650 428614
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424338 -6774 424894
rect -6218 424338 27266 424894
rect 27822 424338 63266 424894
rect 63822 424338 99266 424894
rect 99822 424338 135266 424894
rect 135822 424338 171266 424894
rect 171822 424338 207266 424894
rect 207822 424338 423266 424894
rect 423822 424338 459266 424894
rect 459822 424338 495266 424894
rect 495822 424338 531266 424894
rect 531822 424338 567266 424894
rect 567822 424338 590142 424894
rect 590698 424338 590730 424894
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420618 -4854 421174
rect -4298 420618 23546 421174
rect 24102 420618 59546 421174
rect 60102 420618 95546 421174
rect 96102 420618 131546 421174
rect 132102 420618 167546 421174
rect 168102 420618 203546 421174
rect 204102 420618 419546 421174
rect 420102 420618 455546 421174
rect 456102 420618 491546 421174
rect 492102 420618 527546 421174
rect 528102 420618 563546 421174
rect 564102 420618 588222 421174
rect 588778 420618 588810 421174
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 416898 -2934 417454
rect -2378 416898 19826 417454
rect 20382 416898 55826 417454
rect 56382 416898 91826 417454
rect 92382 416898 127826 417454
rect 128382 416898 163826 417454
rect 164382 416898 199826 417454
rect 200382 417218 254610 417454
rect 254846 417218 285330 417454
rect 285566 417218 316050 417454
rect 316286 417218 346770 417454
rect 347006 417218 377490 417454
rect 377726 417218 408210 417454
rect 408446 417218 451826 417454
rect 200382 417134 451826 417218
rect 200382 416898 254610 417134
rect 254846 416898 285330 417134
rect 285566 416898 316050 417134
rect 316286 416898 346770 417134
rect 347006 416898 377490 417134
rect 377726 416898 408210 417134
rect 408446 416898 451826 417134
rect 452382 416898 487826 417454
rect 488382 416898 523826 417454
rect 524382 416898 559826 417454
rect 560382 416898 586302 417454
rect 586858 416898 586890 417454
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410058 -7734 410614
rect -7178 410058 12986 410614
rect 13542 410058 48986 410614
rect 49542 410058 84986 410614
rect 85542 410058 120986 410614
rect 121542 410058 156986 410614
rect 157542 410058 192986 410614
rect 193542 410058 228986 410614
rect 229542 410058 444986 410614
rect 445542 410058 480986 410614
rect 481542 410058 516986 410614
rect 517542 410058 552986 410614
rect 553542 410058 591102 410614
rect 591658 410058 592650 410614
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406338 -5814 406894
rect -5258 406338 9266 406894
rect 9822 406338 45266 406894
rect 45822 406338 81266 406894
rect 81822 406338 117266 406894
rect 117822 406338 153266 406894
rect 153822 406338 189266 406894
rect 189822 406338 225266 406894
rect 225822 406338 441266 406894
rect 441822 406338 477266 406894
rect 477822 406338 513266 406894
rect 513822 406338 549266 406894
rect 549822 406338 589182 406894
rect 589738 406338 590730 406894
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402618 -3894 403174
rect -3338 402618 5546 403174
rect 6102 402618 41546 403174
rect 42102 402618 77546 403174
rect 78102 402618 113546 403174
rect 114102 402618 149546 403174
rect 150102 402618 185546 403174
rect 186102 402618 221546 403174
rect 222102 402618 437546 403174
rect 438102 402618 473546 403174
rect 474102 402618 509546 403174
rect 510102 402618 545546 403174
rect 546102 402618 581546 403174
rect 582102 402618 587262 403174
rect 587818 402618 588810 403174
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 398898 -1974 399454
rect -1418 398898 1826 399454
rect 2382 398898 37826 399454
rect 38382 398898 73826 399454
rect 74382 398898 109826 399454
rect 110382 398898 145826 399454
rect 146382 398898 181826 399454
rect 182382 398898 217826 399454
rect 218382 399218 239250 399454
rect 239486 399218 269970 399454
rect 270206 399218 300690 399454
rect 300926 399218 331410 399454
rect 331646 399218 362130 399454
rect 362366 399218 392850 399454
rect 393086 399218 433826 399454
rect 218382 399134 433826 399218
rect 218382 398898 239250 399134
rect 239486 398898 269970 399134
rect 270206 398898 300690 399134
rect 300926 398898 331410 399134
rect 331646 398898 362130 399134
rect 362366 398898 392850 399134
rect 393086 398898 433826 399134
rect 434382 398898 469826 399454
rect 470382 398898 505826 399454
rect 506382 398898 541826 399454
rect 542382 398898 577826 399454
rect 578382 398898 585342 399454
rect 585898 398898 586890 399454
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392058 -8694 392614
rect -8138 392058 30986 392614
rect 31542 392058 66986 392614
rect 67542 392058 102986 392614
rect 103542 392058 138986 392614
rect 139542 392058 174986 392614
rect 175542 392058 210986 392614
rect 211542 392058 426986 392614
rect 427542 392058 462986 392614
rect 463542 392058 498986 392614
rect 499542 392058 534986 392614
rect 535542 392058 570986 392614
rect 571542 392058 592062 392614
rect 592618 392058 592650 392614
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388338 -6774 388894
rect -6218 388338 27266 388894
rect 27822 388338 63266 388894
rect 63822 388338 99266 388894
rect 99822 388338 135266 388894
rect 135822 388338 171266 388894
rect 171822 388338 207266 388894
rect 207822 388338 423266 388894
rect 423822 388338 459266 388894
rect 459822 388338 495266 388894
rect 495822 388338 531266 388894
rect 531822 388338 567266 388894
rect 567822 388338 590142 388894
rect 590698 388338 590730 388894
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384618 -4854 385174
rect -4298 384618 23546 385174
rect 24102 384618 59546 385174
rect 60102 384618 95546 385174
rect 96102 384618 131546 385174
rect 132102 384618 167546 385174
rect 168102 384618 203546 385174
rect 204102 384618 419546 385174
rect 420102 384618 455546 385174
rect 456102 384618 491546 385174
rect 492102 384618 527546 385174
rect 528102 384618 563546 385174
rect 564102 384618 588222 385174
rect 588778 384618 588810 385174
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 380898 -2934 381454
rect -2378 380898 19826 381454
rect 20382 380898 55826 381454
rect 56382 380898 91826 381454
rect 92382 380898 127826 381454
rect 128382 380898 163826 381454
rect 164382 380898 199826 381454
rect 200382 381218 254610 381454
rect 254846 381218 285330 381454
rect 285566 381218 316050 381454
rect 316286 381218 346770 381454
rect 347006 381218 377490 381454
rect 377726 381218 408210 381454
rect 408446 381218 451826 381454
rect 200382 381134 451826 381218
rect 200382 380898 254610 381134
rect 254846 380898 285330 381134
rect 285566 380898 316050 381134
rect 316286 380898 346770 381134
rect 347006 380898 377490 381134
rect 377726 380898 408210 381134
rect 408446 380898 451826 381134
rect 452382 380898 487826 381454
rect 488382 380898 523826 381454
rect 524382 380898 559826 381454
rect 560382 380898 586302 381454
rect 586858 380898 586890 381454
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374058 -7734 374614
rect -7178 374058 12986 374614
rect 13542 374058 48986 374614
rect 49542 374058 84986 374614
rect 85542 374058 120986 374614
rect 121542 374058 156986 374614
rect 157542 374058 192986 374614
rect 193542 374058 228986 374614
rect 229542 374058 444986 374614
rect 445542 374058 480986 374614
rect 481542 374058 516986 374614
rect 517542 374058 552986 374614
rect 553542 374058 591102 374614
rect 591658 374058 592650 374614
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370338 -5814 370894
rect -5258 370338 9266 370894
rect 9822 370338 45266 370894
rect 45822 370338 81266 370894
rect 81822 370338 117266 370894
rect 117822 370338 153266 370894
rect 153822 370338 189266 370894
rect 189822 370338 225266 370894
rect 225822 370338 441266 370894
rect 441822 370338 477266 370894
rect 477822 370338 513266 370894
rect 513822 370338 549266 370894
rect 549822 370338 589182 370894
rect 589738 370338 590730 370894
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366618 -3894 367174
rect -3338 366618 5546 367174
rect 6102 366618 41546 367174
rect 42102 366618 77546 367174
rect 78102 366618 113546 367174
rect 114102 366618 149546 367174
rect 150102 366618 185546 367174
rect 186102 366618 221546 367174
rect 222102 366618 437546 367174
rect 438102 366618 473546 367174
rect 474102 366618 509546 367174
rect 510102 366618 545546 367174
rect 546102 366618 581546 367174
rect 582102 366618 587262 367174
rect 587818 366618 588810 367174
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 362898 -1974 363454
rect -1418 362898 1826 363454
rect 2382 362898 37826 363454
rect 38382 362898 73826 363454
rect 74382 362898 109826 363454
rect 110382 362898 145826 363454
rect 146382 362898 181826 363454
rect 182382 362898 217826 363454
rect 218382 363218 239250 363454
rect 239486 363218 269970 363454
rect 270206 363218 300690 363454
rect 300926 363218 331410 363454
rect 331646 363218 362130 363454
rect 362366 363218 392850 363454
rect 393086 363218 433826 363454
rect 218382 363134 433826 363218
rect 218382 362898 239250 363134
rect 239486 362898 269970 363134
rect 270206 362898 300690 363134
rect 300926 362898 331410 363134
rect 331646 362898 362130 363134
rect 362366 362898 392850 363134
rect 393086 362898 433826 363134
rect 434382 362898 469826 363454
rect 470382 362898 505826 363454
rect 506382 362898 541826 363454
rect 542382 362898 577826 363454
rect 578382 362898 585342 363454
rect 585898 362898 586890 363454
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356058 -8694 356614
rect -8138 356058 30986 356614
rect 31542 356058 66986 356614
rect 67542 356058 102986 356614
rect 103542 356058 138986 356614
rect 139542 356058 174986 356614
rect 175542 356058 210986 356614
rect 211542 356058 426986 356614
rect 427542 356058 462986 356614
rect 463542 356058 498986 356614
rect 499542 356058 534986 356614
rect 535542 356058 570986 356614
rect 571542 356058 592062 356614
rect 592618 356058 592650 356614
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352338 -6774 352894
rect -6218 352338 27266 352894
rect 27822 352338 63266 352894
rect 63822 352338 99266 352894
rect 99822 352338 135266 352894
rect 135822 352338 171266 352894
rect 171822 352338 207266 352894
rect 207822 352338 423266 352894
rect 423822 352338 459266 352894
rect 459822 352338 495266 352894
rect 495822 352338 531266 352894
rect 531822 352338 567266 352894
rect 567822 352338 590142 352894
rect 590698 352338 590730 352894
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348618 -4854 349174
rect -4298 348618 23546 349174
rect 24102 348618 59546 349174
rect 60102 348618 95546 349174
rect 96102 348618 131546 349174
rect 132102 348618 167546 349174
rect 168102 348618 203546 349174
rect 204102 348618 419546 349174
rect 420102 348618 455546 349174
rect 456102 348618 491546 349174
rect 492102 348618 527546 349174
rect 528102 348618 563546 349174
rect 564102 348618 588222 349174
rect 588778 348618 588810 349174
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 344898 -2934 345454
rect -2378 344898 19826 345454
rect 20382 344898 55826 345454
rect 56382 344898 91826 345454
rect 92382 344898 127826 345454
rect 128382 344898 163826 345454
rect 164382 344898 199826 345454
rect 200382 345218 254610 345454
rect 254846 345218 285330 345454
rect 285566 345218 316050 345454
rect 316286 345218 346770 345454
rect 347006 345218 377490 345454
rect 377726 345218 408210 345454
rect 408446 345218 451826 345454
rect 200382 345134 451826 345218
rect 200382 344898 254610 345134
rect 254846 344898 285330 345134
rect 285566 344898 316050 345134
rect 316286 344898 346770 345134
rect 347006 344898 377490 345134
rect 377726 344898 408210 345134
rect 408446 344898 451826 345134
rect 452382 344898 487826 345454
rect 488382 344898 523826 345454
rect 524382 344898 559826 345454
rect 560382 344898 586302 345454
rect 586858 344898 586890 345454
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338058 -7734 338614
rect -7178 338058 12986 338614
rect 13542 338058 48986 338614
rect 49542 338058 84986 338614
rect 85542 338058 120986 338614
rect 121542 338058 156986 338614
rect 157542 338058 192986 338614
rect 193542 338058 228986 338614
rect 229542 338058 444986 338614
rect 445542 338058 480986 338614
rect 481542 338058 516986 338614
rect 517542 338058 552986 338614
rect 553542 338058 591102 338614
rect 591658 338058 592650 338614
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334338 -5814 334894
rect -5258 334338 9266 334894
rect 9822 334338 45266 334894
rect 45822 334338 81266 334894
rect 81822 334338 117266 334894
rect 117822 334338 153266 334894
rect 153822 334338 189266 334894
rect 189822 334338 225266 334894
rect 225822 334338 261266 334894
rect 261822 334338 297266 334894
rect 297822 334338 333266 334894
rect 333822 334338 369266 334894
rect 369822 334338 405266 334894
rect 405822 334338 441266 334894
rect 441822 334338 477266 334894
rect 477822 334338 513266 334894
rect 513822 334338 549266 334894
rect 549822 334338 589182 334894
rect 589738 334338 590730 334894
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330618 -3894 331174
rect -3338 330618 5546 331174
rect 6102 330618 41546 331174
rect 42102 330618 77546 331174
rect 78102 330618 113546 331174
rect 114102 330618 149546 331174
rect 150102 330618 185546 331174
rect 186102 330618 221546 331174
rect 222102 330618 257546 331174
rect 258102 330618 293546 331174
rect 294102 330618 329546 331174
rect 330102 330618 365546 331174
rect 366102 330618 401546 331174
rect 402102 330618 437546 331174
rect 438102 330618 473546 331174
rect 474102 330618 509546 331174
rect 510102 330618 545546 331174
rect 546102 330618 581546 331174
rect 582102 330618 587262 331174
rect 587818 330618 588810 331174
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 326898 -1974 327454
rect -1418 326898 1826 327454
rect 2382 326898 37826 327454
rect 38382 326898 73826 327454
rect 74382 326898 109826 327454
rect 110382 326898 145826 327454
rect 146382 326898 181826 327454
rect 182382 326898 217826 327454
rect 218382 326898 253826 327454
rect 254382 326898 289826 327454
rect 290382 326898 325826 327454
rect 326382 326898 361826 327454
rect 362382 326898 397826 327454
rect 398382 326898 433826 327454
rect 434382 326898 469826 327454
rect 470382 326898 505826 327454
rect 506382 326898 541826 327454
rect 542382 326898 577826 327454
rect 578382 326898 585342 327454
rect 585898 326898 586890 327454
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320058 -8694 320614
rect -8138 320058 30986 320614
rect 31542 320058 66986 320614
rect 67542 320058 102986 320614
rect 103542 320058 138986 320614
rect 139542 320058 174986 320614
rect 175542 320058 210986 320614
rect 211542 320058 246986 320614
rect 247542 320058 282986 320614
rect 283542 320058 318986 320614
rect 319542 320058 354986 320614
rect 355542 320058 390986 320614
rect 391542 320058 426986 320614
rect 427542 320058 462986 320614
rect 463542 320058 498986 320614
rect 499542 320058 534986 320614
rect 535542 320058 570986 320614
rect 571542 320058 592062 320614
rect 592618 320058 592650 320614
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316338 -6774 316894
rect -6218 316338 27266 316894
rect 27822 316338 63266 316894
rect 63822 316338 99266 316894
rect 99822 316338 135266 316894
rect 135822 316338 171266 316894
rect 171822 316338 207266 316894
rect 207822 316338 243266 316894
rect 243822 316338 279266 316894
rect 279822 316338 315266 316894
rect 315822 316338 351266 316894
rect 351822 316338 387266 316894
rect 387822 316338 423266 316894
rect 423822 316338 459266 316894
rect 459822 316338 495266 316894
rect 495822 316338 531266 316894
rect 531822 316338 567266 316894
rect 567822 316338 590142 316894
rect 590698 316338 590730 316894
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312618 -4854 313174
rect -4298 312618 23546 313174
rect 24102 312618 59546 313174
rect 60102 312618 95546 313174
rect 96102 312618 131546 313174
rect 132102 312618 167546 313174
rect 168102 312618 203546 313174
rect 204102 312618 239546 313174
rect 240102 312618 275546 313174
rect 276102 312618 311546 313174
rect 312102 312618 347546 313174
rect 348102 312618 383546 313174
rect 384102 312618 419546 313174
rect 420102 312618 455546 313174
rect 456102 312618 491546 313174
rect 492102 312618 527546 313174
rect 528102 312618 563546 313174
rect 564102 312618 588222 313174
rect 588778 312618 588810 313174
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 308898 -2934 309454
rect -2378 308898 19826 309454
rect 20382 308898 55826 309454
rect 56382 308898 91826 309454
rect 92382 308898 127826 309454
rect 128382 308898 163826 309454
rect 164382 308898 199826 309454
rect 200382 308898 235826 309454
rect 236382 308898 271826 309454
rect 272382 308898 307826 309454
rect 308382 308898 343826 309454
rect 344382 308898 379826 309454
rect 380382 308898 415826 309454
rect 416382 308898 451826 309454
rect 452382 308898 487826 309454
rect 488382 308898 523826 309454
rect 524382 308898 559826 309454
rect 560382 308898 586302 309454
rect 586858 308898 586890 309454
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302058 -7734 302614
rect -7178 302058 12986 302614
rect 13542 302058 48986 302614
rect 49542 302058 84986 302614
rect 85542 302058 120986 302614
rect 121542 302058 156986 302614
rect 157542 302058 192986 302614
rect 193542 302058 228986 302614
rect 229542 302058 264986 302614
rect 265542 302058 300986 302614
rect 301542 302058 336986 302614
rect 337542 302058 372986 302614
rect 373542 302058 408986 302614
rect 409542 302058 444986 302614
rect 445542 302058 480986 302614
rect 481542 302058 516986 302614
rect 517542 302058 552986 302614
rect 553542 302058 591102 302614
rect 591658 302058 592650 302614
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298338 -5814 298894
rect -5258 298338 9266 298894
rect 9822 298338 45266 298894
rect 45822 298338 81266 298894
rect 81822 298338 117266 298894
rect 117822 298338 153266 298894
rect 153822 298338 189266 298894
rect 189822 298338 225266 298894
rect 225822 298338 261266 298894
rect 261822 298338 297266 298894
rect 297822 298338 333266 298894
rect 333822 298338 369266 298894
rect 369822 298338 405266 298894
rect 405822 298338 441266 298894
rect 441822 298338 477266 298894
rect 477822 298338 513266 298894
rect 513822 298338 549266 298894
rect 549822 298338 589182 298894
rect 589738 298338 590730 298894
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294618 -3894 295174
rect -3338 294618 5546 295174
rect 6102 294618 41546 295174
rect 42102 294618 77546 295174
rect 78102 294618 113546 295174
rect 114102 294618 149546 295174
rect 150102 294618 185546 295174
rect 186102 294618 221546 295174
rect 222102 294618 257546 295174
rect 258102 294618 293546 295174
rect 294102 294618 329546 295174
rect 330102 294618 365546 295174
rect 366102 294618 401546 295174
rect 402102 294618 437546 295174
rect 438102 294618 473546 295174
rect 474102 294618 509546 295174
rect 510102 294618 545546 295174
rect 546102 294618 581546 295174
rect 582102 294618 587262 295174
rect 587818 294618 588810 295174
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 290898 -1974 291454
rect -1418 290898 1826 291454
rect 2382 290898 37826 291454
rect 38382 290898 73826 291454
rect 74382 290898 109826 291454
rect 110382 290898 145826 291454
rect 146382 290898 181826 291454
rect 182382 290898 217826 291454
rect 218382 290898 253826 291454
rect 254382 290898 289826 291454
rect 290382 290898 325826 291454
rect 326382 290898 361826 291454
rect 362382 290898 397826 291454
rect 398382 290898 433826 291454
rect 434382 290898 469826 291454
rect 470382 290898 505826 291454
rect 506382 290898 541826 291454
rect 542382 290898 577826 291454
rect 578382 290898 585342 291454
rect 585898 290898 586890 291454
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284058 -8694 284614
rect -8138 284058 30986 284614
rect 31542 284058 66986 284614
rect 67542 284058 102986 284614
rect 103542 284058 138986 284614
rect 139542 284058 174986 284614
rect 175542 284058 210986 284614
rect 211542 284058 246986 284614
rect 247542 284058 282986 284614
rect 283542 284058 318986 284614
rect 319542 284058 354986 284614
rect 355542 284058 390986 284614
rect 391542 284058 426986 284614
rect 427542 284058 462986 284614
rect 463542 284058 498986 284614
rect 499542 284058 534986 284614
rect 535542 284058 570986 284614
rect 571542 284058 592062 284614
rect 592618 284058 592650 284614
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280338 -6774 280894
rect -6218 280338 27266 280894
rect 27822 280338 63266 280894
rect 63822 280338 99266 280894
rect 99822 280338 135266 280894
rect 135822 280338 171266 280894
rect 171822 280338 207266 280894
rect 207822 280338 243266 280894
rect 243822 280338 279266 280894
rect 279822 280338 315266 280894
rect 315822 280338 351266 280894
rect 351822 280338 387266 280894
rect 387822 280338 423266 280894
rect 423822 280338 459266 280894
rect 459822 280338 495266 280894
rect 495822 280338 531266 280894
rect 531822 280338 567266 280894
rect 567822 280338 590142 280894
rect 590698 280338 590730 280894
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276618 -4854 277174
rect -4298 276618 23546 277174
rect 24102 276618 59546 277174
rect 60102 276618 95546 277174
rect 96102 276618 131546 277174
rect 132102 276618 167546 277174
rect 168102 276618 203546 277174
rect 204102 276618 239546 277174
rect 240102 276618 275546 277174
rect 276102 276618 311546 277174
rect 312102 276618 347546 277174
rect 348102 276618 383546 277174
rect 384102 276618 419546 277174
rect 420102 276618 455546 277174
rect 456102 276618 491546 277174
rect 492102 276618 527546 277174
rect 528102 276618 563546 277174
rect 564102 276618 588222 277174
rect 588778 276618 588810 277174
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 272898 -2934 273454
rect -2378 272898 19826 273454
rect 20382 272898 55826 273454
rect 56382 272898 91826 273454
rect 92382 272898 127826 273454
rect 128382 272898 163826 273454
rect 164382 272898 199826 273454
rect 200382 272898 235826 273454
rect 236382 272898 271826 273454
rect 272382 272898 307826 273454
rect 308382 272898 343826 273454
rect 344382 272898 379826 273454
rect 380382 272898 415826 273454
rect 416382 272898 451826 273454
rect 452382 272898 487826 273454
rect 488382 272898 523826 273454
rect 524382 272898 559826 273454
rect 560382 272898 586302 273454
rect 586858 272898 586890 273454
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266058 -7734 266614
rect -7178 266058 12986 266614
rect 13542 266058 48986 266614
rect 49542 266058 84986 266614
rect 85542 266058 120986 266614
rect 121542 266058 156986 266614
rect 157542 266058 192986 266614
rect 193542 266058 228986 266614
rect 229542 266058 264986 266614
rect 265542 266058 300986 266614
rect 301542 266058 336986 266614
rect 337542 266058 372986 266614
rect 373542 266058 408986 266614
rect 409542 266058 444986 266614
rect 445542 266058 480986 266614
rect 481542 266058 516986 266614
rect 517542 266058 552986 266614
rect 553542 266058 591102 266614
rect 591658 266058 592650 266614
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262338 -5814 262894
rect -5258 262338 9266 262894
rect 9822 262338 45266 262894
rect 45822 262338 81266 262894
rect 81822 262338 117266 262894
rect 117822 262338 153266 262894
rect 153822 262338 189266 262894
rect 189822 262338 225266 262894
rect 225822 262338 261266 262894
rect 261822 262338 297266 262894
rect 297822 262338 333266 262894
rect 333822 262338 369266 262894
rect 369822 262338 405266 262894
rect 405822 262338 441266 262894
rect 441822 262338 477266 262894
rect 477822 262338 513266 262894
rect 513822 262338 549266 262894
rect 549822 262338 589182 262894
rect 589738 262338 590730 262894
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258618 -3894 259174
rect -3338 258618 5546 259174
rect 6102 258618 41546 259174
rect 42102 258618 77546 259174
rect 78102 258618 113546 259174
rect 114102 258618 149546 259174
rect 150102 258618 185546 259174
rect 186102 258618 221546 259174
rect 222102 258618 257546 259174
rect 258102 258618 293546 259174
rect 294102 258618 329546 259174
rect 330102 258618 365546 259174
rect 366102 258618 401546 259174
rect 402102 258618 437546 259174
rect 438102 258618 473546 259174
rect 474102 258618 509546 259174
rect 510102 258618 545546 259174
rect 546102 258618 581546 259174
rect 582102 258618 587262 259174
rect 587818 258618 588810 259174
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 254898 -1974 255454
rect -1418 254898 1826 255454
rect 2382 254898 37826 255454
rect 38382 254898 73826 255454
rect 74382 254898 109826 255454
rect 110382 254898 145826 255454
rect 146382 254898 181826 255454
rect 182382 254898 217826 255454
rect 218382 254898 253826 255454
rect 254382 254898 289826 255454
rect 290382 254898 325826 255454
rect 326382 254898 361826 255454
rect 362382 254898 397826 255454
rect 398382 254898 433826 255454
rect 434382 254898 469826 255454
rect 470382 254898 505826 255454
rect 506382 254898 541826 255454
rect 542382 254898 577826 255454
rect 578382 254898 585342 255454
rect 585898 254898 586890 255454
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248058 -8694 248614
rect -8138 248058 30986 248614
rect 31542 248058 66986 248614
rect 67542 248058 102986 248614
rect 103542 248058 138986 248614
rect 139542 248058 174986 248614
rect 175542 248058 210986 248614
rect 211542 248058 246986 248614
rect 247542 248058 282986 248614
rect 283542 248058 318986 248614
rect 319542 248058 354986 248614
rect 355542 248058 390986 248614
rect 391542 248058 426986 248614
rect 427542 248058 462986 248614
rect 463542 248058 498986 248614
rect 499542 248058 534986 248614
rect 535542 248058 570986 248614
rect 571542 248058 592062 248614
rect 592618 248058 592650 248614
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244338 -6774 244894
rect -6218 244338 27266 244894
rect 27822 244338 63266 244894
rect 63822 244338 99266 244894
rect 99822 244338 135266 244894
rect 135822 244338 171266 244894
rect 171822 244338 207266 244894
rect 207822 244338 243266 244894
rect 243822 244338 279266 244894
rect 279822 244338 315266 244894
rect 315822 244338 351266 244894
rect 351822 244338 387266 244894
rect 387822 244338 423266 244894
rect 423822 244338 459266 244894
rect 459822 244338 495266 244894
rect 495822 244338 531266 244894
rect 531822 244338 567266 244894
rect 567822 244338 590142 244894
rect 590698 244338 590730 244894
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240618 -4854 241174
rect -4298 240618 23546 241174
rect 24102 240618 59546 241174
rect 60102 240618 95546 241174
rect 96102 240618 131546 241174
rect 132102 240618 167546 241174
rect 168102 240618 203546 241174
rect 204102 240618 239546 241174
rect 240102 240618 275546 241174
rect 276102 240618 311546 241174
rect 312102 240618 347546 241174
rect 348102 240618 383546 241174
rect 384102 240618 419546 241174
rect 420102 240618 455546 241174
rect 456102 240618 491546 241174
rect 492102 240618 527546 241174
rect 528102 240618 563546 241174
rect 564102 240618 588222 241174
rect 588778 240618 588810 241174
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 236898 -2934 237454
rect -2378 236898 19826 237454
rect 20382 236898 55826 237454
rect 56382 236898 91826 237454
rect 92382 236898 127826 237454
rect 128382 236898 163826 237454
rect 164382 236898 199826 237454
rect 200382 236898 235826 237454
rect 236382 236898 271826 237454
rect 272382 236898 307826 237454
rect 308382 236898 343826 237454
rect 344382 236898 379826 237454
rect 380382 236898 415826 237454
rect 416382 236898 451826 237454
rect 452382 236898 487826 237454
rect 488382 236898 523826 237454
rect 524382 236898 559826 237454
rect 560382 236898 586302 237454
rect 586858 236898 586890 237454
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230058 -7734 230614
rect -7178 230058 12986 230614
rect 13542 230058 48986 230614
rect 49542 230058 84986 230614
rect 85542 230058 120986 230614
rect 121542 230058 156986 230614
rect 157542 230058 192986 230614
rect 193542 230058 228986 230614
rect 229542 230058 264986 230614
rect 265542 230058 300986 230614
rect 301542 230058 336986 230614
rect 337542 230058 372986 230614
rect 373542 230058 408986 230614
rect 409542 230058 444986 230614
rect 445542 230058 480986 230614
rect 481542 230058 516986 230614
rect 517542 230058 552986 230614
rect 553542 230058 591102 230614
rect 591658 230058 592650 230614
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226338 -5814 226894
rect -5258 226338 9266 226894
rect 9822 226338 45266 226894
rect 45822 226338 81266 226894
rect 81822 226338 117266 226894
rect 117822 226338 153266 226894
rect 153822 226338 189266 226894
rect 189822 226338 225266 226894
rect 225822 226338 261266 226894
rect 261822 226338 297266 226894
rect 297822 226338 333266 226894
rect 333822 226338 369266 226894
rect 369822 226338 405266 226894
rect 405822 226338 441266 226894
rect 441822 226338 477266 226894
rect 477822 226338 513266 226894
rect 513822 226338 549266 226894
rect 549822 226338 589182 226894
rect 589738 226338 590730 226894
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222618 -3894 223174
rect -3338 222618 5546 223174
rect 6102 222618 41546 223174
rect 42102 222618 77546 223174
rect 78102 222618 113546 223174
rect 114102 222618 149546 223174
rect 150102 222618 185546 223174
rect 186102 222618 221546 223174
rect 222102 222618 257546 223174
rect 258102 222618 293546 223174
rect 294102 222618 329546 223174
rect 330102 222618 365546 223174
rect 366102 222618 401546 223174
rect 402102 222618 437546 223174
rect 438102 222618 473546 223174
rect 474102 222618 509546 223174
rect 510102 222618 545546 223174
rect 546102 222618 581546 223174
rect 582102 222618 587262 223174
rect 587818 222618 588810 223174
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 218898 -1974 219454
rect -1418 218898 1826 219454
rect 2382 218898 37826 219454
rect 38382 218898 73826 219454
rect 74382 218898 109826 219454
rect 110382 218898 145826 219454
rect 146382 218898 181826 219454
rect 182382 218898 217826 219454
rect 218382 218898 253826 219454
rect 254382 218898 289826 219454
rect 290382 218898 325826 219454
rect 326382 218898 361826 219454
rect 362382 218898 397826 219454
rect 398382 218898 433826 219454
rect 434382 218898 469826 219454
rect 470382 218898 505826 219454
rect 506382 218898 541826 219454
rect 542382 218898 577826 219454
rect 578382 218898 585342 219454
rect 585898 218898 586890 219454
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212058 -8694 212614
rect -8138 212058 30986 212614
rect 31542 212058 66986 212614
rect 67542 212058 102986 212614
rect 103542 212058 138986 212614
rect 139542 212058 174986 212614
rect 175542 212058 210986 212614
rect 211542 212058 246986 212614
rect 247542 212058 282986 212614
rect 283542 212058 318986 212614
rect 319542 212058 354986 212614
rect 355542 212058 390986 212614
rect 391542 212058 426986 212614
rect 427542 212058 462986 212614
rect 463542 212058 498986 212614
rect 499542 212058 534986 212614
rect 535542 212058 570986 212614
rect 571542 212058 592062 212614
rect 592618 212058 592650 212614
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208338 -6774 208894
rect -6218 208338 27266 208894
rect 27822 208338 63266 208894
rect 63822 208338 99266 208894
rect 99822 208338 135266 208894
rect 135822 208338 171266 208894
rect 171822 208338 207266 208894
rect 207822 208338 243266 208894
rect 243822 208338 279266 208894
rect 279822 208338 315266 208894
rect 315822 208338 351266 208894
rect 351822 208338 387266 208894
rect 387822 208338 423266 208894
rect 423822 208338 459266 208894
rect 459822 208338 495266 208894
rect 495822 208338 531266 208894
rect 531822 208338 567266 208894
rect 567822 208338 590142 208894
rect 590698 208338 590730 208894
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204618 -4854 205174
rect -4298 204618 23546 205174
rect 24102 204618 59546 205174
rect 60102 204618 95546 205174
rect 96102 204618 131546 205174
rect 132102 204618 167546 205174
rect 168102 204618 203546 205174
rect 204102 204618 239546 205174
rect 240102 204618 275546 205174
rect 276102 204618 311546 205174
rect 312102 204618 347546 205174
rect 348102 204618 383546 205174
rect 384102 204618 419546 205174
rect 420102 204618 455546 205174
rect 456102 204618 491546 205174
rect 492102 204618 527546 205174
rect 528102 204618 563546 205174
rect 564102 204618 588222 205174
rect 588778 204618 588810 205174
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 200898 -2934 201454
rect -2378 200898 19826 201454
rect 20382 200898 55826 201454
rect 56382 200898 91826 201454
rect 92382 200898 127826 201454
rect 128382 200898 163826 201454
rect 164382 200898 199826 201454
rect 200382 200898 235826 201454
rect 236382 200898 271826 201454
rect 272382 200898 307826 201454
rect 308382 200898 343826 201454
rect 344382 200898 379826 201454
rect 380382 200898 415826 201454
rect 416382 200898 451826 201454
rect 452382 200898 487826 201454
rect 488382 200898 523826 201454
rect 524382 200898 559826 201454
rect 560382 200898 586302 201454
rect 586858 200898 586890 201454
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194058 -7734 194614
rect -7178 194058 12986 194614
rect 13542 194058 48986 194614
rect 49542 194058 84986 194614
rect 85542 194058 120986 194614
rect 121542 194058 156986 194614
rect 157542 194058 192986 194614
rect 193542 194058 228986 194614
rect 229542 194058 264986 194614
rect 265542 194058 300986 194614
rect 301542 194058 336986 194614
rect 337542 194058 372986 194614
rect 373542 194058 408986 194614
rect 409542 194058 444986 194614
rect 445542 194058 480986 194614
rect 481542 194058 516986 194614
rect 517542 194058 552986 194614
rect 553542 194058 591102 194614
rect 591658 194058 592650 194614
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190338 -5814 190894
rect -5258 190338 9266 190894
rect 9822 190338 45266 190894
rect 45822 190338 81266 190894
rect 81822 190338 117266 190894
rect 117822 190338 153266 190894
rect 153822 190338 189266 190894
rect 189822 190338 225266 190894
rect 225822 190338 261266 190894
rect 261822 190338 297266 190894
rect 297822 190338 333266 190894
rect 333822 190338 369266 190894
rect 369822 190338 405266 190894
rect 405822 190338 441266 190894
rect 441822 190338 477266 190894
rect 477822 190338 513266 190894
rect 513822 190338 549266 190894
rect 549822 190338 589182 190894
rect 589738 190338 590730 190894
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186618 -3894 187174
rect -3338 186618 5546 187174
rect 6102 186618 41546 187174
rect 42102 186618 77546 187174
rect 78102 186618 113546 187174
rect 114102 186618 149546 187174
rect 150102 186618 185546 187174
rect 186102 186618 221546 187174
rect 222102 186618 257546 187174
rect 258102 186618 293546 187174
rect 294102 186618 329546 187174
rect 330102 186618 365546 187174
rect 366102 186618 401546 187174
rect 402102 186618 437546 187174
rect 438102 186618 473546 187174
rect 474102 186618 509546 187174
rect 510102 186618 545546 187174
rect 546102 186618 581546 187174
rect 582102 186618 587262 187174
rect 587818 186618 588810 187174
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 182898 -1974 183454
rect -1418 182898 1826 183454
rect 2382 182898 37826 183454
rect 38382 182898 73826 183454
rect 74382 182898 109826 183454
rect 110382 182898 145826 183454
rect 146382 182898 181826 183454
rect 182382 182898 217826 183454
rect 218382 182898 253826 183454
rect 254382 182898 289826 183454
rect 290382 182898 325826 183454
rect 326382 182898 361826 183454
rect 362382 182898 397826 183454
rect 398382 182898 433826 183454
rect 434382 182898 469826 183454
rect 470382 182898 505826 183454
rect 506382 182898 541826 183454
rect 542382 182898 577826 183454
rect 578382 182898 585342 183454
rect 585898 182898 586890 183454
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176058 -8694 176614
rect -8138 176058 30986 176614
rect 31542 176058 66986 176614
rect 67542 176058 102986 176614
rect 103542 176058 138986 176614
rect 139542 176058 174986 176614
rect 175542 176058 210986 176614
rect 211542 176058 246986 176614
rect 247542 176058 282986 176614
rect 283542 176058 318986 176614
rect 319542 176058 354986 176614
rect 355542 176058 390986 176614
rect 391542 176058 426986 176614
rect 427542 176058 462986 176614
rect 463542 176058 498986 176614
rect 499542 176058 534986 176614
rect 535542 176058 570986 176614
rect 571542 176058 592062 176614
rect 592618 176058 592650 176614
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172338 -6774 172894
rect -6218 172338 27266 172894
rect 27822 172338 63266 172894
rect 63822 172338 99266 172894
rect 99822 172338 135266 172894
rect 135822 172338 171266 172894
rect 171822 172338 207266 172894
rect 207822 172338 243266 172894
rect 243822 172338 279266 172894
rect 279822 172338 315266 172894
rect 315822 172338 351266 172894
rect 351822 172338 387266 172894
rect 387822 172338 423266 172894
rect 423822 172338 459266 172894
rect 459822 172338 495266 172894
rect 495822 172338 531266 172894
rect 531822 172338 567266 172894
rect 567822 172338 590142 172894
rect 590698 172338 590730 172894
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168618 -4854 169174
rect -4298 168618 23546 169174
rect 24102 168618 59546 169174
rect 60102 168618 95546 169174
rect 96102 168618 131546 169174
rect 132102 168618 167546 169174
rect 168102 168618 203546 169174
rect 204102 168618 239546 169174
rect 240102 168618 275546 169174
rect 276102 168618 311546 169174
rect 312102 168618 347546 169174
rect 348102 168618 383546 169174
rect 384102 168618 419546 169174
rect 420102 168618 455546 169174
rect 456102 168618 491546 169174
rect 492102 168618 527546 169174
rect 528102 168618 563546 169174
rect 564102 168618 588222 169174
rect 588778 168618 588810 169174
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 164898 -2934 165454
rect -2378 164898 19826 165454
rect 20382 164898 55826 165454
rect 56382 164898 91826 165454
rect 92382 164898 127826 165454
rect 128382 164898 163826 165454
rect 164382 164898 199826 165454
rect 200382 164898 235826 165454
rect 236382 164898 271826 165454
rect 272382 164898 307826 165454
rect 308382 164898 343826 165454
rect 344382 164898 379826 165454
rect 380382 164898 415826 165454
rect 416382 164898 451826 165454
rect 452382 164898 487826 165454
rect 488382 164898 523826 165454
rect 524382 164898 559826 165454
rect 560382 164898 586302 165454
rect 586858 164898 586890 165454
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158058 -7734 158614
rect -7178 158058 12986 158614
rect 13542 158058 48986 158614
rect 49542 158058 84986 158614
rect 85542 158058 120986 158614
rect 121542 158058 156986 158614
rect 157542 158058 192986 158614
rect 193542 158058 228986 158614
rect 229542 158058 264986 158614
rect 265542 158058 300986 158614
rect 301542 158058 336986 158614
rect 337542 158058 372986 158614
rect 373542 158058 408986 158614
rect 409542 158058 444986 158614
rect 445542 158058 480986 158614
rect 481542 158058 516986 158614
rect 517542 158058 552986 158614
rect 553542 158058 591102 158614
rect 591658 158058 592650 158614
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154338 -5814 154894
rect -5258 154338 9266 154894
rect 9822 154338 45266 154894
rect 45822 154338 81266 154894
rect 81822 154338 117266 154894
rect 117822 154338 153266 154894
rect 153822 154338 189266 154894
rect 189822 154338 225266 154894
rect 225822 154338 261266 154894
rect 261822 154338 297266 154894
rect 297822 154338 333266 154894
rect 333822 154338 369266 154894
rect 369822 154338 405266 154894
rect 405822 154338 441266 154894
rect 441822 154338 477266 154894
rect 477822 154338 513266 154894
rect 513822 154338 549266 154894
rect 549822 154338 589182 154894
rect 589738 154338 590730 154894
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150618 -3894 151174
rect -3338 150618 5546 151174
rect 6102 150618 41546 151174
rect 42102 150618 77546 151174
rect 78102 150618 113546 151174
rect 114102 150618 149546 151174
rect 150102 150618 185546 151174
rect 186102 150618 221546 151174
rect 222102 150618 257546 151174
rect 258102 150618 293546 151174
rect 294102 150618 329546 151174
rect 330102 150618 365546 151174
rect 366102 150618 401546 151174
rect 402102 150618 437546 151174
rect 438102 150618 473546 151174
rect 474102 150618 509546 151174
rect 510102 150618 545546 151174
rect 546102 150618 581546 151174
rect 582102 150618 587262 151174
rect 587818 150618 588810 151174
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 146898 -1974 147454
rect -1418 146898 1826 147454
rect 2382 146898 37826 147454
rect 38382 146898 73826 147454
rect 74382 146898 109826 147454
rect 110382 146898 145826 147454
rect 146382 146898 181826 147454
rect 182382 146898 217826 147454
rect 218382 146898 253826 147454
rect 254382 146898 289826 147454
rect 290382 146898 325826 147454
rect 326382 146898 361826 147454
rect 362382 146898 397826 147454
rect 398382 146898 433826 147454
rect 434382 146898 469826 147454
rect 470382 146898 505826 147454
rect 506382 146898 541826 147454
rect 542382 146898 577826 147454
rect 578382 146898 585342 147454
rect 585898 146898 586890 147454
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140058 -8694 140614
rect -8138 140058 30986 140614
rect 31542 140058 66986 140614
rect 67542 140058 102986 140614
rect 103542 140058 138986 140614
rect 139542 140058 174986 140614
rect 175542 140058 210986 140614
rect 211542 140058 246986 140614
rect 247542 140058 282986 140614
rect 283542 140058 318986 140614
rect 319542 140058 354986 140614
rect 355542 140058 390986 140614
rect 391542 140058 426986 140614
rect 427542 140058 462986 140614
rect 463542 140058 498986 140614
rect 499542 140058 534986 140614
rect 535542 140058 570986 140614
rect 571542 140058 592062 140614
rect 592618 140058 592650 140614
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136338 -6774 136894
rect -6218 136338 27266 136894
rect 27822 136338 63266 136894
rect 63822 136338 99266 136894
rect 99822 136338 135266 136894
rect 135822 136338 171266 136894
rect 171822 136338 207266 136894
rect 207822 136338 243266 136894
rect 243822 136338 279266 136894
rect 279822 136338 315266 136894
rect 315822 136338 351266 136894
rect 351822 136338 387266 136894
rect 387822 136338 423266 136894
rect 423822 136338 459266 136894
rect 459822 136338 495266 136894
rect 495822 136338 531266 136894
rect 531822 136338 567266 136894
rect 567822 136338 590142 136894
rect 590698 136338 590730 136894
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132618 -4854 133174
rect -4298 132618 23546 133174
rect 24102 132618 59546 133174
rect 60102 132618 95546 133174
rect 96102 132618 131546 133174
rect 132102 132618 167546 133174
rect 168102 132618 203546 133174
rect 204102 132618 239546 133174
rect 240102 132618 275546 133174
rect 276102 132618 311546 133174
rect 312102 132618 347546 133174
rect 348102 132618 383546 133174
rect 384102 132618 419546 133174
rect 420102 132618 455546 133174
rect 456102 132618 491546 133174
rect 492102 132618 527546 133174
rect 528102 132618 563546 133174
rect 564102 132618 588222 133174
rect 588778 132618 588810 133174
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 128898 -2934 129454
rect -2378 128898 19826 129454
rect 20382 128898 55826 129454
rect 56382 128898 91826 129454
rect 92382 128898 127826 129454
rect 128382 128898 163826 129454
rect 164382 128898 199826 129454
rect 200382 128898 235826 129454
rect 236382 128898 271826 129454
rect 272382 128898 307826 129454
rect 308382 128898 343826 129454
rect 344382 128898 379826 129454
rect 380382 128898 415826 129454
rect 416382 128898 451826 129454
rect 452382 128898 487826 129454
rect 488382 128898 523826 129454
rect 524382 128898 559826 129454
rect 560382 128898 586302 129454
rect 586858 128898 586890 129454
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122058 -7734 122614
rect -7178 122058 12986 122614
rect 13542 122058 48986 122614
rect 49542 122058 84986 122614
rect 85542 122058 120986 122614
rect 121542 122058 156986 122614
rect 157542 122058 192986 122614
rect 193542 122058 228986 122614
rect 229542 122058 264986 122614
rect 265542 122058 300986 122614
rect 301542 122058 336986 122614
rect 337542 122058 372986 122614
rect 373542 122058 408986 122614
rect 409542 122058 444986 122614
rect 445542 122058 480986 122614
rect 481542 122058 516986 122614
rect 517542 122058 552986 122614
rect 553542 122058 591102 122614
rect 591658 122058 592650 122614
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118338 -5814 118894
rect -5258 118338 9266 118894
rect 9822 118338 45266 118894
rect 45822 118338 81266 118894
rect 81822 118338 117266 118894
rect 117822 118338 153266 118894
rect 153822 118338 189266 118894
rect 189822 118338 225266 118894
rect 225822 118338 261266 118894
rect 261822 118338 297266 118894
rect 297822 118338 333266 118894
rect 333822 118338 369266 118894
rect 369822 118338 405266 118894
rect 405822 118338 441266 118894
rect 441822 118338 477266 118894
rect 477822 118338 513266 118894
rect 513822 118338 549266 118894
rect 549822 118338 589182 118894
rect 589738 118338 590730 118894
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114618 -3894 115174
rect -3338 114618 5546 115174
rect 6102 114618 41546 115174
rect 42102 114618 77546 115174
rect 78102 114618 113546 115174
rect 114102 114618 149546 115174
rect 150102 114618 185546 115174
rect 186102 114618 221546 115174
rect 222102 114618 257546 115174
rect 258102 114618 293546 115174
rect 294102 114618 329546 115174
rect 330102 114618 365546 115174
rect 366102 114618 401546 115174
rect 402102 114618 437546 115174
rect 438102 114618 473546 115174
rect 474102 114618 509546 115174
rect 510102 114618 545546 115174
rect 546102 114618 581546 115174
rect 582102 114618 587262 115174
rect 587818 114618 588810 115174
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 110898 -1974 111454
rect -1418 110898 1826 111454
rect 2382 110898 37826 111454
rect 38382 110898 73826 111454
rect 74382 110898 109826 111454
rect 110382 110898 145826 111454
rect 146382 110898 181826 111454
rect 182382 110898 217826 111454
rect 218382 110898 253826 111454
rect 254382 110898 289826 111454
rect 290382 110898 325826 111454
rect 326382 110898 361826 111454
rect 362382 110898 397826 111454
rect 398382 110898 433826 111454
rect 434382 110898 469826 111454
rect 470382 110898 505826 111454
rect 506382 110898 541826 111454
rect 542382 110898 577826 111454
rect 578382 110898 585342 111454
rect 585898 110898 586890 111454
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104058 -8694 104614
rect -8138 104058 30986 104614
rect 31542 104058 66986 104614
rect 67542 104058 102986 104614
rect 103542 104058 138986 104614
rect 139542 104058 174986 104614
rect 175542 104058 210986 104614
rect 211542 104058 246986 104614
rect 247542 104058 282986 104614
rect 283542 104058 318986 104614
rect 319542 104058 354986 104614
rect 355542 104058 390986 104614
rect 391542 104058 426986 104614
rect 427542 104058 462986 104614
rect 463542 104058 498986 104614
rect 499542 104058 534986 104614
rect 535542 104058 570986 104614
rect 571542 104058 592062 104614
rect 592618 104058 592650 104614
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100338 -6774 100894
rect -6218 100338 27266 100894
rect 27822 100338 63266 100894
rect 63822 100338 99266 100894
rect 99822 100338 135266 100894
rect 135822 100338 171266 100894
rect 171822 100338 207266 100894
rect 207822 100338 243266 100894
rect 243822 100338 279266 100894
rect 279822 100338 315266 100894
rect 315822 100338 351266 100894
rect 351822 100338 387266 100894
rect 387822 100338 423266 100894
rect 423822 100338 459266 100894
rect 459822 100338 495266 100894
rect 495822 100338 531266 100894
rect 531822 100338 567266 100894
rect 567822 100338 590142 100894
rect 590698 100338 590730 100894
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96618 -4854 97174
rect -4298 96618 23546 97174
rect 24102 96618 59546 97174
rect 60102 96618 95546 97174
rect 96102 96618 131546 97174
rect 132102 96618 167546 97174
rect 168102 96618 203546 97174
rect 204102 96618 239546 97174
rect 240102 96618 275546 97174
rect 276102 96618 311546 97174
rect 312102 96618 347546 97174
rect 348102 96618 383546 97174
rect 384102 96618 419546 97174
rect 420102 96618 455546 97174
rect 456102 96618 491546 97174
rect 492102 96618 527546 97174
rect 528102 96618 563546 97174
rect 564102 96618 588222 97174
rect 588778 96618 588810 97174
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 92898 -2934 93454
rect -2378 92898 19826 93454
rect 20382 92898 55826 93454
rect 56382 92898 91826 93454
rect 92382 92898 127826 93454
rect 128382 92898 163826 93454
rect 164382 92898 199826 93454
rect 200382 92898 235826 93454
rect 236382 92898 271826 93454
rect 272382 92898 307826 93454
rect 308382 92898 343826 93454
rect 344382 92898 379826 93454
rect 380382 92898 415826 93454
rect 416382 92898 451826 93454
rect 452382 92898 487826 93454
rect 488382 92898 523826 93454
rect 524382 92898 559826 93454
rect 560382 92898 586302 93454
rect 586858 92898 586890 93454
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86058 -7734 86614
rect -7178 86058 12986 86614
rect 13542 86058 48986 86614
rect 49542 86058 84986 86614
rect 85542 86058 120986 86614
rect 121542 86058 156986 86614
rect 157542 86058 192986 86614
rect 193542 86058 228986 86614
rect 229542 86058 264986 86614
rect 265542 86058 300986 86614
rect 301542 86058 336986 86614
rect 337542 86058 372986 86614
rect 373542 86058 408986 86614
rect 409542 86058 444986 86614
rect 445542 86058 480986 86614
rect 481542 86058 516986 86614
rect 517542 86058 552986 86614
rect 553542 86058 591102 86614
rect 591658 86058 592650 86614
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82338 -5814 82894
rect -5258 82338 9266 82894
rect 9822 82338 45266 82894
rect 45822 82338 81266 82894
rect 81822 82338 117266 82894
rect 117822 82338 153266 82894
rect 153822 82338 189266 82894
rect 189822 82338 225266 82894
rect 225822 82338 261266 82894
rect 261822 82338 297266 82894
rect 297822 82338 333266 82894
rect 333822 82338 369266 82894
rect 369822 82338 405266 82894
rect 405822 82338 441266 82894
rect 441822 82338 477266 82894
rect 477822 82338 513266 82894
rect 513822 82338 549266 82894
rect 549822 82338 589182 82894
rect 589738 82338 590730 82894
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78618 -3894 79174
rect -3338 78618 5546 79174
rect 6102 78618 41546 79174
rect 42102 78618 77546 79174
rect 78102 78618 113546 79174
rect 114102 78618 149546 79174
rect 150102 78618 185546 79174
rect 186102 78618 221546 79174
rect 222102 78618 257546 79174
rect 258102 78618 293546 79174
rect 294102 78618 329546 79174
rect 330102 78618 365546 79174
rect 366102 78618 401546 79174
rect 402102 78618 437546 79174
rect 438102 78618 473546 79174
rect 474102 78618 509546 79174
rect 510102 78618 545546 79174
rect 546102 78618 581546 79174
rect 582102 78618 587262 79174
rect 587818 78618 588810 79174
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 74898 -1974 75454
rect -1418 74898 1826 75454
rect 2382 74898 37826 75454
rect 38382 74898 73826 75454
rect 74382 74898 109826 75454
rect 110382 74898 145826 75454
rect 146382 74898 181826 75454
rect 182382 74898 217826 75454
rect 218382 74898 253826 75454
rect 254382 74898 289826 75454
rect 290382 74898 325826 75454
rect 326382 74898 361826 75454
rect 362382 74898 397826 75454
rect 398382 74898 433826 75454
rect 434382 74898 469826 75454
rect 470382 74898 505826 75454
rect 506382 74898 541826 75454
rect 542382 74898 577826 75454
rect 578382 74898 585342 75454
rect 585898 74898 586890 75454
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68058 -8694 68614
rect -8138 68058 30986 68614
rect 31542 68058 66986 68614
rect 67542 68058 102986 68614
rect 103542 68058 138986 68614
rect 139542 68058 174986 68614
rect 175542 68058 210986 68614
rect 211542 68058 246986 68614
rect 247542 68058 282986 68614
rect 283542 68058 318986 68614
rect 319542 68058 354986 68614
rect 355542 68058 390986 68614
rect 391542 68058 426986 68614
rect 427542 68058 462986 68614
rect 463542 68058 498986 68614
rect 499542 68058 534986 68614
rect 535542 68058 570986 68614
rect 571542 68058 592062 68614
rect 592618 68058 592650 68614
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64338 -6774 64894
rect -6218 64338 27266 64894
rect 27822 64338 63266 64894
rect 63822 64338 99266 64894
rect 99822 64338 135266 64894
rect 135822 64338 171266 64894
rect 171822 64338 207266 64894
rect 207822 64338 243266 64894
rect 243822 64338 279266 64894
rect 279822 64338 315266 64894
rect 315822 64338 351266 64894
rect 351822 64338 387266 64894
rect 387822 64338 423266 64894
rect 423822 64338 459266 64894
rect 459822 64338 495266 64894
rect 495822 64338 531266 64894
rect 531822 64338 567266 64894
rect 567822 64338 590142 64894
rect 590698 64338 590730 64894
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60618 -4854 61174
rect -4298 60618 23546 61174
rect 24102 60618 59546 61174
rect 60102 60618 95546 61174
rect 96102 60618 131546 61174
rect 132102 60618 167546 61174
rect 168102 60618 203546 61174
rect 204102 60618 239546 61174
rect 240102 60618 275546 61174
rect 276102 60618 311546 61174
rect 312102 60618 347546 61174
rect 348102 60618 383546 61174
rect 384102 60618 419546 61174
rect 420102 60618 455546 61174
rect 456102 60618 491546 61174
rect 492102 60618 527546 61174
rect 528102 60618 563546 61174
rect 564102 60618 588222 61174
rect 588778 60618 588810 61174
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 56898 -2934 57454
rect -2378 56898 19826 57454
rect 20382 56898 55826 57454
rect 56382 56898 91826 57454
rect 92382 56898 127826 57454
rect 128382 56898 163826 57454
rect 164382 56898 199826 57454
rect 200382 56898 235826 57454
rect 236382 56898 271826 57454
rect 272382 56898 307826 57454
rect 308382 56898 343826 57454
rect 344382 56898 379826 57454
rect 380382 56898 415826 57454
rect 416382 56898 451826 57454
rect 452382 56898 487826 57454
rect 488382 56898 523826 57454
rect 524382 56898 559826 57454
rect 560382 56898 586302 57454
rect 586858 56898 586890 57454
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50058 -7734 50614
rect -7178 50058 12986 50614
rect 13542 50058 48986 50614
rect 49542 50058 84986 50614
rect 85542 50058 120986 50614
rect 121542 50058 156986 50614
rect 157542 50058 192986 50614
rect 193542 50058 228986 50614
rect 229542 50058 264986 50614
rect 265542 50058 300986 50614
rect 301542 50058 336986 50614
rect 337542 50058 372986 50614
rect 373542 50058 408986 50614
rect 409542 50058 444986 50614
rect 445542 50058 480986 50614
rect 481542 50058 516986 50614
rect 517542 50058 552986 50614
rect 553542 50058 591102 50614
rect 591658 50058 592650 50614
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46338 -5814 46894
rect -5258 46338 9266 46894
rect 9822 46338 45266 46894
rect 45822 46338 81266 46894
rect 81822 46338 117266 46894
rect 117822 46338 153266 46894
rect 153822 46338 189266 46894
rect 189822 46338 225266 46894
rect 225822 46338 261266 46894
rect 261822 46338 297266 46894
rect 297822 46338 333266 46894
rect 333822 46338 369266 46894
rect 369822 46338 405266 46894
rect 405822 46338 441266 46894
rect 441822 46338 477266 46894
rect 477822 46338 513266 46894
rect 513822 46338 549266 46894
rect 549822 46338 589182 46894
rect 589738 46338 590730 46894
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42618 -3894 43174
rect -3338 42618 5546 43174
rect 6102 42618 41546 43174
rect 42102 42618 77546 43174
rect 78102 42618 113546 43174
rect 114102 42618 149546 43174
rect 150102 42618 185546 43174
rect 186102 42618 221546 43174
rect 222102 42618 257546 43174
rect 258102 42618 293546 43174
rect 294102 42618 329546 43174
rect 330102 42618 365546 43174
rect 366102 42618 401546 43174
rect 402102 42618 437546 43174
rect 438102 42618 473546 43174
rect 474102 42618 509546 43174
rect 510102 42618 545546 43174
rect 546102 42618 581546 43174
rect 582102 42618 587262 43174
rect 587818 42618 588810 43174
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 38898 -1974 39454
rect -1418 38898 1826 39454
rect 2382 38898 37826 39454
rect 38382 38898 73826 39454
rect 74382 38898 109826 39454
rect 110382 38898 145826 39454
rect 146382 38898 181826 39454
rect 182382 38898 217826 39454
rect 218382 38898 253826 39454
rect 254382 38898 289826 39454
rect 290382 38898 325826 39454
rect 326382 38898 361826 39454
rect 362382 38898 397826 39454
rect 398382 38898 433826 39454
rect 434382 38898 469826 39454
rect 470382 38898 505826 39454
rect 506382 38898 541826 39454
rect 542382 38898 577826 39454
rect 578382 38898 585342 39454
rect 585898 38898 586890 39454
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32058 -8694 32614
rect -8138 32058 30986 32614
rect 31542 32058 66986 32614
rect 67542 32058 102986 32614
rect 103542 32058 138986 32614
rect 139542 32058 174986 32614
rect 175542 32058 210986 32614
rect 211542 32058 246986 32614
rect 247542 32058 282986 32614
rect 283542 32058 318986 32614
rect 319542 32058 354986 32614
rect 355542 32058 390986 32614
rect 391542 32058 426986 32614
rect 427542 32058 462986 32614
rect 463542 32058 498986 32614
rect 499542 32058 534986 32614
rect 535542 32058 570986 32614
rect 571542 32058 592062 32614
rect 592618 32058 592650 32614
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28338 -6774 28894
rect -6218 28338 27266 28894
rect 27822 28338 63266 28894
rect 63822 28338 99266 28894
rect 99822 28338 135266 28894
rect 135822 28338 171266 28894
rect 171822 28338 207266 28894
rect 207822 28338 243266 28894
rect 243822 28338 279266 28894
rect 279822 28338 315266 28894
rect 315822 28338 351266 28894
rect 351822 28338 387266 28894
rect 387822 28338 423266 28894
rect 423822 28338 459266 28894
rect 459822 28338 495266 28894
rect 495822 28338 531266 28894
rect 531822 28338 567266 28894
rect 567822 28338 590142 28894
rect 590698 28338 590730 28894
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24618 -4854 25174
rect -4298 24618 23546 25174
rect 24102 24618 59546 25174
rect 60102 24618 95546 25174
rect 96102 24618 131546 25174
rect 132102 24618 167546 25174
rect 168102 24618 203546 25174
rect 204102 24618 239546 25174
rect 240102 24618 275546 25174
rect 276102 24618 311546 25174
rect 312102 24618 347546 25174
rect 348102 24618 383546 25174
rect 384102 24618 419546 25174
rect 420102 24618 455546 25174
rect 456102 24618 491546 25174
rect 492102 24618 527546 25174
rect 528102 24618 563546 25174
rect 564102 24618 588222 25174
rect 588778 24618 588810 25174
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 20898 -2934 21454
rect -2378 20898 19826 21454
rect 20382 20898 55826 21454
rect 56382 20898 91826 21454
rect 92382 20898 127826 21454
rect 128382 20898 163826 21454
rect 164382 20898 199826 21454
rect 200382 20898 235826 21454
rect 236382 20898 271826 21454
rect 272382 20898 307826 21454
rect 308382 20898 343826 21454
rect 344382 20898 379826 21454
rect 380382 20898 415826 21454
rect 416382 20898 451826 21454
rect 452382 20898 487826 21454
rect 488382 20898 523826 21454
rect 524382 20898 559826 21454
rect 560382 20898 586302 21454
rect 586858 20898 586890 21454
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14058 -7734 14614
rect -7178 14058 12986 14614
rect 13542 14058 48986 14614
rect 49542 14058 84986 14614
rect 85542 14058 120986 14614
rect 121542 14058 156986 14614
rect 157542 14058 192986 14614
rect 193542 14058 228986 14614
rect 229542 14058 264986 14614
rect 265542 14058 300986 14614
rect 301542 14058 336986 14614
rect 337542 14058 372986 14614
rect 373542 14058 408986 14614
rect 409542 14058 444986 14614
rect 445542 14058 480986 14614
rect 481542 14058 516986 14614
rect 517542 14058 552986 14614
rect 553542 14058 591102 14614
rect 591658 14058 592650 14614
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10338 -5814 10894
rect -5258 10338 9266 10894
rect 9822 10338 45266 10894
rect 45822 10338 81266 10894
rect 81822 10338 117266 10894
rect 117822 10338 153266 10894
rect 153822 10338 189266 10894
rect 189822 10338 225266 10894
rect 225822 10338 261266 10894
rect 261822 10338 297266 10894
rect 297822 10338 333266 10894
rect 333822 10338 369266 10894
rect 369822 10338 405266 10894
rect 405822 10338 441266 10894
rect 441822 10338 477266 10894
rect 477822 10338 513266 10894
rect 513822 10338 549266 10894
rect 549822 10338 589182 10894
rect 589738 10338 590730 10894
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6618 -3894 7174
rect -3338 6618 5546 7174
rect 6102 6618 41546 7174
rect 42102 6618 77546 7174
rect 78102 6618 113546 7174
rect 114102 6618 149546 7174
rect 150102 6618 185546 7174
rect 186102 6618 221546 7174
rect 222102 6618 257546 7174
rect 258102 6618 293546 7174
rect 294102 6618 329546 7174
rect 330102 6618 365546 7174
rect 366102 6618 401546 7174
rect 402102 6618 437546 7174
rect 438102 6618 473546 7174
rect 474102 6618 509546 7174
rect 510102 6618 545546 7174
rect 546102 6618 581546 7174
rect 582102 6618 587262 7174
rect 587818 6618 588810 7174
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 2898 -1974 3454
rect -1418 2898 1826 3454
rect 2382 2898 37826 3454
rect 38382 2898 73826 3454
rect 74382 2898 109826 3454
rect 110382 2898 145826 3454
rect 146382 2898 181826 3454
rect 182382 2898 217826 3454
rect 218382 2898 253826 3454
rect 254382 2898 289826 3454
rect 290382 2898 325826 3454
rect 326382 2898 361826 3454
rect 362382 2898 397826 3454
rect 398382 2898 433826 3454
rect 434382 2898 469826 3454
rect 470382 2898 505826 3454
rect 506382 2898 541826 3454
rect 542382 2898 577826 3454
rect 578382 2898 585342 3454
rect 585898 2898 586890 3454
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -902 -1974 -346
rect -1418 -902 1826 -346
rect 2382 -902 37826 -346
rect 38382 -902 73826 -346
rect 74382 -902 109826 -346
rect 110382 -902 145826 -346
rect 146382 -902 181826 -346
rect 182382 -902 217826 -346
rect 218382 -902 253826 -346
rect 254382 -902 289826 -346
rect 290382 -902 325826 -346
rect 326382 -902 361826 -346
rect 362382 -902 397826 -346
rect 398382 -902 433826 -346
rect 434382 -902 469826 -346
rect 470382 -902 505826 -346
rect 506382 -902 541826 -346
rect 542382 -902 577826 -346
rect 578382 -902 585342 -346
rect 585898 -902 585930 -346
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1862 -2934 -1306
rect -2378 -1862 19826 -1306
rect 20382 -1862 55826 -1306
rect 56382 -1862 91826 -1306
rect 92382 -1862 127826 -1306
rect 128382 -1862 163826 -1306
rect 164382 -1862 199826 -1306
rect 200382 -1862 235826 -1306
rect 236382 -1862 271826 -1306
rect 272382 -1862 307826 -1306
rect 308382 -1862 343826 -1306
rect 344382 -1862 379826 -1306
rect 380382 -1862 415826 -1306
rect 416382 -1862 451826 -1306
rect 452382 -1862 487826 -1306
rect 488382 -1862 523826 -1306
rect 524382 -1862 559826 -1306
rect 560382 -1862 586302 -1306
rect 586858 -1862 586890 -1306
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2822 -3894 -2266
rect -3338 -2822 5546 -2266
rect 6102 -2822 41546 -2266
rect 42102 -2822 77546 -2266
rect 78102 -2822 113546 -2266
rect 114102 -2822 149546 -2266
rect 150102 -2822 185546 -2266
rect 186102 -2822 221546 -2266
rect 222102 -2822 257546 -2266
rect 258102 -2822 293546 -2266
rect 294102 -2822 329546 -2266
rect 330102 -2822 365546 -2266
rect 366102 -2822 401546 -2266
rect 402102 -2822 437546 -2266
rect 438102 -2822 473546 -2266
rect 474102 -2822 509546 -2266
rect 510102 -2822 545546 -2266
rect 546102 -2822 581546 -2266
rect 582102 -2822 587262 -2266
rect 587818 -2822 587850 -2266
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3782 -4854 -3226
rect -4298 -3782 23546 -3226
rect 24102 -3782 59546 -3226
rect 60102 -3782 95546 -3226
rect 96102 -3782 131546 -3226
rect 132102 -3782 167546 -3226
rect 168102 -3782 203546 -3226
rect 204102 -3782 239546 -3226
rect 240102 -3782 275546 -3226
rect 276102 -3782 311546 -3226
rect 312102 -3782 347546 -3226
rect 348102 -3782 383546 -3226
rect 384102 -3782 419546 -3226
rect 420102 -3782 455546 -3226
rect 456102 -3782 491546 -3226
rect 492102 -3782 527546 -3226
rect 528102 -3782 563546 -3226
rect 564102 -3782 588222 -3226
rect 588778 -3782 588810 -3226
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4742 -5814 -4186
rect -5258 -4742 9266 -4186
rect 9822 -4742 45266 -4186
rect 45822 -4742 81266 -4186
rect 81822 -4742 117266 -4186
rect 117822 -4742 153266 -4186
rect 153822 -4742 189266 -4186
rect 189822 -4742 225266 -4186
rect 225822 -4742 261266 -4186
rect 261822 -4742 297266 -4186
rect 297822 -4742 333266 -4186
rect 333822 -4742 369266 -4186
rect 369822 -4742 405266 -4186
rect 405822 -4742 441266 -4186
rect 441822 -4742 477266 -4186
rect 477822 -4742 513266 -4186
rect 513822 -4742 549266 -4186
rect 549822 -4742 589182 -4186
rect 589738 -4742 589770 -4186
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5702 -6774 -5146
rect -6218 -5702 27266 -5146
rect 27822 -5702 63266 -5146
rect 63822 -5702 99266 -5146
rect 99822 -5702 135266 -5146
rect 135822 -5702 171266 -5146
rect 171822 -5702 207266 -5146
rect 207822 -5702 243266 -5146
rect 243822 -5702 279266 -5146
rect 279822 -5702 315266 -5146
rect 315822 -5702 351266 -5146
rect 351822 -5702 387266 -5146
rect 387822 -5702 423266 -5146
rect 423822 -5702 459266 -5146
rect 459822 -5702 495266 -5146
rect 495822 -5702 531266 -5146
rect 531822 -5702 567266 -5146
rect 567822 -5702 590142 -5146
rect 590698 -5702 590730 -5146
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6662 -7734 -6106
rect -7178 -6662 12986 -6106
rect 13542 -6662 48986 -6106
rect 49542 -6662 84986 -6106
rect 85542 -6662 120986 -6106
rect 121542 -6662 156986 -6106
rect 157542 -6662 192986 -6106
rect 193542 -6662 228986 -6106
rect 229542 -6662 264986 -6106
rect 265542 -6662 300986 -6106
rect 301542 -6662 336986 -6106
rect 337542 -6662 372986 -6106
rect 373542 -6662 408986 -6106
rect 409542 -6662 444986 -6106
rect 445542 -6662 480986 -6106
rect 481542 -6662 516986 -6106
rect 517542 -6662 552986 -6106
rect 553542 -6662 591102 -6106
rect 591658 -6662 591690 -6106
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7622 -8694 -7066
rect -8138 -7622 30986 -7066
rect 31542 -7622 66986 -7066
rect 67542 -7622 102986 -7066
rect 103542 -7622 138986 -7066
rect 139542 -7622 174986 -7066
rect 175542 -7622 210986 -7066
rect 211542 -7622 246986 -7066
rect 247542 -7622 282986 -7066
rect 283542 -7622 318986 -7066
rect 319542 -7622 354986 -7066
rect 355542 -7622 390986 -7066
rect 391542 -7622 426986 -7066
rect 427542 -7622 462986 -7066
rect 463542 -7622 498986 -7066
rect 499542 -7622 534986 -7066
rect 535542 -7622 570986 -7066
rect 571542 -7622 592062 -7066
rect 592618 -7622 592650 -7066
rect -8726 -7654 592650 -7622
use user_proj_example  mprj
timestamp 0
transform 1 0 235000 0 1 338000
box 105 0 179846 120000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 4 analog_io[0]
port 1 nsew
rlabel metal2 s 446098 703520 446210 704960 4 analog_io[10]
port 2 nsew
rlabel metal2 s 381146 703520 381258 704960 4 analog_io[11]
port 3 nsew
rlabel metal2 s 316286 703520 316398 704960 4 analog_io[12]
port 4 nsew
rlabel metal2 s 251426 703520 251538 704960 4 analog_io[13]
port 5 nsew
rlabel metal2 s 186474 703520 186586 704960 4 analog_io[14]
port 6 nsew
rlabel metal2 s 121614 703520 121726 704960 4 analog_io[15]
port 7 nsew
rlabel metal2 s 56754 703520 56866 704960 4 analog_io[16]
port 8 nsew
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 9 nsew
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 10 nsew
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 11 nsew
rlabel metal3 s 583520 338452 584960 338692 4 analog_io[1]
port 12 nsew
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 13 nsew
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 14 nsew
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 15 nsew
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 16 nsew
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 17 nsew
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 18 nsew
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 19 nsew
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 20 nsew
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 21 nsew
rlabel metal3 s 583520 391628 584960 391868 4 analog_io[2]
port 22 nsew
rlabel metal3 s 583520 444668 584960 444908 4 analog_io[3]
port 23 nsew
rlabel metal3 s 583520 497844 584960 498084 4 analog_io[4]
port 24 nsew
rlabel metal3 s 583520 551020 584960 551260 4 analog_io[5]
port 25 nsew
rlabel metal3 s 583520 604060 584960 604300 4 analog_io[6]
port 26 nsew
rlabel metal3 s 583520 657236 584960 657476 4 analog_io[7]
port 27 nsew
rlabel metal2 s 575818 703520 575930 704960 4 analog_io[8]
port 28 nsew
rlabel metal2 s 510958 703520 511070 704960 4 analog_io[9]
port 29 nsew
rlabel metal3 s 583520 6476 584960 6716 4 io_in[0]
port 30 nsew
rlabel metal3 s 583520 457996 584960 458236 4 io_in[10]
port 31 nsew
rlabel metal3 s 583520 511172 584960 511412 4 io_in[11]
port 32 nsew
rlabel metal3 s 583520 564212 584960 564452 4 io_in[12]
port 33 nsew
rlabel metal3 s 583520 617388 584960 617628 4 io_in[13]
port 34 nsew
rlabel metal3 s 583520 670564 584960 670804 4 io_in[14]
port 35 nsew
rlabel metal2 s 559626 703520 559738 704960 4 io_in[15]
port 36 nsew
rlabel metal2 s 494766 703520 494878 704960 4 io_in[16]
port 37 nsew
rlabel metal2 s 429814 703520 429926 704960 4 io_in[17]
port 38 nsew
rlabel metal2 s 364954 703520 365066 704960 4 io_in[18]
port 39 nsew
rlabel metal2 s 300094 703520 300206 704960 4 io_in[19]
port 40 nsew
rlabel metal3 s 583520 46188 584960 46428 4 io_in[1]
port 41 nsew
rlabel metal2 s 235142 703520 235254 704960 4 io_in[20]
port 42 nsew
rlabel metal2 s 170282 703520 170394 704960 4 io_in[21]
port 43 nsew
rlabel metal2 s 105422 703520 105534 704960 4 io_in[22]
port 44 nsew
rlabel metal2 s 40470 703520 40582 704960 4 io_in[23]
port 45 nsew
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 46 nsew
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 47 nsew
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 48 nsew
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 49 nsew
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 50 nsew
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 51 nsew
rlabel metal3 s 583520 86036 584960 86276 4 io_in[2]
port 52 nsew
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 53 nsew
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 54 nsew
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 55 nsew
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 56 nsew
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 57 nsew
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 58 nsew
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 59 nsew
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 60 nsew
rlabel metal3 s 583520 125884 584960 126124 4 io_in[3]
port 61 nsew
rlabel metal3 s 583520 165732 584960 165972 4 io_in[4]
port 62 nsew
rlabel metal3 s 583520 205580 584960 205820 4 io_in[5]
port 63 nsew
rlabel metal3 s 583520 245428 584960 245668 4 io_in[6]
port 64 nsew
rlabel metal3 s 583520 298604 584960 298844 4 io_in[7]
port 65 nsew
rlabel metal3 s 583520 351780 584960 352020 4 io_in[8]
port 66 nsew
rlabel metal3 s 583520 404820 584960 405060 4 io_in[9]
port 67 nsew
rlabel metal3 s 583520 32996 584960 33236 4 io_oeb[0]
port 68 nsew
rlabel metal3 s 583520 484516 584960 484756 4 io_oeb[10]
port 69 nsew
rlabel metal3 s 583520 537692 584960 537932 4 io_oeb[11]
port 70 nsew
rlabel metal3 s 583520 590868 584960 591108 4 io_oeb[12]
port 71 nsew
rlabel metal3 s 583520 643908 584960 644148 4 io_oeb[13]
port 72 nsew
rlabel metal3 s 583520 697084 584960 697324 4 io_oeb[14]
port 73 nsew
rlabel metal2 s 527150 703520 527262 704960 4 io_oeb[15]
port 74 nsew
rlabel metal2 s 462290 703520 462402 704960 4 io_oeb[16]
port 75 nsew
rlabel metal2 s 397430 703520 397542 704960 4 io_oeb[17]
port 76 nsew
rlabel metal2 s 332478 703520 332590 704960 4 io_oeb[18]
port 77 nsew
rlabel metal2 s 267618 703520 267730 704960 4 io_oeb[19]
port 78 nsew
rlabel metal3 s 583520 72844 584960 73084 4 io_oeb[1]
port 79 nsew
rlabel metal2 s 202758 703520 202870 704960 4 io_oeb[20]
port 80 nsew
rlabel metal2 s 137806 703520 137918 704960 4 io_oeb[21]
port 81 nsew
rlabel metal2 s 72946 703520 73058 704960 4 io_oeb[22]
port 82 nsew
rlabel metal2 s 8086 703520 8198 704960 4 io_oeb[23]
port 83 nsew
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 84 nsew
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 85 nsew
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 86 nsew
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 87 nsew
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 88 nsew
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 89 nsew
rlabel metal3 s 583520 112692 584960 112932 4 io_oeb[2]
port 90 nsew
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 91 nsew
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 92 nsew
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 93 nsew
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 94 nsew
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 95 nsew
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 96 nsew
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 97 nsew
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 98 nsew
rlabel metal3 s 583520 152540 584960 152780 4 io_oeb[3]
port 99 nsew
rlabel metal3 s 583520 192388 584960 192628 4 io_oeb[4]
port 100 nsew
rlabel metal3 s 583520 232236 584960 232476 4 io_oeb[5]
port 101 nsew
rlabel metal3 s 583520 272084 584960 272324 4 io_oeb[6]
port 102 nsew
rlabel metal3 s 583520 325124 584960 325364 4 io_oeb[7]
port 103 nsew
rlabel metal3 s 583520 378300 584960 378540 4 io_oeb[8]
port 104 nsew
rlabel metal3 s 583520 431476 584960 431716 4 io_oeb[9]
port 105 nsew
rlabel metal3 s 583520 19668 584960 19908 4 io_out[0]
port 106 nsew
rlabel metal3 s 583520 471324 584960 471564 4 io_out[10]
port 107 nsew
rlabel metal3 s 583520 524364 584960 524604 4 io_out[11]
port 108 nsew
rlabel metal3 s 583520 577540 584960 577780 4 io_out[12]
port 109 nsew
rlabel metal3 s 583520 630716 584960 630956 4 io_out[13]
port 110 nsew
rlabel metal3 s 583520 683756 584960 683996 4 io_out[14]
port 111 nsew
rlabel metal2 s 543434 703520 543546 704960 4 io_out[15]
port 112 nsew
rlabel metal2 s 478482 703520 478594 704960 4 io_out[16]
port 113 nsew
rlabel metal2 s 413622 703520 413734 704960 4 io_out[17]
port 114 nsew
rlabel metal2 s 348762 703520 348874 704960 4 io_out[18]
port 115 nsew
rlabel metal2 s 283810 703520 283922 704960 4 io_out[19]
port 116 nsew
rlabel metal3 s 583520 59516 584960 59756 4 io_out[1]
port 117 nsew
rlabel metal2 s 218950 703520 219062 704960 4 io_out[20]
port 118 nsew
rlabel metal2 s 154090 703520 154202 704960 4 io_out[21]
port 119 nsew
rlabel metal2 s 89138 703520 89250 704960 4 io_out[22]
port 120 nsew
rlabel metal2 s 24278 703520 24390 704960 4 io_out[23]
port 121 nsew
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 122 nsew
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 123 nsew
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 124 nsew
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 125 nsew
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 126 nsew
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 127 nsew
rlabel metal3 s 583520 99364 584960 99604 4 io_out[2]
port 128 nsew
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 129 nsew
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 130 nsew
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 131 nsew
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 132 nsew
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 133 nsew
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 134 nsew
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 135 nsew
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 136 nsew
rlabel metal3 s 583520 139212 584960 139452 4 io_out[3]
port 137 nsew
rlabel metal3 s 583520 179060 584960 179300 4 io_out[4]
port 138 nsew
rlabel metal3 s 583520 218908 584960 219148 4 io_out[5]
port 139 nsew
rlabel metal3 s 583520 258756 584960 258996 4 io_out[6]
port 140 nsew
rlabel metal3 s 583520 311932 584960 312172 4 io_out[7]
port 141 nsew
rlabel metal3 s 583520 364972 584960 365212 4 io_out[8]
port 142 nsew
rlabel metal3 s 583520 418148 584960 418388 4 io_out[9]
port 143 nsew
rlabel metal2 s 125846 -960 125958 480 4 la_data_in[0]
port 144 nsew
rlabel metal2 s 480506 -960 480618 480 4 la_data_in[100]
port 145 nsew
rlabel metal2 s 484002 -960 484114 480 4 la_data_in[101]
port 146 nsew
rlabel metal2 s 487590 -960 487702 480 4 la_data_in[102]
port 147 nsew
rlabel metal2 s 491086 -960 491198 480 4 la_data_in[103]
port 148 nsew
rlabel metal2 s 494674 -960 494786 480 4 la_data_in[104]
port 149 nsew
rlabel metal2 s 498170 -960 498282 480 4 la_data_in[105]
port 150 nsew
rlabel metal2 s 501758 -960 501870 480 4 la_data_in[106]
port 151 nsew
rlabel metal2 s 505346 -960 505458 480 4 la_data_in[107]
port 152 nsew
rlabel metal2 s 508842 -960 508954 480 4 la_data_in[108]
port 153 nsew
rlabel metal2 s 512430 -960 512542 480 4 la_data_in[109]
port 154 nsew
rlabel metal2 s 161266 -960 161378 480 4 la_data_in[10]
port 155 nsew
rlabel metal2 s 515926 -960 516038 480 4 la_data_in[110]
port 156 nsew
rlabel metal2 s 519514 -960 519626 480 4 la_data_in[111]
port 157 nsew
rlabel metal2 s 523010 -960 523122 480 4 la_data_in[112]
port 158 nsew
rlabel metal2 s 526598 -960 526710 480 4 la_data_in[113]
port 159 nsew
rlabel metal2 s 530094 -960 530206 480 4 la_data_in[114]
port 160 nsew
rlabel metal2 s 533682 -960 533794 480 4 la_data_in[115]
port 161 nsew
rlabel metal2 s 537178 -960 537290 480 4 la_data_in[116]
port 162 nsew
rlabel metal2 s 540766 -960 540878 480 4 la_data_in[117]
port 163 nsew
rlabel metal2 s 544354 -960 544466 480 4 la_data_in[118]
port 164 nsew
rlabel metal2 s 547850 -960 547962 480 4 la_data_in[119]
port 165 nsew
rlabel metal2 s 164854 -960 164966 480 4 la_data_in[11]
port 166 nsew
rlabel metal2 s 551438 -960 551550 480 4 la_data_in[120]
port 167 nsew
rlabel metal2 s 554934 -960 555046 480 4 la_data_in[121]
port 168 nsew
rlabel metal2 s 558522 -960 558634 480 4 la_data_in[122]
port 169 nsew
rlabel metal2 s 562018 -960 562130 480 4 la_data_in[123]
port 170 nsew
rlabel metal2 s 565606 -960 565718 480 4 la_data_in[124]
port 171 nsew
rlabel metal2 s 569102 -960 569214 480 4 la_data_in[125]
port 172 nsew
rlabel metal2 s 572690 -960 572802 480 4 la_data_in[126]
port 173 nsew
rlabel metal2 s 576278 -960 576390 480 4 la_data_in[127]
port 174 nsew
rlabel metal2 s 168350 -960 168462 480 4 la_data_in[12]
port 175 nsew
rlabel metal2 s 171938 -960 172050 480 4 la_data_in[13]
port 176 nsew
rlabel metal2 s 175434 -960 175546 480 4 la_data_in[14]
port 177 nsew
rlabel metal2 s 179022 -960 179134 480 4 la_data_in[15]
port 178 nsew
rlabel metal2 s 182518 -960 182630 480 4 la_data_in[16]
port 179 nsew
rlabel metal2 s 186106 -960 186218 480 4 la_data_in[17]
port 180 nsew
rlabel metal2 s 189694 -960 189806 480 4 la_data_in[18]
port 181 nsew
rlabel metal2 s 193190 -960 193302 480 4 la_data_in[19]
port 182 nsew
rlabel metal2 s 129342 -960 129454 480 4 la_data_in[1]
port 183 nsew
rlabel metal2 s 196778 -960 196890 480 4 la_data_in[20]
port 184 nsew
rlabel metal2 s 200274 -960 200386 480 4 la_data_in[21]
port 185 nsew
rlabel metal2 s 203862 -960 203974 480 4 la_data_in[22]
port 186 nsew
rlabel metal2 s 207358 -960 207470 480 4 la_data_in[23]
port 187 nsew
rlabel metal2 s 210946 -960 211058 480 4 la_data_in[24]
port 188 nsew
rlabel metal2 s 214442 -960 214554 480 4 la_data_in[25]
port 189 nsew
rlabel metal2 s 218030 -960 218142 480 4 la_data_in[26]
port 190 nsew
rlabel metal2 s 221526 -960 221638 480 4 la_data_in[27]
port 191 nsew
rlabel metal2 s 225114 -960 225226 480 4 la_data_in[28]
port 192 nsew
rlabel metal2 s 228702 -960 228814 480 4 la_data_in[29]
port 193 nsew
rlabel metal2 s 132930 -960 133042 480 4 la_data_in[2]
port 194 nsew
rlabel metal2 s 232198 -960 232310 480 4 la_data_in[30]
port 195 nsew
rlabel metal2 s 235786 -960 235898 480 4 la_data_in[31]
port 196 nsew
rlabel metal2 s 239282 -960 239394 480 4 la_data_in[32]
port 197 nsew
rlabel metal2 s 242870 -960 242982 480 4 la_data_in[33]
port 198 nsew
rlabel metal2 s 246366 -960 246478 480 4 la_data_in[34]
port 199 nsew
rlabel metal2 s 249954 -960 250066 480 4 la_data_in[35]
port 200 nsew
rlabel metal2 s 253450 -960 253562 480 4 la_data_in[36]
port 201 nsew
rlabel metal2 s 257038 -960 257150 480 4 la_data_in[37]
port 202 nsew
rlabel metal2 s 260626 -960 260738 480 4 la_data_in[38]
port 203 nsew
rlabel metal2 s 264122 -960 264234 480 4 la_data_in[39]
port 204 nsew
rlabel metal2 s 136426 -960 136538 480 4 la_data_in[3]
port 205 nsew
rlabel metal2 s 267710 -960 267822 480 4 la_data_in[40]
port 206 nsew
rlabel metal2 s 271206 -960 271318 480 4 la_data_in[41]
port 207 nsew
rlabel metal2 s 274794 -960 274906 480 4 la_data_in[42]
port 208 nsew
rlabel metal2 s 278290 -960 278402 480 4 la_data_in[43]
port 209 nsew
rlabel metal2 s 281878 -960 281990 480 4 la_data_in[44]
port 210 nsew
rlabel metal2 s 285374 -960 285486 480 4 la_data_in[45]
port 211 nsew
rlabel metal2 s 288962 -960 289074 480 4 la_data_in[46]
port 212 nsew
rlabel metal2 s 292550 -960 292662 480 4 la_data_in[47]
port 213 nsew
rlabel metal2 s 296046 -960 296158 480 4 la_data_in[48]
port 214 nsew
rlabel metal2 s 299634 -960 299746 480 4 la_data_in[49]
port 215 nsew
rlabel metal2 s 140014 -960 140126 480 4 la_data_in[4]
port 216 nsew
rlabel metal2 s 303130 -960 303242 480 4 la_data_in[50]
port 217 nsew
rlabel metal2 s 306718 -960 306830 480 4 la_data_in[51]
port 218 nsew
rlabel metal2 s 310214 -960 310326 480 4 la_data_in[52]
port 219 nsew
rlabel metal2 s 313802 -960 313914 480 4 la_data_in[53]
port 220 nsew
rlabel metal2 s 317298 -960 317410 480 4 la_data_in[54]
port 221 nsew
rlabel metal2 s 320886 -960 320998 480 4 la_data_in[55]
port 222 nsew
rlabel metal2 s 324382 -960 324494 480 4 la_data_in[56]
port 223 nsew
rlabel metal2 s 327970 -960 328082 480 4 la_data_in[57]
port 224 nsew
rlabel metal2 s 331558 -960 331670 480 4 la_data_in[58]
port 225 nsew
rlabel metal2 s 335054 -960 335166 480 4 la_data_in[59]
port 226 nsew
rlabel metal2 s 143510 -960 143622 480 4 la_data_in[5]
port 227 nsew
rlabel metal2 s 338642 -960 338754 480 4 la_data_in[60]
port 228 nsew
rlabel metal2 s 342138 -960 342250 480 4 la_data_in[61]
port 229 nsew
rlabel metal2 s 345726 -960 345838 480 4 la_data_in[62]
port 230 nsew
rlabel metal2 s 349222 -960 349334 480 4 la_data_in[63]
port 231 nsew
rlabel metal2 s 352810 -960 352922 480 4 la_data_in[64]
port 232 nsew
rlabel metal2 s 356306 -960 356418 480 4 la_data_in[65]
port 233 nsew
rlabel metal2 s 359894 -960 360006 480 4 la_data_in[66]
port 234 nsew
rlabel metal2 s 363482 -960 363594 480 4 la_data_in[67]
port 235 nsew
rlabel metal2 s 366978 -960 367090 480 4 la_data_in[68]
port 236 nsew
rlabel metal2 s 370566 -960 370678 480 4 la_data_in[69]
port 237 nsew
rlabel metal2 s 147098 -960 147210 480 4 la_data_in[6]
port 238 nsew
rlabel metal2 s 374062 -960 374174 480 4 la_data_in[70]
port 239 nsew
rlabel metal2 s 377650 -960 377762 480 4 la_data_in[71]
port 240 nsew
rlabel metal2 s 381146 -960 381258 480 4 la_data_in[72]
port 241 nsew
rlabel metal2 s 384734 -960 384846 480 4 la_data_in[73]
port 242 nsew
rlabel metal2 s 388230 -960 388342 480 4 la_data_in[74]
port 243 nsew
rlabel metal2 s 391818 -960 391930 480 4 la_data_in[75]
port 244 nsew
rlabel metal2 s 395314 -960 395426 480 4 la_data_in[76]
port 245 nsew
rlabel metal2 s 398902 -960 399014 480 4 la_data_in[77]
port 246 nsew
rlabel metal2 s 402490 -960 402602 480 4 la_data_in[78]
port 247 nsew
rlabel metal2 s 405986 -960 406098 480 4 la_data_in[79]
port 248 nsew
rlabel metal2 s 150594 -960 150706 480 4 la_data_in[7]
port 249 nsew
rlabel metal2 s 409574 -960 409686 480 4 la_data_in[80]
port 250 nsew
rlabel metal2 s 413070 -960 413182 480 4 la_data_in[81]
port 251 nsew
rlabel metal2 s 416658 -960 416770 480 4 la_data_in[82]
port 252 nsew
rlabel metal2 s 420154 -960 420266 480 4 la_data_in[83]
port 253 nsew
rlabel metal2 s 423742 -960 423854 480 4 la_data_in[84]
port 254 nsew
rlabel metal2 s 427238 -960 427350 480 4 la_data_in[85]
port 255 nsew
rlabel metal2 s 430826 -960 430938 480 4 la_data_in[86]
port 256 nsew
rlabel metal2 s 434414 -960 434526 480 4 la_data_in[87]
port 257 nsew
rlabel metal2 s 437910 -960 438022 480 4 la_data_in[88]
port 258 nsew
rlabel metal2 s 441498 -960 441610 480 4 la_data_in[89]
port 259 nsew
rlabel metal2 s 154182 -960 154294 480 4 la_data_in[8]
port 260 nsew
rlabel metal2 s 444994 -960 445106 480 4 la_data_in[90]
port 261 nsew
rlabel metal2 s 448582 -960 448694 480 4 la_data_in[91]
port 262 nsew
rlabel metal2 s 452078 -960 452190 480 4 la_data_in[92]
port 263 nsew
rlabel metal2 s 455666 -960 455778 480 4 la_data_in[93]
port 264 nsew
rlabel metal2 s 459162 -960 459274 480 4 la_data_in[94]
port 265 nsew
rlabel metal2 s 462750 -960 462862 480 4 la_data_in[95]
port 266 nsew
rlabel metal2 s 466246 -960 466358 480 4 la_data_in[96]
port 267 nsew
rlabel metal2 s 469834 -960 469946 480 4 la_data_in[97]
port 268 nsew
rlabel metal2 s 473422 -960 473534 480 4 la_data_in[98]
port 269 nsew
rlabel metal2 s 476918 -960 477030 480 4 la_data_in[99]
port 270 nsew
rlabel metal2 s 157770 -960 157882 480 4 la_data_in[9]
port 271 nsew
rlabel metal2 s 126950 -960 127062 480 4 la_data_out[0]
port 272 nsew
rlabel metal2 s 481702 -960 481814 480 4 la_data_out[100]
port 273 nsew
rlabel metal2 s 485198 -960 485310 480 4 la_data_out[101]
port 274 nsew
rlabel metal2 s 488786 -960 488898 480 4 la_data_out[102]
port 275 nsew
rlabel metal2 s 492282 -960 492394 480 4 la_data_out[103]
port 276 nsew
rlabel metal2 s 495870 -960 495982 480 4 la_data_out[104]
port 277 nsew
rlabel metal2 s 499366 -960 499478 480 4 la_data_out[105]
port 278 nsew
rlabel metal2 s 502954 -960 503066 480 4 la_data_out[106]
port 279 nsew
rlabel metal2 s 506450 -960 506562 480 4 la_data_out[107]
port 280 nsew
rlabel metal2 s 510038 -960 510150 480 4 la_data_out[108]
port 281 nsew
rlabel metal2 s 513534 -960 513646 480 4 la_data_out[109]
port 282 nsew
rlabel metal2 s 162462 -960 162574 480 4 la_data_out[10]
port 283 nsew
rlabel metal2 s 517122 -960 517234 480 4 la_data_out[110]
port 284 nsew
rlabel metal2 s 520710 -960 520822 480 4 la_data_out[111]
port 285 nsew
rlabel metal2 s 524206 -960 524318 480 4 la_data_out[112]
port 286 nsew
rlabel metal2 s 527794 -960 527906 480 4 la_data_out[113]
port 287 nsew
rlabel metal2 s 531290 -960 531402 480 4 la_data_out[114]
port 288 nsew
rlabel metal2 s 534878 -960 534990 480 4 la_data_out[115]
port 289 nsew
rlabel metal2 s 538374 -960 538486 480 4 la_data_out[116]
port 290 nsew
rlabel metal2 s 541962 -960 542074 480 4 la_data_out[117]
port 291 nsew
rlabel metal2 s 545458 -960 545570 480 4 la_data_out[118]
port 292 nsew
rlabel metal2 s 549046 -960 549158 480 4 la_data_out[119]
port 293 nsew
rlabel metal2 s 166050 -960 166162 480 4 la_data_out[11]
port 294 nsew
rlabel metal2 s 552634 -960 552746 480 4 la_data_out[120]
port 295 nsew
rlabel metal2 s 556130 -960 556242 480 4 la_data_out[121]
port 296 nsew
rlabel metal2 s 559718 -960 559830 480 4 la_data_out[122]
port 297 nsew
rlabel metal2 s 563214 -960 563326 480 4 la_data_out[123]
port 298 nsew
rlabel metal2 s 566802 -960 566914 480 4 la_data_out[124]
port 299 nsew
rlabel metal2 s 570298 -960 570410 480 4 la_data_out[125]
port 300 nsew
rlabel metal2 s 573886 -960 573998 480 4 la_data_out[126]
port 301 nsew
rlabel metal2 s 577382 -960 577494 480 4 la_data_out[127]
port 302 nsew
rlabel metal2 s 169546 -960 169658 480 4 la_data_out[12]
port 303 nsew
rlabel metal2 s 173134 -960 173246 480 4 la_data_out[13]
port 304 nsew
rlabel metal2 s 176630 -960 176742 480 4 la_data_out[14]
port 305 nsew
rlabel metal2 s 180218 -960 180330 480 4 la_data_out[15]
port 306 nsew
rlabel metal2 s 183714 -960 183826 480 4 la_data_out[16]
port 307 nsew
rlabel metal2 s 187302 -960 187414 480 4 la_data_out[17]
port 308 nsew
rlabel metal2 s 190798 -960 190910 480 4 la_data_out[18]
port 309 nsew
rlabel metal2 s 194386 -960 194498 480 4 la_data_out[19]
port 310 nsew
rlabel metal2 s 130538 -960 130650 480 4 la_data_out[1]
port 311 nsew
rlabel metal2 s 197882 -960 197994 480 4 la_data_out[20]
port 312 nsew
rlabel metal2 s 201470 -960 201582 480 4 la_data_out[21]
port 313 nsew
rlabel metal2 s 205058 -960 205170 480 4 la_data_out[22]
port 314 nsew
rlabel metal2 s 208554 -960 208666 480 4 la_data_out[23]
port 315 nsew
rlabel metal2 s 212142 -960 212254 480 4 la_data_out[24]
port 316 nsew
rlabel metal2 s 215638 -960 215750 480 4 la_data_out[25]
port 317 nsew
rlabel metal2 s 219226 -960 219338 480 4 la_data_out[26]
port 318 nsew
rlabel metal2 s 222722 -960 222834 480 4 la_data_out[27]
port 319 nsew
rlabel metal2 s 226310 -960 226422 480 4 la_data_out[28]
port 320 nsew
rlabel metal2 s 229806 -960 229918 480 4 la_data_out[29]
port 321 nsew
rlabel metal2 s 134126 -960 134238 480 4 la_data_out[2]
port 322 nsew
rlabel metal2 s 233394 -960 233506 480 4 la_data_out[30]
port 323 nsew
rlabel metal2 s 236982 -960 237094 480 4 la_data_out[31]
port 324 nsew
rlabel metal2 s 240478 -960 240590 480 4 la_data_out[32]
port 325 nsew
rlabel metal2 s 244066 -960 244178 480 4 la_data_out[33]
port 326 nsew
rlabel metal2 s 247562 -960 247674 480 4 la_data_out[34]
port 327 nsew
rlabel metal2 s 251150 -960 251262 480 4 la_data_out[35]
port 328 nsew
rlabel metal2 s 254646 -960 254758 480 4 la_data_out[36]
port 329 nsew
rlabel metal2 s 258234 -960 258346 480 4 la_data_out[37]
port 330 nsew
rlabel metal2 s 261730 -960 261842 480 4 la_data_out[38]
port 331 nsew
rlabel metal2 s 265318 -960 265430 480 4 la_data_out[39]
port 332 nsew
rlabel metal2 s 137622 -960 137734 480 4 la_data_out[3]
port 333 nsew
rlabel metal2 s 268814 -960 268926 480 4 la_data_out[40]
port 334 nsew
rlabel metal2 s 272402 -960 272514 480 4 la_data_out[41]
port 335 nsew
rlabel metal2 s 275990 -960 276102 480 4 la_data_out[42]
port 336 nsew
rlabel metal2 s 279486 -960 279598 480 4 la_data_out[43]
port 337 nsew
rlabel metal2 s 283074 -960 283186 480 4 la_data_out[44]
port 338 nsew
rlabel metal2 s 286570 -960 286682 480 4 la_data_out[45]
port 339 nsew
rlabel metal2 s 290158 -960 290270 480 4 la_data_out[46]
port 340 nsew
rlabel metal2 s 293654 -960 293766 480 4 la_data_out[47]
port 341 nsew
rlabel metal2 s 297242 -960 297354 480 4 la_data_out[48]
port 342 nsew
rlabel metal2 s 300738 -960 300850 480 4 la_data_out[49]
port 343 nsew
rlabel metal2 s 141210 -960 141322 480 4 la_data_out[4]
port 344 nsew
rlabel metal2 s 304326 -960 304438 480 4 la_data_out[50]
port 345 nsew
rlabel metal2 s 307914 -960 308026 480 4 la_data_out[51]
port 346 nsew
rlabel metal2 s 311410 -960 311522 480 4 la_data_out[52]
port 347 nsew
rlabel metal2 s 314998 -960 315110 480 4 la_data_out[53]
port 348 nsew
rlabel metal2 s 318494 -960 318606 480 4 la_data_out[54]
port 349 nsew
rlabel metal2 s 322082 -960 322194 480 4 la_data_out[55]
port 350 nsew
rlabel metal2 s 325578 -960 325690 480 4 la_data_out[56]
port 351 nsew
rlabel metal2 s 329166 -960 329278 480 4 la_data_out[57]
port 352 nsew
rlabel metal2 s 332662 -960 332774 480 4 la_data_out[58]
port 353 nsew
rlabel metal2 s 336250 -960 336362 480 4 la_data_out[59]
port 354 nsew
rlabel metal2 s 144706 -960 144818 480 4 la_data_out[5]
port 355 nsew
rlabel metal2 s 339838 -960 339950 480 4 la_data_out[60]
port 356 nsew
rlabel metal2 s 343334 -960 343446 480 4 la_data_out[61]
port 357 nsew
rlabel metal2 s 346922 -960 347034 480 4 la_data_out[62]
port 358 nsew
rlabel metal2 s 350418 -960 350530 480 4 la_data_out[63]
port 359 nsew
rlabel metal2 s 354006 -960 354118 480 4 la_data_out[64]
port 360 nsew
rlabel metal2 s 357502 -960 357614 480 4 la_data_out[65]
port 361 nsew
rlabel metal2 s 361090 -960 361202 480 4 la_data_out[66]
port 362 nsew
rlabel metal2 s 364586 -960 364698 480 4 la_data_out[67]
port 363 nsew
rlabel metal2 s 368174 -960 368286 480 4 la_data_out[68]
port 364 nsew
rlabel metal2 s 371670 -960 371782 480 4 la_data_out[69]
port 365 nsew
rlabel metal2 s 148294 -960 148406 480 4 la_data_out[6]
port 366 nsew
rlabel metal2 s 375258 -960 375370 480 4 la_data_out[70]
port 367 nsew
rlabel metal2 s 378846 -960 378958 480 4 la_data_out[71]
port 368 nsew
rlabel metal2 s 382342 -960 382454 480 4 la_data_out[72]
port 369 nsew
rlabel metal2 s 385930 -960 386042 480 4 la_data_out[73]
port 370 nsew
rlabel metal2 s 389426 -960 389538 480 4 la_data_out[74]
port 371 nsew
rlabel metal2 s 393014 -960 393126 480 4 la_data_out[75]
port 372 nsew
rlabel metal2 s 396510 -960 396622 480 4 la_data_out[76]
port 373 nsew
rlabel metal2 s 400098 -960 400210 480 4 la_data_out[77]
port 374 nsew
rlabel metal2 s 403594 -960 403706 480 4 la_data_out[78]
port 375 nsew
rlabel metal2 s 407182 -960 407294 480 4 la_data_out[79]
port 376 nsew
rlabel metal2 s 151790 -960 151902 480 4 la_data_out[7]
port 377 nsew
rlabel metal2 s 410770 -960 410882 480 4 la_data_out[80]
port 378 nsew
rlabel metal2 s 414266 -960 414378 480 4 la_data_out[81]
port 379 nsew
rlabel metal2 s 417854 -960 417966 480 4 la_data_out[82]
port 380 nsew
rlabel metal2 s 421350 -960 421462 480 4 la_data_out[83]
port 381 nsew
rlabel metal2 s 424938 -960 425050 480 4 la_data_out[84]
port 382 nsew
rlabel metal2 s 428434 -960 428546 480 4 la_data_out[85]
port 383 nsew
rlabel metal2 s 432022 -960 432134 480 4 la_data_out[86]
port 384 nsew
rlabel metal2 s 435518 -960 435630 480 4 la_data_out[87]
port 385 nsew
rlabel metal2 s 439106 -960 439218 480 4 la_data_out[88]
port 386 nsew
rlabel metal2 s 442602 -960 442714 480 4 la_data_out[89]
port 387 nsew
rlabel metal2 s 155378 -960 155490 480 4 la_data_out[8]
port 388 nsew
rlabel metal2 s 446190 -960 446302 480 4 la_data_out[90]
port 389 nsew
rlabel metal2 s 449778 -960 449890 480 4 la_data_out[91]
port 390 nsew
rlabel metal2 s 453274 -960 453386 480 4 la_data_out[92]
port 391 nsew
rlabel metal2 s 456862 -960 456974 480 4 la_data_out[93]
port 392 nsew
rlabel metal2 s 460358 -960 460470 480 4 la_data_out[94]
port 393 nsew
rlabel metal2 s 463946 -960 464058 480 4 la_data_out[95]
port 394 nsew
rlabel metal2 s 467442 -960 467554 480 4 la_data_out[96]
port 395 nsew
rlabel metal2 s 471030 -960 471142 480 4 la_data_out[97]
port 396 nsew
rlabel metal2 s 474526 -960 474638 480 4 la_data_out[98]
port 397 nsew
rlabel metal2 s 478114 -960 478226 480 4 la_data_out[99]
port 398 nsew
rlabel metal2 s 158874 -960 158986 480 4 la_data_out[9]
port 399 nsew
rlabel metal2 s 128146 -960 128258 480 4 la_oenb[0]
port 400 nsew
rlabel metal2 s 482806 -960 482918 480 4 la_oenb[100]
port 401 nsew
rlabel metal2 s 486394 -960 486506 480 4 la_oenb[101]
port 402 nsew
rlabel metal2 s 489890 -960 490002 480 4 la_oenb[102]
port 403 nsew
rlabel metal2 s 493478 -960 493590 480 4 la_oenb[103]
port 404 nsew
rlabel metal2 s 497066 -960 497178 480 4 la_oenb[104]
port 405 nsew
rlabel metal2 s 500562 -960 500674 480 4 la_oenb[105]
port 406 nsew
rlabel metal2 s 504150 -960 504262 480 4 la_oenb[106]
port 407 nsew
rlabel metal2 s 507646 -960 507758 480 4 la_oenb[107]
port 408 nsew
rlabel metal2 s 511234 -960 511346 480 4 la_oenb[108]
port 409 nsew
rlabel metal2 s 514730 -960 514842 480 4 la_oenb[109]
port 410 nsew
rlabel metal2 s 163658 -960 163770 480 4 la_oenb[10]
port 411 nsew
rlabel metal2 s 518318 -960 518430 480 4 la_oenb[110]
port 412 nsew
rlabel metal2 s 521814 -960 521926 480 4 la_oenb[111]
port 413 nsew
rlabel metal2 s 525402 -960 525514 480 4 la_oenb[112]
port 414 nsew
rlabel metal2 s 528990 -960 529102 480 4 la_oenb[113]
port 415 nsew
rlabel metal2 s 532486 -960 532598 480 4 la_oenb[114]
port 416 nsew
rlabel metal2 s 536074 -960 536186 480 4 la_oenb[115]
port 417 nsew
rlabel metal2 s 539570 -960 539682 480 4 la_oenb[116]
port 418 nsew
rlabel metal2 s 543158 -960 543270 480 4 la_oenb[117]
port 419 nsew
rlabel metal2 s 546654 -960 546766 480 4 la_oenb[118]
port 420 nsew
rlabel metal2 s 550242 -960 550354 480 4 la_oenb[119]
port 421 nsew
rlabel metal2 s 167154 -960 167266 480 4 la_oenb[11]
port 422 nsew
rlabel metal2 s 553738 -960 553850 480 4 la_oenb[120]
port 423 nsew
rlabel metal2 s 557326 -960 557438 480 4 la_oenb[121]
port 424 nsew
rlabel metal2 s 560822 -960 560934 480 4 la_oenb[122]
port 425 nsew
rlabel metal2 s 564410 -960 564522 480 4 la_oenb[123]
port 426 nsew
rlabel metal2 s 567998 -960 568110 480 4 la_oenb[124]
port 427 nsew
rlabel metal2 s 571494 -960 571606 480 4 la_oenb[125]
port 428 nsew
rlabel metal2 s 575082 -960 575194 480 4 la_oenb[126]
port 429 nsew
rlabel metal2 s 578578 -960 578690 480 4 la_oenb[127]
port 430 nsew
rlabel metal2 s 170742 -960 170854 480 4 la_oenb[12]
port 431 nsew
rlabel metal2 s 174238 -960 174350 480 4 la_oenb[13]
port 432 nsew
rlabel metal2 s 177826 -960 177938 480 4 la_oenb[14]
port 433 nsew
rlabel metal2 s 181414 -960 181526 480 4 la_oenb[15]
port 434 nsew
rlabel metal2 s 184910 -960 185022 480 4 la_oenb[16]
port 435 nsew
rlabel metal2 s 188498 -960 188610 480 4 la_oenb[17]
port 436 nsew
rlabel metal2 s 191994 -960 192106 480 4 la_oenb[18]
port 437 nsew
rlabel metal2 s 195582 -960 195694 480 4 la_oenb[19]
port 438 nsew
rlabel metal2 s 131734 -960 131846 480 4 la_oenb[1]
port 439 nsew
rlabel metal2 s 199078 -960 199190 480 4 la_oenb[20]
port 440 nsew
rlabel metal2 s 202666 -960 202778 480 4 la_oenb[21]
port 441 nsew
rlabel metal2 s 206162 -960 206274 480 4 la_oenb[22]
port 442 nsew
rlabel metal2 s 209750 -960 209862 480 4 la_oenb[23]
port 443 nsew
rlabel metal2 s 213338 -960 213450 480 4 la_oenb[24]
port 444 nsew
rlabel metal2 s 216834 -960 216946 480 4 la_oenb[25]
port 445 nsew
rlabel metal2 s 220422 -960 220534 480 4 la_oenb[26]
port 446 nsew
rlabel metal2 s 223918 -960 224030 480 4 la_oenb[27]
port 447 nsew
rlabel metal2 s 227506 -960 227618 480 4 la_oenb[28]
port 448 nsew
rlabel metal2 s 231002 -960 231114 480 4 la_oenb[29]
port 449 nsew
rlabel metal2 s 135230 -960 135342 480 4 la_oenb[2]
port 450 nsew
rlabel metal2 s 234590 -960 234702 480 4 la_oenb[30]
port 451 nsew
rlabel metal2 s 238086 -960 238198 480 4 la_oenb[31]
port 452 nsew
rlabel metal2 s 241674 -960 241786 480 4 la_oenb[32]
port 453 nsew
rlabel metal2 s 245170 -960 245282 480 4 la_oenb[33]
port 454 nsew
rlabel metal2 s 248758 -960 248870 480 4 la_oenb[34]
port 455 nsew
rlabel metal2 s 252346 -960 252458 480 4 la_oenb[35]
port 456 nsew
rlabel metal2 s 255842 -960 255954 480 4 la_oenb[36]
port 457 nsew
rlabel metal2 s 259430 -960 259542 480 4 la_oenb[37]
port 458 nsew
rlabel metal2 s 262926 -960 263038 480 4 la_oenb[38]
port 459 nsew
rlabel metal2 s 266514 -960 266626 480 4 la_oenb[39]
port 460 nsew
rlabel metal2 s 138818 -960 138930 480 4 la_oenb[3]
port 461 nsew
rlabel metal2 s 270010 -960 270122 480 4 la_oenb[40]
port 462 nsew
rlabel metal2 s 273598 -960 273710 480 4 la_oenb[41]
port 463 nsew
rlabel metal2 s 277094 -960 277206 480 4 la_oenb[42]
port 464 nsew
rlabel metal2 s 280682 -960 280794 480 4 la_oenb[43]
port 465 nsew
rlabel metal2 s 284270 -960 284382 480 4 la_oenb[44]
port 466 nsew
rlabel metal2 s 287766 -960 287878 480 4 la_oenb[45]
port 467 nsew
rlabel metal2 s 291354 -960 291466 480 4 la_oenb[46]
port 468 nsew
rlabel metal2 s 294850 -960 294962 480 4 la_oenb[47]
port 469 nsew
rlabel metal2 s 298438 -960 298550 480 4 la_oenb[48]
port 470 nsew
rlabel metal2 s 301934 -960 302046 480 4 la_oenb[49]
port 471 nsew
rlabel metal2 s 142406 -960 142518 480 4 la_oenb[4]
port 472 nsew
rlabel metal2 s 305522 -960 305634 480 4 la_oenb[50]
port 473 nsew
rlabel metal2 s 309018 -960 309130 480 4 la_oenb[51]
port 474 nsew
rlabel metal2 s 312606 -960 312718 480 4 la_oenb[52]
port 475 nsew
rlabel metal2 s 316194 -960 316306 480 4 la_oenb[53]
port 476 nsew
rlabel metal2 s 319690 -960 319802 480 4 la_oenb[54]
port 477 nsew
rlabel metal2 s 323278 -960 323390 480 4 la_oenb[55]
port 478 nsew
rlabel metal2 s 326774 -960 326886 480 4 la_oenb[56]
port 479 nsew
rlabel metal2 s 330362 -960 330474 480 4 la_oenb[57]
port 480 nsew
rlabel metal2 s 333858 -960 333970 480 4 la_oenb[58]
port 481 nsew
rlabel metal2 s 337446 -960 337558 480 4 la_oenb[59]
port 482 nsew
rlabel metal2 s 145902 -960 146014 480 4 la_oenb[5]
port 483 nsew
rlabel metal2 s 340942 -960 341054 480 4 la_oenb[60]
port 484 nsew
rlabel metal2 s 344530 -960 344642 480 4 la_oenb[61]
port 485 nsew
rlabel metal2 s 348026 -960 348138 480 4 la_oenb[62]
port 486 nsew
rlabel metal2 s 351614 -960 351726 480 4 la_oenb[63]
port 487 nsew
rlabel metal2 s 355202 -960 355314 480 4 la_oenb[64]
port 488 nsew
rlabel metal2 s 358698 -960 358810 480 4 la_oenb[65]
port 489 nsew
rlabel metal2 s 362286 -960 362398 480 4 la_oenb[66]
port 490 nsew
rlabel metal2 s 365782 -960 365894 480 4 la_oenb[67]
port 491 nsew
rlabel metal2 s 369370 -960 369482 480 4 la_oenb[68]
port 492 nsew
rlabel metal2 s 372866 -960 372978 480 4 la_oenb[69]
port 493 nsew
rlabel metal2 s 149490 -960 149602 480 4 la_oenb[6]
port 494 nsew
rlabel metal2 s 376454 -960 376566 480 4 la_oenb[70]
port 495 nsew
rlabel metal2 s 379950 -960 380062 480 4 la_oenb[71]
port 496 nsew
rlabel metal2 s 383538 -960 383650 480 4 la_oenb[72]
port 497 nsew
rlabel metal2 s 387126 -960 387238 480 4 la_oenb[73]
port 498 nsew
rlabel metal2 s 390622 -960 390734 480 4 la_oenb[74]
port 499 nsew
rlabel metal2 s 394210 -960 394322 480 4 la_oenb[75]
port 500 nsew
rlabel metal2 s 397706 -960 397818 480 4 la_oenb[76]
port 501 nsew
rlabel metal2 s 401294 -960 401406 480 4 la_oenb[77]
port 502 nsew
rlabel metal2 s 404790 -960 404902 480 4 la_oenb[78]
port 503 nsew
rlabel metal2 s 408378 -960 408490 480 4 la_oenb[79]
port 504 nsew
rlabel metal2 s 152986 -960 153098 480 4 la_oenb[7]
port 505 nsew
rlabel metal2 s 411874 -960 411986 480 4 la_oenb[80]
port 506 nsew
rlabel metal2 s 415462 -960 415574 480 4 la_oenb[81]
port 507 nsew
rlabel metal2 s 418958 -960 419070 480 4 la_oenb[82]
port 508 nsew
rlabel metal2 s 422546 -960 422658 480 4 la_oenb[83]
port 509 nsew
rlabel metal2 s 426134 -960 426246 480 4 la_oenb[84]
port 510 nsew
rlabel metal2 s 429630 -960 429742 480 4 la_oenb[85]
port 511 nsew
rlabel metal2 s 433218 -960 433330 480 4 la_oenb[86]
port 512 nsew
rlabel metal2 s 436714 -960 436826 480 4 la_oenb[87]
port 513 nsew
rlabel metal2 s 440302 -960 440414 480 4 la_oenb[88]
port 514 nsew
rlabel metal2 s 443798 -960 443910 480 4 la_oenb[89]
port 515 nsew
rlabel metal2 s 156574 -960 156686 480 4 la_oenb[8]
port 516 nsew
rlabel metal2 s 447386 -960 447498 480 4 la_oenb[90]
port 517 nsew
rlabel metal2 s 450882 -960 450994 480 4 la_oenb[91]
port 518 nsew
rlabel metal2 s 454470 -960 454582 480 4 la_oenb[92]
port 519 nsew
rlabel metal2 s 458058 -960 458170 480 4 la_oenb[93]
port 520 nsew
rlabel metal2 s 461554 -960 461666 480 4 la_oenb[94]
port 521 nsew
rlabel metal2 s 465142 -960 465254 480 4 la_oenb[95]
port 522 nsew
rlabel metal2 s 468638 -960 468750 480 4 la_oenb[96]
port 523 nsew
rlabel metal2 s 472226 -960 472338 480 4 la_oenb[97]
port 524 nsew
rlabel metal2 s 475722 -960 475834 480 4 la_oenb[98]
port 525 nsew
rlabel metal2 s 479310 -960 479422 480 4 la_oenb[99]
port 526 nsew
rlabel metal2 s 160070 -960 160182 480 4 la_oenb[9]
port 527 nsew
rlabel metal2 s 579774 -960 579886 480 4 user_clock2
port 528 nsew
rlabel metal2 s 580970 -960 581082 480 4 user_irq[0]
port 529 nsew
rlabel metal2 s 582166 -960 582278 480 4 user_irq[1]
port 530 nsew
rlabel metal2 s 583362 -960 583474 480 4 user_irq[2]
port 531 nsew
rlabel metal5 s -2006 -934 585930 -314 4 vccd1
port 532 nsew
rlabel metal5 s -2966 2866 586890 3486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 38866 586890 39486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 74866 586890 75486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 110866 586890 111486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 146866 586890 147486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 182866 586890 183486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 218866 586890 219486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 254866 586890 255486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 290866 586890 291486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 326866 586890 327486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 362866 586890 363486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 398866 586890 399486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 434866 586890 435486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 470866 586890 471486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 506866 586890 507486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 542866 586890 543486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 578866 586890 579486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 614866 586890 615486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 650866 586890 651486 4 vccd1
port 532 nsew
rlabel metal5 s -2966 686866 586890 687486 4 vccd1
port 532 nsew
rlabel metal5 s -2006 704250 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 253794 -1894 254414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 289794 -1894 290414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 325794 -1894 326414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 361794 -1894 362414 336000 4 vccd1
port 532 nsew
rlabel metal4 s 397794 -1894 398414 336000 4 vccd1
port 532 nsew
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 532 nsew
rlabel metal4 s 585310 -934 585930 704870 4 vccd1
port 532 nsew
rlabel metal4 s 1794 -1894 2414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 37794 -1894 38414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 73794 -1894 74414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 109794 -1894 110414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 145794 -1894 146414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 181794 -1894 182414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 217794 -1894 218414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 253794 460000 254414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 289794 460000 290414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 325794 460000 326414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 361794 460000 362414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 397794 460000 398414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 433794 -1894 434414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 469794 -1894 470414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 505794 -1894 506414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 541794 -1894 542414 705830 4 vccd1
port 532 nsew
rlabel metal4 s 577794 -1894 578414 705830 4 vccd1
port 532 nsew
rlabel metal5 s -3926 -2854 587850 -2234 4 vccd2
port 533 nsew
rlabel metal5 s -4886 6586 588810 7206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 42586 588810 43206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 78586 588810 79206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 114586 588810 115206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 150586 588810 151206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 186586 588810 187206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 222586 588810 223206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 258586 588810 259206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 294586 588810 295206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 330586 588810 331206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 366586 588810 367206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 402586 588810 403206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 438586 588810 439206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 474586 588810 475206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 510586 588810 511206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 546586 588810 547206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 582586 588810 583206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 618586 588810 619206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 654586 588810 655206 4 vccd2
port 533 nsew
rlabel metal5 s -4886 690586 588810 691206 4 vccd2
port 533 nsew
rlabel metal5 s -3926 706170 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 257514 -3814 258134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 293514 -3814 294134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 329514 -3814 330134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 365514 -3814 366134 336000 4 vccd2
port 533 nsew
rlabel metal4 s 401514 -3814 402134 336000 4 vccd2
port 533 nsew
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 533 nsew
rlabel metal4 s 587230 -2854 587850 706790 4 vccd2
port 533 nsew
rlabel metal4 s 5514 -3814 6134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 41514 -3814 42134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 77514 -3814 78134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 113514 -3814 114134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 149514 -3814 150134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 185514 -3814 186134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 221514 -3814 222134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 257514 460000 258134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 293514 460000 294134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 329514 460000 330134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 365514 460000 366134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 401514 460000 402134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 437514 -3814 438134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 473514 -3814 474134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 509514 -3814 510134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 545514 -3814 546134 707750 4 vccd2
port 533 nsew
rlabel metal4 s 581514 -3814 582134 707750 4 vccd2
port 533 nsew
rlabel metal5 s -5846 -4774 589770 -4154 4 vdda1
port 534 nsew
rlabel metal5 s -6806 10306 590730 10926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 46306 590730 46926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 82306 590730 82926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 118306 590730 118926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 154306 590730 154926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 190306 590730 190926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 226306 590730 226926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 262306 590730 262926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 298306 590730 298926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 334306 590730 334926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 370306 590730 370926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 406306 590730 406926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 442306 590730 442926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 478306 590730 478926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 514306 590730 514926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 550306 590730 550926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 586306 590730 586926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 622306 590730 622926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 658306 590730 658926 4 vdda1
port 534 nsew
rlabel metal5 s -6806 694306 590730 694926 4 vdda1
port 534 nsew
rlabel metal5 s -5846 708090 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 261234 -5734 261854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 297234 -5734 297854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 333234 -5734 333854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 369234 -5734 369854 336000 4 vdda1
port 534 nsew
rlabel metal4 s 405234 -5734 405854 336000 4 vdda1
port 534 nsew
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 534 nsew
rlabel metal4 s 589150 -4774 589770 708710 4 vdda1
port 534 nsew
rlabel metal4 s 9234 -5734 9854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 45234 -5734 45854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 81234 -5734 81854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 117234 -5734 117854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 153234 -5734 153854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 189234 -5734 189854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 225234 -5734 225854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 261234 460000 261854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 297234 460000 297854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 333234 460000 333854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 369234 460000 369854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 405234 460000 405854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 441234 -5734 441854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 477234 -5734 477854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 513234 -5734 513854 709670 4 vdda1
port 534 nsew
rlabel metal4 s 549234 -5734 549854 709670 4 vdda1
port 534 nsew
rlabel metal5 s -7766 -6694 591690 -6074 4 vdda2
port 535 nsew
rlabel metal5 s -8726 14026 592650 14646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 50026 592650 50646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 86026 592650 86646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 122026 592650 122646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 158026 592650 158646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 194026 592650 194646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 230026 592650 230646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 266026 592650 266646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 302026 592650 302646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 338026 592650 338646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 374026 592650 374646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 410026 592650 410646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 446026 592650 446646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 482026 592650 482646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 518026 592650 518646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 554026 592650 554646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 590026 592650 590646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 626026 592650 626646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 662026 592650 662646 4 vdda2
port 535 nsew
rlabel metal5 s -8726 698026 592650 698646 4 vdda2
port 535 nsew
rlabel metal5 s -7766 710010 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 264954 -7654 265574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 300954 -7654 301574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 336954 -7654 337574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 372954 -7654 373574 336000 4 vdda2
port 535 nsew
rlabel metal4 s 408954 -7654 409574 336000 4 vdda2
port 535 nsew
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 535 nsew
rlabel metal4 s 591070 -6694 591690 710630 4 vdda2
port 535 nsew
rlabel metal4 s 12954 -7654 13574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 48954 -7654 49574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 84954 -7654 85574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 120954 -7654 121574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 156954 -7654 157574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 192954 -7654 193574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 228954 -7654 229574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 264954 460000 265574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 300954 460000 301574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 336954 460000 337574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 372954 460000 373574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 408954 460000 409574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 444954 -7654 445574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 480954 -7654 481574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 516954 -7654 517574 711590 4 vdda2
port 535 nsew
rlabel metal4 s 552954 -7654 553574 711590 4 vdda2
port 535 nsew
rlabel metal5 s -6806 -5734 590730 -5114 4 vssa1
port 536 nsew
rlabel metal5 s -6806 28306 590730 28926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 64306 590730 64926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 100306 590730 100926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 136306 590730 136926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 172306 590730 172926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 208306 590730 208926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 244306 590730 244926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 280306 590730 280926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 316306 590730 316926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 352306 590730 352926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 388306 590730 388926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 424306 590730 424926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 460306 590730 460926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 496306 590730 496926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 532306 590730 532926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 568306 590730 568926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 604306 590730 604926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 640306 590730 640926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 676306 590730 676926 4 vssa1
port 536 nsew
rlabel metal5 s -6806 709050 590730 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 -5734 243854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 279234 -5734 279854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 315234 -5734 315854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 351234 -5734 351854 336000 4 vssa1
port 536 nsew
rlabel metal4 s 387234 -5734 387854 336000 4 vssa1
port 536 nsew
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 536 nsew
rlabel metal4 s 27234 -5734 27854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 63234 -5734 63854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 99234 -5734 99854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 135234 -5734 135854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 171234 -5734 171854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 207234 -5734 207854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 243234 460000 243854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 279234 460000 279854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 315234 460000 315854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 351234 460000 351854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 387234 460000 387854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 423234 -5734 423854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 459234 -5734 459854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 495234 -5734 495854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 531234 -5734 531854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 567234 -5734 567854 709670 4 vssa1
port 536 nsew
rlabel metal4 s 590110 -5734 590730 709670 4 vssa1
port 536 nsew
rlabel metal5 s -8726 -7654 592650 -7034 4 vssa2
port 537 nsew
rlabel metal5 s -8726 32026 592650 32646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 68026 592650 68646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 104026 592650 104646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 140026 592650 140646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 176026 592650 176646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 212026 592650 212646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 248026 592650 248646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 284026 592650 284646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 320026 592650 320646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 356026 592650 356646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 392026 592650 392646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 428026 592650 428646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 464026 592650 464646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 500026 592650 500646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 536026 592650 536646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 572026 592650 572646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 608026 592650 608646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 644026 592650 644646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 680026 592650 680646 4 vssa2
port 537 nsew
rlabel metal5 s -8726 710970 592650 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 -7654 247574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 282954 -7654 283574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 318954 -7654 319574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 354954 -7654 355574 336000 4 vssa2
port 537 nsew
rlabel metal4 s 390954 -7654 391574 336000 4 vssa2
port 537 nsew
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 537 nsew
rlabel metal4 s 30954 -7654 31574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 66954 -7654 67574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 102954 -7654 103574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 138954 -7654 139574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 174954 -7654 175574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 210954 -7654 211574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 246954 460000 247574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 282954 460000 283574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 318954 460000 319574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 354954 460000 355574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 390954 460000 391574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 426954 -7654 427574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 462954 -7654 463574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 498954 -7654 499574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 534954 -7654 535574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 570954 -7654 571574 711590 4 vssa2
port 537 nsew
rlabel metal4 s 592030 -7654 592650 711590 4 vssa2
port 537 nsew
rlabel metal5 s -2966 -1894 586890 -1274 4 vssd1
port 538 nsew
rlabel metal5 s -2966 20866 586890 21486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 56866 586890 57486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 92866 586890 93486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 128866 586890 129486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 164866 586890 165486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 200866 586890 201486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 236866 586890 237486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 272866 586890 273486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 308866 586890 309486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 344866 586890 345486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 380866 586890 381486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 416866 586890 417486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 452866 586890 453486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 488866 586890 489486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 524866 586890 525486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 560866 586890 561486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 596866 586890 597486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 632866 586890 633486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 668866 586890 669486 4 vssd1
port 538 nsew
rlabel metal5 s -2966 705210 586890 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 -1894 236414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 271794 -1894 272414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 307794 -1894 308414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 343794 -1894 344414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 379794 -1894 380414 336000 4 vssd1
port 538 nsew
rlabel metal4 s 415794 -1894 416414 336000 4 vssd1
port 538 nsew
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 538 nsew
rlabel metal4 s 19794 -1894 20414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 55794 -1894 56414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 91794 -1894 92414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 127794 -1894 128414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 163794 -1894 164414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 199794 -1894 200414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 235794 460000 236414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 271794 460000 272414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 307794 460000 308414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 343794 460000 344414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 379794 460000 380414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 415794 460000 416414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 451794 -1894 452414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 487794 -1894 488414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 523794 -1894 524414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 559794 -1894 560414 705830 4 vssd1
port 538 nsew
rlabel metal4 s 586270 -1894 586890 705830 4 vssd1
port 538 nsew
rlabel metal5 s -4886 -3814 588810 -3194 4 vssd2
port 539 nsew
rlabel metal5 s -4886 24586 588810 25206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 60586 588810 61206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 96586 588810 97206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 132586 588810 133206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 168586 588810 169206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 204586 588810 205206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 240586 588810 241206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 276586 588810 277206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 312586 588810 313206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 348586 588810 349206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 384586 588810 385206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 420586 588810 421206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 456586 588810 457206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 492586 588810 493206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 528586 588810 529206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 564586 588810 565206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 600586 588810 601206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 636586 588810 637206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 672586 588810 673206 4 vssd2
port 539 nsew
rlabel metal5 s -4886 707130 588810 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 -3814 240134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 275514 -3814 276134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 311514 -3814 312134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 347514 -3814 348134 336000 4 vssd2
port 539 nsew
rlabel metal4 s 383514 -3814 384134 336000 4 vssd2
port 539 nsew
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 539 nsew
rlabel metal4 s 23514 -3814 24134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 59514 -3814 60134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 95514 -3814 96134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 131514 -3814 132134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 167514 -3814 168134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 203514 -3814 204134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 239514 460000 240134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 275514 460000 276134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 311514 460000 312134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 347514 460000 348134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 383514 460000 384134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 419514 -3814 420134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 455514 -3814 456134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 491514 -3814 492134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 527514 -3814 528134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 563514 -3814 564134 707750 4 vssd2
port 539 nsew
rlabel metal4 s 588190 -3814 588810 707750 4 vssd2
port 539 nsew
rlabel metal2 s 542 -960 654 480 4 wb_clk_i
port 540 nsew
rlabel metal2 s 1646 -960 1758 480 4 wb_rst_i
port 541 nsew
rlabel metal2 s 2842 -960 2954 480 4 wbs_ack_o
port 542 nsew
rlabel metal2 s 7626 -960 7738 480 4 wbs_adr_i[0]
port 543 nsew
rlabel metal2 s 47830 -960 47942 480 4 wbs_adr_i[10]
port 544 nsew
rlabel metal2 s 51326 -960 51438 480 4 wbs_adr_i[11]
port 545 nsew
rlabel metal2 s 54914 -960 55026 480 4 wbs_adr_i[12]
port 546 nsew
rlabel metal2 s 58410 -960 58522 480 4 wbs_adr_i[13]
port 547 nsew
rlabel metal2 s 61998 -960 62110 480 4 wbs_adr_i[14]
port 548 nsew
rlabel metal2 s 65494 -960 65606 480 4 wbs_adr_i[15]
port 549 nsew
rlabel metal2 s 69082 -960 69194 480 4 wbs_adr_i[16]
port 550 nsew
rlabel metal2 s 72578 -960 72690 480 4 wbs_adr_i[17]
port 551 nsew
rlabel metal2 s 76166 -960 76278 480 4 wbs_adr_i[18]
port 552 nsew
rlabel metal2 s 79662 -960 79774 480 4 wbs_adr_i[19]
port 553 nsew
rlabel metal2 s 12318 -960 12430 480 4 wbs_adr_i[1]
port 554 nsew
rlabel metal2 s 83250 -960 83362 480 4 wbs_adr_i[20]
port 555 nsew
rlabel metal2 s 86838 -960 86950 480 4 wbs_adr_i[21]
port 556 nsew
rlabel metal2 s 90334 -960 90446 480 4 wbs_adr_i[22]
port 557 nsew
rlabel metal2 s 93922 -960 94034 480 4 wbs_adr_i[23]
port 558 nsew
rlabel metal2 s 97418 -960 97530 480 4 wbs_adr_i[24]
port 559 nsew
rlabel metal2 s 101006 -960 101118 480 4 wbs_adr_i[25]
port 560 nsew
rlabel metal2 s 104502 -960 104614 480 4 wbs_adr_i[26]
port 561 nsew
rlabel metal2 s 108090 -960 108202 480 4 wbs_adr_i[27]
port 562 nsew
rlabel metal2 s 111586 -960 111698 480 4 wbs_adr_i[28]
port 563 nsew
rlabel metal2 s 115174 -960 115286 480 4 wbs_adr_i[29]
port 564 nsew
rlabel metal2 s 17010 -960 17122 480 4 wbs_adr_i[2]
port 565 nsew
rlabel metal2 s 118762 -960 118874 480 4 wbs_adr_i[30]
port 566 nsew
rlabel metal2 s 122258 -960 122370 480 4 wbs_adr_i[31]
port 567 nsew
rlabel metal2 s 21794 -960 21906 480 4 wbs_adr_i[3]
port 568 nsew
rlabel metal2 s 26486 -960 26598 480 4 wbs_adr_i[4]
port 569 nsew
rlabel metal2 s 30074 -960 30186 480 4 wbs_adr_i[5]
port 570 nsew
rlabel metal2 s 33570 -960 33682 480 4 wbs_adr_i[6]
port 571 nsew
rlabel metal2 s 37158 -960 37270 480 4 wbs_adr_i[7]
port 572 nsew
rlabel metal2 s 40654 -960 40766 480 4 wbs_adr_i[8]
port 573 nsew
rlabel metal2 s 44242 -960 44354 480 4 wbs_adr_i[9]
port 574 nsew
rlabel metal2 s 4038 -960 4150 480 4 wbs_cyc_i
port 575 nsew
rlabel metal2 s 8730 -960 8842 480 4 wbs_dat_i[0]
port 576 nsew
rlabel metal2 s 48934 -960 49046 480 4 wbs_dat_i[10]
port 577 nsew
rlabel metal2 s 52522 -960 52634 480 4 wbs_dat_i[11]
port 578 nsew
rlabel metal2 s 56018 -960 56130 480 4 wbs_dat_i[12]
port 579 nsew
rlabel metal2 s 59606 -960 59718 480 4 wbs_dat_i[13]
port 580 nsew
rlabel metal2 s 63194 -960 63306 480 4 wbs_dat_i[14]
port 581 nsew
rlabel metal2 s 66690 -960 66802 480 4 wbs_dat_i[15]
port 582 nsew
rlabel metal2 s 70278 -960 70390 480 4 wbs_dat_i[16]
port 583 nsew
rlabel metal2 s 73774 -960 73886 480 4 wbs_dat_i[17]
port 584 nsew
rlabel metal2 s 77362 -960 77474 480 4 wbs_dat_i[18]
port 585 nsew
rlabel metal2 s 80858 -960 80970 480 4 wbs_dat_i[19]
port 586 nsew
rlabel metal2 s 13514 -960 13626 480 4 wbs_dat_i[1]
port 587 nsew
rlabel metal2 s 84446 -960 84558 480 4 wbs_dat_i[20]
port 588 nsew
rlabel metal2 s 87942 -960 88054 480 4 wbs_dat_i[21]
port 589 nsew
rlabel metal2 s 91530 -960 91642 480 4 wbs_dat_i[22]
port 590 nsew
rlabel metal2 s 95118 -960 95230 480 4 wbs_dat_i[23]
port 591 nsew
rlabel metal2 s 98614 -960 98726 480 4 wbs_dat_i[24]
port 592 nsew
rlabel metal2 s 102202 -960 102314 480 4 wbs_dat_i[25]
port 593 nsew
rlabel metal2 s 105698 -960 105810 480 4 wbs_dat_i[26]
port 594 nsew
rlabel metal2 s 109286 -960 109398 480 4 wbs_dat_i[27]
port 595 nsew
rlabel metal2 s 112782 -960 112894 480 4 wbs_dat_i[28]
port 596 nsew
rlabel metal2 s 116370 -960 116482 480 4 wbs_dat_i[29]
port 597 nsew
rlabel metal2 s 18206 -960 18318 480 4 wbs_dat_i[2]
port 598 nsew
rlabel metal2 s 119866 -960 119978 480 4 wbs_dat_i[30]
port 599 nsew
rlabel metal2 s 123454 -960 123566 480 4 wbs_dat_i[31]
port 600 nsew
rlabel metal2 s 22990 -960 23102 480 4 wbs_dat_i[3]
port 601 nsew
rlabel metal2 s 27682 -960 27794 480 4 wbs_dat_i[4]
port 602 nsew
rlabel metal2 s 31270 -960 31382 480 4 wbs_dat_i[5]
port 603 nsew
rlabel metal2 s 34766 -960 34878 480 4 wbs_dat_i[6]
port 604 nsew
rlabel metal2 s 38354 -960 38466 480 4 wbs_dat_i[7]
port 605 nsew
rlabel metal2 s 41850 -960 41962 480 4 wbs_dat_i[8]
port 606 nsew
rlabel metal2 s 45438 -960 45550 480 4 wbs_dat_i[9]
port 607 nsew
rlabel metal2 s 9926 -960 10038 480 4 wbs_dat_o[0]
port 608 nsew
rlabel metal2 s 50130 -960 50242 480 4 wbs_dat_o[10]
port 609 nsew
rlabel metal2 s 53718 -960 53830 480 4 wbs_dat_o[11]
port 610 nsew
rlabel metal2 s 57214 -960 57326 480 4 wbs_dat_o[12]
port 611 nsew
rlabel metal2 s 60802 -960 60914 480 4 wbs_dat_o[13]
port 612 nsew
rlabel metal2 s 64298 -960 64410 480 4 wbs_dat_o[14]
port 613 nsew
rlabel metal2 s 67886 -960 67998 480 4 wbs_dat_o[15]
port 614 nsew
rlabel metal2 s 71474 -960 71586 480 4 wbs_dat_o[16]
port 615 nsew
rlabel metal2 s 74970 -960 75082 480 4 wbs_dat_o[17]
port 616 nsew
rlabel metal2 s 78558 -960 78670 480 4 wbs_dat_o[18]
port 617 nsew
rlabel metal2 s 82054 -960 82166 480 4 wbs_dat_o[19]
port 618 nsew
rlabel metal2 s 14710 -960 14822 480 4 wbs_dat_o[1]
port 619 nsew
rlabel metal2 s 85642 -960 85754 480 4 wbs_dat_o[20]
port 620 nsew
rlabel metal2 s 89138 -960 89250 480 4 wbs_dat_o[21]
port 621 nsew
rlabel metal2 s 92726 -960 92838 480 4 wbs_dat_o[22]
port 622 nsew
rlabel metal2 s 96222 -960 96334 480 4 wbs_dat_o[23]
port 623 nsew
rlabel metal2 s 99810 -960 99922 480 4 wbs_dat_o[24]
port 624 nsew
rlabel metal2 s 103306 -960 103418 480 4 wbs_dat_o[25]
port 625 nsew
rlabel metal2 s 106894 -960 107006 480 4 wbs_dat_o[26]
port 626 nsew
rlabel metal2 s 110482 -960 110594 480 4 wbs_dat_o[27]
port 627 nsew
rlabel metal2 s 113978 -960 114090 480 4 wbs_dat_o[28]
port 628 nsew
rlabel metal2 s 117566 -960 117678 480 4 wbs_dat_o[29]
port 629 nsew
rlabel metal2 s 19402 -960 19514 480 4 wbs_dat_o[2]
port 630 nsew
rlabel metal2 s 121062 -960 121174 480 4 wbs_dat_o[30]
port 631 nsew
rlabel metal2 s 124650 -960 124762 480 4 wbs_dat_o[31]
port 632 nsew
rlabel metal2 s 24186 -960 24298 480 4 wbs_dat_o[3]
port 633 nsew
rlabel metal2 s 28878 -960 28990 480 4 wbs_dat_o[4]
port 634 nsew
rlabel metal2 s 32374 -960 32486 480 4 wbs_dat_o[5]
port 635 nsew
rlabel metal2 s 35962 -960 36074 480 4 wbs_dat_o[6]
port 636 nsew
rlabel metal2 s 39550 -960 39662 480 4 wbs_dat_o[7]
port 637 nsew
rlabel metal2 s 43046 -960 43158 480 4 wbs_dat_o[8]
port 638 nsew
rlabel metal2 s 46634 -960 46746 480 4 wbs_dat_o[9]
port 639 nsew
rlabel metal2 s 11122 -960 11234 480 4 wbs_sel_i[0]
port 640 nsew
rlabel metal2 s 15906 -960 16018 480 4 wbs_sel_i[1]
port 641 nsew
rlabel metal2 s 20598 -960 20710 480 4 wbs_sel_i[2]
port 642 nsew
rlabel metal2 s 25290 -960 25402 480 4 wbs_sel_i[3]
port 643 nsew
rlabel metal2 s 5234 -960 5346 480 4 wbs_stb_i
port 644 nsew
rlabel metal2 s 6430 -960 6542 480 4 wbs_we_i
port 645 nsew
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
