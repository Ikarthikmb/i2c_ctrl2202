/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/rf_npn_05v5/sky130_fd_pr__rf_npn_05v5_W2p00L2p00.spice