/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/open_pdks/sources/sky130_sram_macros/sram_1rw1r_32_256_8_sky130/sram_1rw1r_32_256_8_sky130.lef