magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< poly >>
rect 12348 115 12535 148
rect 12348 81 12365 115
rect 12399 81 12433 115
rect 12467 81 12501 115
rect 12348 48 12535 81
rect 14575 115 14762 148
rect 14609 81 14643 115
rect 14677 81 14711 115
rect 14745 81 14762 115
rect 14575 48 14762 81
<< polycont >>
rect 12365 81 12399 115
rect 12433 81 12467 115
rect 12501 81 12535 115
rect 14575 81 14609 115
rect 14643 81 14677 115
rect 14711 81 14745 115
<< npolyres >>
rect 12535 48 14575 148
<< locali >>
rect 1455 4502 3752 4670
rect 4434 4498 8283 4670
rect 8788 4498 9770 4670
rect 10371 4516 11334 4670
rect 11736 4498 12770 4670
rect 14251 4498 14626 4670
rect 11902 605 11941 639
rect 11975 605 12014 639
rect 12048 605 12087 639
rect 12121 605 12160 639
rect 12194 605 12233 639
rect 12267 605 12306 639
rect 12340 605 12379 639
rect 12413 605 12452 639
rect 12486 605 12525 639
rect 12559 605 12598 639
rect 12632 605 12671 639
rect 12705 605 12744 639
rect 12778 605 12817 639
rect 12851 605 12890 639
rect 12924 605 12963 639
rect 12997 605 13036 639
rect 13070 605 13109 639
rect 13143 605 13182 639
rect 13216 605 13255 639
rect 13289 605 13328 639
rect 13362 605 13401 639
rect 13435 605 13474 639
rect 13508 605 13547 639
rect 13581 605 13620 639
rect 13654 605 13693 639
rect 13727 605 13766 639
rect 13800 605 13839 639
rect 13873 605 13913 639
rect 13947 605 13987 639
rect 14021 605 14061 639
rect 14095 605 14135 639
rect 14169 605 14209 639
rect 14243 605 14283 639
rect 14317 605 14357 639
rect 14391 605 14431 639
rect 14465 605 14505 639
rect 14539 605 14579 639
rect 14613 605 14653 639
rect 14687 605 14727 639
rect 14761 605 14801 639
rect 14835 605 14875 639
rect 11868 567 14909 605
rect 11902 533 11941 567
rect 11975 533 12014 567
rect 12048 533 12087 567
rect 12121 533 12160 567
rect 12194 533 12233 567
rect 12267 533 12306 567
rect 12340 533 12379 567
rect 12413 533 12452 567
rect 12486 533 12525 567
rect 12559 533 12598 567
rect 12632 533 12671 567
rect 12705 533 12744 567
rect 12778 533 12817 567
rect 12851 533 12890 567
rect 12924 533 12963 567
rect 12997 533 13036 567
rect 13070 533 13109 567
rect 13143 533 13182 567
rect 13216 533 13255 567
rect 13289 533 13328 567
rect 13362 533 13401 567
rect 13435 533 13474 567
rect 13508 533 13547 567
rect 13581 533 13620 567
rect 13654 533 13693 567
rect 13727 533 13766 567
rect 13800 533 13839 567
rect 13873 533 13913 567
rect 13947 533 13987 567
rect 14021 533 14061 567
rect 14095 533 14135 567
rect 14169 533 14209 567
rect 14243 533 14283 567
rect 14317 533 14357 567
rect 14391 533 14431 567
rect 14465 533 14505 567
rect 14539 533 14579 567
rect 14613 533 14653 567
rect 14687 533 14727 567
rect 14761 533 14801 567
rect 14835 533 14875 567
rect 11868 495 14909 533
rect 11902 461 11941 495
rect 11975 461 12014 495
rect 12048 461 12087 495
rect 12121 461 12160 495
rect 12194 461 12233 495
rect 12267 461 12306 495
rect 12340 461 12379 495
rect 12413 461 12452 495
rect 12486 461 12525 495
rect 12559 461 12598 495
rect 12632 461 12671 495
rect 12705 461 12744 495
rect 12778 461 12817 495
rect 12851 461 12890 495
rect 12924 461 12963 495
rect 12997 461 13036 495
rect 13070 461 13109 495
rect 13143 461 13182 495
rect 13216 461 13255 495
rect 13289 461 13328 495
rect 13362 461 13401 495
rect 13435 461 13474 495
rect 13508 461 13547 495
rect 13581 461 13620 495
rect 13654 461 13693 495
rect 13727 461 13766 495
rect 13800 461 13839 495
rect 13873 461 13913 495
rect 13947 461 13987 495
rect 14021 461 14061 495
rect 14095 461 14135 495
rect 14169 461 14209 495
rect 14243 461 14283 495
rect 14317 461 14357 495
rect 14391 461 14431 495
rect 14465 461 14505 495
rect 14539 461 14579 495
rect 14613 461 14653 495
rect 14687 461 14727 495
rect 14761 461 14801 495
rect 14835 461 14875 495
rect 14559 162 14761 168
rect 12349 115 12551 131
rect 12349 105 12365 115
rect 12349 71 12362 105
rect 12399 81 12433 115
rect 12467 105 12501 115
rect 12535 111 12551 115
rect 14559 128 14571 162
rect 14605 128 14643 162
rect 14677 128 14715 162
rect 14749 128 14761 162
rect 14559 115 14761 128
rect 12535 105 12552 111
rect 12468 81 12501 105
rect 12396 71 12434 81
rect 12468 71 12506 81
rect 12540 71 12552 105
rect 12349 65 12552 71
rect 14559 81 14575 115
rect 14609 81 14643 115
rect 14677 81 14711 115
rect 14745 81 14761 115
rect 14559 80 14761 81
rect 14559 46 14571 80
rect 14605 46 14643 80
rect 14677 46 14715 80
rect 14749 46 14761 80
rect 14559 40 14761 46
<< viali >>
rect 11868 605 11902 639
rect 11941 605 11975 639
rect 12014 605 12048 639
rect 12087 605 12121 639
rect 12160 605 12194 639
rect 12233 605 12267 639
rect 12306 605 12340 639
rect 12379 605 12413 639
rect 12452 605 12486 639
rect 12525 605 12559 639
rect 12598 605 12632 639
rect 12671 605 12705 639
rect 12744 605 12778 639
rect 12817 605 12851 639
rect 12890 605 12924 639
rect 12963 605 12997 639
rect 13036 605 13070 639
rect 13109 605 13143 639
rect 13182 605 13216 639
rect 13255 605 13289 639
rect 13328 605 13362 639
rect 13401 605 13435 639
rect 13474 605 13508 639
rect 13547 605 13581 639
rect 13620 605 13654 639
rect 13693 605 13727 639
rect 13766 605 13800 639
rect 13839 605 13873 639
rect 13913 605 13947 639
rect 13987 605 14021 639
rect 14061 605 14095 639
rect 14135 605 14169 639
rect 14209 605 14243 639
rect 14283 605 14317 639
rect 14357 605 14391 639
rect 14431 605 14465 639
rect 14505 605 14539 639
rect 14579 605 14613 639
rect 14653 605 14687 639
rect 14727 605 14761 639
rect 14801 605 14835 639
rect 14875 605 14909 639
rect 11868 533 11902 567
rect 11941 533 11975 567
rect 12014 533 12048 567
rect 12087 533 12121 567
rect 12160 533 12194 567
rect 12233 533 12267 567
rect 12306 533 12340 567
rect 12379 533 12413 567
rect 12452 533 12486 567
rect 12525 533 12559 567
rect 12598 533 12632 567
rect 12671 533 12705 567
rect 12744 533 12778 567
rect 12817 533 12851 567
rect 12890 533 12924 567
rect 12963 533 12997 567
rect 13036 533 13070 567
rect 13109 533 13143 567
rect 13182 533 13216 567
rect 13255 533 13289 567
rect 13328 533 13362 567
rect 13401 533 13435 567
rect 13474 533 13508 567
rect 13547 533 13581 567
rect 13620 533 13654 567
rect 13693 533 13727 567
rect 13766 533 13800 567
rect 13839 533 13873 567
rect 13913 533 13947 567
rect 13987 533 14021 567
rect 14061 533 14095 567
rect 14135 533 14169 567
rect 14209 533 14243 567
rect 14283 533 14317 567
rect 14357 533 14391 567
rect 14431 533 14465 567
rect 14505 533 14539 567
rect 14579 533 14613 567
rect 14653 533 14687 567
rect 14727 533 14761 567
rect 14801 533 14835 567
rect 14875 533 14909 567
rect 11868 461 11902 495
rect 11941 461 11975 495
rect 12014 461 12048 495
rect 12087 461 12121 495
rect 12160 461 12194 495
rect 12233 461 12267 495
rect 12306 461 12340 495
rect 12379 461 12413 495
rect 12452 461 12486 495
rect 12525 461 12559 495
rect 12598 461 12632 495
rect 12671 461 12705 495
rect 12744 461 12778 495
rect 12817 461 12851 495
rect 12890 461 12924 495
rect 12963 461 12997 495
rect 13036 461 13070 495
rect 13109 461 13143 495
rect 13182 461 13216 495
rect 13255 461 13289 495
rect 13328 461 13362 495
rect 13401 461 13435 495
rect 13474 461 13508 495
rect 13547 461 13581 495
rect 13620 461 13654 495
rect 13693 461 13727 495
rect 13766 461 13800 495
rect 13839 461 13873 495
rect 13913 461 13947 495
rect 13987 461 14021 495
rect 14061 461 14095 495
rect 14135 461 14169 495
rect 14209 461 14243 495
rect 14283 461 14317 495
rect 14357 461 14391 495
rect 14431 461 14465 495
rect 14505 461 14539 495
rect 14579 461 14613 495
rect 14653 461 14687 495
rect 14727 461 14761 495
rect 14801 461 14835 495
rect 14875 461 14909 495
rect 12362 81 12365 105
rect 12365 81 12396 105
rect 14571 128 14605 162
rect 14643 128 14677 162
rect 14715 128 14749 162
rect 12434 81 12467 105
rect 12467 81 12468 105
rect 12506 81 12535 105
rect 12535 81 12540 105
rect 12362 71 12396 81
rect 12434 71 12468 81
rect 12506 71 12540 81
rect 14571 46 14605 80
rect 14643 46 14677 80
rect 14715 46 14749 80
<< metal1 >>
rect 1427 1478 2325 1608
rect 2455 1478 2755 1608
rect 2885 1602 3747 1608
rect 2885 1550 3593 1602
rect 3645 1550 3671 1602
rect 3723 1550 3747 1602
rect 2885 1536 3747 1550
rect 2885 1484 3593 1536
rect 3645 1484 3671 1536
rect 3723 1484 3747 1536
rect 2885 1478 3747 1484
rect 4439 1478 5301 1608
rect 5431 1478 7285 1608
rect 7367 1556 8282 1608
rect 8334 1556 8349 1608
rect 8401 1556 8407 1608
rect 7367 1530 8407 1556
rect 7367 1478 8282 1530
rect 8334 1478 8349 1530
rect 8401 1478 8407 1530
rect 8837 1556 9132 1608
rect 9184 1556 9199 1608
rect 9251 1556 9267 1608
rect 9319 1556 9335 1608
rect 9387 1556 9403 1608
rect 9455 1556 9471 1608
rect 9523 1556 9539 1608
rect 9591 1556 9607 1608
rect 9659 1556 9675 1608
rect 9727 1556 9733 1608
rect 8837 1530 9733 1556
rect 8837 1478 9132 1530
rect 9184 1478 9199 1530
rect 9251 1478 9267 1530
rect 9319 1478 9335 1530
rect 9387 1478 9403 1530
rect 9455 1478 9471 1530
rect 9523 1478 9539 1530
rect 9591 1478 9607 1530
rect 9659 1478 9675 1530
rect 9727 1478 9733 1530
rect 10391 1556 10950 1608
rect 11002 1556 11025 1608
rect 11077 1556 11100 1608
rect 11152 1556 11175 1608
rect 11227 1556 11250 1608
rect 11302 1556 11325 1608
rect 11377 1556 11383 1608
rect 10391 1530 11383 1556
rect 10391 1478 10950 1530
rect 11002 1478 11025 1530
rect 11077 1478 11100 1530
rect 11152 1478 11175 1530
rect 11227 1478 11250 1530
rect 11302 1478 11325 1530
rect 11377 1478 11383 1530
rect 11745 1556 12273 1608
rect 12325 1556 12339 1608
rect 12391 1556 12405 1608
rect 12457 1556 12472 1608
rect 12524 1556 12539 1608
rect 12591 1556 12606 1608
rect 12658 1556 12673 1608
rect 12725 1556 12731 1608
rect 11745 1530 12731 1556
rect 11745 1478 12273 1530
rect 12325 1478 12339 1530
rect 12391 1478 12405 1530
rect 12457 1478 12472 1530
rect 12524 1478 12539 1530
rect 12591 1478 12606 1530
rect 12658 1478 12673 1530
rect 12725 1478 12731 1530
rect 13237 1601 13367 1608
rect 13237 1549 13243 1601
rect 13295 1549 13309 1601
rect 13361 1549 13367 1601
rect 13237 1537 13367 1549
rect 13237 1485 13243 1537
rect 13295 1485 13309 1537
rect 13361 1485 13367 1537
rect 13237 1478 13367 1485
rect 13667 1601 13797 1608
rect 13667 1549 13673 1601
rect 13725 1549 13739 1601
rect 13791 1549 13797 1601
rect 13667 1537 13797 1549
rect 13667 1485 13673 1537
rect 13725 1485 13739 1537
rect 13791 1485 13797 1537
rect 13667 1478 13797 1485
rect 14229 1601 14587 1608
rect 14229 1549 14235 1601
rect 14287 1549 14301 1601
rect 14353 1549 14587 1601
rect 14229 1537 14587 1549
rect 14229 1485 14235 1537
rect 14287 1485 14301 1537
rect 14353 1485 14587 1537
rect 14229 1478 14587 1485
rect 12712 661 12811 745
rect 11856 639 14921 645
rect 11856 605 11868 639
rect 11902 605 11941 639
rect 11975 605 12014 639
rect 12048 605 12087 639
rect 12121 605 12160 639
rect 12194 605 12233 639
rect 12267 605 12306 639
rect 12340 605 12379 639
rect 12413 605 12452 639
rect 12486 605 12525 639
rect 12559 605 12598 639
rect 12632 605 12671 639
rect 12705 605 12744 639
rect 12778 605 12817 639
rect 12851 605 12890 639
rect 12924 605 12963 639
rect 12997 605 13036 639
rect 13070 605 13109 639
rect 13143 605 13182 639
rect 13216 605 13255 639
rect 13289 605 13328 639
rect 13362 605 13401 639
rect 13435 605 13474 639
rect 13508 605 13547 639
rect 13581 605 13620 639
rect 13654 605 13693 639
rect 13727 605 13766 639
rect 13800 605 13839 639
rect 13873 605 13913 639
rect 13947 605 13987 639
rect 14021 605 14061 639
rect 14095 605 14135 639
rect 14169 605 14209 639
rect 14243 605 14283 639
rect 14317 605 14357 639
rect 14391 605 14431 639
rect 14465 605 14505 639
rect 14539 605 14579 639
rect 14613 605 14653 639
rect 14687 605 14727 639
rect 14761 605 14801 639
rect 14835 605 14875 639
rect 14909 605 14921 639
rect 11856 567 14921 605
rect 11856 533 11868 567
rect 11902 533 11941 567
rect 11975 533 12014 567
rect 12048 533 12087 567
rect 12121 533 12160 567
rect 12194 533 12233 567
rect 12267 533 12306 567
rect 12340 533 12379 567
rect 12413 533 12452 567
rect 12486 533 12525 567
rect 12559 533 12598 567
rect 12632 533 12671 567
rect 12705 533 12744 567
rect 12778 533 12817 567
rect 12851 533 12890 567
rect 12924 533 12963 567
rect 12997 533 13036 567
rect 13070 533 13109 567
rect 13143 533 13182 567
rect 13216 533 13255 567
rect 13289 533 13328 567
rect 13362 533 13401 567
rect 13435 533 13474 567
rect 13508 533 13547 567
rect 13581 533 13620 567
rect 13654 533 13693 567
rect 13727 533 13766 567
rect 13800 533 13839 567
rect 13873 533 13913 567
rect 13947 533 13987 567
rect 14021 533 14061 567
rect 14095 533 14135 567
rect 14169 533 14209 567
rect 14243 533 14283 567
rect 14317 533 14357 567
rect 14391 533 14431 567
rect 14465 533 14505 567
rect 14539 533 14579 567
rect 14613 533 14653 567
rect 14687 533 14727 567
rect 14761 533 14801 567
rect 14835 533 14875 567
rect 14909 533 14921 567
rect 11856 495 14921 533
rect 11856 461 11868 495
rect 11902 461 11941 495
rect 11975 461 12014 495
rect 12048 461 12087 495
rect 12121 461 12160 495
rect 12194 461 12233 495
rect 12267 461 12306 495
rect 12340 461 12379 495
rect 12413 461 12452 495
rect 12486 461 12525 495
rect 12559 461 12598 495
rect 12632 461 12671 495
rect 12705 461 12744 495
rect 12778 461 12817 495
rect 12851 461 12890 495
rect 12924 461 12963 495
rect 12997 461 13036 495
rect 13070 461 13109 495
rect 13143 461 13182 495
rect 13216 461 13255 495
rect 13289 461 13328 495
rect 13362 461 13401 495
rect 13435 461 13474 495
rect 13508 461 13547 495
rect 13581 461 13620 495
rect 13654 461 13693 495
rect 13727 461 13766 495
rect 13800 461 13839 495
rect 13873 461 13913 495
rect 13947 461 13987 495
rect 14021 461 14061 495
rect 14095 461 14135 495
rect 14169 461 14209 495
rect 14243 461 14283 495
rect 14317 461 14357 495
rect 14391 461 14431 495
rect 14465 461 14505 495
rect 14539 461 14579 495
rect 14613 461 14653 495
rect 14687 461 14727 495
rect 14761 461 14801 495
rect 14835 461 14875 495
rect 14909 461 14921 495
rect 11856 455 14921 461
rect 11936 232 11942 284
rect 11994 232 12015 284
rect 12067 232 12087 284
rect 12139 232 14108 284
rect 11936 204 14108 232
rect 11936 152 11942 204
rect 11994 152 12015 204
rect 12067 152 12087 204
rect 12139 168 14108 204
tri 14108 168 14224 284 sw
rect 12139 162 14761 168
rect 12139 152 14571 162
tri 14058 128 14082 152 ne
rect 14082 128 14571 152
rect 14605 128 14643 162
rect 14677 128 14715 162
rect 14749 128 14761 162
tri 14082 111 14099 128 ne
rect 14099 111 14761 128
rect 12003 59 12009 111
rect 12061 59 12073 111
rect 12125 105 12552 111
rect 12125 71 12362 105
rect 12396 71 12434 105
rect 12468 71 12506 105
rect 12540 71 12552 105
tri 14099 80 14130 111 ne
rect 14130 80 14761 111
rect 12125 59 12552 71
tri 14130 65 14145 80 ne
rect 14145 65 14571 80
tri 14145 59 14151 65 ne
rect 14151 59 14571 65
tri 14151 46 14164 59 ne
rect 14164 46 14571 59
rect 14605 46 14643 80
rect 14677 46 14715 80
rect 14749 46 14761 80
tri 14164 40 14170 46 ne
rect 14170 40 14761 46
tri 14471 -317 14498 -290 se
rect 14498 -317 14725 -290
tri 8008 -369 8060 -317 se
rect 8060 -369 9847 -317
rect 9899 -369 9911 -317
rect 9963 -369 11429 -317
rect 11481 -369 11493 -317
rect 11545 -369 12758 -317
rect 12810 -369 12822 -317
rect 12874 -369 13141 -317
rect 13193 -369 13207 -317
rect 13259 -369 14082 -317
rect 14134 -369 14146 -317
rect 14198 -342 14725 -317
rect 14777 -342 14789 -290
rect 14841 -342 14853 -290
rect 14905 -342 14917 -290
rect 14969 -342 14975 -290
rect 14198 -369 14550 -342
tri 14550 -369 14577 -342 nw
tri 7986 -391 8008 -369 se
rect 8008 -391 8060 -369
tri 8060 -391 8082 -369 nw
tri 14613 -391 14629 -375 se
rect 14629 -391 14905 -375
tri 7975 -402 7986 -391 se
rect 7986 -402 8049 -391
tri 8049 -402 8060 -391 nw
tri 14602 -402 14613 -391 se
rect 14613 -402 14905 -391
rect 7615 -454 7621 -402
rect 7673 -454 7685 -402
rect 7737 -454 7997 -402
tri 7997 -454 8049 -402 nw
rect 8246 -454 8252 -402
rect 8304 -454 8360 -402
rect 8412 -454 9612 -402
rect 9664 -454 9676 -402
rect 9728 -454 11194 -402
rect 11246 -454 11258 -402
rect 11310 -454 12517 -402
rect 12569 -454 12581 -402
rect 12633 -454 13845 -402
rect 13897 -454 13909 -402
rect 13961 -454 14539 -402
rect 14591 -454 14603 -402
rect 14655 -427 14905 -402
rect 14957 -427 14970 -375
rect 15022 -427 15028 -375
rect 14655 -454 14665 -427
tri 14665 -454 14692 -427 nw
tri 14689 -482 14716 -455 se
rect 14716 -461 14954 -455
rect 14716 -482 14902 -461
rect 7649 -534 9370 -482
rect 9422 -534 9434 -482
rect 9486 -534 10952 -482
rect 11004 -534 11016 -482
rect 11068 -534 12006 -482
rect 12058 -534 12070 -482
rect 12122 -534 12275 -482
rect 12327 -534 12339 -482
rect 12391 -534 13600 -482
rect 13652 -534 13664 -482
rect 13716 -534 14294 -482
rect 14346 -534 14358 -482
rect 14410 -507 14902 -482
rect 14410 -534 14753 -507
tri 14753 -534 14780 -507 nw
tri 14858 -534 14885 -507 ne
rect 14885 -513 14902 -507
rect 14885 -525 14954 -513
rect 14885 -534 14902 -525
tri 14885 -551 14902 -534 ne
rect 14902 -583 14954 -577
<< via1 >>
rect 3593 1550 3645 1602
rect 3671 1550 3723 1602
rect 3593 1484 3645 1536
rect 3671 1484 3723 1536
rect 8282 1556 8334 1608
rect 8349 1556 8401 1608
rect 8282 1478 8334 1530
rect 8349 1478 8401 1530
rect 9132 1556 9184 1608
rect 9199 1556 9251 1608
rect 9267 1556 9319 1608
rect 9335 1556 9387 1608
rect 9403 1556 9455 1608
rect 9471 1556 9523 1608
rect 9539 1556 9591 1608
rect 9607 1556 9659 1608
rect 9675 1556 9727 1608
rect 9132 1478 9184 1530
rect 9199 1478 9251 1530
rect 9267 1478 9319 1530
rect 9335 1478 9387 1530
rect 9403 1478 9455 1530
rect 9471 1478 9523 1530
rect 9539 1478 9591 1530
rect 9607 1478 9659 1530
rect 9675 1478 9727 1530
rect 10950 1556 11002 1608
rect 11025 1556 11077 1608
rect 11100 1556 11152 1608
rect 11175 1556 11227 1608
rect 11250 1556 11302 1608
rect 11325 1556 11377 1608
rect 10950 1478 11002 1530
rect 11025 1478 11077 1530
rect 11100 1478 11152 1530
rect 11175 1478 11227 1530
rect 11250 1478 11302 1530
rect 11325 1478 11377 1530
rect 12273 1556 12325 1608
rect 12339 1556 12391 1608
rect 12405 1556 12457 1608
rect 12472 1556 12524 1608
rect 12539 1556 12591 1608
rect 12606 1556 12658 1608
rect 12673 1556 12725 1608
rect 12273 1478 12325 1530
rect 12339 1478 12391 1530
rect 12405 1478 12457 1530
rect 12472 1478 12524 1530
rect 12539 1478 12591 1530
rect 12606 1478 12658 1530
rect 12673 1478 12725 1530
rect 13243 1549 13295 1601
rect 13309 1549 13361 1601
rect 13243 1485 13295 1537
rect 13309 1485 13361 1537
rect 13673 1549 13725 1601
rect 13739 1549 13791 1601
rect 13673 1485 13725 1537
rect 13739 1485 13791 1537
rect 14235 1549 14287 1601
rect 14301 1549 14353 1601
rect 14235 1485 14287 1537
rect 14301 1485 14353 1537
rect 11942 232 11994 284
rect 12015 232 12067 284
rect 12087 232 12139 284
rect 11942 152 11994 204
rect 12015 152 12067 204
rect 12087 152 12139 204
rect 12009 59 12061 111
rect 12073 59 12125 111
rect 9847 -369 9899 -317
rect 9911 -369 9963 -317
rect 11429 -369 11481 -317
rect 11493 -369 11545 -317
rect 12758 -369 12810 -317
rect 12822 -369 12874 -317
rect 13141 -369 13193 -317
rect 13207 -369 13259 -317
rect 14082 -369 14134 -317
rect 14146 -369 14198 -317
rect 14725 -342 14777 -290
rect 14789 -342 14841 -290
rect 14853 -342 14905 -290
rect 14917 -342 14969 -290
rect 7621 -454 7673 -402
rect 7685 -454 7737 -402
rect 8252 -454 8304 -402
rect 8360 -454 8412 -402
rect 9612 -454 9664 -402
rect 9676 -454 9728 -402
rect 11194 -454 11246 -402
rect 11258 -454 11310 -402
rect 12517 -454 12569 -402
rect 12581 -454 12633 -402
rect 13845 -454 13897 -402
rect 13909 -454 13961 -402
rect 14539 -454 14591 -402
rect 14603 -454 14655 -402
rect 14905 -427 14957 -375
rect 14970 -427 15022 -375
rect 9370 -534 9422 -482
rect 9434 -534 9486 -482
rect 10952 -534 11004 -482
rect 11016 -534 11068 -482
rect 12006 -534 12058 -482
rect 12070 -534 12122 -482
rect 12275 -534 12327 -482
rect 12339 -534 12391 -482
rect 13600 -534 13652 -482
rect 13664 -534 13716 -482
rect 14294 -534 14346 -482
rect 14358 -534 14410 -482
rect 14902 -513 14954 -461
rect 14902 -577 14954 -525
<< metal2 >>
rect 3593 1602 3723 1608
rect 3645 1550 3671 1602
rect 3593 1536 3723 1550
rect 3645 1484 3671 1536
rect 3593 -328 3723 1484
rect 8246 1556 8282 1608
rect 8334 1556 8349 1608
rect 8401 1556 8418 1608
rect 8246 1530 8418 1556
rect 8246 1478 8282 1530
rect 8334 1478 8349 1530
rect 8401 1478 8418 1530
tri 3593 -369 3634 -328 ne
rect 3634 -369 3723 -328
tri 3723 -369 3771 -321 sw
tri 3634 -375 3640 -369 ne
rect 3640 -375 3771 -369
tri 3771 -375 3777 -369 sw
tri 3640 -402 3667 -375 ne
rect 3667 -402 3777 -375
tri 3777 -402 3804 -375 sw
rect 8246 -402 8418 1478
rect 9126 1556 9132 1608
rect 9184 1556 9199 1608
rect 9251 1556 9267 1608
rect 9319 1556 9335 1608
rect 9387 1556 9403 1608
rect 9455 1556 9471 1608
rect 9523 1556 9539 1608
rect 9591 1556 9607 1608
rect 9659 1556 9675 1608
rect 9727 1556 9733 1608
rect 9126 1530 9733 1556
rect 9126 1478 9132 1530
rect 9184 1478 9199 1530
rect 9251 1478 9267 1530
rect 9319 1478 9335 1530
rect 9387 1478 9403 1530
rect 9455 1478 9471 1530
rect 9523 1478 9539 1530
rect 9591 1478 9607 1530
rect 9659 1478 9675 1530
rect 9727 1478 9733 1530
rect 9126 1457 9697 1478
tri 9126 1442 9141 1457 ne
rect 9141 1442 9697 1457
tri 9697 1442 9733 1478 nw
rect 10944 1556 10950 1608
rect 11002 1556 11025 1608
rect 11077 1556 11100 1608
rect 11152 1556 11175 1608
rect 11227 1556 11250 1608
rect 11302 1556 11325 1608
rect 11377 1556 11383 1608
rect 10944 1530 11383 1556
rect 10944 1478 10950 1530
rect 11002 1478 11025 1530
rect 11077 1478 11100 1530
rect 11152 1478 11175 1530
rect 11227 1478 11250 1530
rect 11302 1478 11325 1530
rect 11377 1478 11383 1530
tri 9141 1221 9362 1442 ne
rect 9362 284 9697 1442
tri 9697 284 9945 532 sw
rect 10944 284 11383 1478
rect 12267 1556 12273 1608
rect 12325 1556 12339 1608
rect 12391 1556 12405 1608
rect 12457 1556 12472 1608
rect 12524 1556 12539 1608
rect 12591 1556 12606 1608
rect 12658 1556 12673 1608
rect 12725 1556 12731 1608
tri 13198 1601 13205 1608 se
rect 13205 1601 13367 1608
rect 12267 1530 12731 1556
tri 13146 1549 13198 1601 se
rect 13198 1549 13243 1601
rect 13295 1549 13309 1601
rect 13361 1549 13367 1601
rect 12267 1478 12273 1530
rect 12325 1478 12339 1530
rect 12391 1478 12405 1530
rect 12457 1478 12472 1530
rect 12524 1478 12539 1530
rect 12591 1478 12606 1530
rect 12658 1478 12673 1530
rect 12725 1478 12731 1530
tri 11383 284 11527 428 sw
rect 11931 351 11940 407
rect 11996 351 12064 407
rect 12120 351 12145 407
rect 11931 321 12145 351
rect 9362 260 9945 284
tri 9945 260 9969 284 sw
rect 9362 146 9969 260
rect 9362 94 9492 146
tri 9492 114 9524 146 nw
tri 9571 114 9603 146 ne
rect 9603 114 9734 146
tri 9734 114 9766 146 nw
tri 9805 114 9837 146 ne
rect 9837 114 9969 146
tri 9603 113 9604 114 ne
rect 9363 92 9491 93
rect 9604 94 9734 114
tri 9837 112 9839 114 ne
rect 9605 92 9733 93
rect 9839 94 9969 114
rect 9840 92 9968 93
rect 10944 260 11527 284
tri 11527 260 11551 284 sw
rect 10944 146 11551 260
rect 11931 265 11940 321
rect 11996 284 12064 321
rect 12120 284 12145 321
rect 11996 265 12015 284
rect 11931 232 11942 265
rect 11994 232 12015 265
rect 12067 232 12087 265
rect 12139 232 12145 284
rect 11931 204 12145 232
rect 11931 152 11942 204
rect 11994 152 12015 204
rect 12067 152 12087 204
rect 12139 152 12145 204
rect 12267 189 12731 1478
tri 13135 1538 13146 1549 se
rect 13146 1538 13367 1549
rect 13135 1537 13367 1538
rect 13135 1485 13243 1537
rect 13295 1485 13309 1537
rect 13361 1485 13367 1537
rect 13135 1478 13367 1485
rect 13667 1601 13797 1608
rect 13667 1549 13673 1601
rect 13725 1549 13739 1601
rect 13791 1549 13797 1601
rect 13667 1537 13797 1549
rect 13667 1485 13673 1537
rect 13725 1485 13739 1537
rect 13791 1485 13797 1537
tri 12731 189 12880 338 sw
rect 10944 94 11074 146
tri 11074 114 11106 146 nw
tri 11153 114 11185 146 ne
rect 11185 114 11316 146
tri 11316 114 11348 146 nw
tri 11387 114 11419 146 ne
rect 11419 114 11551 146
tri 11185 113 11186 114 ne
rect 10945 92 11073 93
rect 11186 94 11316 114
tri 11419 113 11420 114 ne
rect 11420 113 11551 114
tri 11420 112 11421 113 ne
rect 11187 92 11315 93
rect 11421 94 11551 113
rect 11422 92 11550 93
rect 9839 -208 9969 92
rect 11186 -208 11316 92
rect 12003 59 12009 111
rect 12061 59 12073 111
rect 12125 59 12131 111
tri 12003 41 12021 59 ne
rect 12021 41 12113 59
tri 12113 41 12131 59 nw
rect 12267 75 12880 189
tri 12021 21 12041 41 ne
tri 3667 -454 3719 -402 ne
rect 3719 -454 7621 -402
rect 7673 -454 7685 -402
rect 7737 -454 7743 -402
rect 8246 -454 8252 -402
rect 8304 -454 8360 -402
rect 8412 -454 8418 -402
rect 9363 -209 9491 -208
rect 9362 -482 9492 -210
rect 9605 -209 9733 -208
rect 9604 -402 9734 -210
rect 9840 -209 9968 -208
rect 9839 -317 9969 -210
rect 9839 -369 9847 -317
rect 9899 -369 9911 -317
rect 9963 -369 9969 -317
rect 10945 -209 11073 -208
rect 9604 -454 9612 -402
rect 9664 -454 9676 -402
rect 9728 -454 9734 -402
rect 9362 -534 9370 -482
rect 9422 -534 9434 -482
rect 9486 -534 9492 -482
rect 10944 -482 11074 -210
rect 11187 -209 11315 -208
rect 11186 -402 11316 -210
rect 11422 -209 11550 -208
rect 11421 -317 11551 -210
rect 11421 -369 11429 -317
rect 11481 -369 11493 -317
rect 11545 -369 11551 -317
rect 11186 -454 11194 -402
rect 11246 -454 11258 -402
rect 11310 -454 11316 -402
tri 12028 -454 12041 -441 se
rect 12041 -454 12093 41
tri 12093 21 12113 41 nw
rect 12267 23 12397 75
tri 12397 41 12431 75 nw
tri 12475 41 12509 75 ne
rect 12268 21 12396 22
rect 12509 23 12639 75
tri 12639 41 12673 75 nw
tri 12716 41 12750 75 ne
rect 12510 21 12638 22
rect 12750 23 12880 75
rect 12751 21 12879 22
rect 12267 -279 12397 21
rect 12268 -280 12396 -279
tri 12093 -454 12100 -447 sw
tri 12021 -461 12028 -454 se
rect 12028 -461 12100 -454
tri 12100 -461 12107 -454 sw
rect 10944 -534 10952 -482
rect 11004 -534 11016 -482
rect 11068 -534 11074 -482
tri 12000 -482 12021 -461 se
rect 12021 -482 12107 -461
tri 12107 -482 12128 -461 sw
rect 12000 -534 12006 -482
rect 12058 -534 12070 -482
rect 12122 -534 12128 -482
rect 12267 -482 12397 -281
rect 12510 -280 12638 -279
rect 12509 -402 12639 -281
rect 12751 -280 12879 -279
rect 12750 -317 12880 -281
rect 12750 -369 12758 -317
rect 12810 -369 12822 -317
rect 12874 -369 12880 -317
rect 13135 -317 13265 1478
tri 13265 1408 13335 1478 nw
tri 13592 1147 13667 1222 se
rect 13667 1147 13797 1485
rect 14229 1601 14359 1608
rect 14229 1549 14235 1601
rect 14287 1549 14301 1601
rect 14353 1549 14359 1601
rect 14229 1537 14359 1549
rect 14229 1485 14235 1537
rect 14287 1485 14301 1537
rect 14353 1485 14359 1537
rect 14229 1357 14359 1485
tri 14229 1328 14258 1357 ne
rect 14258 1328 14359 1357
tri 14359 1328 14442 1411 sw
tri 14258 1300 14286 1328 ne
rect 13592 1126 13797 1147
tri 13797 1126 13893 1222 sw
rect 14286 1126 14442 1328
tri 14442 1126 14563 1247 sw
rect 13592 1012 14204 1126
rect 13592 960 13722 1012
tri 13722 978 13756 1012 nw
tri 13803 978 13837 1012 ne
rect 13593 958 13721 959
rect 13837 960 13967 1012
tri 13967 978 14001 1012 nw
tri 14040 978 14074 1012 ne
rect 13838 958 13966 959
rect 14074 960 14204 1012
rect 14075 958 14203 959
rect 14286 1012 14898 1126
rect 14286 960 14416 1012
tri 14416 978 14450 1012 nw
tri 14497 978 14531 1012 ne
rect 14287 958 14415 959
rect 14531 960 14661 1012
tri 14661 978 14695 1012 nw
tri 14734 978 14768 1012 ne
rect 14532 958 14660 959
rect 14768 960 14898 1012
rect 14769 958 14897 959
rect 13837 658 13967 958
rect 14286 658 14416 958
rect 13135 -369 13141 -317
rect 13193 -369 13207 -317
rect 13259 -369 13265 -317
rect 13593 657 13721 658
rect 12509 -454 12517 -402
rect 12569 -454 12581 -402
rect 12633 -454 12639 -402
rect 12267 -534 12275 -482
rect 12327 -534 12339 -482
rect 12391 -534 12397 -482
rect 13592 -482 13722 656
rect 13838 657 13966 658
rect 13837 -402 13967 656
rect 14075 657 14203 658
rect 14074 -317 14204 656
rect 14074 -369 14082 -317
rect 14134 -369 14146 -317
rect 14198 -369 14204 -317
rect 14287 657 14415 658
rect 13837 -454 13845 -402
rect 13897 -454 13909 -402
rect 13961 -454 13967 -402
rect 13592 -534 13600 -482
rect 13652 -534 13664 -482
rect 13716 -534 13722 -482
rect 14286 -482 14416 656
rect 14532 657 14660 658
rect 14531 -402 14661 656
rect 14769 657 14897 658
tri 14740 -262 14768 -234 se
rect 14768 -262 14898 656
tri 14712 -290 14740 -262 se
rect 14740 -290 14898 -262
tri 14898 -290 14972 -216 sw
rect 14712 -342 14725 -290
rect 14777 -342 14789 -290
rect 14841 -342 14853 -290
rect 14905 -342 14917 -290
rect 14969 -342 14975 -290
rect 14531 -454 14539 -402
rect 14591 -454 14603 -402
rect 14655 -454 14661 -402
rect 14899 -427 14905 -375
rect 14957 -427 14970 -375
rect 15022 -427 15028 -375
rect 14286 -534 14294 -482
rect 14346 -534 14358 -482
rect 14410 -534 14416 -482
rect 14902 -461 14954 -455
rect 14902 -525 14954 -513
rect 14902 -583 14954 -577
<< rmetal2 >>
rect 9362 93 9492 94
rect 9362 92 9363 93
rect 9491 92 9492 93
rect 9604 93 9734 94
rect 9604 92 9605 93
rect 9733 92 9734 93
rect 9839 93 9969 94
rect 9839 92 9840 93
rect 9968 92 9969 93
rect 10944 93 11074 94
rect 10944 92 10945 93
rect 11073 92 11074 93
rect 11186 93 11316 94
rect 11186 92 11187 93
rect 11315 92 11316 93
rect 11421 93 11551 94
rect 11421 92 11422 93
rect 11550 92 11551 93
rect 9362 -209 9363 -208
rect 9491 -209 9492 -208
rect 9362 -210 9492 -209
rect 9604 -209 9605 -208
rect 9733 -209 9734 -208
rect 9604 -210 9734 -209
rect 9839 -209 9840 -208
rect 9968 -209 9969 -208
rect 9839 -210 9969 -209
rect 10944 -209 10945 -208
rect 11073 -209 11074 -208
rect 10944 -210 11074 -209
rect 11186 -209 11187 -208
rect 11315 -209 11316 -208
rect 11186 -210 11316 -209
rect 11421 -209 11422 -208
rect 11550 -209 11551 -208
rect 11421 -210 11551 -209
rect 12267 22 12397 23
rect 12267 21 12268 22
rect 12396 21 12397 22
rect 12509 22 12639 23
rect 12509 21 12510 22
rect 12638 21 12639 22
rect 12750 22 12880 23
rect 12750 21 12751 22
rect 12879 21 12880 22
rect 12267 -280 12268 -279
rect 12396 -280 12397 -279
rect 12267 -281 12397 -280
rect 12509 -280 12510 -279
rect 12638 -280 12639 -279
rect 12509 -281 12639 -280
rect 12750 -280 12751 -279
rect 12879 -280 12880 -279
rect 12750 -281 12880 -280
rect 13592 959 13722 960
rect 13592 958 13593 959
rect 13721 958 13722 959
rect 13837 959 13967 960
rect 13837 958 13838 959
rect 13966 958 13967 959
rect 14074 959 14204 960
rect 14074 958 14075 959
rect 14203 958 14204 959
rect 14286 959 14416 960
rect 14286 958 14287 959
rect 14415 958 14416 959
rect 14531 959 14661 960
rect 14531 958 14532 959
rect 14660 958 14661 959
rect 14768 959 14898 960
rect 14768 958 14769 959
rect 14897 958 14898 959
rect 13592 657 13593 658
rect 13721 657 13722 658
rect 13592 656 13722 657
rect 13837 657 13838 658
rect 13966 657 13967 658
rect 13837 656 13967 657
rect 14074 657 14075 658
rect 14203 657 14204 658
rect 14074 656 14204 657
rect 14286 657 14287 658
rect 14415 657 14416 658
rect 14286 656 14416 657
rect 14531 657 14532 658
rect 14660 657 14661 658
rect 14531 656 14661 657
rect 14768 657 14769 658
rect 14897 657 14898 658
rect 14768 656 14898 657
<< via2 >>
rect 11940 351 11996 407
rect 12064 351 12120 407
rect 11940 284 11996 321
rect 12064 284 12120 321
rect 11940 265 11942 284
rect 11942 265 11994 284
rect 11994 265 11996 284
rect 12064 265 12067 284
rect 12067 265 12087 284
rect 12087 265 12120 284
<< metal3 >>
rect 11935 407 12125 412
rect 11935 351 11940 407
rect 11996 351 12064 407
rect 12120 351 12125 407
rect 11935 321 12125 351
rect 11935 265 11940 321
rect 11996 265 12064 321
rect 12120 265 12125 321
rect 11935 260 12125 265
use sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2  sky130_fd_io__pfet_con_diff_wo_abt_270_xres4v2_0
timestamp 1644511149
transform 1 0 457 0 1 346
box 15 283 15097 5150
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_0
timestamp 1644511149
transform 0 1 14074 1 0 604
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_1
timestamp 1644511149
transform 0 1 14531 1 0 604
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_2
timestamp 1644511149
transform 0 1 13592 1 0 604
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_3
timestamp 1644511149
transform 0 1 9362 1 0 -262
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_4
timestamp 1644511149
transform 0 1 9604 1 0 -262
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_5
timestamp 1644511149
transform 0 1 11421 1 0 -262
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_6
timestamp 1644511149
transform 0 1 10944 1 0 -262
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_7
timestamp 1644511149
transform 0 1 12750 1 0 -333
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_8
timestamp 1644511149
transform 0 1 14768 1 0 604
box 0 24 408 28
use sky130_fd_io__tk_em2o_cdns_55959141808653  sky130_fd_io__tk_em2o_cdns_55959141808653_9
timestamp 1644511149
transform 0 1 12509 1 0 -333
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_0
timestamp 1644511149
transform 0 1 14286 1 0 604
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_1
timestamp 1644511149
transform 0 1 13837 1 0 604
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_2
timestamp 1644511149
transform 0 1 9839 1 0 -262
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_3
timestamp 1644511149
transform 0 1 11186 1 0 -262
box 0 24 408 28
use sky130_fd_io__tk_em2s_cdns_55959141808652  sky130_fd_io__tk_em2s_cdns_55959141808652_4
timestamp 1644511149
transform 0 1 12267 1 0 -333
box 0 24 408 28
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_0
timestamp 1644511149
transform 1 0 12535 0 1 48
box 15 17 2025 18
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_0
timestamp 1644511149
transform -1 0 14660 0 -1 98
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_1
timestamp 1644511149
transform 1 0 12450 0 -1 98
box 0 0 1 1
<< labels >>
flabel comment s 13504 107 13504 107 0 FreeSans 440 0 0 0 LEAKER
flabel metal1 s 10483 -454 10635 -402 0 FreeSans 400 180 0 0 PU_H_N[3]
port 1 nsew
flabel metal1 s 10299 -369 10384 -317 0 FreeSans 400 180 0 0 PU_H_N[2]
port 2 nsew
flabel metal1 s 9905 -508 9905 -508 0 FreeSans 400 180 0 0 TIE_HI_ESD
port 3 nsew
flabel metal1 s 12712 661 12811 745 3 FreeSans 520 0 0 0 VNB
port 4 nsew
<< properties >>
string GDS_END 30610258
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 30581732
<< end >>
