magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< dnwell >>
rect 214 214 1978 2378
<< nwell >>
rect 134 2098 2058 2458
rect 134 494 494 2098
rect 1698 494 2058 2098
rect 134 134 2058 494
<< pwell >>
rect 0 2458 2192 2592
rect 0 134 134 2458
rect 628 628 1564 1964
rect 2058 134 2192 2458
rect 0 0 2192 134
<< ndiff >>
rect 896 1653 1296 1696
rect 896 939 909 1653
rect 1283 939 1296 1653
rect 896 896 1296 939
<< ndiffc >>
rect 909 939 1283 1653
<< psubdiff >>
rect 26 2542 2166 2566
rect 26 2508 50 2542
rect 84 2508 127 2542
rect 161 2508 195 2542
rect 229 2508 263 2542
rect 297 2508 331 2542
rect 365 2508 399 2542
rect 433 2508 467 2542
rect 501 2508 535 2542
rect 569 2508 603 2542
rect 637 2508 671 2542
rect 705 2508 739 2542
rect 773 2508 807 2542
rect 841 2508 875 2542
rect 909 2508 943 2542
rect 977 2508 1011 2542
rect 1045 2508 1079 2542
rect 1113 2508 1147 2542
rect 1181 2508 1215 2542
rect 1249 2508 1283 2542
rect 1317 2508 1351 2542
rect 1385 2508 1419 2542
rect 1453 2508 1487 2542
rect 1521 2508 1555 2542
rect 1589 2508 1623 2542
rect 1657 2508 1691 2542
rect 1725 2508 1759 2542
rect 1793 2508 1827 2542
rect 1861 2508 1895 2542
rect 1929 2508 1963 2542
rect 1997 2508 2031 2542
rect 2065 2508 2108 2542
rect 2142 2508 2166 2542
rect 26 2484 2166 2508
rect 26 2469 108 2484
rect 26 2435 50 2469
rect 84 2435 108 2469
rect 26 2401 108 2435
rect 26 2367 50 2401
rect 84 2367 108 2401
rect 26 2333 108 2367
rect 2084 2469 2166 2484
rect 2084 2435 2108 2469
rect 2142 2435 2166 2469
rect 2084 2401 2166 2435
rect 2084 2367 2108 2401
rect 2142 2367 2166 2401
rect 26 2299 50 2333
rect 84 2299 108 2333
rect 26 2265 108 2299
rect 26 2231 50 2265
rect 84 2231 108 2265
rect 26 2197 108 2231
rect 26 2163 50 2197
rect 84 2163 108 2197
rect 26 2129 108 2163
rect 26 2095 50 2129
rect 84 2095 108 2129
rect 26 2061 108 2095
rect 26 2027 50 2061
rect 84 2027 108 2061
rect 26 1993 108 2027
rect 26 1959 50 1993
rect 84 1959 108 1993
rect 26 1925 108 1959
rect 26 1891 50 1925
rect 84 1891 108 1925
rect 26 1857 108 1891
rect 26 1823 50 1857
rect 84 1823 108 1857
rect 26 1789 108 1823
rect 26 1755 50 1789
rect 84 1755 108 1789
rect 26 1721 108 1755
rect 26 1687 50 1721
rect 84 1687 108 1721
rect 26 1653 108 1687
rect 26 1619 50 1653
rect 84 1619 108 1653
rect 26 1585 108 1619
rect 26 1551 50 1585
rect 84 1551 108 1585
rect 26 1517 108 1551
rect 26 1483 50 1517
rect 84 1483 108 1517
rect 26 1449 108 1483
rect 26 1415 50 1449
rect 84 1415 108 1449
rect 26 1381 108 1415
rect 26 1347 50 1381
rect 84 1347 108 1381
rect 26 1313 108 1347
rect 26 1279 50 1313
rect 84 1279 108 1313
rect 26 1245 108 1279
rect 26 1211 50 1245
rect 84 1211 108 1245
rect 26 1177 108 1211
rect 26 1143 50 1177
rect 84 1143 108 1177
rect 26 1109 108 1143
rect 26 1075 50 1109
rect 84 1075 108 1109
rect 26 1041 108 1075
rect 26 1007 50 1041
rect 84 1007 108 1041
rect 26 973 108 1007
rect 26 939 50 973
rect 84 939 108 973
rect 26 905 108 939
rect 26 871 50 905
rect 84 871 108 905
rect 26 837 108 871
rect 26 803 50 837
rect 84 803 108 837
rect 26 769 108 803
rect 26 735 50 769
rect 84 735 108 769
rect 26 701 108 735
rect 26 667 50 701
rect 84 667 108 701
rect 26 633 108 667
rect 26 599 50 633
rect 84 599 108 633
rect 26 565 108 599
rect 26 531 50 565
rect 84 531 108 565
rect 26 497 108 531
rect 26 463 50 497
rect 84 463 108 497
rect 26 429 108 463
rect 26 395 50 429
rect 84 395 108 429
rect 26 361 108 395
rect 26 327 50 361
rect 84 327 108 361
rect 26 293 108 327
rect 26 259 50 293
rect 84 259 108 293
rect 26 225 108 259
rect 654 1914 1538 1938
rect 654 1880 678 1914
rect 712 1880 773 1914
rect 807 1880 841 1914
rect 875 1880 909 1914
rect 943 1880 977 1914
rect 1011 1880 1045 1914
rect 1079 1880 1113 1914
rect 1147 1880 1181 1914
rect 1215 1880 1249 1914
rect 1283 1880 1317 1914
rect 1351 1880 1385 1914
rect 1419 1880 1480 1914
rect 1514 1880 1538 1914
rect 654 1856 1538 1880
rect 654 1823 736 1856
rect 654 1789 678 1823
rect 712 1789 736 1823
rect 654 1755 736 1789
rect 654 1721 678 1755
rect 712 1721 736 1755
rect 654 1687 736 1721
rect 1456 1823 1538 1856
rect 1456 1789 1480 1823
rect 1514 1789 1538 1823
rect 1456 1755 1538 1789
rect 1456 1721 1480 1755
rect 1514 1721 1538 1755
rect 654 1653 678 1687
rect 712 1653 736 1687
rect 654 1619 736 1653
rect 654 1585 678 1619
rect 712 1585 736 1619
rect 654 1551 736 1585
rect 654 1517 678 1551
rect 712 1517 736 1551
rect 654 1483 736 1517
rect 654 1449 678 1483
rect 712 1449 736 1483
rect 654 1415 736 1449
rect 654 1381 678 1415
rect 712 1381 736 1415
rect 654 1347 736 1381
rect 654 1313 678 1347
rect 712 1313 736 1347
rect 654 1279 736 1313
rect 654 1245 678 1279
rect 712 1245 736 1279
rect 654 1211 736 1245
rect 654 1177 678 1211
rect 712 1177 736 1211
rect 654 1143 736 1177
rect 654 1109 678 1143
rect 712 1109 736 1143
rect 654 1075 736 1109
rect 654 1041 678 1075
rect 712 1041 736 1075
rect 654 1007 736 1041
rect 654 973 678 1007
rect 712 973 736 1007
rect 654 939 736 973
rect 654 905 678 939
rect 712 905 736 939
rect 654 871 736 905
rect 1456 1687 1538 1721
rect 1456 1653 1480 1687
rect 1514 1653 1538 1687
rect 1456 1619 1538 1653
rect 1456 1585 1480 1619
rect 1514 1585 1538 1619
rect 1456 1551 1538 1585
rect 1456 1517 1480 1551
rect 1514 1517 1538 1551
rect 1456 1483 1538 1517
rect 1456 1449 1480 1483
rect 1514 1449 1538 1483
rect 1456 1415 1538 1449
rect 1456 1381 1480 1415
rect 1514 1381 1538 1415
rect 1456 1347 1538 1381
rect 1456 1313 1480 1347
rect 1514 1313 1538 1347
rect 1456 1279 1538 1313
rect 1456 1245 1480 1279
rect 1514 1245 1538 1279
rect 1456 1211 1538 1245
rect 1456 1177 1480 1211
rect 1514 1177 1538 1211
rect 1456 1143 1538 1177
rect 1456 1109 1480 1143
rect 1514 1109 1538 1143
rect 1456 1075 1538 1109
rect 1456 1041 1480 1075
rect 1514 1041 1538 1075
rect 1456 1007 1538 1041
rect 1456 973 1480 1007
rect 1514 973 1538 1007
rect 1456 939 1538 973
rect 1456 905 1480 939
rect 1514 905 1538 939
rect 654 837 678 871
rect 712 837 736 871
rect 654 803 736 837
rect 654 769 678 803
rect 712 769 736 803
rect 654 736 736 769
rect 1456 871 1538 905
rect 1456 837 1480 871
rect 1514 837 1538 871
rect 1456 803 1538 837
rect 1456 769 1480 803
rect 1514 769 1538 803
rect 1456 736 1538 769
rect 654 712 1538 736
rect 654 678 678 712
rect 712 678 773 712
rect 807 678 841 712
rect 875 678 909 712
rect 943 678 977 712
rect 1011 678 1045 712
rect 1079 678 1113 712
rect 1147 678 1181 712
rect 1215 678 1249 712
rect 1283 678 1317 712
rect 1351 678 1385 712
rect 1419 678 1480 712
rect 1514 678 1538 712
rect 654 654 1538 678
rect 2084 2333 2166 2367
rect 2084 2299 2108 2333
rect 2142 2299 2166 2333
rect 2084 2265 2166 2299
rect 2084 2231 2108 2265
rect 2142 2231 2166 2265
rect 2084 2197 2166 2231
rect 2084 2163 2108 2197
rect 2142 2163 2166 2197
rect 2084 2129 2166 2163
rect 2084 2095 2108 2129
rect 2142 2095 2166 2129
rect 2084 2061 2166 2095
rect 2084 2027 2108 2061
rect 2142 2027 2166 2061
rect 2084 1993 2166 2027
rect 2084 1959 2108 1993
rect 2142 1959 2166 1993
rect 2084 1925 2166 1959
rect 2084 1891 2108 1925
rect 2142 1891 2166 1925
rect 2084 1857 2166 1891
rect 2084 1823 2108 1857
rect 2142 1823 2166 1857
rect 2084 1789 2166 1823
rect 2084 1755 2108 1789
rect 2142 1755 2166 1789
rect 2084 1721 2166 1755
rect 2084 1687 2108 1721
rect 2142 1687 2166 1721
rect 2084 1653 2166 1687
rect 2084 1619 2108 1653
rect 2142 1619 2166 1653
rect 2084 1585 2166 1619
rect 2084 1551 2108 1585
rect 2142 1551 2166 1585
rect 2084 1517 2166 1551
rect 2084 1483 2108 1517
rect 2142 1483 2166 1517
rect 2084 1449 2166 1483
rect 2084 1415 2108 1449
rect 2142 1415 2166 1449
rect 2084 1381 2166 1415
rect 2084 1347 2108 1381
rect 2142 1347 2166 1381
rect 2084 1313 2166 1347
rect 2084 1279 2108 1313
rect 2142 1279 2166 1313
rect 2084 1245 2166 1279
rect 2084 1211 2108 1245
rect 2142 1211 2166 1245
rect 2084 1177 2166 1211
rect 2084 1143 2108 1177
rect 2142 1143 2166 1177
rect 2084 1109 2166 1143
rect 2084 1075 2108 1109
rect 2142 1075 2166 1109
rect 2084 1041 2166 1075
rect 2084 1007 2108 1041
rect 2142 1007 2166 1041
rect 2084 973 2166 1007
rect 2084 939 2108 973
rect 2142 939 2166 973
rect 2084 905 2166 939
rect 2084 871 2108 905
rect 2142 871 2166 905
rect 2084 837 2166 871
rect 2084 803 2108 837
rect 2142 803 2166 837
rect 2084 769 2166 803
rect 2084 735 2108 769
rect 2142 735 2166 769
rect 2084 701 2166 735
rect 2084 667 2108 701
rect 2142 667 2166 701
rect 2084 633 2166 667
rect 2084 599 2108 633
rect 2142 599 2166 633
rect 2084 565 2166 599
rect 2084 531 2108 565
rect 2142 531 2166 565
rect 2084 497 2166 531
rect 2084 463 2108 497
rect 2142 463 2166 497
rect 2084 429 2166 463
rect 2084 395 2108 429
rect 2142 395 2166 429
rect 2084 361 2166 395
rect 2084 327 2108 361
rect 2142 327 2166 361
rect 2084 293 2166 327
rect 2084 259 2108 293
rect 2142 259 2166 293
rect 26 191 50 225
rect 84 191 108 225
rect 26 157 108 191
rect 26 123 50 157
rect 84 123 108 157
rect 26 108 108 123
rect 2084 225 2166 259
rect 2084 191 2108 225
rect 2142 191 2166 225
rect 2084 157 2166 191
rect 2084 123 2108 157
rect 2142 123 2166 157
rect 2084 108 2166 123
rect 26 84 2166 108
rect 26 50 50 84
rect 84 50 127 84
rect 161 50 195 84
rect 229 50 263 84
rect 297 50 331 84
rect 365 50 399 84
rect 433 50 467 84
rect 501 50 535 84
rect 569 50 603 84
rect 637 50 671 84
rect 705 50 739 84
rect 773 50 807 84
rect 841 50 875 84
rect 909 50 943 84
rect 977 50 1011 84
rect 1045 50 1079 84
rect 1113 50 1147 84
rect 1181 50 1215 84
rect 1249 50 1283 84
rect 1317 50 1351 84
rect 1385 50 1419 84
rect 1453 50 1487 84
rect 1521 50 1555 84
rect 1589 50 1623 84
rect 1657 50 1691 84
rect 1725 50 1759 84
rect 1793 50 1827 84
rect 1861 50 1895 84
rect 1929 50 1963 84
rect 1997 50 2031 84
rect 2065 50 2108 84
rect 2142 50 2166 84
rect 26 26 2166 50
<< nsubdiff >>
rect 252 2316 1940 2340
rect 252 2282 276 2316
rect 310 2282 365 2316
rect 399 2282 433 2316
rect 467 2282 501 2316
rect 535 2282 569 2316
rect 603 2282 637 2316
rect 671 2282 705 2316
rect 739 2282 773 2316
rect 807 2282 841 2316
rect 875 2282 909 2316
rect 943 2282 977 2316
rect 1011 2282 1045 2316
rect 1079 2282 1113 2316
rect 1147 2282 1181 2316
rect 1215 2282 1249 2316
rect 1283 2282 1317 2316
rect 1351 2282 1385 2316
rect 1419 2282 1453 2316
rect 1487 2282 1521 2316
rect 1555 2282 1589 2316
rect 1623 2282 1657 2316
rect 1691 2282 1725 2316
rect 1759 2282 1793 2316
rect 1827 2282 1882 2316
rect 1916 2282 1940 2316
rect 252 2258 1940 2282
rect 252 2231 334 2258
rect 252 2197 276 2231
rect 310 2197 334 2231
rect 252 2163 334 2197
rect 252 2129 276 2163
rect 310 2129 334 2163
rect 252 2095 334 2129
rect 252 2061 276 2095
rect 310 2061 334 2095
rect 252 2027 334 2061
rect 252 1993 276 2027
rect 310 1993 334 2027
rect 252 1959 334 1993
rect 252 1925 276 1959
rect 310 1925 334 1959
rect 1858 2231 1940 2258
rect 1858 2197 1882 2231
rect 1916 2197 1940 2231
rect 1858 2163 1940 2197
rect 1858 2129 1882 2163
rect 1916 2129 1940 2163
rect 1858 2095 1940 2129
rect 1858 2061 1882 2095
rect 1916 2061 1940 2095
rect 1858 2027 1940 2061
rect 1858 1993 1882 2027
rect 1916 1993 1940 2027
rect 1858 1959 1940 1993
rect 252 1891 334 1925
rect 252 1857 276 1891
rect 310 1857 334 1891
rect 252 1823 334 1857
rect 252 1789 276 1823
rect 310 1789 334 1823
rect 252 1755 334 1789
rect 252 1721 276 1755
rect 310 1721 334 1755
rect 252 1687 334 1721
rect 252 1653 276 1687
rect 310 1653 334 1687
rect 252 1619 334 1653
rect 252 1585 276 1619
rect 310 1585 334 1619
rect 252 1551 334 1585
rect 252 1517 276 1551
rect 310 1517 334 1551
rect 252 1483 334 1517
rect 252 1449 276 1483
rect 310 1449 334 1483
rect 252 1415 334 1449
rect 252 1381 276 1415
rect 310 1381 334 1415
rect 252 1347 334 1381
rect 252 1313 276 1347
rect 310 1313 334 1347
rect 252 1279 334 1313
rect 252 1245 276 1279
rect 310 1245 334 1279
rect 252 1211 334 1245
rect 252 1177 276 1211
rect 310 1177 334 1211
rect 252 1143 334 1177
rect 252 1109 276 1143
rect 310 1109 334 1143
rect 252 1075 334 1109
rect 252 1041 276 1075
rect 310 1041 334 1075
rect 252 1007 334 1041
rect 252 973 276 1007
rect 310 973 334 1007
rect 252 939 334 973
rect 252 905 276 939
rect 310 905 334 939
rect 252 871 334 905
rect 252 837 276 871
rect 310 837 334 871
rect 252 803 334 837
rect 252 769 276 803
rect 310 769 334 803
rect 252 735 334 769
rect 252 701 276 735
rect 310 701 334 735
rect 252 667 334 701
rect 252 633 276 667
rect 310 633 334 667
rect 1858 1925 1882 1959
rect 1916 1925 1940 1959
rect 1858 1891 1940 1925
rect 1858 1857 1882 1891
rect 1916 1857 1940 1891
rect 1858 1823 1940 1857
rect 1858 1789 1882 1823
rect 1916 1789 1940 1823
rect 1858 1755 1940 1789
rect 1858 1721 1882 1755
rect 1916 1721 1940 1755
rect 1858 1687 1940 1721
rect 1858 1653 1882 1687
rect 1916 1653 1940 1687
rect 1858 1619 1940 1653
rect 1858 1585 1882 1619
rect 1916 1585 1940 1619
rect 1858 1551 1940 1585
rect 1858 1517 1882 1551
rect 1916 1517 1940 1551
rect 1858 1483 1940 1517
rect 1858 1449 1882 1483
rect 1916 1449 1940 1483
rect 1858 1415 1940 1449
rect 1858 1381 1882 1415
rect 1916 1381 1940 1415
rect 1858 1347 1940 1381
rect 1858 1313 1882 1347
rect 1916 1313 1940 1347
rect 1858 1279 1940 1313
rect 1858 1245 1882 1279
rect 1916 1245 1940 1279
rect 1858 1211 1940 1245
rect 1858 1177 1882 1211
rect 1916 1177 1940 1211
rect 1858 1143 1940 1177
rect 1858 1109 1882 1143
rect 1916 1109 1940 1143
rect 1858 1075 1940 1109
rect 1858 1041 1882 1075
rect 1916 1041 1940 1075
rect 1858 1007 1940 1041
rect 1858 973 1882 1007
rect 1916 973 1940 1007
rect 1858 939 1940 973
rect 1858 905 1882 939
rect 1916 905 1940 939
rect 1858 871 1940 905
rect 1858 837 1882 871
rect 1916 837 1940 871
rect 1858 803 1940 837
rect 1858 769 1882 803
rect 1916 769 1940 803
rect 1858 735 1940 769
rect 1858 701 1882 735
rect 1916 701 1940 735
rect 1858 667 1940 701
rect 252 599 334 633
rect 252 565 276 599
rect 310 565 334 599
rect 252 531 334 565
rect 252 497 276 531
rect 310 497 334 531
rect 252 463 334 497
rect 252 429 276 463
rect 310 429 334 463
rect 252 395 334 429
rect 252 361 276 395
rect 310 361 334 395
rect 252 334 334 361
rect 1858 633 1882 667
rect 1916 633 1940 667
rect 1858 599 1940 633
rect 1858 565 1882 599
rect 1916 565 1940 599
rect 1858 531 1940 565
rect 1858 497 1882 531
rect 1916 497 1940 531
rect 1858 463 1940 497
rect 1858 429 1882 463
rect 1916 429 1940 463
rect 1858 395 1940 429
rect 1858 361 1882 395
rect 1916 361 1940 395
rect 1858 334 1940 361
rect 252 310 1940 334
rect 252 276 276 310
rect 310 276 365 310
rect 399 276 433 310
rect 467 276 501 310
rect 535 276 569 310
rect 603 276 637 310
rect 671 276 705 310
rect 739 276 773 310
rect 807 276 841 310
rect 875 276 909 310
rect 943 276 977 310
rect 1011 276 1045 310
rect 1079 276 1113 310
rect 1147 276 1181 310
rect 1215 276 1249 310
rect 1283 276 1317 310
rect 1351 276 1385 310
rect 1419 276 1453 310
rect 1487 276 1521 310
rect 1555 276 1589 310
rect 1623 276 1657 310
rect 1691 276 1725 310
rect 1759 276 1793 310
rect 1827 276 1882 310
rect 1916 276 1940 310
rect 252 252 1940 276
<< psubdiffcont >>
rect 50 2508 84 2542
rect 127 2508 161 2542
rect 195 2508 229 2542
rect 263 2508 297 2542
rect 331 2508 365 2542
rect 399 2508 433 2542
rect 467 2508 501 2542
rect 535 2508 569 2542
rect 603 2508 637 2542
rect 671 2508 705 2542
rect 739 2508 773 2542
rect 807 2508 841 2542
rect 875 2508 909 2542
rect 943 2508 977 2542
rect 1011 2508 1045 2542
rect 1079 2508 1113 2542
rect 1147 2508 1181 2542
rect 1215 2508 1249 2542
rect 1283 2508 1317 2542
rect 1351 2508 1385 2542
rect 1419 2508 1453 2542
rect 1487 2508 1521 2542
rect 1555 2508 1589 2542
rect 1623 2508 1657 2542
rect 1691 2508 1725 2542
rect 1759 2508 1793 2542
rect 1827 2508 1861 2542
rect 1895 2508 1929 2542
rect 1963 2508 1997 2542
rect 2031 2508 2065 2542
rect 2108 2508 2142 2542
rect 50 2435 84 2469
rect 50 2367 84 2401
rect 2108 2435 2142 2469
rect 2108 2367 2142 2401
rect 50 2299 84 2333
rect 50 2231 84 2265
rect 50 2163 84 2197
rect 50 2095 84 2129
rect 50 2027 84 2061
rect 50 1959 84 1993
rect 50 1891 84 1925
rect 50 1823 84 1857
rect 50 1755 84 1789
rect 50 1687 84 1721
rect 50 1619 84 1653
rect 50 1551 84 1585
rect 50 1483 84 1517
rect 50 1415 84 1449
rect 50 1347 84 1381
rect 50 1279 84 1313
rect 50 1211 84 1245
rect 50 1143 84 1177
rect 50 1075 84 1109
rect 50 1007 84 1041
rect 50 939 84 973
rect 50 871 84 905
rect 50 803 84 837
rect 50 735 84 769
rect 50 667 84 701
rect 50 599 84 633
rect 50 531 84 565
rect 50 463 84 497
rect 50 395 84 429
rect 50 327 84 361
rect 50 259 84 293
rect 678 1880 712 1914
rect 773 1880 807 1914
rect 841 1880 875 1914
rect 909 1880 943 1914
rect 977 1880 1011 1914
rect 1045 1880 1079 1914
rect 1113 1880 1147 1914
rect 1181 1880 1215 1914
rect 1249 1880 1283 1914
rect 1317 1880 1351 1914
rect 1385 1880 1419 1914
rect 1480 1880 1514 1914
rect 678 1789 712 1823
rect 678 1721 712 1755
rect 1480 1789 1514 1823
rect 1480 1721 1514 1755
rect 678 1653 712 1687
rect 678 1585 712 1619
rect 678 1517 712 1551
rect 678 1449 712 1483
rect 678 1381 712 1415
rect 678 1313 712 1347
rect 678 1245 712 1279
rect 678 1177 712 1211
rect 678 1109 712 1143
rect 678 1041 712 1075
rect 678 973 712 1007
rect 678 905 712 939
rect 1480 1653 1514 1687
rect 1480 1585 1514 1619
rect 1480 1517 1514 1551
rect 1480 1449 1514 1483
rect 1480 1381 1514 1415
rect 1480 1313 1514 1347
rect 1480 1245 1514 1279
rect 1480 1177 1514 1211
rect 1480 1109 1514 1143
rect 1480 1041 1514 1075
rect 1480 973 1514 1007
rect 1480 905 1514 939
rect 678 837 712 871
rect 678 769 712 803
rect 1480 837 1514 871
rect 1480 769 1514 803
rect 678 678 712 712
rect 773 678 807 712
rect 841 678 875 712
rect 909 678 943 712
rect 977 678 1011 712
rect 1045 678 1079 712
rect 1113 678 1147 712
rect 1181 678 1215 712
rect 1249 678 1283 712
rect 1317 678 1351 712
rect 1385 678 1419 712
rect 1480 678 1514 712
rect 2108 2299 2142 2333
rect 2108 2231 2142 2265
rect 2108 2163 2142 2197
rect 2108 2095 2142 2129
rect 2108 2027 2142 2061
rect 2108 1959 2142 1993
rect 2108 1891 2142 1925
rect 2108 1823 2142 1857
rect 2108 1755 2142 1789
rect 2108 1687 2142 1721
rect 2108 1619 2142 1653
rect 2108 1551 2142 1585
rect 2108 1483 2142 1517
rect 2108 1415 2142 1449
rect 2108 1347 2142 1381
rect 2108 1279 2142 1313
rect 2108 1211 2142 1245
rect 2108 1143 2142 1177
rect 2108 1075 2142 1109
rect 2108 1007 2142 1041
rect 2108 939 2142 973
rect 2108 871 2142 905
rect 2108 803 2142 837
rect 2108 735 2142 769
rect 2108 667 2142 701
rect 2108 599 2142 633
rect 2108 531 2142 565
rect 2108 463 2142 497
rect 2108 395 2142 429
rect 2108 327 2142 361
rect 2108 259 2142 293
rect 50 191 84 225
rect 50 123 84 157
rect 2108 191 2142 225
rect 2108 123 2142 157
rect 50 50 84 84
rect 127 50 161 84
rect 195 50 229 84
rect 263 50 297 84
rect 331 50 365 84
rect 399 50 433 84
rect 467 50 501 84
rect 535 50 569 84
rect 603 50 637 84
rect 671 50 705 84
rect 739 50 773 84
rect 807 50 841 84
rect 875 50 909 84
rect 943 50 977 84
rect 1011 50 1045 84
rect 1079 50 1113 84
rect 1147 50 1181 84
rect 1215 50 1249 84
rect 1283 50 1317 84
rect 1351 50 1385 84
rect 1419 50 1453 84
rect 1487 50 1521 84
rect 1555 50 1589 84
rect 1623 50 1657 84
rect 1691 50 1725 84
rect 1759 50 1793 84
rect 1827 50 1861 84
rect 1895 50 1929 84
rect 1963 50 1997 84
rect 2031 50 2065 84
rect 2108 50 2142 84
<< nsubdiffcont >>
rect 276 2282 310 2316
rect 365 2282 399 2316
rect 433 2282 467 2316
rect 501 2282 535 2316
rect 569 2282 603 2316
rect 637 2282 671 2316
rect 705 2282 739 2316
rect 773 2282 807 2316
rect 841 2282 875 2316
rect 909 2282 943 2316
rect 977 2282 1011 2316
rect 1045 2282 1079 2316
rect 1113 2282 1147 2316
rect 1181 2282 1215 2316
rect 1249 2282 1283 2316
rect 1317 2282 1351 2316
rect 1385 2282 1419 2316
rect 1453 2282 1487 2316
rect 1521 2282 1555 2316
rect 1589 2282 1623 2316
rect 1657 2282 1691 2316
rect 1725 2282 1759 2316
rect 1793 2282 1827 2316
rect 1882 2282 1916 2316
rect 276 2197 310 2231
rect 276 2129 310 2163
rect 276 2061 310 2095
rect 276 1993 310 2027
rect 276 1925 310 1959
rect 1882 2197 1916 2231
rect 1882 2129 1916 2163
rect 1882 2061 1916 2095
rect 1882 1993 1916 2027
rect 276 1857 310 1891
rect 276 1789 310 1823
rect 276 1721 310 1755
rect 276 1653 310 1687
rect 276 1585 310 1619
rect 276 1517 310 1551
rect 276 1449 310 1483
rect 276 1381 310 1415
rect 276 1313 310 1347
rect 276 1245 310 1279
rect 276 1177 310 1211
rect 276 1109 310 1143
rect 276 1041 310 1075
rect 276 973 310 1007
rect 276 905 310 939
rect 276 837 310 871
rect 276 769 310 803
rect 276 701 310 735
rect 276 633 310 667
rect 1882 1925 1916 1959
rect 1882 1857 1916 1891
rect 1882 1789 1916 1823
rect 1882 1721 1916 1755
rect 1882 1653 1916 1687
rect 1882 1585 1916 1619
rect 1882 1517 1916 1551
rect 1882 1449 1916 1483
rect 1882 1381 1916 1415
rect 1882 1313 1916 1347
rect 1882 1245 1916 1279
rect 1882 1177 1916 1211
rect 1882 1109 1916 1143
rect 1882 1041 1916 1075
rect 1882 973 1916 1007
rect 1882 905 1916 939
rect 1882 837 1916 871
rect 1882 769 1916 803
rect 1882 701 1916 735
rect 276 565 310 599
rect 276 497 310 531
rect 276 429 310 463
rect 276 361 310 395
rect 1882 633 1916 667
rect 1882 565 1916 599
rect 1882 497 1916 531
rect 1882 429 1916 463
rect 1882 361 1916 395
rect 276 276 310 310
rect 365 276 399 310
rect 433 276 467 310
rect 501 276 535 310
rect 569 276 603 310
rect 637 276 671 310
rect 705 276 739 310
rect 773 276 807 310
rect 841 276 875 310
rect 909 276 943 310
rect 977 276 1011 310
rect 1045 276 1079 310
rect 1113 276 1147 310
rect 1181 276 1215 310
rect 1249 276 1283 310
rect 1317 276 1351 310
rect 1385 276 1419 310
rect 1453 276 1487 310
rect 1521 276 1555 310
rect 1589 276 1623 310
rect 1657 276 1691 310
rect 1725 276 1759 310
rect 1793 276 1827 310
rect 1882 276 1916 310
<< locali >>
rect 34 2542 2158 2558
rect 34 2508 50 2542
rect 84 2508 127 2542
rect 177 2508 195 2542
rect 249 2508 263 2542
rect 321 2508 331 2542
rect 393 2508 399 2542
rect 465 2508 467 2542
rect 501 2508 503 2542
rect 569 2508 575 2542
rect 637 2508 647 2542
rect 705 2508 719 2542
rect 773 2508 791 2542
rect 841 2508 863 2542
rect 909 2508 935 2542
rect 977 2508 1007 2542
rect 1045 2508 1079 2542
rect 1113 2508 1147 2542
rect 1185 2508 1215 2542
rect 1257 2508 1283 2542
rect 1329 2508 1351 2542
rect 1401 2508 1419 2542
rect 1473 2508 1487 2542
rect 1545 2508 1555 2542
rect 1617 2508 1623 2542
rect 1689 2508 1691 2542
rect 1725 2508 1727 2542
rect 1793 2508 1799 2542
rect 1861 2508 1871 2542
rect 1929 2508 1943 2542
rect 1997 2508 2015 2542
rect 2065 2508 2108 2542
rect 2142 2508 2158 2542
rect 34 2492 2158 2508
rect 34 2469 100 2492
rect 34 2431 50 2469
rect 84 2431 100 2469
rect 34 2401 100 2431
rect 34 2359 50 2401
rect 84 2359 100 2401
rect 34 2333 100 2359
rect 34 2287 50 2333
rect 84 2287 100 2333
rect 2092 2469 2158 2492
rect 2092 2431 2108 2469
rect 2142 2431 2158 2469
rect 2092 2401 2158 2431
rect 2092 2359 2108 2401
rect 2142 2359 2158 2401
rect 2092 2333 2158 2359
rect 34 2265 100 2287
rect 34 2215 50 2265
rect 84 2215 100 2265
rect 34 2197 100 2215
rect 34 2143 50 2197
rect 84 2143 100 2197
rect 34 2129 100 2143
rect 34 2071 50 2129
rect 84 2071 100 2129
rect 34 2061 100 2071
rect 34 1999 50 2061
rect 84 1999 100 2061
rect 34 1993 100 1999
rect 34 1927 50 1993
rect 84 1927 100 1993
rect 34 1925 100 1927
rect 34 1891 50 1925
rect 84 1891 100 1925
rect 34 1889 100 1891
rect 34 1823 50 1889
rect 84 1823 100 1889
rect 34 1817 100 1823
rect 34 1755 50 1817
rect 84 1755 100 1817
rect 34 1745 100 1755
rect 34 1687 50 1745
rect 84 1687 100 1745
rect 34 1673 100 1687
rect 34 1619 50 1673
rect 84 1619 100 1673
rect 34 1601 100 1619
rect 34 1551 50 1601
rect 84 1551 100 1601
rect 34 1529 100 1551
rect 34 1483 50 1529
rect 84 1483 100 1529
rect 34 1457 100 1483
rect 34 1415 50 1457
rect 84 1415 100 1457
rect 34 1385 100 1415
rect 34 1347 50 1385
rect 84 1347 100 1385
rect 34 1313 100 1347
rect 34 1279 50 1313
rect 84 1279 100 1313
rect 34 1245 100 1279
rect 34 1207 50 1245
rect 84 1207 100 1245
rect 34 1177 100 1207
rect 34 1135 50 1177
rect 84 1135 100 1177
rect 34 1109 100 1135
rect 34 1063 50 1109
rect 84 1063 100 1109
rect 34 1041 100 1063
rect 34 991 50 1041
rect 84 991 100 1041
rect 34 973 100 991
rect 34 919 50 973
rect 84 919 100 973
rect 34 905 100 919
rect 34 847 50 905
rect 84 847 100 905
rect 34 837 100 847
rect 34 775 50 837
rect 84 775 100 837
rect 34 769 100 775
rect 34 703 50 769
rect 84 703 100 769
rect 34 701 100 703
rect 34 667 50 701
rect 84 667 100 701
rect 34 665 100 667
rect 34 599 50 665
rect 84 599 100 665
rect 34 593 100 599
rect 34 531 50 593
rect 84 531 100 593
rect 34 521 100 531
rect 34 463 50 521
rect 84 463 100 521
rect 34 449 100 463
rect 34 395 50 449
rect 84 395 100 449
rect 34 377 100 395
rect 34 327 50 377
rect 84 327 100 377
rect 34 305 100 327
rect 34 259 50 305
rect 84 259 100 305
rect 260 2316 1932 2332
rect 260 2282 276 2316
rect 310 2282 359 2316
rect 399 2282 431 2316
rect 467 2282 501 2316
rect 537 2282 569 2316
rect 609 2282 637 2316
rect 681 2282 705 2316
rect 753 2282 773 2316
rect 825 2282 841 2316
rect 897 2282 909 2316
rect 969 2282 977 2316
rect 1041 2282 1045 2316
rect 1147 2282 1151 2316
rect 1215 2282 1223 2316
rect 1283 2282 1295 2316
rect 1351 2282 1367 2316
rect 1419 2282 1439 2316
rect 1487 2282 1511 2316
rect 1555 2282 1583 2316
rect 1623 2282 1655 2316
rect 1691 2282 1725 2316
rect 1761 2282 1793 2316
rect 1833 2282 1882 2316
rect 1916 2282 1932 2316
rect 260 2266 1932 2282
rect 260 2231 326 2266
rect 260 2179 276 2231
rect 310 2179 326 2231
rect 260 2163 326 2179
rect 260 2107 276 2163
rect 310 2107 326 2163
rect 260 2095 326 2107
rect 260 2035 276 2095
rect 310 2035 326 2095
rect 260 2027 326 2035
rect 260 1963 276 2027
rect 310 1963 326 2027
rect 260 1959 326 1963
rect 260 1857 276 1959
rect 310 1857 326 1959
rect 1866 2231 1932 2266
rect 1866 2179 1882 2231
rect 1916 2179 1932 2231
rect 1866 2163 1932 2179
rect 1866 2107 1882 2163
rect 1916 2107 1932 2163
rect 1866 2095 1932 2107
rect 1866 2035 1882 2095
rect 1916 2035 1932 2095
rect 1866 2027 1932 2035
rect 1866 1963 1882 2027
rect 1916 1963 1932 2027
rect 1866 1959 1932 1963
rect 260 1853 326 1857
rect 260 1789 276 1853
rect 310 1789 326 1853
rect 260 1781 326 1789
rect 260 1721 276 1781
rect 310 1721 326 1781
rect 260 1709 326 1721
rect 260 1653 276 1709
rect 310 1653 326 1709
rect 260 1637 326 1653
rect 260 1585 276 1637
rect 310 1585 326 1637
rect 260 1565 326 1585
rect 260 1517 276 1565
rect 310 1517 326 1565
rect 260 1493 326 1517
rect 260 1449 276 1493
rect 310 1449 326 1493
rect 260 1421 326 1449
rect 260 1381 276 1421
rect 310 1381 326 1421
rect 260 1349 326 1381
rect 260 1313 276 1349
rect 310 1313 326 1349
rect 260 1279 326 1313
rect 260 1243 276 1279
rect 310 1243 326 1279
rect 260 1211 326 1243
rect 260 1171 276 1211
rect 310 1171 326 1211
rect 260 1143 326 1171
rect 260 1099 276 1143
rect 310 1099 326 1143
rect 260 1075 326 1099
rect 260 1027 276 1075
rect 310 1027 326 1075
rect 260 1007 326 1027
rect 260 955 276 1007
rect 310 955 326 1007
rect 260 939 326 955
rect 260 883 276 939
rect 310 883 326 939
rect 260 871 326 883
rect 260 811 276 871
rect 310 811 326 871
rect 260 803 326 811
rect 260 739 276 803
rect 310 739 326 803
rect 260 735 326 739
rect 260 633 276 735
rect 310 633 326 735
rect 662 1914 1530 1930
rect 662 1880 678 1914
rect 712 1880 755 1914
rect 807 1880 827 1914
rect 875 1880 899 1914
rect 943 1880 971 1914
rect 1011 1880 1043 1914
rect 1079 1880 1113 1914
rect 1149 1880 1181 1914
rect 1221 1880 1249 1914
rect 1293 1880 1317 1914
rect 1365 1880 1385 1914
rect 1437 1880 1480 1914
rect 1514 1880 1530 1914
rect 662 1864 1530 1880
rect 662 1823 728 1864
rect 662 1783 678 1823
rect 712 1783 728 1823
rect 662 1755 728 1783
rect 662 1711 678 1755
rect 712 1711 728 1755
rect 662 1687 728 1711
rect 1464 1823 1530 1864
rect 1464 1783 1480 1823
rect 1514 1783 1530 1823
rect 1464 1755 1530 1783
rect 1464 1711 1480 1755
rect 1514 1711 1530 1755
rect 662 1639 678 1687
rect 712 1639 728 1687
rect 662 1619 728 1639
rect 662 1567 678 1619
rect 712 1567 728 1619
rect 662 1551 728 1567
rect 662 1495 678 1551
rect 712 1495 728 1551
rect 662 1483 728 1495
rect 662 1423 678 1483
rect 712 1423 728 1483
rect 662 1415 728 1423
rect 662 1351 678 1415
rect 712 1351 728 1415
rect 662 1347 728 1351
rect 662 1245 678 1347
rect 712 1245 728 1347
rect 662 1241 728 1245
rect 662 1177 678 1241
rect 712 1177 728 1241
rect 662 1169 728 1177
rect 662 1109 678 1169
rect 712 1109 728 1169
rect 662 1097 728 1109
rect 662 1041 678 1097
rect 712 1041 728 1097
rect 662 1025 728 1041
rect 662 973 678 1025
rect 712 973 728 1025
rect 662 953 728 973
rect 662 905 678 953
rect 712 905 728 953
rect 662 881 728 905
rect 893 1653 1299 1699
rect 893 939 909 1653
rect 1283 939 1299 1653
rect 893 893 1299 939
rect 1464 1687 1530 1711
rect 1464 1639 1480 1687
rect 1514 1639 1530 1687
rect 1464 1619 1530 1639
rect 1464 1567 1480 1619
rect 1514 1567 1530 1619
rect 1464 1551 1530 1567
rect 1464 1495 1480 1551
rect 1514 1495 1530 1551
rect 1464 1483 1530 1495
rect 1464 1423 1480 1483
rect 1514 1423 1530 1483
rect 1464 1415 1530 1423
rect 1464 1351 1480 1415
rect 1514 1351 1530 1415
rect 1464 1347 1530 1351
rect 1464 1245 1480 1347
rect 1514 1245 1530 1347
rect 1464 1241 1530 1245
rect 1464 1177 1480 1241
rect 1514 1177 1530 1241
rect 1464 1169 1530 1177
rect 1464 1109 1480 1169
rect 1514 1109 1530 1169
rect 1464 1097 1530 1109
rect 1464 1041 1480 1097
rect 1514 1041 1530 1097
rect 1464 1025 1530 1041
rect 1464 973 1480 1025
rect 1514 973 1530 1025
rect 1464 953 1530 973
rect 1464 905 1480 953
rect 1514 905 1530 953
rect 662 837 678 881
rect 712 837 728 881
rect 662 809 728 837
rect 662 769 678 809
rect 712 769 728 809
rect 662 728 728 769
rect 1464 881 1530 905
rect 1464 837 1480 881
rect 1514 837 1530 881
rect 1464 809 1530 837
rect 1464 769 1480 809
rect 1514 769 1530 809
rect 1464 728 1530 769
rect 662 712 1530 728
rect 662 678 678 712
rect 712 678 755 712
rect 807 678 827 712
rect 875 678 899 712
rect 943 678 971 712
rect 1011 678 1043 712
rect 1079 678 1113 712
rect 1149 678 1181 712
rect 1221 678 1249 712
rect 1293 678 1317 712
rect 1365 678 1385 712
rect 1437 678 1480 712
rect 1514 678 1530 712
rect 662 662 1530 678
rect 1866 1857 1882 1959
rect 1916 1857 1932 1959
rect 1866 1853 1932 1857
rect 1866 1789 1882 1853
rect 1916 1789 1932 1853
rect 1866 1781 1932 1789
rect 1866 1721 1882 1781
rect 1916 1721 1932 1781
rect 1866 1709 1932 1721
rect 1866 1653 1882 1709
rect 1916 1653 1932 1709
rect 1866 1637 1932 1653
rect 1866 1585 1882 1637
rect 1916 1585 1932 1637
rect 1866 1565 1932 1585
rect 1866 1517 1882 1565
rect 1916 1517 1932 1565
rect 1866 1493 1932 1517
rect 1866 1449 1882 1493
rect 1916 1449 1932 1493
rect 1866 1421 1932 1449
rect 1866 1381 1882 1421
rect 1916 1381 1932 1421
rect 1866 1349 1932 1381
rect 1866 1313 1882 1349
rect 1916 1313 1932 1349
rect 1866 1279 1932 1313
rect 1866 1243 1882 1279
rect 1916 1243 1932 1279
rect 1866 1211 1932 1243
rect 1866 1171 1882 1211
rect 1916 1171 1932 1211
rect 1866 1143 1932 1171
rect 1866 1099 1882 1143
rect 1916 1099 1932 1143
rect 1866 1075 1932 1099
rect 1866 1027 1882 1075
rect 1916 1027 1932 1075
rect 1866 1007 1932 1027
rect 1866 955 1882 1007
rect 1916 955 1932 1007
rect 1866 939 1932 955
rect 1866 883 1882 939
rect 1916 883 1932 939
rect 1866 871 1932 883
rect 1866 811 1882 871
rect 1916 811 1932 871
rect 1866 803 1932 811
rect 1866 739 1882 803
rect 1916 739 1932 803
rect 1866 735 1932 739
rect 260 629 326 633
rect 260 565 276 629
rect 310 565 326 629
rect 260 557 326 565
rect 260 497 276 557
rect 310 497 326 557
rect 260 485 326 497
rect 260 429 276 485
rect 310 429 326 485
rect 260 413 326 429
rect 260 361 276 413
rect 310 361 326 413
rect 260 326 326 361
rect 1866 633 1882 735
rect 1916 633 1932 735
rect 1866 629 1932 633
rect 1866 565 1882 629
rect 1916 565 1932 629
rect 1866 557 1932 565
rect 1866 497 1882 557
rect 1916 497 1932 557
rect 1866 485 1932 497
rect 1866 429 1882 485
rect 1916 429 1932 485
rect 1866 413 1932 429
rect 1866 361 1882 413
rect 1916 361 1932 413
rect 1866 326 1932 361
rect 260 310 1932 326
rect 260 276 276 310
rect 310 276 359 310
rect 399 276 431 310
rect 467 276 501 310
rect 537 276 569 310
rect 609 276 637 310
rect 681 276 705 310
rect 753 276 773 310
rect 825 276 841 310
rect 897 276 909 310
rect 969 276 977 310
rect 1041 276 1045 310
rect 1147 276 1151 310
rect 1215 276 1223 310
rect 1283 276 1295 310
rect 1351 276 1367 310
rect 1419 276 1439 310
rect 1487 276 1511 310
rect 1555 276 1583 310
rect 1623 276 1655 310
rect 1691 276 1725 310
rect 1761 276 1793 310
rect 1833 276 1882 310
rect 1916 276 1932 310
rect 260 260 1932 276
rect 2092 2287 2108 2333
rect 2142 2287 2158 2333
rect 2092 2265 2158 2287
rect 2092 2215 2108 2265
rect 2142 2215 2158 2265
rect 2092 2197 2158 2215
rect 2092 2143 2108 2197
rect 2142 2143 2158 2197
rect 2092 2129 2158 2143
rect 2092 2071 2108 2129
rect 2142 2071 2158 2129
rect 2092 2061 2158 2071
rect 2092 1999 2108 2061
rect 2142 1999 2158 2061
rect 2092 1993 2158 1999
rect 2092 1927 2108 1993
rect 2142 1927 2158 1993
rect 2092 1925 2158 1927
rect 2092 1891 2108 1925
rect 2142 1891 2158 1925
rect 2092 1889 2158 1891
rect 2092 1823 2108 1889
rect 2142 1823 2158 1889
rect 2092 1817 2158 1823
rect 2092 1755 2108 1817
rect 2142 1755 2158 1817
rect 2092 1745 2158 1755
rect 2092 1687 2108 1745
rect 2142 1687 2158 1745
rect 2092 1673 2158 1687
rect 2092 1619 2108 1673
rect 2142 1619 2158 1673
rect 2092 1601 2158 1619
rect 2092 1551 2108 1601
rect 2142 1551 2158 1601
rect 2092 1529 2158 1551
rect 2092 1483 2108 1529
rect 2142 1483 2158 1529
rect 2092 1457 2158 1483
rect 2092 1415 2108 1457
rect 2142 1415 2158 1457
rect 2092 1385 2158 1415
rect 2092 1347 2108 1385
rect 2142 1347 2158 1385
rect 2092 1313 2158 1347
rect 2092 1279 2108 1313
rect 2142 1279 2158 1313
rect 2092 1245 2158 1279
rect 2092 1207 2108 1245
rect 2142 1207 2158 1245
rect 2092 1177 2158 1207
rect 2092 1135 2108 1177
rect 2142 1135 2158 1177
rect 2092 1109 2158 1135
rect 2092 1063 2108 1109
rect 2142 1063 2158 1109
rect 2092 1041 2158 1063
rect 2092 991 2108 1041
rect 2142 991 2158 1041
rect 2092 973 2158 991
rect 2092 919 2108 973
rect 2142 919 2158 973
rect 2092 905 2158 919
rect 2092 847 2108 905
rect 2142 847 2158 905
rect 2092 837 2158 847
rect 2092 775 2108 837
rect 2142 775 2158 837
rect 2092 769 2158 775
rect 2092 703 2108 769
rect 2142 703 2158 769
rect 2092 701 2158 703
rect 2092 667 2108 701
rect 2142 667 2158 701
rect 2092 665 2158 667
rect 2092 599 2108 665
rect 2142 599 2158 665
rect 2092 593 2158 599
rect 2092 531 2108 593
rect 2142 531 2158 593
rect 2092 521 2158 531
rect 2092 463 2108 521
rect 2142 463 2158 521
rect 2092 449 2158 463
rect 2092 395 2108 449
rect 2142 395 2158 449
rect 2092 377 2158 395
rect 2092 327 2108 377
rect 2142 327 2158 377
rect 2092 305 2158 327
rect 34 233 100 259
rect 34 191 50 233
rect 84 191 100 233
rect 34 161 100 191
rect 34 123 50 161
rect 84 123 100 161
rect 34 100 100 123
rect 2092 259 2108 305
rect 2142 259 2158 305
rect 2092 233 2158 259
rect 2092 191 2108 233
rect 2142 191 2158 233
rect 2092 161 2158 191
rect 2092 123 2108 161
rect 2142 123 2158 161
rect 2092 100 2158 123
rect 34 84 2158 100
rect 34 50 50 84
rect 84 50 127 84
rect 177 50 195 84
rect 249 50 263 84
rect 321 50 331 84
rect 393 50 399 84
rect 465 50 467 84
rect 501 50 503 84
rect 569 50 575 84
rect 637 50 647 84
rect 705 50 719 84
rect 773 50 791 84
rect 841 50 863 84
rect 909 50 935 84
rect 977 50 1007 84
rect 1045 50 1079 84
rect 1113 50 1147 84
rect 1185 50 1215 84
rect 1257 50 1283 84
rect 1329 50 1351 84
rect 1401 50 1419 84
rect 1473 50 1487 84
rect 1545 50 1555 84
rect 1617 50 1623 84
rect 1689 50 1691 84
rect 1725 50 1727 84
rect 1793 50 1799 84
rect 1861 50 1871 84
rect 1929 50 1943 84
rect 1997 50 2015 84
rect 2065 50 2108 84
rect 2142 50 2158 84
rect 34 34 2158 50
<< viali >>
rect 50 2508 84 2542
rect 143 2508 161 2542
rect 161 2508 177 2542
rect 215 2508 229 2542
rect 229 2508 249 2542
rect 287 2508 297 2542
rect 297 2508 321 2542
rect 359 2508 365 2542
rect 365 2508 393 2542
rect 431 2508 433 2542
rect 433 2508 465 2542
rect 503 2508 535 2542
rect 535 2508 537 2542
rect 575 2508 603 2542
rect 603 2508 609 2542
rect 647 2508 671 2542
rect 671 2508 681 2542
rect 719 2508 739 2542
rect 739 2508 753 2542
rect 791 2508 807 2542
rect 807 2508 825 2542
rect 863 2508 875 2542
rect 875 2508 897 2542
rect 935 2508 943 2542
rect 943 2508 969 2542
rect 1007 2508 1011 2542
rect 1011 2508 1041 2542
rect 1079 2508 1113 2542
rect 1151 2508 1181 2542
rect 1181 2508 1185 2542
rect 1223 2508 1249 2542
rect 1249 2508 1257 2542
rect 1295 2508 1317 2542
rect 1317 2508 1329 2542
rect 1367 2508 1385 2542
rect 1385 2508 1401 2542
rect 1439 2508 1453 2542
rect 1453 2508 1473 2542
rect 1511 2508 1521 2542
rect 1521 2508 1545 2542
rect 1583 2508 1589 2542
rect 1589 2508 1617 2542
rect 1655 2508 1657 2542
rect 1657 2508 1689 2542
rect 1727 2508 1759 2542
rect 1759 2508 1761 2542
rect 1799 2508 1827 2542
rect 1827 2508 1833 2542
rect 1871 2508 1895 2542
rect 1895 2508 1905 2542
rect 1943 2508 1963 2542
rect 1963 2508 1977 2542
rect 2015 2508 2031 2542
rect 2031 2508 2049 2542
rect 2108 2508 2142 2542
rect 50 2435 84 2465
rect 50 2431 84 2435
rect 50 2367 84 2393
rect 50 2359 84 2367
rect 50 2299 84 2321
rect 50 2287 84 2299
rect 2108 2435 2142 2465
rect 2108 2431 2142 2435
rect 2108 2367 2142 2393
rect 2108 2359 2142 2367
rect 50 2231 84 2249
rect 50 2215 84 2231
rect 50 2163 84 2177
rect 50 2143 84 2163
rect 50 2095 84 2105
rect 50 2071 84 2095
rect 50 2027 84 2033
rect 50 1999 84 2027
rect 50 1959 84 1961
rect 50 1927 84 1959
rect 50 1857 84 1889
rect 50 1855 84 1857
rect 50 1789 84 1817
rect 50 1783 84 1789
rect 50 1721 84 1745
rect 50 1711 84 1721
rect 50 1653 84 1673
rect 50 1639 84 1653
rect 50 1585 84 1601
rect 50 1567 84 1585
rect 50 1517 84 1529
rect 50 1495 84 1517
rect 50 1449 84 1457
rect 50 1423 84 1449
rect 50 1381 84 1385
rect 50 1351 84 1381
rect 50 1279 84 1313
rect 50 1211 84 1241
rect 50 1207 84 1211
rect 50 1143 84 1169
rect 50 1135 84 1143
rect 50 1075 84 1097
rect 50 1063 84 1075
rect 50 1007 84 1025
rect 50 991 84 1007
rect 50 939 84 953
rect 50 919 84 939
rect 50 871 84 881
rect 50 847 84 871
rect 50 803 84 809
rect 50 775 84 803
rect 50 735 84 737
rect 50 703 84 735
rect 50 633 84 665
rect 50 631 84 633
rect 50 565 84 593
rect 50 559 84 565
rect 50 497 84 521
rect 50 487 84 497
rect 50 429 84 449
rect 50 415 84 429
rect 50 361 84 377
rect 50 343 84 361
rect 50 293 84 305
rect 50 271 84 293
rect 276 2282 310 2316
rect 359 2282 365 2316
rect 365 2282 393 2316
rect 431 2282 433 2316
rect 433 2282 465 2316
rect 503 2282 535 2316
rect 535 2282 537 2316
rect 575 2282 603 2316
rect 603 2282 609 2316
rect 647 2282 671 2316
rect 671 2282 681 2316
rect 719 2282 739 2316
rect 739 2282 753 2316
rect 791 2282 807 2316
rect 807 2282 825 2316
rect 863 2282 875 2316
rect 875 2282 897 2316
rect 935 2282 943 2316
rect 943 2282 969 2316
rect 1007 2282 1011 2316
rect 1011 2282 1041 2316
rect 1079 2282 1113 2316
rect 1151 2282 1181 2316
rect 1181 2282 1185 2316
rect 1223 2282 1249 2316
rect 1249 2282 1257 2316
rect 1295 2282 1317 2316
rect 1317 2282 1329 2316
rect 1367 2282 1385 2316
rect 1385 2282 1401 2316
rect 1439 2282 1453 2316
rect 1453 2282 1473 2316
rect 1511 2282 1521 2316
rect 1521 2282 1545 2316
rect 1583 2282 1589 2316
rect 1589 2282 1617 2316
rect 1655 2282 1657 2316
rect 1657 2282 1689 2316
rect 1727 2282 1759 2316
rect 1759 2282 1761 2316
rect 1799 2282 1827 2316
rect 1827 2282 1833 2316
rect 1882 2282 1916 2316
rect 276 2197 310 2213
rect 276 2179 310 2197
rect 276 2129 310 2141
rect 276 2107 310 2129
rect 276 2061 310 2069
rect 276 2035 310 2061
rect 276 1993 310 1997
rect 276 1963 310 1993
rect 276 1891 310 1925
rect 1882 2197 1916 2213
rect 1882 2179 1916 2197
rect 1882 2129 1916 2141
rect 1882 2107 1916 2129
rect 1882 2061 1916 2069
rect 1882 2035 1916 2061
rect 1882 1993 1916 1997
rect 1882 1963 1916 1993
rect 276 1823 310 1853
rect 276 1819 310 1823
rect 276 1755 310 1781
rect 276 1747 310 1755
rect 276 1687 310 1709
rect 276 1675 310 1687
rect 276 1619 310 1637
rect 276 1603 310 1619
rect 276 1551 310 1565
rect 276 1531 310 1551
rect 276 1483 310 1493
rect 276 1459 310 1483
rect 276 1415 310 1421
rect 276 1387 310 1415
rect 276 1347 310 1349
rect 276 1315 310 1347
rect 276 1245 310 1277
rect 276 1243 310 1245
rect 276 1177 310 1205
rect 276 1171 310 1177
rect 276 1109 310 1133
rect 276 1099 310 1109
rect 276 1041 310 1061
rect 276 1027 310 1041
rect 276 973 310 989
rect 276 955 310 973
rect 276 905 310 917
rect 276 883 310 905
rect 276 837 310 845
rect 276 811 310 837
rect 276 769 310 773
rect 276 739 310 769
rect 276 667 310 701
rect 678 1880 712 1914
rect 755 1880 773 1914
rect 773 1880 789 1914
rect 827 1880 841 1914
rect 841 1880 861 1914
rect 899 1880 909 1914
rect 909 1880 933 1914
rect 971 1880 977 1914
rect 977 1880 1005 1914
rect 1043 1880 1045 1914
rect 1045 1880 1077 1914
rect 1115 1880 1147 1914
rect 1147 1880 1149 1914
rect 1187 1880 1215 1914
rect 1215 1880 1221 1914
rect 1259 1880 1283 1914
rect 1283 1880 1293 1914
rect 1331 1880 1351 1914
rect 1351 1880 1365 1914
rect 1403 1880 1419 1914
rect 1419 1880 1437 1914
rect 1480 1880 1514 1914
rect 678 1789 712 1817
rect 678 1783 712 1789
rect 678 1721 712 1745
rect 678 1711 712 1721
rect 1480 1789 1514 1817
rect 1480 1783 1514 1789
rect 1480 1721 1514 1745
rect 1480 1711 1514 1721
rect 678 1653 712 1673
rect 678 1639 712 1653
rect 678 1585 712 1601
rect 678 1567 712 1585
rect 678 1517 712 1529
rect 678 1495 712 1517
rect 678 1449 712 1457
rect 678 1423 712 1449
rect 678 1381 712 1385
rect 678 1351 712 1381
rect 678 1279 712 1313
rect 678 1211 712 1241
rect 678 1207 712 1211
rect 678 1143 712 1169
rect 678 1135 712 1143
rect 678 1075 712 1097
rect 678 1063 712 1075
rect 678 1007 712 1025
rect 678 991 712 1007
rect 678 939 712 953
rect 678 919 712 939
rect 935 955 1257 1637
rect 1480 1653 1514 1673
rect 1480 1639 1514 1653
rect 1480 1585 1514 1601
rect 1480 1567 1514 1585
rect 1480 1517 1514 1529
rect 1480 1495 1514 1517
rect 1480 1449 1514 1457
rect 1480 1423 1514 1449
rect 1480 1381 1514 1385
rect 1480 1351 1514 1381
rect 1480 1279 1514 1313
rect 1480 1211 1514 1241
rect 1480 1207 1514 1211
rect 1480 1143 1514 1169
rect 1480 1135 1514 1143
rect 1480 1075 1514 1097
rect 1480 1063 1514 1075
rect 1480 1007 1514 1025
rect 1480 991 1514 1007
rect 1480 939 1514 953
rect 1480 919 1514 939
rect 678 871 712 881
rect 678 847 712 871
rect 678 803 712 809
rect 678 775 712 803
rect 1480 871 1514 881
rect 1480 847 1514 871
rect 1480 803 1514 809
rect 1480 775 1514 803
rect 678 678 712 712
rect 755 678 773 712
rect 773 678 789 712
rect 827 678 841 712
rect 841 678 861 712
rect 899 678 909 712
rect 909 678 933 712
rect 971 678 977 712
rect 977 678 1005 712
rect 1043 678 1045 712
rect 1045 678 1077 712
rect 1115 678 1147 712
rect 1147 678 1149 712
rect 1187 678 1215 712
rect 1215 678 1221 712
rect 1259 678 1283 712
rect 1283 678 1293 712
rect 1331 678 1351 712
rect 1351 678 1365 712
rect 1403 678 1419 712
rect 1419 678 1437 712
rect 1480 678 1514 712
rect 1882 1891 1916 1925
rect 1882 1823 1916 1853
rect 1882 1819 1916 1823
rect 1882 1755 1916 1781
rect 1882 1747 1916 1755
rect 1882 1687 1916 1709
rect 1882 1675 1916 1687
rect 1882 1619 1916 1637
rect 1882 1603 1916 1619
rect 1882 1551 1916 1565
rect 1882 1531 1916 1551
rect 1882 1483 1916 1493
rect 1882 1459 1916 1483
rect 1882 1415 1916 1421
rect 1882 1387 1916 1415
rect 1882 1347 1916 1349
rect 1882 1315 1916 1347
rect 1882 1245 1916 1277
rect 1882 1243 1916 1245
rect 1882 1177 1916 1205
rect 1882 1171 1916 1177
rect 1882 1109 1916 1133
rect 1882 1099 1916 1109
rect 1882 1041 1916 1061
rect 1882 1027 1916 1041
rect 1882 973 1916 989
rect 1882 955 1916 973
rect 1882 905 1916 917
rect 1882 883 1916 905
rect 1882 837 1916 845
rect 1882 811 1916 837
rect 1882 769 1916 773
rect 1882 739 1916 769
rect 276 599 310 629
rect 276 595 310 599
rect 276 531 310 557
rect 276 523 310 531
rect 276 463 310 485
rect 276 451 310 463
rect 276 395 310 413
rect 276 379 310 395
rect 1882 667 1916 701
rect 1882 599 1916 629
rect 1882 595 1916 599
rect 1882 531 1916 557
rect 1882 523 1916 531
rect 1882 463 1916 485
rect 1882 451 1916 463
rect 1882 395 1916 413
rect 1882 379 1916 395
rect 276 276 310 310
rect 359 276 365 310
rect 365 276 393 310
rect 431 276 433 310
rect 433 276 465 310
rect 503 276 535 310
rect 535 276 537 310
rect 575 276 603 310
rect 603 276 609 310
rect 647 276 671 310
rect 671 276 681 310
rect 719 276 739 310
rect 739 276 753 310
rect 791 276 807 310
rect 807 276 825 310
rect 863 276 875 310
rect 875 276 897 310
rect 935 276 943 310
rect 943 276 969 310
rect 1007 276 1011 310
rect 1011 276 1041 310
rect 1079 276 1113 310
rect 1151 276 1181 310
rect 1181 276 1185 310
rect 1223 276 1249 310
rect 1249 276 1257 310
rect 1295 276 1317 310
rect 1317 276 1329 310
rect 1367 276 1385 310
rect 1385 276 1401 310
rect 1439 276 1453 310
rect 1453 276 1473 310
rect 1511 276 1521 310
rect 1521 276 1545 310
rect 1583 276 1589 310
rect 1589 276 1617 310
rect 1655 276 1657 310
rect 1657 276 1689 310
rect 1727 276 1759 310
rect 1759 276 1761 310
rect 1799 276 1827 310
rect 1827 276 1833 310
rect 1882 276 1916 310
rect 2108 2299 2142 2321
rect 2108 2287 2142 2299
rect 2108 2231 2142 2249
rect 2108 2215 2142 2231
rect 2108 2163 2142 2177
rect 2108 2143 2142 2163
rect 2108 2095 2142 2105
rect 2108 2071 2142 2095
rect 2108 2027 2142 2033
rect 2108 1999 2142 2027
rect 2108 1959 2142 1961
rect 2108 1927 2142 1959
rect 2108 1857 2142 1889
rect 2108 1855 2142 1857
rect 2108 1789 2142 1817
rect 2108 1783 2142 1789
rect 2108 1721 2142 1745
rect 2108 1711 2142 1721
rect 2108 1653 2142 1673
rect 2108 1639 2142 1653
rect 2108 1585 2142 1601
rect 2108 1567 2142 1585
rect 2108 1517 2142 1529
rect 2108 1495 2142 1517
rect 2108 1449 2142 1457
rect 2108 1423 2142 1449
rect 2108 1381 2142 1385
rect 2108 1351 2142 1381
rect 2108 1279 2142 1313
rect 2108 1211 2142 1241
rect 2108 1207 2142 1211
rect 2108 1143 2142 1169
rect 2108 1135 2142 1143
rect 2108 1075 2142 1097
rect 2108 1063 2142 1075
rect 2108 1007 2142 1025
rect 2108 991 2142 1007
rect 2108 939 2142 953
rect 2108 919 2142 939
rect 2108 871 2142 881
rect 2108 847 2142 871
rect 2108 803 2142 809
rect 2108 775 2142 803
rect 2108 735 2142 737
rect 2108 703 2142 735
rect 2108 633 2142 665
rect 2108 631 2142 633
rect 2108 565 2142 593
rect 2108 559 2142 565
rect 2108 497 2142 521
rect 2108 487 2142 497
rect 2108 429 2142 449
rect 2108 415 2142 429
rect 2108 361 2142 377
rect 2108 343 2142 361
rect 50 225 84 233
rect 50 199 84 225
rect 50 157 84 161
rect 50 127 84 157
rect 2108 293 2142 305
rect 2108 271 2142 293
rect 2108 225 2142 233
rect 2108 199 2142 225
rect 2108 157 2142 161
rect 2108 127 2142 157
rect 50 50 84 84
rect 143 50 161 84
rect 161 50 177 84
rect 215 50 229 84
rect 229 50 249 84
rect 287 50 297 84
rect 297 50 321 84
rect 359 50 365 84
rect 365 50 393 84
rect 431 50 433 84
rect 433 50 465 84
rect 503 50 535 84
rect 535 50 537 84
rect 575 50 603 84
rect 603 50 609 84
rect 647 50 671 84
rect 671 50 681 84
rect 719 50 739 84
rect 739 50 753 84
rect 791 50 807 84
rect 807 50 825 84
rect 863 50 875 84
rect 875 50 897 84
rect 935 50 943 84
rect 943 50 969 84
rect 1007 50 1011 84
rect 1011 50 1041 84
rect 1079 50 1113 84
rect 1151 50 1181 84
rect 1181 50 1185 84
rect 1223 50 1249 84
rect 1249 50 1257 84
rect 1295 50 1317 84
rect 1317 50 1329 84
rect 1367 50 1385 84
rect 1385 50 1401 84
rect 1439 50 1453 84
rect 1453 50 1473 84
rect 1511 50 1521 84
rect 1521 50 1545 84
rect 1583 50 1589 84
rect 1589 50 1617 84
rect 1655 50 1657 84
rect 1657 50 1689 84
rect 1727 50 1759 84
rect 1759 50 1761 84
rect 1799 50 1827 84
rect 1827 50 1833 84
rect 1871 50 1895 84
rect 1895 50 1905 84
rect 1943 50 1963 84
rect 1963 50 1977 84
rect 2015 50 2031 84
rect 2031 50 2049 84
rect 2108 50 2142 84
<< metal1 >>
rect 38 2542 2154 2554
rect 38 2508 50 2542
rect 84 2508 143 2542
rect 177 2508 215 2542
rect 249 2508 287 2542
rect 321 2508 359 2542
rect 393 2508 431 2542
rect 465 2508 503 2542
rect 537 2508 575 2542
rect 609 2508 647 2542
rect 681 2508 719 2542
rect 753 2508 791 2542
rect 825 2508 863 2542
rect 897 2508 935 2542
rect 969 2508 1007 2542
rect 1041 2508 1079 2542
rect 1113 2508 1151 2542
rect 1185 2508 1223 2542
rect 1257 2508 1295 2542
rect 1329 2508 1367 2542
rect 1401 2508 1439 2542
rect 1473 2508 1511 2542
rect 1545 2508 1583 2542
rect 1617 2508 1655 2542
rect 1689 2508 1727 2542
rect 1761 2508 1799 2542
rect 1833 2508 1871 2542
rect 1905 2508 1943 2542
rect 1977 2508 2015 2542
rect 2049 2508 2108 2542
rect 2142 2508 2154 2542
rect 38 2496 2154 2508
rect 38 2465 96 2496
rect 38 2431 50 2465
rect 84 2431 96 2465
rect 38 2393 96 2431
rect 38 2359 50 2393
rect 84 2359 96 2393
rect 38 2321 96 2359
rect 2096 2465 2154 2496
rect 2096 2431 2108 2465
rect 2142 2431 2154 2465
rect 2096 2393 2154 2431
rect 2096 2359 2108 2393
rect 2142 2359 2154 2393
rect 38 2287 50 2321
rect 84 2287 96 2321
rect 38 2249 96 2287
rect 38 2215 50 2249
rect 84 2215 96 2249
rect 38 2177 96 2215
rect 38 2143 50 2177
rect 84 2143 96 2177
rect 38 2105 96 2143
rect 38 2071 50 2105
rect 84 2071 96 2105
rect 38 2033 96 2071
rect 38 1999 50 2033
rect 84 1999 96 2033
rect 38 1961 96 1999
rect 38 1927 50 1961
rect 84 1927 96 1961
rect 38 1889 96 1927
rect 38 1855 50 1889
rect 84 1855 96 1889
rect 38 1817 96 1855
rect 38 1783 50 1817
rect 84 1783 96 1817
rect 38 1745 96 1783
rect 38 1711 50 1745
rect 84 1711 96 1745
rect 38 1673 96 1711
rect 38 1639 50 1673
rect 84 1639 96 1673
rect 38 1601 96 1639
rect 38 1567 50 1601
rect 84 1567 96 1601
rect 38 1529 96 1567
rect 38 1495 50 1529
rect 84 1495 96 1529
rect 38 1457 96 1495
rect 38 1423 50 1457
rect 84 1423 96 1457
rect 38 1385 96 1423
rect 38 1351 50 1385
rect 84 1351 96 1385
rect 38 1313 96 1351
rect 38 1279 50 1313
rect 84 1279 96 1313
rect 38 1241 96 1279
rect 38 1207 50 1241
rect 84 1207 96 1241
rect 38 1169 96 1207
rect 38 1135 50 1169
rect 84 1135 96 1169
rect 38 1097 96 1135
rect 38 1063 50 1097
rect 84 1063 96 1097
rect 38 1025 96 1063
rect 38 991 50 1025
rect 84 991 96 1025
rect 38 953 96 991
rect 38 919 50 953
rect 84 919 96 953
rect 38 881 96 919
rect 38 847 50 881
rect 84 847 96 881
rect 38 809 96 847
rect 38 775 50 809
rect 84 775 96 809
rect 38 737 96 775
rect 38 703 50 737
rect 84 703 96 737
rect 38 665 96 703
rect 38 631 50 665
rect 84 631 96 665
rect 38 593 96 631
rect 38 559 50 593
rect 84 559 96 593
rect 38 521 96 559
rect 38 487 50 521
rect 84 487 96 521
rect 38 449 96 487
rect 38 415 50 449
rect 84 415 96 449
rect 38 377 96 415
rect 38 343 50 377
rect 84 343 96 377
rect 38 305 96 343
rect 38 271 50 305
rect 84 271 96 305
rect 38 233 96 271
rect 264 2316 1928 2328
rect 264 2282 276 2316
rect 310 2282 359 2316
rect 393 2282 431 2316
rect 465 2282 503 2316
rect 537 2282 575 2316
rect 609 2282 647 2316
rect 681 2282 719 2316
rect 753 2282 791 2316
rect 825 2282 863 2316
rect 897 2282 935 2316
rect 969 2282 1007 2316
rect 1041 2282 1079 2316
rect 1113 2282 1151 2316
rect 1185 2282 1223 2316
rect 1257 2282 1295 2316
rect 1329 2282 1367 2316
rect 1401 2282 1439 2316
rect 1473 2282 1511 2316
rect 1545 2282 1583 2316
rect 1617 2282 1655 2316
rect 1689 2282 1727 2316
rect 1761 2282 1799 2316
rect 1833 2282 1882 2316
rect 1916 2282 1928 2316
rect 264 2270 1928 2282
rect 264 2213 322 2270
rect 264 2179 276 2213
rect 310 2179 322 2213
rect 264 2141 322 2179
rect 264 2107 276 2141
rect 310 2107 322 2141
rect 264 2069 322 2107
rect 264 2035 276 2069
rect 310 2035 322 2069
rect 264 1997 322 2035
rect 264 1963 276 1997
rect 310 1963 322 1997
rect 264 1925 322 1963
rect 1870 2213 1928 2270
rect 1870 2179 1882 2213
rect 1916 2179 1928 2213
rect 1870 2141 1928 2179
rect 1870 2107 1882 2141
rect 1916 2107 1928 2141
rect 1870 2069 1928 2107
rect 1870 2035 1882 2069
rect 1916 2035 1928 2069
rect 1870 1997 1928 2035
rect 1870 1963 1882 1997
rect 1916 1963 1928 1997
rect 264 1891 276 1925
rect 310 1891 322 1925
rect 264 1853 322 1891
rect 264 1819 276 1853
rect 310 1819 322 1853
rect 264 1781 322 1819
rect 264 1747 276 1781
rect 310 1747 322 1781
rect 264 1709 322 1747
rect 264 1675 276 1709
rect 310 1675 322 1709
rect 264 1637 322 1675
rect 264 1603 276 1637
rect 310 1603 322 1637
rect 264 1565 322 1603
rect 264 1531 276 1565
rect 310 1531 322 1565
rect 264 1493 322 1531
rect 264 1459 276 1493
rect 310 1459 322 1493
rect 264 1421 322 1459
rect 264 1387 276 1421
rect 310 1387 322 1421
rect 264 1349 322 1387
rect 264 1315 276 1349
rect 310 1315 322 1349
rect 264 1277 322 1315
rect 264 1243 276 1277
rect 310 1243 322 1277
rect 264 1205 322 1243
rect 264 1171 276 1205
rect 310 1171 322 1205
rect 264 1133 322 1171
rect 264 1099 276 1133
rect 310 1099 322 1133
rect 264 1061 322 1099
rect 264 1027 276 1061
rect 310 1027 322 1061
rect 264 989 322 1027
rect 264 955 276 989
rect 310 955 322 989
rect 264 917 322 955
rect 264 883 276 917
rect 310 883 322 917
rect 264 845 322 883
rect 264 811 276 845
rect 310 811 322 845
rect 264 773 322 811
rect 264 739 276 773
rect 310 739 322 773
rect 264 701 322 739
rect 264 667 276 701
rect 310 667 322 701
rect 264 629 322 667
rect 666 1914 1526 1926
rect 666 1880 678 1914
rect 712 1880 755 1914
rect 789 1880 827 1914
rect 861 1880 899 1914
rect 933 1880 971 1914
rect 1005 1880 1043 1914
rect 1077 1880 1115 1914
rect 1149 1880 1187 1914
rect 1221 1880 1259 1914
rect 1293 1880 1331 1914
rect 1365 1880 1403 1914
rect 1437 1880 1480 1914
rect 1514 1880 1526 1914
rect 666 1868 1526 1880
rect 666 1817 724 1868
rect 666 1783 678 1817
rect 712 1783 724 1817
rect 666 1745 724 1783
rect 666 1711 678 1745
rect 712 1711 724 1745
rect 666 1673 724 1711
rect 666 1639 678 1673
rect 712 1639 724 1673
rect 1468 1817 1526 1868
rect 1468 1783 1480 1817
rect 1514 1783 1526 1817
rect 1468 1745 1526 1783
rect 1468 1711 1480 1745
rect 1514 1711 1526 1745
rect 1468 1673 1526 1711
rect 666 1601 724 1639
rect 666 1567 678 1601
rect 712 1567 724 1601
rect 666 1529 724 1567
rect 666 1495 678 1529
rect 712 1495 724 1529
rect 666 1457 724 1495
rect 666 1423 678 1457
rect 712 1423 724 1457
rect 666 1385 724 1423
rect 666 1351 678 1385
rect 712 1351 724 1385
rect 666 1313 724 1351
rect 666 1279 678 1313
rect 712 1279 724 1313
rect 666 1241 724 1279
rect 666 1207 678 1241
rect 712 1207 724 1241
rect 666 1169 724 1207
rect 666 1135 678 1169
rect 712 1135 724 1169
rect 666 1097 724 1135
rect 666 1063 678 1097
rect 712 1063 724 1097
rect 666 1025 724 1063
rect 666 991 678 1025
rect 712 991 724 1025
rect 666 953 724 991
rect 666 919 678 953
rect 712 919 724 953
rect 923 1637 1269 1649
rect 923 955 935 1637
rect 1257 955 1269 1637
rect 923 943 1269 955
rect 1468 1639 1480 1673
rect 1514 1639 1526 1673
rect 1468 1601 1526 1639
rect 1468 1567 1480 1601
rect 1514 1567 1526 1601
rect 1468 1529 1526 1567
rect 1468 1495 1480 1529
rect 1514 1495 1526 1529
rect 1468 1457 1526 1495
rect 1468 1423 1480 1457
rect 1514 1423 1526 1457
rect 1468 1385 1526 1423
rect 1468 1351 1480 1385
rect 1514 1351 1526 1385
rect 1468 1313 1526 1351
rect 1468 1279 1480 1313
rect 1514 1279 1526 1313
rect 1468 1241 1526 1279
rect 1468 1207 1480 1241
rect 1514 1207 1526 1241
rect 1468 1169 1526 1207
rect 1468 1135 1480 1169
rect 1514 1135 1526 1169
rect 1468 1097 1526 1135
rect 1468 1063 1480 1097
rect 1514 1063 1526 1097
rect 1468 1025 1526 1063
rect 1468 991 1480 1025
rect 1514 991 1526 1025
rect 1468 953 1526 991
rect 666 881 724 919
rect 666 847 678 881
rect 712 847 724 881
rect 666 809 724 847
rect 666 775 678 809
rect 712 775 724 809
rect 666 724 724 775
rect 1468 919 1480 953
rect 1514 919 1526 953
rect 1468 881 1526 919
rect 1468 847 1480 881
rect 1514 847 1526 881
rect 1468 809 1526 847
rect 1468 775 1480 809
rect 1514 775 1526 809
rect 1468 724 1526 775
rect 666 712 1526 724
rect 666 678 678 712
rect 712 678 755 712
rect 789 678 827 712
rect 861 678 899 712
rect 933 678 971 712
rect 1005 678 1043 712
rect 1077 678 1115 712
rect 1149 678 1187 712
rect 1221 678 1259 712
rect 1293 678 1331 712
rect 1365 678 1403 712
rect 1437 678 1480 712
rect 1514 678 1526 712
rect 666 666 1526 678
rect 1870 1925 1928 1963
rect 1870 1891 1882 1925
rect 1916 1891 1928 1925
rect 1870 1853 1928 1891
rect 1870 1819 1882 1853
rect 1916 1819 1928 1853
rect 1870 1781 1928 1819
rect 1870 1747 1882 1781
rect 1916 1747 1928 1781
rect 1870 1709 1928 1747
rect 1870 1675 1882 1709
rect 1916 1675 1928 1709
rect 1870 1637 1928 1675
rect 1870 1603 1882 1637
rect 1916 1603 1928 1637
rect 1870 1565 1928 1603
rect 1870 1531 1882 1565
rect 1916 1531 1928 1565
rect 1870 1493 1928 1531
rect 1870 1459 1882 1493
rect 1916 1459 1928 1493
rect 1870 1421 1928 1459
rect 1870 1387 1882 1421
rect 1916 1387 1928 1421
rect 1870 1349 1928 1387
rect 1870 1315 1882 1349
rect 1916 1315 1928 1349
rect 1870 1277 1928 1315
rect 1870 1243 1882 1277
rect 1916 1243 1928 1277
rect 1870 1205 1928 1243
rect 1870 1171 1882 1205
rect 1916 1171 1928 1205
rect 1870 1133 1928 1171
rect 1870 1099 1882 1133
rect 1916 1099 1928 1133
rect 1870 1061 1928 1099
rect 1870 1027 1882 1061
rect 1916 1027 1928 1061
rect 1870 989 1928 1027
rect 1870 955 1882 989
rect 1916 955 1928 989
rect 1870 917 1928 955
rect 1870 883 1882 917
rect 1916 883 1928 917
rect 1870 845 1928 883
rect 1870 811 1882 845
rect 1916 811 1928 845
rect 1870 773 1928 811
rect 1870 739 1882 773
rect 1916 739 1928 773
rect 1870 701 1928 739
rect 1870 667 1882 701
rect 1916 667 1928 701
rect 264 595 276 629
rect 310 595 322 629
rect 264 557 322 595
rect 264 523 276 557
rect 310 523 322 557
rect 264 485 322 523
rect 264 451 276 485
rect 310 451 322 485
rect 264 413 322 451
rect 264 379 276 413
rect 310 379 322 413
rect 264 322 322 379
rect 1870 629 1928 667
rect 1870 595 1882 629
rect 1916 595 1928 629
rect 1870 557 1928 595
rect 1870 523 1882 557
rect 1916 523 1928 557
rect 1870 485 1928 523
rect 1870 451 1882 485
rect 1916 451 1928 485
rect 1870 413 1928 451
rect 1870 379 1882 413
rect 1916 379 1928 413
rect 1870 322 1928 379
rect 264 310 1928 322
rect 264 276 276 310
rect 310 276 359 310
rect 393 276 431 310
rect 465 276 503 310
rect 537 276 575 310
rect 609 276 647 310
rect 681 276 719 310
rect 753 276 791 310
rect 825 276 863 310
rect 897 276 935 310
rect 969 276 1007 310
rect 1041 276 1079 310
rect 1113 276 1151 310
rect 1185 276 1223 310
rect 1257 276 1295 310
rect 1329 276 1367 310
rect 1401 276 1439 310
rect 1473 276 1511 310
rect 1545 276 1583 310
rect 1617 276 1655 310
rect 1689 276 1727 310
rect 1761 276 1799 310
rect 1833 276 1882 310
rect 1916 276 1928 310
rect 264 264 1928 276
rect 2096 2321 2154 2359
rect 2096 2287 2108 2321
rect 2142 2287 2154 2321
rect 2096 2249 2154 2287
rect 2096 2215 2108 2249
rect 2142 2215 2154 2249
rect 2096 2177 2154 2215
rect 2096 2143 2108 2177
rect 2142 2143 2154 2177
rect 2096 2105 2154 2143
rect 2096 2071 2108 2105
rect 2142 2071 2154 2105
rect 2096 2033 2154 2071
rect 2096 1999 2108 2033
rect 2142 1999 2154 2033
rect 2096 1961 2154 1999
rect 2096 1927 2108 1961
rect 2142 1927 2154 1961
rect 2096 1889 2154 1927
rect 2096 1855 2108 1889
rect 2142 1855 2154 1889
rect 2096 1817 2154 1855
rect 2096 1783 2108 1817
rect 2142 1783 2154 1817
rect 2096 1745 2154 1783
rect 2096 1711 2108 1745
rect 2142 1711 2154 1745
rect 2096 1673 2154 1711
rect 2096 1639 2108 1673
rect 2142 1639 2154 1673
rect 2096 1601 2154 1639
rect 2096 1567 2108 1601
rect 2142 1567 2154 1601
rect 2096 1529 2154 1567
rect 2096 1495 2108 1529
rect 2142 1495 2154 1529
rect 2096 1457 2154 1495
rect 2096 1423 2108 1457
rect 2142 1423 2154 1457
rect 2096 1385 2154 1423
rect 2096 1351 2108 1385
rect 2142 1351 2154 1385
rect 2096 1313 2154 1351
rect 2096 1279 2108 1313
rect 2142 1279 2154 1313
rect 2096 1241 2154 1279
rect 2096 1207 2108 1241
rect 2142 1207 2154 1241
rect 2096 1169 2154 1207
rect 2096 1135 2108 1169
rect 2142 1135 2154 1169
rect 2096 1097 2154 1135
rect 2096 1063 2108 1097
rect 2142 1063 2154 1097
rect 2096 1025 2154 1063
rect 2096 991 2108 1025
rect 2142 991 2154 1025
rect 2096 953 2154 991
rect 2096 919 2108 953
rect 2142 919 2154 953
rect 2096 881 2154 919
rect 2096 847 2108 881
rect 2142 847 2154 881
rect 2096 809 2154 847
rect 2096 775 2108 809
rect 2142 775 2154 809
rect 2096 737 2154 775
rect 2096 703 2108 737
rect 2142 703 2154 737
rect 2096 665 2154 703
rect 2096 631 2108 665
rect 2142 631 2154 665
rect 2096 593 2154 631
rect 2096 559 2108 593
rect 2142 559 2154 593
rect 2096 521 2154 559
rect 2096 487 2108 521
rect 2142 487 2154 521
rect 2096 449 2154 487
rect 2096 415 2108 449
rect 2142 415 2154 449
rect 2096 377 2154 415
rect 2096 343 2108 377
rect 2142 343 2154 377
rect 2096 305 2154 343
rect 2096 271 2108 305
rect 2142 271 2154 305
rect 38 199 50 233
rect 84 199 96 233
rect 38 161 96 199
rect 38 127 50 161
rect 84 127 96 161
rect 38 96 96 127
rect 2096 233 2154 271
rect 2096 199 2108 233
rect 2142 199 2154 233
rect 2096 161 2154 199
rect 2096 127 2108 161
rect 2142 127 2154 161
rect 2096 96 2154 127
rect 38 84 2154 96
rect 38 50 50 84
rect 84 50 143 84
rect 177 50 215 84
rect 249 50 287 84
rect 321 50 359 84
rect 393 50 431 84
rect 465 50 503 84
rect 537 50 575 84
rect 609 50 647 84
rect 681 50 719 84
rect 753 50 791 84
rect 825 50 863 84
rect 897 50 935 84
rect 969 50 1007 84
rect 1041 50 1079 84
rect 1113 50 1151 84
rect 1185 50 1223 84
rect 1257 50 1295 84
rect 1329 50 1367 84
rect 1401 50 1439 84
rect 1473 50 1511 84
rect 1545 50 1583 84
rect 1617 50 1655 84
rect 1689 50 1727 84
rect 1761 50 1799 84
rect 1833 50 1871 84
rect 1905 50 1943 84
rect 1977 50 2015 84
rect 2049 50 2108 84
rect 2142 50 2154 84
rect 38 38 2154 50
<< properties >>
string GDS_END 8926674
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8873862
string path 7.850 12.350 7.850 56.950 46.950 56.950 46.950 7.850 3.350 7.850 
<< end >>
