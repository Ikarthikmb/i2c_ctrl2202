magic
tech sky130A
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_0
timestamp 1644511149
transform 1 0 30 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_1
timestamp 1644511149
transform 1 0 116 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_2
timestamp 1644511149
transform 1 0 202 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_3
timestamp 1644511149
transform 1 0 288 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 316 97 316 97 0 FreeSans 300 0 0 0 D
flabel comment s 230 97 230 97 0 FreeSans 300 0 0 0 S
flabel comment s 144 97 144 97 0 FreeSans 300 0 0 0 D
flabel comment s 58 97 58 97 0 FreeSans 300 0 0 0 S
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 6768094
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6765612
<< end >>
