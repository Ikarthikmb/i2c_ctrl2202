magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 2 21 1088 203
rect 29 -17 63 21
<< locali >>
rect 180 370 428 421
rect 25 289 360 336
rect 394 325 428 370
rect 394 289 651 325
rect 25 209 91 289
rect 323 255 360 289
rect 151 215 285 255
rect 323 206 395 255
rect 437 206 571 255
rect 605 169 651 289
rect 693 289 1058 335
rect 693 197 743 289
rect 794 203 945 255
rect 979 199 1058 289
rect 24 161 651 169
rect 24 123 1071 161
rect 24 51 76 123
rect 210 51 259 123
rect 393 51 459 123
rect 593 55 659 123
rect 1004 59 1071 123
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 20 459 597 493
rect 20 455 437 459
rect 20 374 92 455
rect 563 427 597 459
rect 631 419 704 493
rect 738 455 804 527
rect 838 421 880 493
rect 914 455 980 527
rect 1014 421 1080 493
rect 838 419 1080 421
rect 462 393 528 412
rect 631 393 1080 419
rect 462 369 1080 393
rect 462 359 667 369
rect 110 17 176 89
rect 293 17 359 89
rect 493 17 559 89
rect 825 17 891 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
<< metal1 >>
rect 0 561 1104 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1104 561
rect 0 496 1104 527
rect 0 17 1104 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1104 17
rect 0 -48 1104 -17
<< labels >>
rlabel locali s 979 199 1058 289 6 A1
port 1 nsew signal input
rlabel locali s 693 197 743 289 6 A1
port 1 nsew signal input
rlabel locali s 693 289 1058 335 6 A1
port 1 nsew signal input
rlabel locali s 794 203 945 255 6 A2
port 2 nsew signal input
rlabel locali s 437 206 571 255 6 B1
port 3 nsew signal input
rlabel locali s 323 206 395 255 6 C1
port 4 nsew signal input
rlabel locali s 323 255 360 289 6 C1
port 4 nsew signal input
rlabel locali s 25 209 91 289 6 C1
port 4 nsew signal input
rlabel locali s 25 289 360 336 6 C1
port 4 nsew signal input
rlabel locali s 151 215 285 255 6 D1
port 5 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 2 21 1088 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 1004 59 1071 123 6 Y
port 10 nsew signal output
rlabel locali s 593 55 659 123 6 Y
port 10 nsew signal output
rlabel locali s 393 51 459 123 6 Y
port 10 nsew signal output
rlabel locali s 210 51 259 123 6 Y
port 10 nsew signal output
rlabel locali s 24 51 76 123 6 Y
port 10 nsew signal output
rlabel locali s 24 123 1071 161 6 Y
port 10 nsew signal output
rlabel locali s 24 161 651 169 6 Y
port 10 nsew signal output
rlabel locali s 605 169 651 289 6 Y
port 10 nsew signal output
rlabel locali s 394 289 651 325 6 Y
port 10 nsew signal output
rlabel locali s 394 325 428 370 6 Y
port 10 nsew signal output
rlabel locali s 180 370 428 421 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3799438
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3791210
<< end >>
