/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/sky130A/libs.tech/ngspice/corners/ss.spice