magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< metal1 >>
rect 15240 14951 17187 15070
rect 15240 5427 15324 14951
rect 17040 9639 17187 14951
rect 17104 5427 17187 9639
rect 5101 -7 5685 83
rect 4185 -163 11313 -7
rect 15240 -163 17187 5427
rect 4185 -1384 17187 -163
rect 4185 -2184 16387 -1384
tri 16387 -2184 17187 -1384 nw
<< via1 >>
rect 15324 9639 17040 14951
rect 15324 5427 17104 9639
<< metal2 >>
rect 15240 39515 17187 39586
rect 15240 34819 15307 39515
rect 17123 34819 17187 39515
rect 15240 14951 17187 34819
rect 15240 5613 15324 14951
rect 17040 9639 17187 14951
rect 17104 5613 17187 9639
rect 15240 4837 15298 5613
rect 17114 4837 17187 5613
rect 15240 4678 17187 4837
<< via2 >>
rect 15307 34819 17123 39515
rect 15298 5427 15324 5613
rect 15324 5427 17104 5613
rect 17104 5427 17114 5613
rect 15298 4837 17114 5427
<< metal3 >>
rect 15240 39519 17187 39586
rect 15240 34815 15303 39519
rect 17127 34815 17187 39519
rect 15240 34743 17187 34815
rect 15240 5617 17187 5683
rect 15240 4833 15294 5617
rect 17118 4833 17187 5617
rect 15240 4753 17187 4833
<< via3 >>
rect 15303 39515 17127 39519
rect 15303 34819 15307 39515
rect 15307 34819 17123 39515
rect 17123 34819 17127 39515
rect 15303 34815 17127 34819
rect 15294 5613 17118 5617
rect 15294 4837 15298 5613
rect 15298 4837 17114 5613
rect 17114 4837 17118 5613
rect 15294 4833 17118 4837
<< metal4 >>
rect 14957 39519 17187 39586
rect 14957 34815 15303 39519
rect 17127 34815 17187 39519
rect 14957 34743 17187 34815
rect 14987 5617 17187 5683
rect 14987 4833 15294 5617
rect 17118 4833 17187 5617
rect 14987 4753 17187 4833
<< properties >>
string FIXED_BBOX 0 -7 15000 39593
string GDS_END 465730
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_ef_io.gds
string GDS_START 134
<< end >>
