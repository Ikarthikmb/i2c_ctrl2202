magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 1 21 1491 203
rect 30 -17 64 21
<< locali >>
rect 119 349 153 493
rect 287 349 321 493
rect 30 315 321 349
rect 30 161 64 315
rect 427 215 629 256
rect 679 215 813 259
rect 855 215 995 257
rect 1031 215 1237 259
rect 1299 215 1501 259
rect 30 127 321 161
rect 119 51 153 127
rect 287 51 321 127
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 19 383 85 527
rect 187 383 253 527
rect 355 383 425 527
rect 475 459 681 493
rect 475 359 509 459
rect 543 391 609 425
rect 559 325 593 391
rect 355 291 593 325
rect 647 341 681 459
rect 715 383 781 527
rect 815 341 849 493
rect 883 383 949 527
rect 987 341 1021 493
rect 1069 383 1207 527
rect 1255 341 1289 493
rect 1323 383 1389 527
rect 1423 341 1457 493
rect 647 307 1474 341
rect 355 249 389 291
rect 98 215 389 249
rect 355 163 389 215
rect 355 129 781 163
rect 815 129 1033 163
rect 1071 129 1457 163
rect 19 17 85 93
rect 187 17 253 93
rect 355 17 425 93
rect 459 51 493 129
rect 815 93 849 129
rect 527 17 593 93
rect 631 59 849 93
rect 883 59 1221 93
rect 1323 17 1389 93
rect 1423 51 1457 129
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
rlabel locali s 679 215 813 259 6 A1
port 1 nsew signal input
rlabel locali s 855 215 995 257 6 A2
port 2 nsew signal input
rlabel locali s 1031 215 1237 259 6 A3
port 3 nsew signal input
rlabel locali s 1299 215 1501 259 6 A4
port 4 nsew signal input
rlabel locali s 427 215 629 256 6 B1
port 5 nsew signal input
rlabel metal1 s 0 -48 1564 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1491 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1602 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1564 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 287 51 321 127 6 X
port 10 nsew signal output
rlabel locali s 119 51 153 127 6 X
port 10 nsew signal output
rlabel locali s 30 127 321 161 6 X
port 10 nsew signal output
rlabel locali s 30 161 64 315 6 X
port 10 nsew signal output
rlabel locali s 30 315 321 349 6 X
port 10 nsew signal output
rlabel locali s 287 349 321 493 6 X
port 10 nsew signal output
rlabel locali s 119 349 153 493 6 X
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1564 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3542148
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3529682
<< end >>
