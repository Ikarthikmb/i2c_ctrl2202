magic
tech sky130A
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_0
timestamp 1644511149
transform -1 0 -40 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_1
timestamp 1644511149
transform 1 0 314 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_2
timestamp 1644511149
transform 1 0 868 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_3
timestamp 1644511149
transform 1 0 1422 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_4
timestamp 1644511149
transform 1 0 1976 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_5
timestamp 1644511149
transform 1 0 2530 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_6
timestamp 1644511149
transform 1 0 3084 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_7
timestamp 1644511149
transform 1 0 3638 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_8
timestamp 1644511149
transform 1 0 4192 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_9
timestamp 1644511149
transform 1 0 4746 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_10
timestamp 1644511149
transform 1 0 5300 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_11
timestamp 1644511149
transform 1 0 5854 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_12
timestamp 1644511149
transform 1 0 6408 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_13
timestamp 1644511149
transform 1 0 6962 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_14
timestamp 1644511149
transform 1 0 7516 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_15
timestamp 1644511149
transform 1 0 8070 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_16
timestamp 1644511149
transform 1 0 8624 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_17
timestamp 1644511149
transform 1 0 9178 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_18
timestamp 1644511149
transform 1 0 9732 0 1 0
box 0 0 1 1
use sky130_fd_pr__dftpl1s2__example_55959141808694  sky130_fd_pr__dftpl1s2__example_55959141808694_19
timestamp 1644511149
transform 1 0 10286 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 10386 471 10386 471 0 FreeSans 300 0 0 0 S
flabel comment s 10109 500 10109 500 0 FreeSans 300 0 0 0 D
flabel comment s 9832 471 9832 471 0 FreeSans 300 0 0 0 S
flabel comment s 9555 500 9555 500 0 FreeSans 300 0 0 0 D
flabel comment s 9278 471 9278 471 0 FreeSans 300 0 0 0 S
flabel comment s 9001 500 9001 500 0 FreeSans 300 0 0 0 D
flabel comment s 8724 471 8724 471 0 FreeSans 300 0 0 0 S
flabel comment s 8447 500 8447 500 0 FreeSans 300 0 0 0 D
flabel comment s 8170 471 8170 471 0 FreeSans 300 0 0 0 S
flabel comment s 7893 500 7893 500 0 FreeSans 300 0 0 0 D
flabel comment s 7616 471 7616 471 0 FreeSans 300 0 0 0 S
flabel comment s 7339 500 7339 500 0 FreeSans 300 0 0 0 D
flabel comment s 7062 471 7062 471 0 FreeSans 300 0 0 0 S
flabel comment s 6785 500 6785 500 0 FreeSans 300 0 0 0 D
flabel comment s 6508 471 6508 471 0 FreeSans 300 0 0 0 S
flabel comment s 6231 500 6231 500 0 FreeSans 300 0 0 0 D
flabel comment s 5954 471 5954 471 0 FreeSans 300 0 0 0 S
flabel comment s 5677 500 5677 500 0 FreeSans 300 0 0 0 D
flabel comment s 5400 471 5400 471 0 FreeSans 300 0 0 0 S
flabel comment s 5123 500 5123 500 0 FreeSans 300 0 0 0 D
flabel comment s 4846 471 4846 471 0 FreeSans 300 0 0 0 S
flabel comment s 4569 500 4569 500 0 FreeSans 300 0 0 0 D
flabel comment s 4292 471 4292 471 0 FreeSans 300 0 0 0 S
flabel comment s 4015 500 4015 500 0 FreeSans 300 0 0 0 D
flabel comment s 3738 471 3738 471 0 FreeSans 300 0 0 0 S
flabel comment s 3461 500 3461 500 0 FreeSans 300 0 0 0 D
flabel comment s 3184 471 3184 471 0 FreeSans 300 0 0 0 S
flabel comment s 2907 500 2907 500 0 FreeSans 300 0 0 0 D
flabel comment s 2630 471 2630 471 0 FreeSans 300 0 0 0 S
flabel comment s 2353 500 2353 500 0 FreeSans 300 0 0 0 D
flabel comment s 2076 471 2076 471 0 FreeSans 300 0 0 0 S
flabel comment s 1799 500 1799 500 0 FreeSans 300 0 0 0 D
flabel comment s 1522 471 1522 471 0 FreeSans 300 0 0 0 S
flabel comment s 1245 500 1245 500 0 FreeSans 300 0 0 0 D
flabel comment s 968 471 968 471 0 FreeSans 300 0 0 0 S
flabel comment s 691 500 691 500 0 FreeSans 300 0 0 0 D
flabel comment s 414 471 414 471 0 FreeSans 300 0 0 0 S
flabel comment s 137 500 137 500 0 FreeSans 300 0 0 0 D
flabel comment s -140 471 -140 471 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 15462022
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15442182
<< end >>
