magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< obsli1 >>
rect 98 1119 368 1135
rect 98 1085 108 1119
rect 142 1085 180 1119
rect 214 1085 252 1119
rect 286 1085 324 1119
rect 358 1085 368 1119
rect 98 1067 368 1085
rect 44 983 78 1021
rect 44 911 78 949
rect 44 839 78 877
rect 44 767 78 805
rect 44 695 78 733
rect 44 623 78 661
rect 44 551 78 589
rect 44 479 78 517
rect 44 407 78 445
rect 44 335 78 373
rect 44 263 78 301
rect 44 191 78 229
rect 44 119 78 157
rect 44 51 78 85
rect 130 51 164 1021
rect 216 983 250 1021
rect 216 911 250 949
rect 216 839 250 877
rect 216 767 250 805
rect 216 695 250 733
rect 216 623 250 661
rect 216 551 250 589
rect 216 479 250 517
rect 216 407 250 445
rect 216 335 250 373
rect 216 263 250 301
rect 216 191 250 229
rect 216 119 250 157
rect 216 51 250 85
rect 302 51 336 1021
rect 388 983 422 1021
rect 388 911 422 949
rect 388 839 422 877
rect 388 767 422 805
rect 388 695 422 733
rect 388 623 422 661
rect 388 551 422 589
rect 388 479 422 517
rect 388 407 422 445
rect 388 335 422 373
rect 388 263 422 301
rect 388 191 422 229
rect 388 119 422 157
rect 388 51 422 85
<< obsli1c >>
rect 108 1085 142 1119
rect 180 1085 214 1119
rect 252 1085 286 1119
rect 324 1085 358 1119
rect 44 949 78 983
rect 44 877 78 911
rect 44 805 78 839
rect 44 733 78 767
rect 44 661 78 695
rect 44 589 78 623
rect 44 517 78 551
rect 44 445 78 479
rect 44 373 78 407
rect 44 301 78 335
rect 44 229 78 263
rect 44 157 78 191
rect 44 85 78 119
rect 216 949 250 983
rect 216 877 250 911
rect 216 805 250 839
rect 216 733 250 767
rect 216 661 250 695
rect 216 589 250 623
rect 216 517 250 551
rect 216 445 250 479
rect 216 373 250 407
rect 216 301 250 335
rect 216 229 250 263
rect 216 157 250 191
rect 216 85 250 119
rect 388 949 422 983
rect 388 877 422 911
rect 388 805 422 839
rect 388 733 422 767
rect 388 661 422 695
rect 388 589 422 623
rect 388 517 422 551
rect 388 445 422 479
rect 388 373 422 407
rect 388 301 422 335
rect 388 229 422 263
rect 388 157 422 191
rect 388 85 422 119
<< metal1 >>
rect 96 1119 370 1131
rect 96 1085 108 1119
rect 142 1085 180 1119
rect 214 1085 252 1119
rect 286 1085 324 1119
rect 358 1085 370 1119
rect 96 1073 370 1085
rect 38 983 84 1021
rect 38 949 44 983
rect 78 949 84 983
rect 38 911 84 949
rect 38 877 44 911
rect 78 877 84 911
rect 38 839 84 877
rect 38 805 44 839
rect 78 805 84 839
rect 38 767 84 805
rect 38 733 44 767
rect 78 733 84 767
rect 38 695 84 733
rect 38 661 44 695
rect 78 661 84 695
rect 38 623 84 661
rect 38 589 44 623
rect 78 589 84 623
rect 38 551 84 589
rect 38 517 44 551
rect 78 517 84 551
rect 38 479 84 517
rect 38 445 44 479
rect 78 445 84 479
rect 38 407 84 445
rect 38 373 44 407
rect 78 373 84 407
rect 38 335 84 373
rect 38 301 44 335
rect 78 301 84 335
rect 38 263 84 301
rect 38 229 44 263
rect 78 229 84 263
rect 38 191 84 229
rect 38 157 44 191
rect 78 157 84 191
rect 38 119 84 157
rect 38 85 44 119
rect 78 85 84 119
rect 38 -45 84 85
rect 210 983 256 1021
rect 210 949 216 983
rect 250 949 256 983
rect 210 911 256 949
rect 210 877 216 911
rect 250 877 256 911
rect 210 839 256 877
rect 210 805 216 839
rect 250 805 256 839
rect 210 767 256 805
rect 210 733 216 767
rect 250 733 256 767
rect 210 695 256 733
rect 210 661 216 695
rect 250 661 256 695
rect 210 623 256 661
rect 210 589 216 623
rect 250 589 256 623
rect 210 551 256 589
rect 210 517 216 551
rect 250 517 256 551
rect 210 479 256 517
rect 210 445 216 479
rect 250 445 256 479
rect 210 407 256 445
rect 210 373 216 407
rect 250 373 256 407
rect 210 335 256 373
rect 210 301 216 335
rect 250 301 256 335
rect 210 263 256 301
rect 210 229 216 263
rect 250 229 256 263
rect 210 191 256 229
rect 210 157 216 191
rect 250 157 256 191
rect 210 119 256 157
rect 210 85 216 119
rect 250 85 256 119
rect 210 -45 256 85
rect 382 983 428 1021
rect 382 949 388 983
rect 422 949 428 983
rect 382 911 428 949
rect 382 877 388 911
rect 422 877 428 911
rect 382 839 428 877
rect 382 805 388 839
rect 422 805 428 839
rect 382 767 428 805
rect 382 733 388 767
rect 422 733 428 767
rect 382 695 428 733
rect 382 661 388 695
rect 422 661 428 695
rect 382 623 428 661
rect 382 589 388 623
rect 422 589 428 623
rect 382 551 428 589
rect 382 517 388 551
rect 422 517 428 551
rect 382 479 428 517
rect 382 445 388 479
rect 422 445 428 479
rect 382 407 428 445
rect 382 373 388 407
rect 422 373 428 407
rect 382 335 428 373
rect 382 301 388 335
rect 422 301 428 335
rect 382 263 428 301
rect 382 229 388 263
rect 422 229 428 263
rect 382 191 428 229
rect 382 157 388 191
rect 422 157 428 191
rect 382 119 428 157
rect 382 85 388 119
rect 422 85 428 119
rect 382 -45 428 85
rect 38 -97 428 -45
<< obsm1 >>
rect 121 51 173 1021
rect 293 51 345 1021
<< obsm2 >>
rect 114 875 180 1029
rect 286 875 352 1029
<< metal3 >>
rect 114 963 352 1029
rect 114 875 180 963
rect 286 875 352 963
<< labels >>
rlabel metal3 s 286 875 352 963 6 DRAIN
port 1 nsew
rlabel metal3 s 114 963 352 1029 6 DRAIN
port 1 nsew
rlabel metal3 s 114 875 180 963 6 DRAIN
port 1 nsew
rlabel metal1 s 96 1073 370 1131 6 GATE
port 2 nsew
rlabel metal1 s 382 -45 428 1021 6 SOURCE
port 3 nsew
rlabel metal1 s 210 -45 256 1021 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -45 84 1021 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -97 428 -45 8 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 -97 466 1135
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9269534
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9255814
<< end >>
