/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/open_pdks/sky130/custom/sky130_fd_io/spice/sky130_fd_io.spice