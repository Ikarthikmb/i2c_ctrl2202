/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/res_high_po/sky130_fd_pr__res_high_po_0p35.model.spice