magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1326 582
<< pwell >>
rect 79 21 1287 203
rect 29 -17 63 17
<< scnmos >>
rect 158 47 188 177
rect 244 47 274 177
rect 330 47 360 177
rect 419 47 449 177
rect 506 47 536 177
rect 600 47 630 177
rect 697 47 727 177
rect 805 47 835 177
rect 921 47 951 177
rect 1007 47 1037 177
rect 1093 47 1123 177
rect 1179 47 1209 177
<< scpmoshvt >>
rect 79 297 109 497
rect 165 297 195 497
rect 251 297 281 497
rect 337 297 367 497
rect 525 297 555 497
rect 611 297 641 497
rect 697 297 727 497
rect 791 297 821 497
rect 899 297 929 497
rect 1007 297 1037 497
rect 1093 297 1123 497
rect 1179 297 1209 497
<< ndiff >>
rect 105 93 158 177
rect 105 59 113 93
rect 147 59 158 93
rect 105 47 158 59
rect 188 101 244 177
rect 188 67 199 101
rect 233 67 244 101
rect 188 47 244 67
rect 274 89 330 177
rect 274 55 285 89
rect 319 55 330 89
rect 274 47 330 55
rect 360 101 419 177
rect 360 67 371 101
rect 405 67 419 101
rect 360 47 419 67
rect 449 89 506 177
rect 449 55 461 89
rect 495 55 506 89
rect 449 47 506 55
rect 536 114 600 177
rect 536 80 547 114
rect 581 80 600 114
rect 536 47 600 80
rect 630 89 697 177
rect 630 55 644 89
rect 678 55 697 89
rect 630 47 697 55
rect 727 161 805 177
rect 727 127 750 161
rect 784 127 805 161
rect 727 93 805 127
rect 727 59 750 93
rect 784 59 805 93
rect 727 47 805 59
rect 835 89 921 177
rect 835 55 854 89
rect 888 55 921 89
rect 835 47 921 55
rect 951 47 1007 177
rect 1037 157 1093 177
rect 1037 123 1048 157
rect 1082 123 1093 157
rect 1037 89 1093 123
rect 1037 55 1048 89
rect 1082 55 1093 89
rect 1037 47 1093 55
rect 1123 47 1179 177
rect 1209 161 1261 177
rect 1209 127 1219 161
rect 1253 127 1261 161
rect 1209 93 1261 127
rect 1209 59 1219 93
rect 1253 59 1261 93
rect 1209 47 1261 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 409 79 451
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 477 165 497
rect 109 443 120 477
rect 154 443 165 477
rect 109 388 165 443
rect 109 354 120 388
rect 154 354 165 388
rect 109 297 165 354
rect 195 485 251 497
rect 195 451 206 485
rect 240 451 251 485
rect 195 409 251 451
rect 195 375 206 409
rect 240 375 251 409
rect 195 297 251 375
rect 281 477 337 497
rect 281 443 292 477
rect 326 443 337 477
rect 281 388 337 443
rect 281 354 292 388
rect 326 354 337 388
rect 281 297 337 354
rect 367 485 419 497
rect 367 451 377 485
rect 411 451 419 485
rect 367 417 419 451
rect 367 383 377 417
rect 411 383 419 417
rect 367 297 419 383
rect 473 485 525 497
rect 473 451 481 485
rect 515 451 525 485
rect 473 297 525 451
rect 555 297 611 497
rect 641 408 697 497
rect 641 374 652 408
rect 686 374 697 408
rect 641 297 697 374
rect 727 297 791 497
rect 821 485 899 497
rect 821 451 840 485
rect 874 451 899 485
rect 821 417 899 451
rect 821 383 840 417
rect 874 383 899 417
rect 821 297 899 383
rect 929 489 1007 497
rect 929 455 940 489
rect 974 455 1007 489
rect 929 297 1007 455
rect 1037 477 1093 497
rect 1037 443 1048 477
rect 1082 443 1093 477
rect 1037 297 1093 443
rect 1123 489 1179 497
rect 1123 455 1134 489
rect 1168 455 1179 489
rect 1123 297 1179 455
rect 1209 477 1261 497
rect 1209 443 1219 477
rect 1253 443 1261 477
rect 1209 343 1261 443
rect 1209 309 1219 343
rect 1253 309 1261 343
rect 1209 297 1261 309
<< ndiffc >>
rect 113 59 147 93
rect 199 67 233 101
rect 285 55 319 89
rect 371 67 405 101
rect 461 55 495 89
rect 547 80 581 114
rect 644 55 678 89
rect 750 127 784 161
rect 750 59 784 93
rect 854 55 888 89
rect 1048 123 1082 157
rect 1048 55 1082 89
rect 1219 127 1253 161
rect 1219 59 1253 93
<< pdiffc >>
rect 35 451 69 485
rect 35 375 69 409
rect 120 443 154 477
rect 120 354 154 388
rect 206 451 240 485
rect 206 375 240 409
rect 292 443 326 477
rect 292 354 326 388
rect 377 451 411 485
rect 377 383 411 417
rect 481 451 515 485
rect 652 374 686 408
rect 840 451 874 485
rect 840 383 874 417
rect 940 455 974 489
rect 1048 443 1082 477
rect 1134 455 1168 489
rect 1219 443 1253 477
rect 1219 309 1253 343
<< poly >>
rect 79 497 109 523
rect 165 497 195 523
rect 251 497 281 523
rect 337 497 367 523
rect 525 497 555 523
rect 611 497 641 523
rect 697 497 727 523
rect 791 497 821 523
rect 899 497 929 523
rect 1007 497 1037 523
rect 1093 497 1123 523
rect 1179 497 1209 523
rect 79 270 109 297
rect 165 270 195 297
rect 251 270 281 297
rect 337 270 367 297
rect 525 270 555 297
rect 611 271 641 297
rect 697 271 727 297
rect 79 249 449 270
rect 79 215 131 249
rect 165 215 199 249
rect 233 215 267 249
rect 301 215 335 249
rect 369 215 449 249
rect 79 204 449 215
rect 492 249 558 270
rect 492 215 508 249
rect 542 215 558 249
rect 492 204 558 215
rect 600 249 727 271
rect 791 270 821 297
rect 899 280 929 297
rect 600 215 611 249
rect 645 215 679 249
rect 713 215 727 249
rect 158 177 188 204
rect 244 177 274 204
rect 330 177 360 204
rect 419 177 449 204
rect 506 177 536 204
rect 600 198 727 215
rect 600 177 630 198
rect 697 177 727 198
rect 769 249 835 270
rect 769 215 785 249
rect 819 215 835 249
rect 769 197 835 215
rect 899 249 965 280
rect 899 215 915 249
rect 949 215 965 249
rect 899 204 965 215
rect 1007 270 1037 297
rect 1093 270 1123 297
rect 1007 249 1123 270
rect 1007 215 1023 249
rect 1057 215 1123 249
rect 1007 204 1123 215
rect 805 177 835 197
rect 921 177 951 204
rect 1007 177 1037 204
rect 1093 177 1123 204
rect 1179 270 1209 297
rect 1179 249 1245 270
rect 1179 215 1195 249
rect 1229 215 1245 249
rect 1179 202 1245 215
rect 1179 177 1209 202
rect 158 21 188 47
rect 244 21 274 47
rect 330 21 360 47
rect 419 21 449 47
rect 506 21 536 47
rect 600 21 630 47
rect 697 21 727 47
rect 805 21 835 47
rect 921 21 951 47
rect 1007 21 1037 47
rect 1093 21 1123 47
rect 1179 21 1209 47
<< polycont >>
rect 131 215 165 249
rect 199 215 233 249
rect 267 215 301 249
rect 335 215 369 249
rect 508 215 542 249
rect 611 215 645 249
rect 679 215 713 249
rect 785 215 819 249
rect 915 215 949 249
rect 1023 215 1057 249
rect 1195 215 1229 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 18 485 85 527
rect 18 451 35 485
rect 69 451 85 485
rect 18 409 85 451
rect 18 375 35 409
rect 69 375 85 409
rect 119 477 156 493
rect 119 443 120 477
rect 154 443 156 477
rect 119 388 156 443
rect 119 354 120 388
rect 154 354 156 388
rect 190 485 256 527
rect 190 451 206 485
rect 240 451 256 485
rect 190 409 256 451
rect 190 375 206 409
rect 240 375 256 409
rect 290 477 328 493
rect 290 443 292 477
rect 326 443 328 477
rect 290 388 328 443
rect 119 341 156 354
rect 290 354 292 388
rect 326 354 328 388
rect 362 485 412 527
rect 362 451 377 485
rect 411 451 412 485
rect 362 417 412 451
rect 464 485 890 493
rect 464 451 481 485
rect 515 451 840 485
rect 874 451 890 485
rect 924 489 990 527
rect 924 455 940 489
rect 974 455 990 489
rect 1032 477 1084 493
rect 464 442 890 451
rect 362 383 377 417
rect 411 383 412 417
rect 824 421 890 442
rect 1032 443 1048 477
rect 1082 443 1084 477
rect 1118 489 1184 527
rect 1118 455 1134 489
rect 1168 455 1184 489
rect 1218 477 1269 493
rect 1032 421 1084 443
rect 1218 443 1219 477
rect 1253 443 1269 477
rect 1218 421 1269 443
rect 824 417 1269 421
rect 362 367 412 383
rect 456 374 652 408
rect 686 374 702 408
rect 824 383 840 417
rect 874 383 1269 417
rect 824 376 1269 383
rect 290 341 328 354
rect 17 299 328 341
rect 456 335 491 374
rect 1203 343 1269 376
rect 437 301 491 335
rect 17 175 68 299
rect 437 265 474 301
rect 525 289 835 340
rect 525 265 561 289
rect 105 249 474 265
rect 105 215 131 249
rect 165 215 199 249
rect 233 215 267 249
rect 301 215 335 249
rect 369 215 474 249
rect 105 209 474 215
rect 17 127 405 175
rect 197 123 405 127
rect 439 161 474 209
rect 508 249 561 265
rect 542 215 561 249
rect 508 197 561 215
rect 595 249 729 255
rect 595 215 611 249
rect 645 215 679 249
rect 713 215 729 249
rect 595 197 729 215
rect 769 249 835 289
rect 769 215 785 249
rect 819 215 835 249
rect 769 197 835 215
rect 899 302 1169 340
rect 1203 309 1219 343
rect 1253 309 1269 343
rect 1203 307 1269 309
rect 899 249 965 302
rect 899 215 915 249
rect 949 215 965 249
rect 899 204 965 215
rect 1007 249 1076 266
rect 1007 215 1023 249
rect 1057 215 1076 249
rect 1007 204 1076 215
rect 1127 264 1169 302
rect 1127 249 1245 264
rect 1127 215 1195 249
rect 1229 215 1245 249
rect 1127 204 1245 215
rect 439 127 750 161
rect 784 157 1098 161
rect 784 127 1048 157
rect 439 123 1048 127
rect 1082 123 1098 157
rect 197 101 235 123
rect 97 59 113 93
rect 147 59 163 93
rect 97 17 163 59
rect 197 67 199 101
rect 233 67 235 101
rect 369 101 405 123
rect 197 51 235 67
rect 269 55 285 89
rect 319 55 335 89
rect 269 17 335 55
rect 369 67 371 101
rect 545 114 594 123
rect 369 51 405 67
rect 444 55 461 89
rect 495 55 511 89
rect 444 17 511 55
rect 545 80 547 114
rect 581 80 594 114
rect 728 93 804 123
rect 545 51 594 80
rect 628 55 644 89
rect 678 55 694 89
rect 628 17 694 55
rect 728 59 750 93
rect 784 59 804 93
rect 1032 89 1098 123
rect 728 51 804 59
rect 838 55 854 89
rect 888 55 912 89
rect 1032 55 1048 89
rect 1082 55 1098 89
rect 1203 127 1219 161
rect 1253 127 1269 161
rect 1203 93 1269 127
rect 1203 59 1219 93
rect 1253 59 1269 93
rect 838 17 912 55
rect 1203 17 1269 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
<< metal1 >>
rect 0 561 1288 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1288 561
rect 0 496 1288 527
rect 0 17 1288 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1288 17
rect 0 -48 1288 -17
<< labels >>
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 674 221 708 255 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 766 289 800 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 29 153 63 187 0 FreeSans 340 0 0 0 X
port 9 nsew signal output
flabel locali s 1134 289 1168 323 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 1042 221 1076 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
rlabel comment s 0 0 0 0 4 a211o_4
rlabel metal1 s 0 -48 1288 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1288 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1288 544
string GDS_END 3621678
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3612618
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 32.200 13.600 
<< end >>
