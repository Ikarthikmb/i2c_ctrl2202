magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< poly >>
rect 17980 33806 18080 33823
rect 17980 33772 18013 33806
rect 18047 33772 18080 33806
rect 17980 33738 18080 33772
rect 17980 33704 18013 33738
rect 18047 33704 18080 33738
rect 17980 33670 18080 33704
rect 17980 33636 18013 33670
rect 18047 33636 18080 33670
rect 4262 33100 4396 33116
rect 4262 33066 4278 33100
rect 4312 33066 4346 33100
rect 4380 33066 4396 33100
rect 4262 33050 4396 33066
rect 5554 33100 5688 33116
rect 5554 33066 5570 33100
rect 5604 33066 5638 33100
rect 5672 33066 5688 33100
rect 5554 33050 5688 33066
rect 7550 33100 7684 33116
rect 7550 33066 7566 33100
rect 7600 33066 7634 33100
rect 7668 33066 7684 33100
rect 7550 33050 7684 33066
rect 8844 33100 8978 33116
rect 8844 33066 8860 33100
rect 8894 33066 8928 33100
rect 8962 33066 8978 33100
rect 8844 33050 8978 33066
rect 9356 33100 9490 33116
rect 9356 33066 9372 33100
rect 9406 33066 9440 33100
rect 9474 33066 9490 33100
rect 9356 33050 9490 33066
rect 10646 33100 10780 33116
rect 10646 33066 10662 33100
rect 10696 33066 10730 33100
rect 10764 33066 10780 33100
rect 10646 33050 10780 33066
rect 11161 33100 11295 33116
rect 11161 33066 11177 33100
rect 11211 33066 11245 33100
rect 11279 33066 11295 33100
rect 11161 33050 11295 33066
rect 12455 33100 12589 33116
rect 12455 33066 12471 33100
rect 12505 33066 12539 33100
rect 12573 33066 12589 33100
rect 12455 33050 12589 33066
rect 12962 33100 13096 33116
rect 12962 33066 12978 33100
rect 13012 33066 13046 33100
rect 13080 33066 13096 33100
rect 12962 33050 13096 33066
rect 14256 33100 14390 33116
rect 14256 33066 14272 33100
rect 14306 33066 14340 33100
rect 14374 33066 14390 33100
rect 14256 33050 14390 33066
rect 14770 33100 14904 33116
rect 14770 33066 14786 33100
rect 14820 33066 14854 33100
rect 14888 33066 14904 33100
rect 14770 33050 14904 33066
rect 16060 33100 16194 33116
rect 16060 33066 16076 33100
rect 16110 33066 16144 33100
rect 16178 33066 16194 33100
rect 16060 33050 16194 33066
rect 17980 31562 18013 31596
rect 18047 31562 18080 31596
rect 17980 31528 18080 31562
rect 17980 31494 18013 31528
rect 18047 31494 18080 31528
rect 17980 31460 18080 31494
rect 17980 31426 18013 31460
rect 18047 31426 18080 31460
rect 17980 31409 18080 31426
<< polycont >>
rect 18013 33772 18047 33806
rect 18013 33704 18047 33738
rect 18013 33636 18047 33670
rect 4278 33066 4312 33100
rect 4346 33066 4380 33100
rect 5570 33066 5604 33100
rect 5638 33066 5672 33100
rect 7566 33066 7600 33100
rect 7634 33066 7668 33100
rect 8860 33066 8894 33100
rect 8928 33066 8962 33100
rect 9372 33066 9406 33100
rect 9440 33066 9474 33100
rect 10662 33066 10696 33100
rect 10730 33066 10764 33100
rect 11177 33066 11211 33100
rect 11245 33066 11279 33100
rect 12471 33066 12505 33100
rect 12539 33066 12573 33100
rect 12978 33066 13012 33100
rect 13046 33066 13080 33100
rect 14272 33066 14306 33100
rect 14340 33066 14374 33100
rect 14786 33066 14820 33100
rect 14854 33066 14888 33100
rect 16076 33066 16110 33100
rect 16144 33066 16178 33100
rect 18013 31562 18047 31596
rect 18013 31494 18047 31528
rect 18013 31426 18047 31460
<< npolyres >>
rect 17980 31596 18080 33636
<< locali >>
rect 17997 33810 18063 33822
rect 17997 33776 18005 33810
rect 18039 33806 18063 33810
rect 17997 33772 18013 33776
rect 18047 33772 18063 33806
rect 17997 33738 18063 33772
rect 17997 33704 18005 33738
rect 18047 33704 18063 33738
rect 17997 33670 18063 33704
rect 17997 33666 18013 33670
rect 17997 33632 18005 33666
rect 18047 33636 18063 33670
rect 18039 33632 18063 33636
rect 17997 33620 18063 33632
rect 4262 33404 4396 33418
rect 4262 33370 4274 33404
rect 4308 33370 4350 33404
rect 4384 33370 4396 33404
rect 4262 33100 4396 33370
rect 4262 33073 4278 33100
rect 4312 33066 4346 33100
rect 4380 33073 4396 33100
rect 5554 33404 5688 33418
rect 5554 33370 5566 33404
rect 5600 33370 5642 33404
rect 5676 33370 5688 33404
rect 5554 33100 5688 33370
rect 5554 33073 5570 33100
rect 4278 33050 4380 33066
rect 5604 33066 5638 33100
rect 5672 33073 5688 33100
rect 7550 33404 7684 33418
rect 7550 33370 7562 33404
rect 7596 33370 7638 33404
rect 7672 33370 7684 33404
rect 7550 33100 7684 33370
rect 7550 33073 7566 33100
rect 5570 33050 5672 33066
rect 7600 33066 7634 33100
rect 7668 33073 7684 33100
rect 8844 33404 8978 33418
rect 8844 33370 8856 33404
rect 8890 33370 8932 33404
rect 8966 33370 8978 33404
rect 8844 33100 8978 33370
rect 8844 33073 8860 33100
rect 7566 33050 7668 33066
rect 8894 33066 8928 33100
rect 8962 33073 8978 33100
rect 9356 33404 9490 33418
rect 9356 33370 9368 33404
rect 9402 33370 9444 33404
rect 9478 33370 9490 33404
rect 9356 33100 9490 33370
rect 9356 33073 9372 33100
rect 8860 33050 8962 33066
rect 9406 33066 9440 33100
rect 9474 33073 9490 33100
rect 10646 33404 10780 33418
rect 10646 33370 10658 33404
rect 10692 33370 10734 33404
rect 10768 33370 10780 33404
rect 10646 33100 10780 33370
rect 10646 33073 10662 33100
rect 9372 33050 9474 33066
rect 10696 33066 10730 33100
rect 10764 33073 10780 33100
rect 11161 33404 11295 33418
rect 11161 33370 11173 33404
rect 11207 33370 11249 33404
rect 11283 33370 11295 33404
rect 11161 33100 11295 33370
rect 11161 33073 11177 33100
rect 10662 33050 10764 33066
rect 11211 33066 11245 33100
rect 11279 33073 11295 33100
rect 12455 33404 12589 33418
rect 12455 33370 12467 33404
rect 12501 33370 12543 33404
rect 12577 33370 12589 33404
rect 12455 33100 12589 33370
rect 12455 33073 12471 33100
rect 11177 33050 11279 33066
rect 12505 33066 12539 33100
rect 12573 33073 12589 33100
rect 12962 33404 13096 33418
rect 12962 33370 12974 33404
rect 13008 33370 13050 33404
rect 13084 33370 13096 33404
rect 12962 33100 13096 33370
rect 12962 33073 12978 33100
rect 12471 33050 12573 33066
rect 13012 33066 13046 33100
rect 13080 33073 13096 33100
rect 14256 33404 14390 33418
rect 14256 33370 14268 33404
rect 14302 33370 14344 33404
rect 14378 33370 14390 33404
rect 14256 33100 14390 33370
rect 14256 33073 14272 33100
rect 12978 33050 13080 33066
rect 14306 33066 14340 33100
rect 14374 33073 14390 33100
rect 14770 33404 14904 33418
rect 14770 33370 14782 33404
rect 14816 33370 14858 33404
rect 14892 33370 14904 33404
rect 14770 33100 14904 33370
rect 14770 33073 14786 33100
rect 14272 33050 14374 33066
rect 14820 33066 14854 33100
rect 14888 33073 14904 33100
rect 16060 33404 16194 33418
rect 16060 33370 16072 33404
rect 16106 33370 16148 33404
rect 16182 33370 16194 33404
rect 16060 33100 16194 33370
rect 14786 33050 14888 33066
rect 16060 33066 16076 33100
rect 16110 33066 16144 33100
rect 16178 33066 16194 33100
rect 16060 33050 16194 33066
rect 18009 31612 18055 31613
rect 17997 31601 18063 31612
rect 17997 31596 18015 31601
rect 17997 31562 18013 31596
rect 18049 31567 18063 31601
rect 18047 31562 18063 31567
rect 17997 31529 18063 31562
rect 17997 31528 18015 31529
rect 17997 31494 18013 31528
rect 18049 31495 18063 31529
rect 18047 31494 18063 31495
rect 17997 31460 18063 31494
rect 17997 31426 18013 31460
rect 18047 31457 18063 31460
rect 17997 31423 18015 31426
rect 18049 31423 18063 31457
rect 17997 31410 18063 31423
<< viali >>
rect 18005 33806 18039 33810
rect 18005 33776 18013 33806
rect 18013 33776 18039 33806
rect 18005 33704 18013 33738
rect 18013 33704 18039 33738
rect 18005 33636 18013 33666
rect 18013 33636 18039 33666
rect 18005 33632 18039 33636
rect 4274 33370 4308 33404
rect 4350 33370 4384 33404
rect 5566 33370 5600 33404
rect 5642 33370 5676 33404
rect 7562 33370 7596 33404
rect 7638 33370 7672 33404
rect 8856 33370 8890 33404
rect 8932 33370 8966 33404
rect 9368 33370 9402 33404
rect 9444 33370 9478 33404
rect 10658 33370 10692 33404
rect 10734 33370 10768 33404
rect 11173 33370 11207 33404
rect 11249 33370 11283 33404
rect 12467 33370 12501 33404
rect 12543 33370 12577 33404
rect 12974 33370 13008 33404
rect 13050 33370 13084 33404
rect 14268 33370 14302 33404
rect 14344 33370 14378 33404
rect 14782 33370 14816 33404
rect 14858 33370 14892 33404
rect 16072 33370 16106 33404
rect 16148 33370 16182 33404
rect 18015 31596 18049 31601
rect 18015 31567 18047 31596
rect 18047 31567 18049 31596
rect 18015 31528 18049 31529
rect 18015 31495 18047 31528
rect 18047 31495 18049 31528
rect 18015 31426 18047 31457
rect 18047 31426 18049 31457
rect 18015 31423 18049 31426
<< metal1 >>
rect 17996 33837 18048 33843
rect 17996 33776 18005 33785
rect 18039 33776 18048 33785
rect 17996 33769 18048 33776
rect 17996 33704 18005 33717
rect 18039 33704 18048 33717
rect 17996 33701 18048 33704
rect 17996 33632 18005 33649
rect 18039 33632 18048 33649
rect 17996 33620 18048 33632
rect 3687 33404 5688 33433
rect 3687 33370 4274 33404
rect 4308 33370 4350 33404
rect 4384 33370 5566 33404
rect 5600 33370 5642 33404
rect 5676 33370 5688 33404
rect 3687 33355 5688 33370
rect 7549 33421 9498 33433
rect 7549 33420 8766 33421
rect 7549 33368 7555 33420
rect 7607 33368 7619 33420
rect 7671 33404 8766 33420
rect 7672 33370 8766 33404
rect 7671 33369 8766 33370
rect 8818 33369 8830 33421
rect 8882 33404 9362 33421
rect 8890 33370 8932 33404
rect 8966 33370 9362 33404
rect 8882 33369 9362 33370
rect 9414 33369 9426 33421
rect 9478 33369 9498 33421
rect 10648 33420 16381 33433
rect 10648 33418 16130 33420
rect 7671 33368 9498 33369
rect 7549 33355 9498 33368
rect 10646 33404 16130 33418
rect 10646 33370 10658 33404
rect 10692 33370 10734 33404
rect 10768 33370 11173 33404
rect 11207 33370 11249 33404
rect 11283 33370 12467 33404
rect 12501 33370 12543 33404
rect 12577 33370 12974 33404
rect 13008 33370 13050 33404
rect 13084 33370 14268 33404
rect 14302 33370 14344 33404
rect 14378 33370 14782 33404
rect 14816 33370 14858 33404
rect 14892 33370 16072 33404
rect 16106 33370 16130 33404
rect 10646 33368 16130 33370
rect 16182 33368 16195 33420
rect 16247 33368 16259 33420
rect 16311 33368 16323 33420
rect 16375 33368 16381 33420
rect 10646 33356 16381 33368
rect 10648 33355 16381 33356
rect 17962 31607 18083 31613
rect 17962 31555 17967 31607
rect 18019 31601 18031 31607
rect 18019 31555 18031 31567
rect 17962 31538 18083 31555
rect 17962 31486 17967 31538
rect 18019 31529 18031 31538
rect 18019 31486 18031 31495
rect 17962 31468 18083 31486
rect 17962 31416 17967 31468
rect 18019 31457 18031 31468
rect 18019 31416 18031 31423
rect 17962 31410 18083 31416
rect 5837 24643 5972 24745
rect 3101 23975 3213 24075
<< via1 >>
rect 17996 33810 18048 33837
rect 17996 33785 18005 33810
rect 18005 33785 18039 33810
rect 18039 33785 18048 33810
rect 17996 33738 18048 33769
rect 17996 33717 18005 33738
rect 18005 33717 18039 33738
rect 18039 33717 18048 33738
rect 17996 33666 18048 33701
rect 17996 33649 18005 33666
rect 18005 33649 18039 33666
rect 18039 33649 18048 33666
rect 7555 33404 7607 33420
rect 7555 33370 7562 33404
rect 7562 33370 7596 33404
rect 7596 33370 7607 33404
rect 7555 33368 7607 33370
rect 7619 33404 7671 33420
rect 7619 33370 7638 33404
rect 7638 33370 7671 33404
rect 7619 33368 7671 33370
rect 8766 33369 8818 33421
rect 8830 33404 8882 33421
rect 9362 33404 9414 33421
rect 8830 33370 8856 33404
rect 8856 33370 8882 33404
rect 9362 33370 9368 33404
rect 9368 33370 9402 33404
rect 9402 33370 9414 33404
rect 8830 33369 8882 33370
rect 9362 33369 9414 33370
rect 9426 33404 9478 33421
rect 9426 33370 9444 33404
rect 9444 33370 9478 33404
rect 9426 33369 9478 33370
rect 16130 33404 16182 33420
rect 16130 33370 16148 33404
rect 16148 33370 16182 33404
rect 16130 33368 16182 33370
rect 16195 33368 16247 33420
rect 16259 33368 16311 33420
rect 16323 33368 16375 33420
rect 17967 31601 18019 31607
rect 18031 31601 18083 31607
rect 17967 31567 18015 31601
rect 18015 31567 18019 31601
rect 18031 31567 18049 31601
rect 18049 31567 18083 31601
rect 17967 31555 18019 31567
rect 18031 31555 18083 31567
rect 17967 31529 18019 31538
rect 18031 31529 18083 31538
rect 17967 31495 18015 31529
rect 18015 31495 18019 31529
rect 18031 31495 18049 31529
rect 18049 31495 18083 31529
rect 17967 31486 18019 31495
rect 18031 31486 18083 31495
rect 17967 31457 18019 31468
rect 18031 31457 18083 31468
rect 17967 31423 18015 31457
rect 18015 31423 18019 31457
rect 18031 31423 18049 31457
rect 18049 31423 18083 31457
rect 17967 31416 18019 31423
rect 18031 31416 18083 31423
<< metal2 >>
rect 7549 34022 17952 34074
rect 7549 33420 7677 34022
tri 7677 33997 7702 34022 nw
rect 10636 33957 18007 33989
tri 17966 33948 17975 33957 ne
rect 17975 33948 18007 33957
tri 18007 33948 18048 33989 sw
tri 17975 33927 17996 33948 ne
rect 17996 33837 18048 33948
rect 17996 33769 18048 33785
rect 17996 33701 18048 33717
rect 17996 33643 18048 33649
rect 7549 33368 7555 33420
rect 7607 33368 7619 33420
rect 7671 33368 7677 33420
rect 8760 33369 8766 33421
rect 8818 33369 8830 33421
rect 8882 33369 8888 33421
rect 9356 33369 9362 33421
rect 9414 33369 9426 33421
rect 9478 33369 9484 33421
rect 16124 33420 18191 33433
rect 7549 33355 7677 33368
rect 16124 33368 16130 33420
rect 16182 33368 16195 33420
rect 16247 33368 16259 33420
rect 16311 33368 16323 33420
rect 16375 33368 18191 33420
rect 16124 33355 18191 33368
tri 16686 31613 16774 31701 sw
rect 16686 31607 18083 31613
rect 16686 31555 17967 31607
rect 18019 31555 18031 31607
rect 16686 31538 18083 31555
rect 16686 31486 17967 31538
rect 18019 31486 18031 31538
rect 16686 31468 18083 31486
rect 16686 31416 17967 31468
rect 18019 31416 18031 31468
rect 16686 31410 18083 31416
tri 16686 31325 16771 31410 nw
<< metal3 >>
rect 3777 34055 4373 36549
rect 5579 35290 6175 36515
rect 4683 24636 5275 33634
rect 7066 32939 7658 39298
rect 7968 24620 8560 33634
rect 8870 32930 9462 39298
rect 9772 24620 10364 33634
rect 10674 32939 11266 39298
rect 11576 24620 12168 33634
rect 12478 32930 13070 38307
rect 13380 24620 13972 33634
rect 14282 32930 14874 38307
rect 15184 24620 15776 33634
rect 16086 32930 16686 38307
tri 16086 32925 16091 32930 ne
<< metal4 >>
rect 3801 38307 11797 39298
tri 11797 38307 12788 39298 sw
rect 3801 35624 23573 38307
rect 5263 33972 15541 34482
rect 6494 21432 14283 21952
use sky130_fd_io__gpio_ovtv2_esd_signal_40_sym_hv_2k_dnwl_aup1_b  sky130_fd_io__gpio_ovtv2_esd_signal_40_sym_hv_2k_dnwl_aup1_b_0
timestamp 1644511149
transform 1 0 2709 0 1 23956
box 145 -11849 14642 15342
use sky130_fd_pr__res_generic_po__example_5595914180838  sky130_fd_pr__res_generic_po__example_5595914180838_0
timestamp 1644511149
transform 0 -1 18080 -1 0 33636
box 15 17 2025 18
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1644511149
transform 1 0 16060 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1644511149
transform 1 0 9356 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1644511149
transform 1 0 8844 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_3
timestamp 1644511149
transform 1 0 10646 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_4
timestamp 1644511149
transform 1 0 11161 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_5
timestamp 1644511149
transform 1 0 12455 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_6
timestamp 1644511149
transform 1 0 12962 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_7
timestamp 1644511149
transform 1 0 14256 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_8
timestamp 1644511149
transform 1 0 14770 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_9
timestamp 1644511149
transform 1 0 7550 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_10
timestamp 1644511149
transform -1 0 4396 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_11
timestamp 1644511149
transform -1 0 5688 0 1 33050
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_0
timestamp 1644511149
transform 0 1 18030 1 0 31511
box 0 0 1 1
use sky130_fd_pr__via_pol1_centered__example_559591418081  sky130_fd_pr__via_pol1_centered__example_559591418081_1
timestamp 1644511149
transform 0 1 18030 -1 0 33721
box 0 0 1 1
<< labels >>
flabel comment s 658 31742 658 31742 0 FreeSans 400 180 0 0 P1G
flabel comment s 18018 32511 18018 32511 0 FreeSans 440 270 0 0 LEAKER
flabel metal2 s 17422 34022 17614 34074 3 FreeSans 520 0 0 0 PD_H[2]
port 1 nsew
flabel metal2 s 17422 33355 17614 33433 3 FreeSans 520 0 0 0 PD_H[3]
port 2 nsew
flabel metal1 s 18000 33685 18044 33776 0 FreeSans 400 90 0 0 TIE_LO_ESD
port 3 nsew
flabel metal1 s 18001 31480 18073 31532 0 FreeSans 400 180 0 0 VSSIO
port 4 nsew
flabel metal1 s 3701 33371 3893 33411 3 FreeSans 520 0 0 0 PD_CSD
port 5 nsew
flabel metal1 s 5837 24643 5972 24744 3 FreeSans 200 0 0 0 VSSIO_Q
port 6 nsew
flabel metal1 s 3101 23975 3213 24075 3 FreeSans 200 0 0 0 VDDIO
port 7 nsew
flabel metal3 s 16375 35379 16447 35431 0 FreeSans 400 180 0 0 VSSIO
port 4 nsew
flabel metal3 s 15416 33471 15546 33521 0 FreeSans 200 0 0 0 PAD
port 8 nsew
flabel metal3 s 13629 33471 13759 33521 0 FreeSans 200 0 0 0 PAD
port 8 nsew
flabel metal3 s 11792 33471 11922 33521 0 FreeSans 200 0 0 0 PAD
port 8 nsew
flabel metal3 s 10021 33471 10151 33521 0 FreeSans 200 0 0 0 PAD
port 8 nsew
flabel metal3 s 8190 33471 8320 33521 0 FreeSans 200 0 0 0 PAD
port 8 nsew
flabel metal3 s 4944 33471 5074 33521 0 FreeSans 200 0 0 0 PAD
port 8 nsew
flabel metal3 s 5847 35379 5919 35431 0 FreeSans 400 180 0 0 VSSIO
port 4 nsew
flabel metal3 s 4050 35379 4122 35431 0 FreeSans 400 180 0 0 VSSIO
port 4 nsew
flabel metal3 s 9079 35379 9151 35431 0 FreeSans 400 180 0 0 VSSIO
port 4 nsew
flabel metal3 s 7401 35379 7473 35431 0 FreeSans 400 180 0 0 VSSIO
port 4 nsew
flabel metal3 s 12721 35379 12793 35431 0 FreeSans 400 180 0 0 VSSIO
port 4 nsew
flabel metal3 s 10923 35379 10995 35431 0 FreeSans 400 180 0 0 VSSIO
port 4 nsew
flabel metal3 s 14538 35379 14610 35431 0 FreeSans 400 180 0 0 VSSIO
port 4 nsew
<< properties >>
string GDS_END 43302456
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 43289548
<< end >>
