magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 2614 582
<< pwell >>
rect 1930 201 2575 203
rect 784 157 1238 201
rect 1559 157 2575 201
rect 1 21 2575 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 446 47 476 119
rect 554 47 584 119
rect 650 47 680 131
rect 760 47 790 131
rect 860 47 890 175
rect 944 47 974 175
rect 1132 47 1162 175
rect 1227 47 1257 119
rect 1336 47 1366 119
rect 1431 47 1461 131
rect 1517 47 1547 131
rect 1635 47 1665 175
rect 1719 47 1749 175
rect 1911 47 1941 131
rect 2008 47 2038 177
rect 2092 47 2122 177
rect 2288 47 2318 131
rect 2383 47 2413 177
rect 2467 47 2497 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 413 381 497
rect 446 413 476 497
rect 530 413 560 497
rect 650 413 680 497
rect 756 413 786 497
rect 864 329 894 497
rect 944 329 974 497
rect 1085 329 1115 497
rect 1229 413 1259 497
rect 1313 413 1343 497
rect 1431 413 1461 497
rect 1539 413 1569 497
rect 1635 329 1665 497
rect 1707 329 1737 497
rect 1911 301 1941 429
rect 2008 297 2038 497
rect 2092 297 2122 497
rect 2288 353 2318 481
rect 2383 297 2413 497
rect 2467 297 2497 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 93 351 131
rect 299 59 307 93
rect 341 59 351 93
rect 299 47 351 59
rect 381 119 431 131
rect 810 131 860 175
rect 599 119 650 131
rect 381 111 446 119
rect 381 77 391 111
rect 425 77 446 111
rect 381 47 446 77
rect 476 93 554 119
rect 476 59 499 93
rect 533 59 554 93
rect 476 47 554 59
rect 584 47 650 119
rect 680 89 760 131
rect 680 55 716 89
rect 750 55 760 89
rect 680 47 760 55
rect 790 109 860 131
rect 790 75 800 109
rect 834 75 860 109
rect 790 47 860 75
rect 890 153 944 175
rect 890 119 900 153
rect 934 119 944 153
rect 890 47 944 119
rect 974 127 1026 175
rect 974 93 984 127
rect 1018 93 1026 127
rect 974 47 1026 93
rect 1080 93 1132 175
rect 1080 59 1088 93
rect 1122 59 1132 93
rect 1080 47 1132 59
rect 1162 119 1212 175
rect 1585 131 1635 175
rect 1381 119 1431 131
rect 1162 47 1227 119
rect 1257 93 1336 119
rect 1257 59 1282 93
rect 1316 59 1336 93
rect 1257 47 1336 59
rect 1366 47 1431 119
rect 1461 89 1517 131
rect 1461 55 1473 89
rect 1507 55 1517 89
rect 1461 47 1517 55
rect 1547 109 1635 131
rect 1547 75 1575 109
rect 1609 75 1635 109
rect 1547 47 1635 75
rect 1665 153 1719 175
rect 1665 119 1675 153
rect 1709 119 1719 153
rect 1665 47 1719 119
rect 1749 101 1804 175
rect 1956 161 2008 177
rect 1956 131 1964 161
rect 1749 67 1759 101
rect 1793 67 1804 101
rect 1749 47 1804 67
rect 1858 103 1911 131
rect 1858 69 1866 103
rect 1900 69 1911 103
rect 1858 47 1911 69
rect 1941 127 1964 131
rect 1998 127 2008 161
rect 1941 93 2008 127
rect 1941 59 1964 93
rect 1998 59 2008 93
rect 1941 47 2008 59
rect 2038 127 2092 177
rect 2038 93 2048 127
rect 2082 93 2092 127
rect 2038 47 2092 93
rect 2122 161 2182 177
rect 2122 127 2140 161
rect 2174 127 2182 161
rect 2333 131 2383 177
rect 2122 93 2182 127
rect 2122 59 2140 93
rect 2174 59 2182 93
rect 2122 47 2182 59
rect 2236 119 2288 131
rect 2236 85 2244 119
rect 2278 85 2288 119
rect 2236 47 2288 85
rect 2318 93 2383 131
rect 2318 59 2339 93
rect 2373 59 2383 93
rect 2318 47 2383 59
rect 2413 129 2467 177
rect 2413 95 2423 129
rect 2457 95 2467 129
rect 2413 47 2467 95
rect 2497 161 2549 177
rect 2497 127 2507 161
rect 2541 127 2549 161
rect 2497 93 2549 127
rect 2497 59 2507 93
rect 2541 59 2549 93
rect 2497 47 2549 59
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 299 461 351 497
rect 299 427 307 461
rect 341 427 351 461
rect 299 413 351 427
rect 381 477 446 497
rect 381 443 391 477
rect 425 443 446 477
rect 381 413 446 443
rect 476 484 530 497
rect 476 450 486 484
rect 520 450 530 484
rect 476 413 530 450
rect 560 413 650 497
rect 680 475 756 497
rect 680 441 700 475
rect 734 441 756 475
rect 680 413 756 441
rect 786 459 864 497
rect 786 425 820 459
rect 854 425 864 459
rect 786 413 864 425
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 802 391 864 413
rect 802 357 820 391
rect 854 357 864 391
rect 802 329 864 357
rect 894 329 944 497
rect 974 485 1085 497
rect 974 451 994 485
rect 1028 451 1085 485
rect 974 417 1085 451
rect 974 383 994 417
rect 1028 383 1085 417
rect 974 329 1085 383
rect 1115 413 1229 497
rect 1259 484 1313 497
rect 1259 450 1269 484
rect 1303 450 1313 484
rect 1259 413 1313 450
rect 1343 413 1431 497
rect 1461 485 1539 497
rect 1461 451 1483 485
rect 1517 451 1539 485
rect 1461 413 1539 451
rect 1569 459 1635 497
rect 1569 425 1591 459
rect 1625 425 1635 459
rect 1569 413 1635 425
rect 1115 329 1167 413
rect 1584 329 1635 413
rect 1665 329 1707 497
rect 1737 485 1789 497
rect 1737 451 1747 485
rect 1781 451 1789 485
rect 1956 485 2008 497
rect 1737 329 1789 451
rect 1956 451 1964 485
rect 1998 451 2008 485
rect 1956 429 2008 451
rect 1856 349 1911 429
rect 1856 315 1864 349
rect 1898 315 1911 349
rect 1856 301 1911 315
rect 1941 301 2008 429
rect 1956 297 2008 301
rect 2038 448 2092 497
rect 2038 414 2048 448
rect 2082 414 2092 448
rect 2038 380 2092 414
rect 2038 346 2048 380
rect 2082 346 2092 380
rect 2038 297 2092 346
rect 2122 479 2182 497
rect 2333 481 2383 497
rect 2122 445 2140 479
rect 2174 445 2182 479
rect 2122 411 2182 445
rect 2122 377 2140 411
rect 2174 377 2182 411
rect 2122 343 2182 377
rect 2236 467 2288 481
rect 2236 433 2244 467
rect 2278 433 2288 467
rect 2236 399 2288 433
rect 2236 365 2244 399
rect 2278 365 2288 399
rect 2236 353 2288 365
rect 2318 473 2383 481
rect 2318 439 2339 473
rect 2373 439 2383 473
rect 2318 405 2383 439
rect 2318 371 2339 405
rect 2373 371 2383 405
rect 2318 353 2383 371
rect 2122 309 2140 343
rect 2174 309 2182 343
rect 2122 297 2182 309
rect 2333 297 2383 353
rect 2413 449 2467 497
rect 2413 415 2423 449
rect 2457 415 2467 449
rect 2413 381 2467 415
rect 2413 347 2423 381
rect 2457 347 2467 381
rect 2413 297 2467 347
rect 2497 479 2549 497
rect 2497 445 2507 479
rect 2541 445 2549 479
rect 2497 411 2549 445
rect 2497 377 2507 411
rect 2541 377 2549 411
rect 2497 343 2549 377
rect 2497 309 2507 343
rect 2541 309 2549 343
rect 2497 297 2549 309
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 59 341 93
rect 391 77 425 111
rect 499 59 533 93
rect 716 55 750 89
rect 800 75 834 109
rect 900 119 934 153
rect 984 93 1018 127
rect 1088 59 1122 93
rect 1282 59 1316 93
rect 1473 55 1507 89
rect 1575 75 1609 109
rect 1675 119 1709 153
rect 1759 67 1793 101
rect 1866 69 1900 103
rect 1964 127 1998 161
rect 1964 59 1998 93
rect 2048 93 2082 127
rect 2140 127 2174 161
rect 2140 59 2174 93
rect 2244 85 2278 119
rect 2339 59 2373 93
rect 2423 95 2457 129
rect 2507 127 2541 161
rect 2507 59 2541 93
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 307 427 341 461
rect 391 443 425 477
rect 486 450 520 484
rect 700 441 734 475
rect 820 425 854 459
rect 203 375 237 409
rect 820 357 854 391
rect 994 451 1028 485
rect 994 383 1028 417
rect 1269 450 1303 484
rect 1483 451 1517 485
rect 1591 425 1625 459
rect 1747 451 1781 485
rect 1964 451 1998 485
rect 1864 315 1898 349
rect 2048 414 2082 448
rect 2048 346 2082 380
rect 2140 445 2174 479
rect 2140 377 2174 411
rect 2244 433 2278 467
rect 2244 365 2278 399
rect 2339 439 2373 473
rect 2339 371 2373 405
rect 2140 309 2174 343
rect 2423 415 2457 449
rect 2423 347 2457 381
rect 2507 445 2541 479
rect 2507 377 2541 411
rect 2507 309 2541 343
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 446 497 476 523
rect 530 497 560 523
rect 650 497 680 523
rect 756 497 786 523
rect 864 497 894 523
rect 944 497 974 523
rect 1085 497 1115 523
rect 1229 497 1259 523
rect 1313 497 1343 523
rect 1431 497 1461 523
rect 1539 497 1569 523
rect 1635 497 1665 523
rect 1707 497 1737 523
rect 2008 497 2038 523
rect 2092 497 2122 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 351 267 381 413
rect 446 279 476 413
rect 530 375 560 413
rect 650 381 680 413
rect 518 365 584 375
rect 518 331 534 365
rect 568 331 584 365
rect 518 321 584 331
rect 650 365 714 381
rect 650 331 670 365
rect 704 331 714 365
rect 650 315 714 331
rect 118 230 134 264
rect 168 230 193 264
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 342 251 396 267
rect 342 217 352 251
rect 386 217 396 251
rect 446 249 584 279
rect 342 201 396 217
rect 554 219 584 249
rect 351 131 381 201
rect 446 191 512 207
rect 446 157 468 191
rect 502 157 512 191
rect 446 141 512 157
rect 554 203 608 219
rect 554 169 564 203
rect 598 169 608 203
rect 554 153 608 169
rect 446 119 476 141
rect 554 119 584 153
rect 650 131 680 315
rect 756 229 786 413
rect 1229 381 1259 413
rect 1205 365 1259 381
rect 1313 375 1343 413
rect 1431 381 1461 413
rect 1205 331 1215 365
rect 1249 331 1259 365
rect 864 297 894 329
rect 828 281 894 297
rect 828 247 838 281
rect 872 247 894 281
rect 828 231 894 247
rect 944 297 974 329
rect 944 281 1034 297
rect 944 247 990 281
rect 1024 247 1034 281
rect 944 231 1034 247
rect 1085 263 1115 329
rect 1205 315 1259 331
rect 1301 365 1367 375
rect 1301 331 1317 365
rect 1351 331 1367 365
rect 1301 321 1367 331
rect 1431 365 1497 381
rect 1431 331 1453 365
rect 1487 331 1497 365
rect 1229 279 1259 315
rect 1431 315 1497 331
rect 1085 247 1162 263
rect 1229 249 1366 279
rect 1085 233 1118 247
rect 726 213 786 229
rect 726 179 736 213
rect 770 193 786 213
rect 770 179 790 193
rect 726 163 790 179
rect 860 175 890 231
rect 944 175 974 231
rect 1108 213 1118 233
rect 1152 213 1162 247
rect 1108 197 1162 213
rect 1132 175 1162 197
rect 1227 191 1294 207
rect 760 131 790 163
rect 1227 157 1250 191
rect 1284 157 1294 191
rect 1227 141 1294 157
rect 1227 119 1257 141
rect 1336 119 1366 249
rect 1431 131 1461 315
rect 1539 229 1569 413
rect 1911 429 1941 455
rect 1635 281 1665 329
rect 1503 213 1569 229
rect 1611 265 1665 281
rect 1707 297 1737 329
rect 1707 281 1803 297
rect 1707 267 1759 281
rect 1611 231 1621 265
rect 1655 231 1665 265
rect 1611 215 1665 231
rect 1503 179 1513 213
rect 1547 179 1569 213
rect 1503 163 1569 179
rect 1635 175 1665 215
rect 1719 247 1759 267
rect 1793 247 1803 281
rect 1911 269 1941 301
rect 2288 481 2318 507
rect 2383 497 2413 523
rect 2467 497 2497 523
rect 2288 337 2318 353
rect 2262 307 2318 337
rect 1719 231 1803 247
rect 1856 253 1941 269
rect 2008 265 2038 297
rect 1719 175 1749 231
rect 1856 219 1866 253
rect 1900 219 1941 253
rect 1856 203 1941 219
rect 1517 131 1547 163
rect 1911 131 1941 203
rect 1984 259 2038 265
rect 2092 259 2122 297
rect 2262 259 2292 307
rect 2383 265 2413 297
rect 2467 265 2497 297
rect 1984 249 2292 259
rect 1984 215 1994 249
rect 2028 215 2292 249
rect 1984 205 2292 215
rect 1984 199 2038 205
rect 2008 177 2038 199
rect 2092 177 2122 205
rect 2262 176 2292 205
rect 2354 249 2497 265
rect 2354 215 2364 249
rect 2398 215 2497 249
rect 2354 199 2497 215
rect 2383 177 2413 199
rect 2467 177 2497 199
rect 2262 146 2318 176
rect 2288 131 2318 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 446 21 476 47
rect 554 21 584 47
rect 650 21 680 47
rect 760 21 790 47
rect 860 21 890 47
rect 944 21 974 47
rect 1132 21 1162 47
rect 1227 21 1257 47
rect 1336 21 1366 47
rect 1431 21 1461 47
rect 1517 21 1547 47
rect 1635 21 1665 47
rect 1719 21 1749 47
rect 1911 21 1941 47
rect 2008 21 2038 47
rect 2092 21 2122 47
rect 2288 21 2318 47
rect 2383 21 2413 47
rect 2467 21 2497 47
<< polycont >>
rect 32 230 66 264
rect 534 331 568 365
rect 670 331 704 365
rect 134 230 168 264
rect 352 217 386 251
rect 468 157 502 191
rect 564 169 598 203
rect 1215 331 1249 365
rect 838 247 872 281
rect 990 247 1024 281
rect 1317 331 1351 365
rect 1453 331 1487 365
rect 736 179 770 213
rect 1118 213 1152 247
rect 1250 157 1284 191
rect 1621 231 1655 265
rect 1513 179 1547 213
rect 1759 247 1793 281
rect 1866 219 1900 253
rect 1994 215 2028 249
rect 2364 215 2398 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 237 443 248 477
rect 17 375 35 409
rect 203 409 248 443
rect 289 461 357 527
rect 289 427 307 461
rect 341 427 357 461
rect 391 477 425 493
rect 470 450 486 484
rect 520 450 636 484
rect 69 375 168 393
rect 17 359 168 375
rect 17 264 88 325
rect 17 230 32 264
rect 66 230 88 264
rect 17 195 88 230
rect 122 264 168 359
rect 122 230 134 264
rect 122 187 168 230
rect 17 153 122 161
rect 156 153 168 187
rect 17 127 168 153
rect 237 391 248 409
rect 391 393 425 443
rect 203 357 214 375
rect 17 119 69 127
rect 17 85 35 119
rect 203 119 248 357
rect 284 359 425 393
rect 284 165 318 359
rect 468 357 492 391
rect 526 365 568 391
rect 526 357 534 365
rect 468 331 534 357
rect 352 251 434 325
rect 386 217 434 251
rect 352 201 434 217
rect 468 315 568 331
rect 468 191 512 315
rect 602 281 636 450
rect 684 475 760 527
rect 978 485 1044 527
rect 684 441 700 475
rect 734 441 760 475
rect 820 459 854 475
rect 820 407 854 425
rect 978 451 994 485
rect 1028 451 1044 485
rect 1467 485 1543 527
rect 978 417 1044 451
rect 1253 450 1269 484
rect 1303 450 1419 484
rect 1467 451 1483 485
rect 1517 451 1543 485
rect 1731 485 2014 527
rect 1591 459 1625 475
rect 670 391 940 407
rect 670 365 820 391
rect 704 357 820 365
rect 854 357 940 391
rect 978 383 994 417
rect 1028 383 1044 417
rect 1215 391 1262 397
rect 704 331 720 357
rect 670 315 720 331
rect 822 281 872 297
rect 602 247 838 281
rect 602 239 682 247
rect 284 127 425 165
rect 502 157 512 191
rect 468 141 512 157
rect 548 169 564 203
rect 598 187 614 203
rect 548 153 580 169
rect 548 129 614 153
rect 17 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 248 119
rect 391 111 425 127
rect 203 69 248 85
rect 103 17 169 59
rect 289 59 307 93
rect 341 59 357 93
rect 648 93 682 239
rect 828 231 872 247
rect 906 213 940 357
rect 1215 365 1228 391
rect 1249 331 1262 357
rect 974 323 1175 331
rect 974 289 1136 323
rect 1170 289 1175 323
rect 1215 315 1262 331
rect 1310 365 1351 381
rect 1310 331 1317 365
rect 974 283 1175 289
rect 974 281 1040 283
rect 974 247 990 281
rect 1024 247 1040 281
rect 1310 261 1351 331
rect 1227 255 1351 261
rect 1102 213 1118 247
rect 1152 213 1168 247
rect 720 179 736 213
rect 770 193 786 213
rect 770 187 802 193
rect 720 153 768 179
rect 906 179 1168 213
rect 1227 221 1228 255
rect 1262 225 1351 255
rect 1385 281 1419 450
rect 1731 451 1747 485
rect 1781 451 1964 485
rect 1998 451 2014 485
rect 1591 417 1625 425
rect 2048 448 2100 493
rect 1453 383 2014 417
rect 1453 365 1503 383
rect 1487 331 1503 365
rect 1453 315 1503 331
rect 1385 265 1655 281
rect 1385 247 1621 265
rect 1262 221 1284 225
rect 1227 191 1284 221
rect 906 153 950 179
rect 720 147 802 153
rect 884 119 900 153
rect 934 119 950 153
rect 1227 157 1250 191
rect 984 127 1034 143
rect 1227 141 1284 157
rect 391 61 425 77
rect 289 17 357 59
rect 483 59 499 93
rect 533 59 682 93
rect 483 53 682 59
rect 716 89 750 105
rect 716 17 750 55
rect 784 75 800 109
rect 834 85 850 109
rect 1018 93 1034 127
rect 1385 93 1419 247
rect 1611 231 1621 247
rect 1611 215 1655 231
rect 1494 187 1513 213
rect 1494 153 1504 187
rect 1547 179 1569 213
rect 1538 153 1569 179
rect 1689 156 1725 383
rect 1494 147 1569 153
rect 1659 153 1725 156
rect 1659 119 1675 153
rect 1709 119 1725 153
rect 1759 323 1864 349
rect 1759 289 1780 323
rect 1814 315 1864 323
rect 1898 315 1914 349
rect 1759 281 1814 289
rect 1793 247 1814 281
rect 1980 265 2014 383
rect 2082 414 2100 448
rect 2048 380 2100 414
rect 2082 346 2100 380
rect 2048 326 2100 346
rect 1759 185 1814 247
rect 1850 253 1946 265
rect 1850 219 1866 253
rect 1900 219 1946 253
rect 1980 249 2028 265
rect 1980 215 1994 249
rect 1980 199 2028 215
rect 1759 151 1900 185
rect 984 85 1034 93
rect 834 75 1034 85
rect 784 51 1034 75
rect 1072 59 1088 93
rect 1122 59 1138 93
rect 1072 17 1138 59
rect 1266 59 1282 93
rect 1316 59 1419 93
rect 1266 53 1419 59
rect 1455 89 1507 105
rect 1455 55 1473 89
rect 1455 17 1507 55
rect 1559 75 1575 109
rect 1609 85 1625 109
rect 1759 101 1793 117
rect 1609 75 1759 85
rect 1559 67 1759 75
rect 1559 51 1793 67
rect 1856 103 1900 151
rect 1856 69 1866 103
rect 1856 53 1900 69
rect 1948 127 1964 161
rect 1998 127 2014 161
rect 2064 143 2100 326
rect 2136 479 2182 527
rect 2136 445 2140 479
rect 2174 445 2182 479
rect 2136 411 2182 445
rect 2136 377 2140 411
rect 2174 377 2182 411
rect 2136 343 2182 377
rect 2136 309 2140 343
rect 2174 309 2182 343
rect 2136 293 2182 309
rect 2243 467 2294 483
rect 2243 433 2244 467
rect 2278 433 2294 467
rect 2243 399 2294 433
rect 2243 365 2244 399
rect 2278 365 2294 399
rect 2243 265 2294 365
rect 2330 473 2389 527
rect 2330 439 2339 473
rect 2373 439 2389 473
rect 2330 405 2389 439
rect 2330 371 2339 405
rect 2373 371 2389 405
rect 2330 353 2389 371
rect 2423 449 2469 493
rect 2457 415 2469 449
rect 2423 381 2469 415
rect 2457 347 2469 381
rect 2423 289 2469 347
rect 2503 479 2559 527
rect 2503 445 2507 479
rect 2541 445 2559 479
rect 2503 411 2559 445
rect 2503 377 2507 411
rect 2541 377 2559 411
rect 2503 343 2559 377
rect 2503 309 2507 343
rect 2541 309 2559 343
rect 2503 293 2559 309
rect 2243 249 2398 265
rect 2243 215 2364 249
rect 2243 199 2398 215
rect 1948 93 2014 127
rect 1948 59 1964 93
rect 1998 59 2014 93
rect 1948 17 2014 59
rect 2048 127 2100 143
rect 2082 93 2100 127
rect 2048 51 2100 93
rect 2136 161 2182 177
rect 2136 127 2140 161
rect 2174 127 2182 161
rect 2136 93 2182 127
rect 2136 59 2140 93
rect 2174 59 2182 93
rect 2136 17 2182 59
rect 2243 119 2294 199
rect 2432 165 2469 289
rect 2243 85 2244 119
rect 2278 85 2294 119
rect 2423 129 2469 165
rect 2243 51 2294 85
rect 2330 93 2389 109
rect 2330 59 2339 93
rect 2373 59 2389 93
rect 2330 17 2389 59
rect 2457 95 2469 129
rect 2423 51 2469 95
rect 2503 161 2559 177
rect 2503 127 2507 161
rect 2541 127 2559 161
rect 2503 93 2559 127
rect 2503 59 2507 93
rect 2541 59 2559 93
rect 2503 17 2559 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 2421 527 2455 561
rect 2513 527 2547 561
rect 122 153 156 187
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 492 357 526 391
rect 580 169 598 187
rect 598 169 614 187
rect 580 153 614 169
rect 1228 365 1262 391
rect 1228 357 1249 365
rect 1249 357 1262 365
rect 1136 289 1170 323
rect 768 179 770 187
rect 770 179 802 187
rect 768 153 802 179
rect 1228 221 1262 255
rect 1504 179 1513 187
rect 1513 179 1538 187
rect 1504 153 1538 179
rect 1780 289 1814 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
rect 2421 -17 2455 17
rect 2513 -17 2547 17
<< metal1 >>
rect 0 561 2576 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2421 561
rect 2455 527 2513 561
rect 2547 527 2576 561
rect 0 496 2576 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 480 391 538 397
rect 480 388 492 391
rect 248 360 492 388
rect 248 357 260 360
rect 202 351 260 357
rect 480 357 492 360
rect 526 388 538 391
rect 1216 391 1274 397
rect 1216 388 1228 391
rect 526 360 1228 388
rect 526 357 538 360
rect 480 351 538 357
rect 1216 357 1228 360
rect 1262 357 1274 391
rect 1216 351 1274 357
rect 1124 323 1182 329
rect 1124 289 1136 323
rect 1170 320 1182 323
rect 1768 323 1826 329
rect 1768 320 1780 323
rect 1170 292 1780 320
rect 1170 289 1182 292
rect 1124 283 1182 289
rect 1768 289 1780 292
rect 1814 289 1826 323
rect 1768 283 1826 289
rect 1216 255 1274 261
rect 1216 252 1228 255
rect 587 224 1228 252
rect 587 193 626 224
rect 1216 221 1228 224
rect 1262 221 1274 255
rect 1216 215 1274 221
rect 110 187 168 193
rect 110 153 122 187
rect 156 184 168 187
rect 568 187 626 193
rect 568 184 580 187
rect 156 156 580 184
rect 156 153 168 156
rect 110 147 168 153
rect 568 153 580 156
rect 614 153 626 187
rect 568 147 626 153
rect 756 187 814 193
rect 756 153 768 187
rect 802 184 814 187
rect 1492 187 1550 193
rect 1492 184 1504 187
rect 802 156 1504 184
rect 802 153 814 156
rect 756 147 814 153
rect 1492 153 1504 156
rect 1538 153 1550 187
rect 1492 147 1550 153
rect 0 17 2576 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2421 17
rect 2455 -17 2513 17
rect 2547 -17 2576 17
rect 0 -48 2576 -17
<< labels >>
flabel locali s 1872 221 1906 255 0 FreeSans 400 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 30 -17 64 17 3 FreeSans 400 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 CLK_N
port 1 nsew clock input
flabel locali s 768 153 802 187 0 FreeSans 400 0 0 0 SET_B
port 4 nsew signal input
flabel locali s 2428 85 2462 119 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel locali s 2428 357 2462 391 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel locali s 2428 425 2462 459 0 FreeSans 400 0 0 0 Q
port 9 nsew signal output
flabel locali s 30 527 64 561 3 FreeSans 400 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 400 221 434 255 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 400 289 434 323 0 FreeSans 200 0 0 0 D
port 2 nsew signal input
flabel locali s 2056 425 2090 459 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2056 357 2090 391 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 2056 85 2090 119 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 3 FreeSans 400 0 0 0 VPB
port 7 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
port 7 nsew
flabel pwell s 30 -17 64 17 3 FreeSans 400 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
port 6 nsew
rlabel comment s 0 0 0 0 4 dfbbn_2
rlabel locali s 1494 147 1569 213 1 SET_B
port 4 nsew signal input
rlabel metal1 s 1492 184 1550 193 1 SET_B
port 4 nsew signal input
rlabel metal1 s 1492 147 1550 156 1 SET_B
port 4 nsew signal input
rlabel metal1 s 756 184 814 193 1 SET_B
port 4 nsew signal input
rlabel metal1 s 756 156 1550 184 1 SET_B
port 4 nsew signal input
rlabel metal1 s 756 147 814 156 1 SET_B
port 4 nsew signal input
rlabel metal1 s 0 -48 2576 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2576 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2576 544
string GDS_END 3382204
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3362206
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
