magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< pwell >>
rect 0 66 756 1128
<< nmoslvt >>
rect 194 92 244 1102
rect 300 92 350 1102
rect 406 92 456 1102
rect 512 92 562 1102
<< ndiff >>
rect 138 1090 194 1102
rect 138 1056 149 1090
rect 183 1056 194 1090
rect 138 1022 194 1056
rect 138 988 149 1022
rect 183 988 194 1022
rect 138 954 194 988
rect 138 920 149 954
rect 183 920 194 954
rect 138 886 194 920
rect 138 852 149 886
rect 183 852 194 886
rect 138 818 194 852
rect 138 784 149 818
rect 183 784 194 818
rect 138 750 194 784
rect 138 716 149 750
rect 183 716 194 750
rect 138 682 194 716
rect 138 648 149 682
rect 183 648 194 682
rect 138 614 194 648
rect 138 580 149 614
rect 183 580 194 614
rect 138 546 194 580
rect 138 512 149 546
rect 183 512 194 546
rect 138 478 194 512
rect 138 444 149 478
rect 183 444 194 478
rect 138 410 194 444
rect 138 376 149 410
rect 183 376 194 410
rect 138 342 194 376
rect 138 308 149 342
rect 183 308 194 342
rect 138 274 194 308
rect 138 240 149 274
rect 183 240 194 274
rect 138 206 194 240
rect 138 172 149 206
rect 183 172 194 206
rect 138 138 194 172
rect 138 104 149 138
rect 183 104 194 138
rect 138 92 194 104
rect 244 1090 300 1102
rect 244 1056 255 1090
rect 289 1056 300 1090
rect 244 1022 300 1056
rect 244 988 255 1022
rect 289 988 300 1022
rect 244 954 300 988
rect 244 920 255 954
rect 289 920 300 954
rect 244 886 300 920
rect 244 852 255 886
rect 289 852 300 886
rect 244 818 300 852
rect 244 784 255 818
rect 289 784 300 818
rect 244 750 300 784
rect 244 716 255 750
rect 289 716 300 750
rect 244 682 300 716
rect 244 648 255 682
rect 289 648 300 682
rect 244 614 300 648
rect 244 580 255 614
rect 289 580 300 614
rect 244 546 300 580
rect 244 512 255 546
rect 289 512 300 546
rect 244 478 300 512
rect 244 444 255 478
rect 289 444 300 478
rect 244 410 300 444
rect 244 376 255 410
rect 289 376 300 410
rect 244 342 300 376
rect 244 308 255 342
rect 289 308 300 342
rect 244 274 300 308
rect 244 240 255 274
rect 289 240 300 274
rect 244 206 300 240
rect 244 172 255 206
rect 289 172 300 206
rect 244 138 300 172
rect 244 104 255 138
rect 289 104 300 138
rect 244 92 300 104
rect 350 1090 406 1102
rect 350 1056 361 1090
rect 395 1056 406 1090
rect 350 1022 406 1056
rect 350 988 361 1022
rect 395 988 406 1022
rect 350 954 406 988
rect 350 920 361 954
rect 395 920 406 954
rect 350 886 406 920
rect 350 852 361 886
rect 395 852 406 886
rect 350 818 406 852
rect 350 784 361 818
rect 395 784 406 818
rect 350 750 406 784
rect 350 716 361 750
rect 395 716 406 750
rect 350 682 406 716
rect 350 648 361 682
rect 395 648 406 682
rect 350 614 406 648
rect 350 580 361 614
rect 395 580 406 614
rect 350 546 406 580
rect 350 512 361 546
rect 395 512 406 546
rect 350 478 406 512
rect 350 444 361 478
rect 395 444 406 478
rect 350 410 406 444
rect 350 376 361 410
rect 395 376 406 410
rect 350 342 406 376
rect 350 308 361 342
rect 395 308 406 342
rect 350 274 406 308
rect 350 240 361 274
rect 395 240 406 274
rect 350 206 406 240
rect 350 172 361 206
rect 395 172 406 206
rect 350 138 406 172
rect 350 104 361 138
rect 395 104 406 138
rect 350 92 406 104
rect 456 1090 512 1102
rect 456 1056 467 1090
rect 501 1056 512 1090
rect 456 1022 512 1056
rect 456 988 467 1022
rect 501 988 512 1022
rect 456 954 512 988
rect 456 920 467 954
rect 501 920 512 954
rect 456 886 512 920
rect 456 852 467 886
rect 501 852 512 886
rect 456 818 512 852
rect 456 784 467 818
rect 501 784 512 818
rect 456 750 512 784
rect 456 716 467 750
rect 501 716 512 750
rect 456 682 512 716
rect 456 648 467 682
rect 501 648 512 682
rect 456 614 512 648
rect 456 580 467 614
rect 501 580 512 614
rect 456 546 512 580
rect 456 512 467 546
rect 501 512 512 546
rect 456 478 512 512
rect 456 444 467 478
rect 501 444 512 478
rect 456 410 512 444
rect 456 376 467 410
rect 501 376 512 410
rect 456 342 512 376
rect 456 308 467 342
rect 501 308 512 342
rect 456 274 512 308
rect 456 240 467 274
rect 501 240 512 274
rect 456 206 512 240
rect 456 172 467 206
rect 501 172 512 206
rect 456 138 512 172
rect 456 104 467 138
rect 501 104 512 138
rect 456 92 512 104
rect 562 1090 618 1102
rect 562 1056 573 1090
rect 607 1056 618 1090
rect 562 1022 618 1056
rect 562 988 573 1022
rect 607 988 618 1022
rect 562 954 618 988
rect 562 920 573 954
rect 607 920 618 954
rect 562 886 618 920
rect 562 852 573 886
rect 607 852 618 886
rect 562 818 618 852
rect 562 784 573 818
rect 607 784 618 818
rect 562 750 618 784
rect 562 716 573 750
rect 607 716 618 750
rect 562 682 618 716
rect 562 648 573 682
rect 607 648 618 682
rect 562 614 618 648
rect 562 580 573 614
rect 607 580 618 614
rect 562 546 618 580
rect 562 512 573 546
rect 607 512 618 546
rect 562 478 618 512
rect 562 444 573 478
rect 607 444 618 478
rect 562 410 618 444
rect 562 376 573 410
rect 607 376 618 410
rect 562 342 618 376
rect 562 308 573 342
rect 607 308 618 342
rect 562 274 618 308
rect 562 240 573 274
rect 607 240 618 274
rect 562 206 618 240
rect 562 172 573 206
rect 607 172 618 206
rect 562 138 618 172
rect 562 104 573 138
rect 607 104 618 138
rect 562 92 618 104
<< ndiffc >>
rect 149 1056 183 1090
rect 149 988 183 1022
rect 149 920 183 954
rect 149 852 183 886
rect 149 784 183 818
rect 149 716 183 750
rect 149 648 183 682
rect 149 580 183 614
rect 149 512 183 546
rect 149 444 183 478
rect 149 376 183 410
rect 149 308 183 342
rect 149 240 183 274
rect 149 172 183 206
rect 149 104 183 138
rect 255 1056 289 1090
rect 255 988 289 1022
rect 255 920 289 954
rect 255 852 289 886
rect 255 784 289 818
rect 255 716 289 750
rect 255 648 289 682
rect 255 580 289 614
rect 255 512 289 546
rect 255 444 289 478
rect 255 376 289 410
rect 255 308 289 342
rect 255 240 289 274
rect 255 172 289 206
rect 255 104 289 138
rect 361 1056 395 1090
rect 361 988 395 1022
rect 361 920 395 954
rect 361 852 395 886
rect 361 784 395 818
rect 361 716 395 750
rect 361 648 395 682
rect 361 580 395 614
rect 361 512 395 546
rect 361 444 395 478
rect 361 376 395 410
rect 361 308 395 342
rect 361 240 395 274
rect 361 172 395 206
rect 361 104 395 138
rect 467 1056 501 1090
rect 467 988 501 1022
rect 467 920 501 954
rect 467 852 501 886
rect 467 784 501 818
rect 467 716 501 750
rect 467 648 501 682
rect 467 580 501 614
rect 467 512 501 546
rect 467 444 501 478
rect 467 376 501 410
rect 467 308 501 342
rect 467 240 501 274
rect 467 172 501 206
rect 467 104 501 138
rect 573 1056 607 1090
rect 573 988 607 1022
rect 573 920 607 954
rect 573 852 607 886
rect 573 784 607 818
rect 573 716 607 750
rect 573 648 607 682
rect 573 580 607 614
rect 573 512 607 546
rect 573 444 607 478
rect 573 376 607 410
rect 573 308 607 342
rect 573 240 607 274
rect 573 172 607 206
rect 573 104 607 138
<< psubdiff >>
rect 26 1056 84 1102
rect 26 1022 38 1056
rect 72 1022 84 1056
rect 26 988 84 1022
rect 26 954 38 988
rect 72 954 84 988
rect 26 920 84 954
rect 26 886 38 920
rect 72 886 84 920
rect 26 852 84 886
rect 26 818 38 852
rect 72 818 84 852
rect 26 784 84 818
rect 26 750 38 784
rect 72 750 84 784
rect 26 716 84 750
rect 26 682 38 716
rect 72 682 84 716
rect 26 648 84 682
rect 26 614 38 648
rect 72 614 84 648
rect 26 580 84 614
rect 26 546 38 580
rect 72 546 84 580
rect 26 512 84 546
rect 26 478 38 512
rect 72 478 84 512
rect 26 444 84 478
rect 26 410 38 444
rect 72 410 84 444
rect 26 376 84 410
rect 26 342 38 376
rect 72 342 84 376
rect 26 308 84 342
rect 26 274 38 308
rect 72 274 84 308
rect 26 240 84 274
rect 26 206 38 240
rect 72 206 84 240
rect 26 172 84 206
rect 26 138 38 172
rect 72 138 84 172
rect 26 92 84 138
rect 672 1056 730 1102
rect 672 1022 684 1056
rect 718 1022 730 1056
rect 672 988 730 1022
rect 672 954 684 988
rect 718 954 730 988
rect 672 920 730 954
rect 672 886 684 920
rect 718 886 730 920
rect 672 852 730 886
rect 672 818 684 852
rect 718 818 730 852
rect 672 784 730 818
rect 672 750 684 784
rect 718 750 730 784
rect 672 716 730 750
rect 672 682 684 716
rect 718 682 730 716
rect 672 648 730 682
rect 672 614 684 648
rect 718 614 730 648
rect 672 580 730 614
rect 672 546 684 580
rect 718 546 730 580
rect 672 512 730 546
rect 672 478 684 512
rect 718 478 730 512
rect 672 444 730 478
rect 672 410 684 444
rect 718 410 730 444
rect 672 376 730 410
rect 672 342 684 376
rect 718 342 730 376
rect 672 308 730 342
rect 672 274 684 308
rect 718 274 730 308
rect 672 240 730 274
rect 672 206 684 240
rect 718 206 730 240
rect 672 172 730 206
rect 672 138 684 172
rect 718 138 730 172
rect 672 92 730 138
<< psubdiffcont >>
rect 38 1022 72 1056
rect 38 954 72 988
rect 38 886 72 920
rect 38 818 72 852
rect 38 750 72 784
rect 38 682 72 716
rect 38 614 72 648
rect 38 546 72 580
rect 38 478 72 512
rect 38 410 72 444
rect 38 342 72 376
rect 38 274 72 308
rect 38 206 72 240
rect 38 138 72 172
rect 684 1022 718 1056
rect 684 954 718 988
rect 684 886 718 920
rect 684 818 718 852
rect 684 750 718 784
rect 684 682 718 716
rect 684 614 718 648
rect 684 546 718 580
rect 684 478 718 512
rect 684 410 718 444
rect 684 342 718 376
rect 684 274 718 308
rect 684 206 718 240
rect 684 138 718 172
<< poly >>
rect 175 1174 581 1194
rect 175 1140 191 1174
rect 225 1140 259 1174
rect 293 1140 327 1174
rect 361 1140 395 1174
rect 429 1140 463 1174
rect 497 1140 531 1174
rect 565 1140 581 1174
rect 175 1124 581 1140
rect 194 1102 244 1124
rect 300 1102 350 1124
rect 406 1102 456 1124
rect 512 1102 562 1124
rect 194 70 244 92
rect 300 70 350 92
rect 406 70 456 92
rect 512 70 562 92
rect 175 54 581 70
rect 175 20 191 54
rect 225 20 259 54
rect 293 20 327 54
rect 361 20 395 54
rect 429 20 463 54
rect 497 20 531 54
rect 565 20 581 54
rect 175 0 581 20
<< polycont >>
rect 191 1140 225 1174
rect 259 1140 293 1174
rect 327 1140 361 1174
rect 395 1140 429 1174
rect 463 1140 497 1174
rect 531 1140 565 1174
rect 191 20 225 54
rect 259 20 293 54
rect 327 20 361 54
rect 395 20 429 54
rect 463 20 497 54
rect 531 20 565 54
<< locali >>
rect 175 1140 182 1174
rect 225 1140 254 1174
rect 293 1140 326 1174
rect 361 1140 395 1174
rect 432 1140 463 1174
rect 504 1140 531 1174
rect 576 1140 581 1174
rect 149 1090 183 1106
rect 38 1010 72 1022
rect 38 938 72 954
rect 38 866 72 886
rect 38 794 72 818
rect 38 722 72 750
rect 38 650 72 682
rect 38 580 72 614
rect 38 512 72 544
rect 38 444 72 472
rect 38 376 72 400
rect 38 308 72 328
rect 38 240 72 256
rect 38 172 72 184
rect 149 1022 183 1048
rect 149 954 183 976
rect 149 886 183 904
rect 149 818 183 832
rect 149 750 183 760
rect 149 682 183 688
rect 149 614 183 616
rect 149 578 183 580
rect 149 506 183 512
rect 149 434 183 444
rect 149 362 183 376
rect 149 290 183 308
rect 149 218 183 240
rect 149 146 183 172
rect 149 88 183 104
rect 255 1090 289 1106
rect 255 1022 289 1048
rect 255 954 289 976
rect 255 886 289 904
rect 255 818 289 832
rect 255 750 289 760
rect 255 682 289 688
rect 255 614 289 616
rect 255 578 289 580
rect 255 506 289 512
rect 255 434 289 444
rect 255 362 289 376
rect 255 290 289 308
rect 255 218 289 240
rect 255 146 289 172
rect 255 88 289 104
rect 361 1090 395 1106
rect 361 1022 395 1048
rect 361 954 395 976
rect 361 886 395 904
rect 361 818 395 832
rect 361 750 395 760
rect 361 682 395 688
rect 361 614 395 616
rect 361 578 395 580
rect 361 506 395 512
rect 361 434 395 444
rect 361 362 395 376
rect 361 290 395 308
rect 361 218 395 240
rect 361 146 395 172
rect 361 88 395 104
rect 467 1090 501 1106
rect 467 1022 501 1048
rect 467 954 501 976
rect 467 886 501 904
rect 467 818 501 832
rect 467 750 501 760
rect 467 682 501 688
rect 467 614 501 616
rect 467 578 501 580
rect 467 506 501 512
rect 467 434 501 444
rect 467 362 501 376
rect 467 290 501 308
rect 467 218 501 240
rect 467 146 501 172
rect 467 88 501 104
rect 573 1090 607 1106
rect 573 1022 607 1048
rect 573 954 607 976
rect 573 886 607 904
rect 573 818 607 832
rect 573 750 607 760
rect 573 682 607 688
rect 573 614 607 616
rect 573 578 607 580
rect 573 506 607 512
rect 573 434 607 444
rect 573 362 607 376
rect 573 290 607 308
rect 573 218 607 240
rect 573 146 607 172
rect 684 1010 718 1022
rect 684 938 718 954
rect 684 866 718 886
rect 684 794 718 818
rect 684 722 718 750
rect 684 650 718 682
rect 684 580 718 614
rect 684 512 718 544
rect 684 444 718 472
rect 684 376 718 400
rect 684 308 718 328
rect 684 240 718 256
rect 684 172 718 184
rect 573 88 607 104
rect 175 20 182 54
rect 225 20 254 54
rect 293 20 326 54
rect 361 20 395 54
rect 432 20 463 54
rect 504 20 531 54
rect 576 20 581 54
<< viali >>
rect 182 1140 191 1174
rect 191 1140 216 1174
rect 254 1140 259 1174
rect 259 1140 288 1174
rect 326 1140 327 1174
rect 327 1140 360 1174
rect 398 1140 429 1174
rect 429 1140 432 1174
rect 470 1140 497 1174
rect 497 1140 504 1174
rect 542 1140 565 1174
rect 565 1140 576 1174
rect 38 1056 72 1082
rect 38 1048 72 1056
rect 38 988 72 1010
rect 38 976 72 988
rect 38 920 72 938
rect 38 904 72 920
rect 38 852 72 866
rect 38 832 72 852
rect 38 784 72 794
rect 38 760 72 784
rect 38 716 72 722
rect 38 688 72 716
rect 38 648 72 650
rect 38 616 72 648
rect 38 546 72 578
rect 38 544 72 546
rect 38 478 72 506
rect 38 472 72 478
rect 38 410 72 434
rect 38 400 72 410
rect 38 342 72 362
rect 38 328 72 342
rect 38 274 72 290
rect 38 256 72 274
rect 38 206 72 218
rect 38 184 72 206
rect 38 138 72 146
rect 38 112 72 138
rect 149 1056 183 1082
rect 149 1048 183 1056
rect 149 988 183 1010
rect 149 976 183 988
rect 149 920 183 938
rect 149 904 183 920
rect 149 852 183 866
rect 149 832 183 852
rect 149 784 183 794
rect 149 760 183 784
rect 149 716 183 722
rect 149 688 183 716
rect 149 648 183 650
rect 149 616 183 648
rect 149 546 183 578
rect 149 544 183 546
rect 149 478 183 506
rect 149 472 183 478
rect 149 410 183 434
rect 149 400 183 410
rect 149 342 183 362
rect 149 328 183 342
rect 149 274 183 290
rect 149 256 183 274
rect 149 206 183 218
rect 149 184 183 206
rect 149 138 183 146
rect 149 112 183 138
rect 255 1056 289 1082
rect 255 1048 289 1056
rect 255 988 289 1010
rect 255 976 289 988
rect 255 920 289 938
rect 255 904 289 920
rect 255 852 289 866
rect 255 832 289 852
rect 255 784 289 794
rect 255 760 289 784
rect 255 716 289 722
rect 255 688 289 716
rect 255 648 289 650
rect 255 616 289 648
rect 255 546 289 578
rect 255 544 289 546
rect 255 478 289 506
rect 255 472 289 478
rect 255 410 289 434
rect 255 400 289 410
rect 255 342 289 362
rect 255 328 289 342
rect 255 274 289 290
rect 255 256 289 274
rect 255 206 289 218
rect 255 184 289 206
rect 255 138 289 146
rect 255 112 289 138
rect 361 1056 395 1082
rect 361 1048 395 1056
rect 361 988 395 1010
rect 361 976 395 988
rect 361 920 395 938
rect 361 904 395 920
rect 361 852 395 866
rect 361 832 395 852
rect 361 784 395 794
rect 361 760 395 784
rect 361 716 395 722
rect 361 688 395 716
rect 361 648 395 650
rect 361 616 395 648
rect 361 546 395 578
rect 361 544 395 546
rect 361 478 395 506
rect 361 472 395 478
rect 361 410 395 434
rect 361 400 395 410
rect 361 342 395 362
rect 361 328 395 342
rect 361 274 395 290
rect 361 256 395 274
rect 361 206 395 218
rect 361 184 395 206
rect 361 138 395 146
rect 361 112 395 138
rect 467 1056 501 1082
rect 467 1048 501 1056
rect 467 988 501 1010
rect 467 976 501 988
rect 467 920 501 938
rect 467 904 501 920
rect 467 852 501 866
rect 467 832 501 852
rect 467 784 501 794
rect 467 760 501 784
rect 467 716 501 722
rect 467 688 501 716
rect 467 648 501 650
rect 467 616 501 648
rect 467 546 501 578
rect 467 544 501 546
rect 467 478 501 506
rect 467 472 501 478
rect 467 410 501 434
rect 467 400 501 410
rect 467 342 501 362
rect 467 328 501 342
rect 467 274 501 290
rect 467 256 501 274
rect 467 206 501 218
rect 467 184 501 206
rect 467 138 501 146
rect 467 112 501 138
rect 573 1056 607 1082
rect 573 1048 607 1056
rect 573 988 607 1010
rect 573 976 607 988
rect 573 920 607 938
rect 573 904 607 920
rect 573 852 607 866
rect 573 832 607 852
rect 573 784 607 794
rect 573 760 607 784
rect 573 716 607 722
rect 573 688 607 716
rect 573 648 607 650
rect 573 616 607 648
rect 573 546 607 578
rect 573 544 607 546
rect 573 478 607 506
rect 573 472 607 478
rect 573 410 607 434
rect 573 400 607 410
rect 573 342 607 362
rect 573 328 607 342
rect 573 274 607 290
rect 573 256 607 274
rect 573 206 607 218
rect 573 184 607 206
rect 573 138 607 146
rect 573 112 607 138
rect 684 1056 718 1082
rect 684 1048 718 1056
rect 684 988 718 1010
rect 684 976 718 988
rect 684 920 718 938
rect 684 904 718 920
rect 684 852 718 866
rect 684 832 718 852
rect 684 784 718 794
rect 684 760 718 784
rect 684 716 718 722
rect 684 688 718 716
rect 684 648 718 650
rect 684 616 718 648
rect 684 546 718 578
rect 684 544 718 546
rect 684 478 718 506
rect 684 472 718 478
rect 684 410 718 434
rect 684 400 718 410
rect 684 342 718 362
rect 684 328 718 342
rect 684 274 718 290
rect 684 256 718 274
rect 684 206 718 218
rect 684 184 718 206
rect 684 138 718 146
rect 684 112 718 138
rect 182 20 191 54
rect 191 20 216 54
rect 254 20 259 54
rect 259 20 288 54
rect 326 20 327 54
rect 327 20 360 54
rect 398 20 429 54
rect 429 20 432 54
rect 470 20 497 54
rect 497 20 504 54
rect 542 20 565 54
rect 565 20 576 54
<< metal1 >>
rect 170 1174 588 1194
rect 170 1140 182 1174
rect 216 1140 254 1174
rect 288 1140 326 1174
rect 360 1140 398 1174
rect 432 1140 470 1174
rect 504 1140 542 1174
rect 576 1140 588 1174
rect 170 1128 588 1140
rect 26 1082 84 1094
rect 26 1048 38 1082
rect 72 1048 84 1082
rect 26 1010 84 1048
rect 26 976 38 1010
rect 72 976 84 1010
rect 26 938 84 976
rect 26 904 38 938
rect 72 904 84 938
rect 26 866 84 904
rect 26 832 38 866
rect 72 832 84 866
rect 26 794 84 832
rect 26 760 38 794
rect 72 760 84 794
rect 26 722 84 760
rect 26 688 38 722
rect 72 688 84 722
rect 26 650 84 688
rect 26 616 38 650
rect 72 616 84 650
rect 26 578 84 616
rect 26 544 38 578
rect 72 544 84 578
rect 26 506 84 544
rect 26 472 38 506
rect 72 472 84 506
rect 26 434 84 472
rect 26 400 38 434
rect 72 400 84 434
rect 26 362 84 400
rect 26 328 38 362
rect 72 328 84 362
rect 26 290 84 328
rect 26 256 38 290
rect 72 256 84 290
rect 26 218 84 256
rect 26 184 38 218
rect 72 184 84 218
rect 26 146 84 184
rect 26 112 38 146
rect 72 112 84 146
rect 26 100 84 112
rect 140 1082 192 1094
rect 140 1048 149 1082
rect 183 1048 192 1082
rect 140 1010 192 1048
rect 140 976 149 1010
rect 183 976 192 1010
rect 140 938 192 976
rect 140 904 149 938
rect 183 904 192 938
rect 140 866 192 904
rect 140 832 149 866
rect 183 832 192 866
rect 140 794 192 832
rect 140 760 149 794
rect 183 760 192 794
rect 140 722 192 760
rect 140 688 149 722
rect 183 688 192 722
rect 140 650 192 688
rect 140 616 149 650
rect 183 616 192 650
rect 140 578 192 616
rect 140 544 149 578
rect 183 544 192 578
rect 140 542 192 544
rect 140 478 149 490
rect 183 478 192 490
rect 140 414 149 426
rect 183 414 192 426
rect 140 350 149 362
rect 183 350 192 362
rect 140 290 192 298
rect 140 286 149 290
rect 183 286 192 290
rect 140 222 192 234
rect 140 158 192 170
rect 140 100 192 106
rect 246 1088 298 1094
rect 246 1024 298 1036
rect 246 960 298 972
rect 246 904 255 908
rect 289 904 298 908
rect 246 896 298 904
rect 246 832 255 844
rect 289 832 298 844
rect 246 768 255 780
rect 289 768 298 780
rect 246 704 255 716
rect 289 704 298 716
rect 246 650 298 652
rect 246 616 255 650
rect 289 616 298 650
rect 246 578 298 616
rect 246 544 255 578
rect 289 544 298 578
rect 246 506 298 544
rect 246 472 255 506
rect 289 472 298 506
rect 246 434 298 472
rect 246 400 255 434
rect 289 400 298 434
rect 246 362 298 400
rect 246 328 255 362
rect 289 328 298 362
rect 246 290 298 328
rect 246 256 255 290
rect 289 256 298 290
rect 246 218 298 256
rect 246 184 255 218
rect 289 184 298 218
rect 246 146 298 184
rect 246 112 255 146
rect 289 112 298 146
rect 246 100 298 112
rect 352 1082 404 1094
rect 352 1048 361 1082
rect 395 1048 404 1082
rect 352 1010 404 1048
rect 352 976 361 1010
rect 395 976 404 1010
rect 352 938 404 976
rect 352 904 361 938
rect 395 904 404 938
rect 352 866 404 904
rect 352 832 361 866
rect 395 832 404 866
rect 352 794 404 832
rect 352 760 361 794
rect 395 760 404 794
rect 352 722 404 760
rect 352 688 361 722
rect 395 688 404 722
rect 352 650 404 688
rect 352 616 361 650
rect 395 616 404 650
rect 352 578 404 616
rect 352 544 361 578
rect 395 544 404 578
rect 352 542 404 544
rect 352 478 361 490
rect 395 478 404 490
rect 352 414 361 426
rect 395 414 404 426
rect 352 350 361 362
rect 395 350 404 362
rect 352 290 404 298
rect 352 286 361 290
rect 395 286 404 290
rect 352 222 404 234
rect 352 158 404 170
rect 352 100 404 106
rect 458 1088 510 1094
rect 458 1024 510 1036
rect 458 960 510 972
rect 458 904 467 908
rect 501 904 510 908
rect 458 896 510 904
rect 458 832 467 844
rect 501 832 510 844
rect 458 768 467 780
rect 501 768 510 780
rect 458 704 467 716
rect 501 704 510 716
rect 458 650 510 652
rect 458 616 467 650
rect 501 616 510 650
rect 458 578 510 616
rect 458 544 467 578
rect 501 544 510 578
rect 458 506 510 544
rect 458 472 467 506
rect 501 472 510 506
rect 458 434 510 472
rect 458 400 467 434
rect 501 400 510 434
rect 458 362 510 400
rect 458 328 467 362
rect 501 328 510 362
rect 458 290 510 328
rect 458 256 467 290
rect 501 256 510 290
rect 458 218 510 256
rect 458 184 467 218
rect 501 184 510 218
rect 458 146 510 184
rect 458 112 467 146
rect 501 112 510 146
rect 458 100 510 112
rect 564 1082 616 1094
rect 564 1048 573 1082
rect 607 1048 616 1082
rect 564 1010 616 1048
rect 564 976 573 1010
rect 607 976 616 1010
rect 564 938 616 976
rect 564 904 573 938
rect 607 904 616 938
rect 564 866 616 904
rect 564 832 573 866
rect 607 832 616 866
rect 564 794 616 832
rect 564 760 573 794
rect 607 760 616 794
rect 564 722 616 760
rect 564 688 573 722
rect 607 688 616 722
rect 564 650 616 688
rect 564 616 573 650
rect 607 616 616 650
rect 564 578 616 616
rect 564 544 573 578
rect 607 544 616 578
rect 564 542 616 544
rect 564 478 573 490
rect 607 478 616 490
rect 564 414 573 426
rect 607 414 616 426
rect 564 350 573 362
rect 607 350 616 362
rect 564 290 616 298
rect 564 286 573 290
rect 607 286 616 290
rect 564 222 616 234
rect 564 158 616 170
rect 564 100 616 106
rect 672 1082 730 1094
rect 672 1048 684 1082
rect 718 1048 730 1082
rect 672 1010 730 1048
rect 672 976 684 1010
rect 718 976 730 1010
rect 672 938 730 976
rect 672 904 684 938
rect 718 904 730 938
rect 672 866 730 904
rect 672 832 684 866
rect 718 832 730 866
rect 672 794 730 832
rect 672 760 684 794
rect 718 760 730 794
rect 672 722 730 760
rect 672 688 684 722
rect 718 688 730 722
rect 672 650 730 688
rect 672 616 684 650
rect 718 616 730 650
rect 672 578 730 616
rect 672 544 684 578
rect 718 544 730 578
rect 672 506 730 544
rect 672 472 684 506
rect 718 472 730 506
rect 672 434 730 472
rect 672 400 684 434
rect 718 400 730 434
rect 672 362 730 400
rect 672 328 684 362
rect 718 328 730 362
rect 672 290 730 328
rect 672 256 684 290
rect 718 256 730 290
rect 672 218 730 256
rect 672 184 684 218
rect 718 184 730 218
rect 672 146 730 184
rect 672 112 684 146
rect 718 112 730 146
rect 672 100 730 112
rect 170 54 588 66
rect 170 20 182 54
rect 216 20 254 54
rect 288 20 326 54
rect 360 20 398 54
rect 432 20 470 54
rect 504 20 542 54
rect 576 20 588 54
rect 170 0 588 20
<< via1 >>
rect 140 506 192 542
rect 140 490 149 506
rect 149 490 183 506
rect 183 490 192 506
rect 140 472 149 478
rect 149 472 183 478
rect 183 472 192 478
rect 140 434 192 472
rect 140 426 149 434
rect 149 426 183 434
rect 183 426 192 434
rect 140 400 149 414
rect 149 400 183 414
rect 183 400 192 414
rect 140 362 192 400
rect 140 328 149 350
rect 149 328 183 350
rect 183 328 192 350
rect 140 298 192 328
rect 140 256 149 286
rect 149 256 183 286
rect 183 256 192 286
rect 140 234 192 256
rect 140 218 192 222
rect 140 184 149 218
rect 149 184 183 218
rect 183 184 192 218
rect 140 170 192 184
rect 140 146 192 158
rect 140 112 149 146
rect 149 112 183 146
rect 183 112 192 146
rect 140 106 192 112
rect 246 1082 298 1088
rect 246 1048 255 1082
rect 255 1048 289 1082
rect 289 1048 298 1082
rect 246 1036 298 1048
rect 246 1010 298 1024
rect 246 976 255 1010
rect 255 976 289 1010
rect 289 976 298 1010
rect 246 972 298 976
rect 246 938 298 960
rect 246 908 255 938
rect 255 908 289 938
rect 289 908 298 938
rect 246 866 298 896
rect 246 844 255 866
rect 255 844 289 866
rect 289 844 298 866
rect 246 794 298 832
rect 246 780 255 794
rect 255 780 289 794
rect 289 780 298 794
rect 246 760 255 768
rect 255 760 289 768
rect 289 760 298 768
rect 246 722 298 760
rect 246 716 255 722
rect 255 716 289 722
rect 289 716 298 722
rect 246 688 255 704
rect 255 688 289 704
rect 289 688 298 704
rect 246 652 298 688
rect 352 506 404 542
rect 352 490 361 506
rect 361 490 395 506
rect 395 490 404 506
rect 352 472 361 478
rect 361 472 395 478
rect 395 472 404 478
rect 352 434 404 472
rect 352 426 361 434
rect 361 426 395 434
rect 395 426 404 434
rect 352 400 361 414
rect 361 400 395 414
rect 395 400 404 414
rect 352 362 404 400
rect 352 328 361 350
rect 361 328 395 350
rect 395 328 404 350
rect 352 298 404 328
rect 352 256 361 286
rect 361 256 395 286
rect 395 256 404 286
rect 352 234 404 256
rect 352 218 404 222
rect 352 184 361 218
rect 361 184 395 218
rect 395 184 404 218
rect 352 170 404 184
rect 352 146 404 158
rect 352 112 361 146
rect 361 112 395 146
rect 395 112 404 146
rect 352 106 404 112
rect 458 1082 510 1088
rect 458 1048 467 1082
rect 467 1048 501 1082
rect 501 1048 510 1082
rect 458 1036 510 1048
rect 458 1010 510 1024
rect 458 976 467 1010
rect 467 976 501 1010
rect 501 976 510 1010
rect 458 972 510 976
rect 458 938 510 960
rect 458 908 467 938
rect 467 908 501 938
rect 501 908 510 938
rect 458 866 510 896
rect 458 844 467 866
rect 467 844 501 866
rect 501 844 510 866
rect 458 794 510 832
rect 458 780 467 794
rect 467 780 501 794
rect 501 780 510 794
rect 458 760 467 768
rect 467 760 501 768
rect 501 760 510 768
rect 458 722 510 760
rect 458 716 467 722
rect 467 716 501 722
rect 501 716 510 722
rect 458 688 467 704
rect 467 688 501 704
rect 501 688 510 704
rect 458 652 510 688
rect 564 506 616 542
rect 564 490 573 506
rect 573 490 607 506
rect 607 490 616 506
rect 564 472 573 478
rect 573 472 607 478
rect 607 472 616 478
rect 564 434 616 472
rect 564 426 573 434
rect 573 426 607 434
rect 607 426 616 434
rect 564 400 573 414
rect 573 400 607 414
rect 607 400 616 414
rect 564 362 616 400
rect 564 328 573 350
rect 573 328 607 350
rect 607 328 616 350
rect 564 298 616 328
rect 564 256 573 286
rect 573 256 607 286
rect 607 256 616 286
rect 564 234 616 256
rect 564 218 616 222
rect 564 184 573 218
rect 573 184 607 218
rect 607 184 616 218
rect 564 170 616 184
rect 564 146 616 158
rect 564 112 573 146
rect 573 112 607 146
rect 607 112 616 146
rect 564 106 616 112
<< metal2 >>
rect 0 1088 756 1094
rect 0 1036 246 1088
rect 298 1036 458 1088
rect 510 1036 756 1088
rect 0 1024 756 1036
rect 0 972 246 1024
rect 298 972 458 1024
rect 510 972 756 1024
rect 0 960 756 972
rect 0 908 246 960
rect 298 908 458 960
rect 510 908 756 960
rect 0 896 756 908
rect 0 844 246 896
rect 298 844 458 896
rect 510 844 756 896
rect 0 832 756 844
rect 0 780 246 832
rect 298 780 458 832
rect 510 780 756 832
rect 0 768 756 780
rect 0 716 246 768
rect 298 716 458 768
rect 510 716 756 768
rect 0 704 756 716
rect 0 652 246 704
rect 298 652 458 704
rect 510 652 756 704
rect 0 622 756 652
rect 0 542 756 572
rect 0 490 140 542
rect 192 490 352 542
rect 404 490 564 542
rect 616 490 756 542
rect 0 478 756 490
rect 0 426 140 478
rect 192 426 352 478
rect 404 426 564 478
rect 616 426 756 478
rect 0 414 756 426
rect 0 362 140 414
rect 192 362 352 414
rect 404 362 564 414
rect 616 362 756 414
rect 0 350 756 362
rect 0 298 140 350
rect 192 298 352 350
rect 404 298 564 350
rect 616 298 756 350
rect 0 286 756 298
rect 0 234 140 286
rect 192 234 352 286
rect 404 234 564 286
rect 616 234 756 286
rect 0 222 756 234
rect 0 170 140 222
rect 192 170 352 222
rect 404 170 564 222
rect 616 170 756 222
rect 0 158 756 170
rect 0 106 140 158
rect 192 106 352 158
rect 404 106 564 158
rect 616 106 756 158
rect 0 100 756 106
<< labels >>
flabel comment s 166 597 166 597 0 FreeSans 300 0 0 0 S
flabel comment s 166 597 166 597 0 FreeSans 300 0 0 0 S
flabel comment s 272 597 272 597 0 FreeSans 300 0 0 0 S
flabel comment s 272 597 272 597 0 FreeSans 300 0 0 0 D
flabel comment s 378 597 378 597 0 FreeSans 300 0 0 0 S
flabel comment s 378 597 378 597 0 FreeSans 300 0 0 0 S
flabel comment s 484 597 484 597 0 FreeSans 300 0 0 0 S
flabel comment s 484 597 484 597 0 FreeSans 300 0 0 0 D
flabel comment s 590 597 590 597 0 FreeSans 300 0 0 0 S
flabel metal2 s 4 817 22 887 0 FreeSans 300 90 0 0 DRAIN
port 1 nsew
flabel metal2 s 3 312 23 376 0 FreeSans 300 90 0 0 SOURCE
port 3 nsew
flabel metal1 s 338 24 420 49 0 FreeSans 300 0 0 0 GATE
port 2 nsew
flabel metal1 s 51 714 51 714 7 FreeSans 300 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 699 704 699 704 7 FreeSans 300 90 0 0 SUBSTRATE
port 4 nsew
flabel metal1 s 339 1145 421 1170 0 FreeSans 300 0 0 0 GATE
port 2 nsew
<< properties >>
string GDS_END 6246124
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 6223778
<< end >>
