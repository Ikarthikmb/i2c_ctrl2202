magic
tech sky130A
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_0
timestamp 1644511149
transform -1 0 -7 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_1
timestamp 1644511149
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_2
timestamp 1644511149
transform 1 0 263 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_3
timestamp 1644511149
transform 1 0 426 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_4
timestamp 1644511149
transform 1 0 589 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_5
timestamp 1644511149
transform 1 0 752 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_6
timestamp 1644511149
transform 1 0 915 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_7
timestamp 1644511149
transform 1 0 1078 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_8
timestamp 1644511149
transform 1 0 1241 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 1269 675 1269 675 0 FreeSans 300 0 0 0 S
flabel comment s 1106 675 1106 675 0 FreeSans 300 0 0 0 D
flabel comment s 943 675 943 675 0 FreeSans 300 0 0 0 S
flabel comment s 780 675 780 675 0 FreeSans 300 0 0 0 D
flabel comment s 617 675 617 675 0 FreeSans 300 0 0 0 S
flabel comment s 454 675 454 675 0 FreeSans 300 0 0 0 D
flabel comment s 291 675 291 675 0 FreeSans 300 0 0 0 S
flabel comment s 128 675 128 675 0 FreeSans 300 0 0 0 D
flabel comment s -35 675 -35 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 8691024
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8685956
<< end >>
