magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1418 582
<< pwell >>
rect 505 157 712 203
rect 1195 157 1379 203
rect 1 21 1379 157
rect 29 -17 63 21
<< locali >>
rect 17 191 68 333
rect 176 289 247 391
rect 176 265 238 289
rect 170 191 238 265
rect 1306 299 1363 493
rect 942 253 986 265
rect 942 191 1202 253
rect 1329 165 1363 299
rect 1306 51 1363 165
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 17 367 69 527
rect 108 425 251 493
rect 285 425 440 493
rect 108 351 142 425
rect 102 292 142 351
rect 102 157 136 292
rect 281 265 372 391
rect 272 241 372 265
rect 406 275 440 425
rect 474 415 602 527
rect 636 417 680 493
rect 716 451 1098 527
rect 1132 417 1166 493
rect 1206 451 1272 527
rect 636 383 1090 417
rect 636 381 680 383
rect 474 327 680 381
rect 474 315 508 327
rect 406 241 602 275
rect 17 123 238 157
rect 272 141 340 241
rect 374 141 431 207
rect 465 199 602 241
rect 17 51 69 123
rect 103 17 169 89
rect 203 51 238 123
rect 465 107 499 199
rect 272 51 499 107
rect 533 17 602 165
rect 636 51 680 327
rect 716 315 798 349
rect 716 187 750 315
rect 832 299 992 349
rect 1028 321 1090 383
rect 1132 355 1272 417
rect 832 255 893 299
rect 1028 287 1122 321
rect 1156 287 1272 355
rect 1238 265 1272 287
rect 784 221 893 255
rect 716 153 801 187
rect 835 157 893 221
rect 1238 199 1292 265
rect 1238 157 1272 199
rect 716 51 782 153
rect 835 123 966 157
rect 816 17 882 89
rect 916 51 966 123
rect 1002 123 1272 157
rect 1002 51 1054 123
rect 1101 17 1272 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
<< metal1 >>
rect 0 561 1380 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1380 561
rect 0 496 1380 527
rect 0 17 1380 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1380 17
rect 0 -48 1380 -17
<< obsm1 >>
rect 293 320 351 329
rect 847 320 905 329
rect 293 292 905 320
rect 293 283 351 292
rect 847 283 905 292
rect 385 184 443 193
rect 755 184 813 193
rect 385 156 813 184
rect 385 147 443 156
rect 755 147 813 156
<< labels >>
rlabel locali s 942 191 1202 253 6 CLK
port 1 nsew clock input
rlabel locali s 942 253 986 265 6 CLK
port 1 nsew clock input
rlabel locali s 170 191 238 265 6 GATE
port 2 nsew signal input
rlabel locali s 176 265 238 289 6 GATE
port 2 nsew signal input
rlabel locali s 176 289 247 391 6 GATE
port 2 nsew signal input
rlabel locali s 17 191 68 333 6 SCE
port 3 nsew signal input
rlabel metal1 s 0 -48 1380 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 1379 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1195 157 1379 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 505 157 712 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 1418 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 1380 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 1306 51 1363 165 6 GCLK
port 8 nsew signal output
rlabel locali s 1329 165 1363 299 6 GCLK
port 8 nsew signal output
rlabel locali s 1306 299 1363 493 6 GCLK
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1380 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 419710
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 408734
<< end >>
