magic
tech sky130B
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdfm1sd2__example_55959141808765  sky130_fd_pr__hvdfm1sd2__example_55959141808765_0
timestamp 1644511149
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd__example_5595914180835  sky130_fd_pr__hvdfm1sd__example_5595914180835_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 128 265 128 265 0 FreeSans 300 0 0 0 D
flabel comment s -28 265 -28 265 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 27744374
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 27743446
<< end >>
