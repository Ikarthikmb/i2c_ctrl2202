/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/sky130A/libs.tech/ngspice/parasitics/sky130_fd_pr__model__parasitic__diodes_pw2dn.model.spice