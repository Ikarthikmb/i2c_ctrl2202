magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -66 377 834 897
<< pwell >>
rect 502 217 764 283
rect 4 43 764 217
rect -26 -43 794 43
<< locali >>
rect 121 382 307 652
rect 106 216 263 278
rect 383 216 490 278
rect 692 99 743 751
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 324 735 656 751
rect 324 701 334 735
rect 368 701 406 735
rect 440 701 478 735
rect 512 701 550 735
rect 584 701 622 735
rect 324 686 656 701
rect 29 346 79 556
rect 341 435 656 686
rect 585 346 651 387
rect 29 312 651 346
rect 29 99 72 312
rect 313 182 347 312
rect 106 113 277 182
rect 106 79 116 113
rect 150 79 233 113
rect 267 79 277 113
rect 313 99 393 182
rect 524 113 658 265
rect 106 73 277 79
rect 524 79 538 113
rect 572 79 610 113
rect 644 79 658 113
rect 524 73 658 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 334 701 368 735
rect 406 701 440 735
rect 478 701 512 735
rect 550 701 584 735
rect 622 701 656 735
rect 116 79 150 113
rect 233 79 267 113
rect 538 79 572 113
rect 610 79 644 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
<< metal1 >>
rect 0 831 768 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 768 831
rect 0 791 768 797
rect 0 735 768 763
rect 0 701 334 735
rect 368 701 406 735
rect 440 701 478 735
rect 512 701 550 735
rect 584 701 622 735
rect 656 701 768 735
rect 0 689 768 701
rect 0 113 768 125
rect 0 79 116 113
rect 150 79 233 113
rect 267 79 538 113
rect 572 79 610 113
rect 644 79 768 113
rect 0 51 768 79
rect 0 17 768 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 768 17
rect 0 -23 768 -17
<< labels >>
rlabel locali s 383 216 490 278 6 A
port 1 nsew signal input
rlabel locali s 121 382 307 652 6 B
port 2 nsew signal input
rlabel locali s 106 216 263 278 6 C
port 3 nsew signal input
rlabel metal1 s 0 51 768 125 6 VGND
port 4 nsew ground bidirectional
rlabel metal1 s 0 -23 768 23 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s -26 -43 794 43 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 4 43 764 217 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 502 217 764 283 6 VNB
port 5 nsew ground bidirectional
rlabel metal1 s 0 791 768 837 6 VPB
port 6 nsew power bidirectional
rlabel nwell s -66 377 834 897 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 689 768 763 6 VPWR
port 7 nsew power bidirectional
rlabel locali s 692 99 743 751 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 768 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 367552
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 357224
<< end >>
