magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 891 203
rect 30 -17 64 21
<< scnmos >>
rect 83 47 113 177
rect 167 47 197 177
rect 251 47 281 177
rect 335 47 365 177
rect 531 47 561 177
rect 615 47 645 177
rect 699 47 729 177
rect 783 47 813 177
<< scpmoshvt >>
rect 83 297 113 497
rect 167 297 197 497
rect 251 297 281 497
rect 335 297 365 497
rect 531 297 561 497
rect 615 297 645 497
rect 699 297 729 497
rect 783 297 813 497
<< ndiff >>
rect 27 163 83 177
rect 27 129 39 163
rect 73 129 83 163
rect 27 95 83 129
rect 27 61 39 95
rect 73 61 83 95
rect 27 47 83 61
rect 113 163 167 177
rect 113 129 123 163
rect 157 129 167 163
rect 113 47 167 129
rect 197 95 251 177
rect 197 61 207 95
rect 241 61 251 95
rect 197 47 251 61
rect 281 163 335 177
rect 281 129 291 163
rect 325 129 335 163
rect 281 47 335 129
rect 365 95 531 177
rect 365 61 375 95
rect 409 61 486 95
rect 520 61 531 95
rect 365 47 531 61
rect 561 95 615 177
rect 561 61 571 95
rect 605 61 615 95
rect 561 47 615 61
rect 645 163 699 177
rect 645 129 655 163
rect 689 129 699 163
rect 645 95 699 129
rect 645 61 655 95
rect 689 61 699 95
rect 645 47 699 61
rect 729 95 783 177
rect 729 61 739 95
rect 773 61 783 95
rect 729 47 783 61
rect 813 163 865 177
rect 813 129 823 163
rect 857 129 865 163
rect 813 95 865 129
rect 813 61 823 95
rect 857 61 865 95
rect 813 47 865 61
<< pdiff >>
rect 27 477 83 497
rect 27 443 39 477
rect 73 443 83 477
rect 27 409 83 443
rect 27 375 39 409
rect 73 375 83 409
rect 27 341 83 375
rect 27 307 39 341
rect 73 307 83 341
rect 27 297 83 307
rect 113 477 167 497
rect 113 443 123 477
rect 157 443 167 477
rect 113 409 167 443
rect 113 375 123 409
rect 157 375 167 409
rect 113 297 167 375
rect 197 477 251 497
rect 197 443 207 477
rect 241 443 251 477
rect 197 409 251 443
rect 197 375 207 409
rect 241 375 251 409
rect 197 341 251 375
rect 197 307 207 341
rect 241 307 251 341
rect 197 297 251 307
rect 281 409 335 497
rect 281 375 291 409
rect 325 375 335 409
rect 281 341 335 375
rect 281 307 291 341
rect 325 307 335 341
rect 281 297 335 307
rect 365 477 421 497
rect 365 443 375 477
rect 409 443 421 477
rect 365 409 421 443
rect 365 375 375 409
rect 409 375 421 409
rect 365 297 421 375
rect 475 477 531 497
rect 475 443 487 477
rect 521 443 531 477
rect 475 409 531 443
rect 475 375 487 409
rect 521 375 531 409
rect 475 297 531 375
rect 561 409 615 497
rect 561 375 571 409
rect 605 375 615 409
rect 561 341 615 375
rect 561 307 571 341
rect 605 307 615 341
rect 561 297 615 307
rect 645 477 699 497
rect 645 443 655 477
rect 689 443 699 477
rect 645 409 699 443
rect 645 375 655 409
rect 689 375 699 409
rect 645 341 699 375
rect 645 307 655 341
rect 689 307 699 341
rect 645 297 699 307
rect 729 477 783 497
rect 729 443 739 477
rect 773 443 783 477
rect 729 409 783 443
rect 729 375 739 409
rect 773 375 783 409
rect 729 297 783 375
rect 813 477 869 497
rect 813 443 823 477
rect 857 443 869 477
rect 813 409 869 443
rect 813 375 823 409
rect 857 375 869 409
rect 813 341 869 375
rect 813 307 823 341
rect 857 307 869 341
rect 813 297 869 307
<< ndiffc >>
rect 39 129 73 163
rect 39 61 73 95
rect 123 129 157 163
rect 207 61 241 95
rect 291 129 325 163
rect 375 61 409 95
rect 486 61 520 95
rect 571 61 605 95
rect 655 129 689 163
rect 655 61 689 95
rect 739 61 773 95
rect 823 129 857 163
rect 823 61 857 95
<< pdiffc >>
rect 39 443 73 477
rect 39 375 73 409
rect 39 307 73 341
rect 123 443 157 477
rect 123 375 157 409
rect 207 443 241 477
rect 207 375 241 409
rect 207 307 241 341
rect 291 375 325 409
rect 291 307 325 341
rect 375 443 409 477
rect 375 375 409 409
rect 487 443 521 477
rect 487 375 521 409
rect 571 375 605 409
rect 571 307 605 341
rect 655 443 689 477
rect 655 375 689 409
rect 655 307 689 341
rect 739 443 773 477
rect 739 375 773 409
rect 823 443 857 477
rect 823 375 857 409
rect 823 307 857 341
<< poly >>
rect 83 497 113 523
rect 167 497 197 523
rect 251 497 281 523
rect 335 497 365 523
rect 531 497 561 523
rect 615 497 645 523
rect 699 497 729 523
rect 783 497 813 523
rect 83 265 113 297
rect 167 265 197 297
rect 63 249 197 265
rect 63 215 79 249
rect 113 215 147 249
rect 181 215 197 249
rect 63 199 197 215
rect 83 177 113 199
rect 167 177 197 199
rect 251 265 281 297
rect 335 265 365 297
rect 531 265 561 297
rect 615 265 645 297
rect 251 249 385 265
rect 251 215 267 249
rect 301 215 335 249
rect 369 215 385 249
rect 251 199 385 215
rect 511 249 645 265
rect 511 215 527 249
rect 561 215 595 249
rect 629 215 645 249
rect 511 199 645 215
rect 251 177 281 199
rect 335 177 365 199
rect 531 177 561 199
rect 615 177 645 199
rect 699 265 729 297
rect 783 265 813 297
rect 699 249 833 265
rect 699 215 715 249
rect 749 215 783 249
rect 817 215 833 249
rect 699 199 833 215
rect 699 177 729 199
rect 783 177 813 199
rect 83 21 113 47
rect 167 21 197 47
rect 251 21 281 47
rect 335 21 365 47
rect 531 21 561 47
rect 615 21 645 47
rect 699 21 729 47
rect 783 21 813 47
<< polycont >>
rect 79 215 113 249
rect 147 215 181 249
rect 267 215 301 249
rect 335 215 369 249
rect 527 215 561 249
rect 595 215 629 249
rect 715 215 749 249
rect 783 215 817 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 30 477 81 493
rect 30 443 39 477
rect 73 443 81 477
rect 30 409 81 443
rect 30 375 39 409
rect 73 375 81 409
rect 30 341 81 375
rect 115 477 165 527
rect 115 443 123 477
rect 157 443 165 477
rect 115 409 165 443
rect 115 375 123 409
rect 157 375 165 409
rect 115 359 165 375
rect 199 477 417 493
rect 199 443 207 477
rect 241 459 375 477
rect 241 443 249 459
rect 199 409 249 443
rect 367 443 375 459
rect 409 443 417 477
rect 199 375 207 409
rect 241 375 249 409
rect 30 307 39 341
rect 73 325 81 341
rect 199 341 249 375
rect 199 325 207 341
rect 73 307 207 325
rect 241 307 249 341
rect 30 291 249 307
rect 283 409 333 425
rect 283 375 291 409
rect 325 375 333 409
rect 283 341 333 375
rect 367 409 417 443
rect 367 375 375 409
rect 409 375 417 409
rect 367 359 417 375
rect 479 477 697 493
rect 479 443 487 477
rect 521 459 655 477
rect 521 443 529 459
rect 479 409 529 443
rect 647 443 655 459
rect 689 443 697 477
rect 479 375 487 409
rect 521 375 529 409
rect 479 359 529 375
rect 563 409 613 425
rect 563 375 571 409
rect 605 375 613 409
rect 283 307 291 341
rect 325 325 333 341
rect 563 341 613 375
rect 563 325 571 341
rect 325 307 571 325
rect 605 307 613 341
rect 283 289 613 307
rect 647 409 697 443
rect 647 375 655 409
rect 689 375 697 409
rect 647 341 697 375
rect 731 477 781 527
rect 731 443 739 477
rect 773 443 781 477
rect 731 409 781 443
rect 731 375 739 409
rect 773 375 781 409
rect 731 359 781 375
rect 815 477 866 493
rect 815 443 823 477
rect 857 443 866 477
rect 815 409 866 443
rect 815 375 823 409
rect 857 375 866 409
rect 647 307 655 341
rect 689 325 697 341
rect 815 341 866 375
rect 815 325 823 341
rect 689 307 823 325
rect 857 307 866 341
rect 647 291 866 307
rect 40 249 197 257
rect 40 215 79 249
rect 113 215 147 249
rect 181 215 197 249
rect 231 249 385 255
rect 231 215 267 249
rect 301 215 335 249
rect 369 215 385 249
rect 419 181 468 289
rect 511 249 645 255
rect 511 215 527 249
rect 561 215 595 249
rect 629 215 645 249
rect 679 249 833 257
rect 679 215 715 249
rect 749 215 783 249
rect 817 215 833 249
rect 18 163 73 181
rect 18 129 39 163
rect 107 163 468 181
rect 107 129 123 163
rect 157 145 291 163
rect 157 129 173 145
rect 275 129 291 145
rect 325 145 468 163
rect 502 163 873 181
rect 502 145 655 163
rect 325 129 341 145
rect 18 95 73 129
rect 502 95 536 145
rect 639 129 655 145
rect 689 145 823 163
rect 689 129 705 145
rect 18 61 39 95
rect 73 61 207 95
rect 241 61 375 95
rect 409 61 486 95
rect 520 61 536 95
rect 571 95 605 111
rect 571 17 605 61
rect 639 95 705 129
rect 807 129 823 145
rect 857 129 873 163
rect 639 61 655 95
rect 689 61 705 95
rect 639 51 705 61
rect 739 95 773 111
rect 739 17 773 61
rect 807 95 873 129
rect 807 61 823 95
rect 857 61 873 95
rect 807 51 873 61
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 306 221 340 255 0 FreeSans 400 0 0 0 B2
port 4 nsew signal input
flabel locali s 122 221 156 255 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel locali s 398 289 432 323 0 FreeSans 400 0 0 0 Y
port 9 nsew signal output
flabel locali s 770 221 804 255 0 FreeSans 400 0 0 0 A1
port 1 nsew signal input
flabel locali s 586 221 620 255 0 FreeSans 400 0 0 0 A2
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 o22ai_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 1406564
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1398688
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 4.600 0.000 
<< end >>
