magic
tech sky130B
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdfl1sd2__example_55959141808385  sky130_fd_pr__hvdfl1sd2__example_55959141808385_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 145 70 145 70 0 FreeSans 300 0 0 0 D
flabel comment s -28 63 -28 63 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 48781068
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 48780274
<< end >>
