/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/nfet_20v0_nvt_iso/sky130_fd_pr__nfet_20v0_nvt_iso__sf_discrete.corner.spice