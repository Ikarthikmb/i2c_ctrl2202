magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -66 377 1122 897
<< pwell >>
rect 4 43 998 283
rect -26 -43 1082 43
<< mvnmos >>
rect 87 107 187 257
rect 243 107 343 257
rect 517 107 617 257
rect 659 107 759 257
rect 815 107 915 257
<< mvpmos >>
rect 87 443 187 743
rect 229 443 329 743
rect 431 443 531 743
rect 587 443 687 743
rect 869 443 969 743
<< mvndiff >>
rect 30 249 87 257
rect 30 215 42 249
rect 76 215 87 249
rect 30 149 87 215
rect 30 115 42 149
rect 76 115 87 149
rect 30 107 87 115
rect 187 249 243 257
rect 187 215 198 249
rect 232 215 243 249
rect 187 149 243 215
rect 187 115 198 149
rect 232 115 243 149
rect 187 107 243 115
rect 343 249 517 257
rect 343 215 354 249
rect 388 215 517 249
rect 343 149 517 215
rect 343 115 354 149
rect 388 115 517 149
rect 343 107 517 115
rect 617 107 659 257
rect 759 249 815 257
rect 759 215 770 249
rect 804 215 815 249
rect 759 149 815 215
rect 759 115 770 149
rect 804 115 815 149
rect 759 107 815 115
rect 915 249 972 257
rect 915 215 926 249
rect 960 215 972 249
rect 915 149 972 215
rect 915 115 926 149
rect 960 115 972 149
rect 915 107 972 115
<< mvpdiff >>
rect 30 735 87 743
rect 30 701 42 735
rect 76 701 87 735
rect 30 652 87 701
rect 30 618 42 652
rect 76 618 87 652
rect 30 568 87 618
rect 30 534 42 568
rect 76 534 87 568
rect 30 485 87 534
rect 30 451 42 485
rect 76 451 87 485
rect 30 443 87 451
rect 187 443 229 743
rect 329 735 431 743
rect 329 701 340 735
rect 374 701 431 735
rect 329 663 431 701
rect 329 629 340 663
rect 374 629 431 663
rect 329 591 431 629
rect 329 557 340 591
rect 374 557 431 591
rect 329 443 431 557
rect 531 735 587 743
rect 531 701 542 735
rect 576 701 587 735
rect 531 607 587 701
rect 531 573 542 607
rect 576 573 587 607
rect 531 443 587 573
rect 687 715 744 743
rect 687 681 698 715
rect 732 681 744 715
rect 687 443 744 681
rect 812 485 869 743
rect 812 451 824 485
rect 858 451 869 485
rect 812 443 869 451
rect 969 735 1026 743
rect 969 701 980 735
rect 1014 701 1026 735
rect 969 652 1026 701
rect 969 618 980 652
rect 1014 618 1026 652
rect 969 568 1026 618
rect 969 534 980 568
rect 1014 534 1026 568
rect 969 485 1026 534
rect 969 451 980 485
rect 1014 451 1026 485
rect 969 443 1026 451
<< mvndiffc >>
rect 42 215 76 249
rect 42 115 76 149
rect 198 215 232 249
rect 198 115 232 149
rect 354 215 388 249
rect 354 115 388 149
rect 770 215 804 249
rect 770 115 804 149
rect 926 215 960 249
rect 926 115 960 149
<< mvpdiffc >>
rect 42 701 76 735
rect 42 618 76 652
rect 42 534 76 568
rect 42 451 76 485
rect 340 701 374 735
rect 340 629 374 663
rect 340 557 374 591
rect 542 701 576 735
rect 542 573 576 607
rect 698 681 732 715
rect 824 451 858 485
rect 980 701 1014 735
rect 980 618 1014 652
rect 980 534 1014 568
rect 980 451 1014 485
<< mvpsubdiff >>
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< mvnsubdiff >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
<< mvpsubdiffcont >>
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< mvnsubdiffcont >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
<< poly >>
rect 87 743 187 769
rect 229 743 329 769
rect 431 743 531 769
rect 587 743 687 769
rect 869 743 969 769
rect 87 395 187 443
rect 87 361 128 395
rect 162 361 187 395
rect 229 421 329 443
rect 431 421 531 443
rect 229 395 531 421
rect 229 371 451 395
rect 87 257 187 361
rect 243 361 451 371
rect 485 361 531 395
rect 587 421 687 443
rect 869 421 969 443
rect 587 371 759 421
rect 243 329 531 361
rect 659 351 759 371
rect 243 283 617 329
rect 243 257 343 283
rect 431 279 617 283
rect 517 257 617 279
rect 659 317 696 351
rect 730 317 759 351
rect 659 257 759 317
rect 815 383 980 421
rect 815 349 926 383
rect 960 349 980 383
rect 815 321 980 349
rect 815 257 915 321
rect 87 81 187 107
rect 243 81 343 107
rect 517 81 617 107
rect 659 81 759 107
rect 815 81 915 107
<< polycont >>
rect 128 361 162 395
rect 451 361 485 395
rect 696 317 730 351
rect 926 349 960 383
<< locali >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 26 735 76 751
rect 26 701 42 735
rect 26 652 76 701
rect 26 618 42 652
rect 26 568 76 618
rect 26 534 42 568
rect 112 735 506 751
rect 146 701 184 735
rect 218 701 256 735
rect 290 701 328 735
rect 374 701 400 735
rect 434 701 472 735
rect 112 663 506 701
rect 112 629 340 663
rect 374 629 506 663
rect 112 591 506 629
rect 112 557 340 591
rect 374 557 506 591
rect 542 735 576 751
rect 542 625 576 701
rect 612 735 944 751
rect 612 701 617 735
rect 651 701 689 735
rect 723 715 761 735
rect 732 701 761 715
rect 795 701 833 735
rect 867 701 905 735
rect 939 701 944 735
rect 612 681 698 701
rect 732 681 944 701
rect 612 661 944 681
rect 980 735 1030 751
rect 1014 701 1030 735
rect 980 652 1030 701
rect 542 618 980 625
rect 1014 618 1030 652
rect 542 607 1030 618
rect 576 591 1030 607
rect 542 557 576 573
rect 980 568 1030 591
rect 26 521 76 534
rect 612 521 944 555
rect 26 487 646 521
rect 26 485 76 487
rect 26 451 42 485
rect 26 319 76 451
rect 793 451 824 485
rect 858 451 874 485
rect 112 395 302 411
rect 112 361 128 395
rect 162 361 302 395
rect 112 355 302 361
rect 409 395 647 430
rect 409 361 451 395
rect 485 361 647 395
rect 409 355 647 361
rect 268 319 302 355
rect 683 351 743 367
rect 683 319 696 351
rect 26 285 232 319
rect 268 317 696 319
rect 730 317 743 351
rect 268 301 743 317
rect 268 285 717 301
rect 182 249 232 285
rect 793 265 874 451
rect 910 399 944 521
rect 1014 534 1030 568
rect 980 485 1030 534
rect 1014 451 1030 485
rect 980 435 1030 451
rect 910 383 976 399
rect 910 349 926 383
rect 960 349 976 383
rect 910 333 976 349
rect 770 249 874 265
rect 18 215 42 249
rect 76 215 136 249
rect 18 149 136 215
rect 18 115 42 149
rect 76 115 136 149
rect 18 113 136 115
rect 18 79 24 113
rect 58 79 96 113
rect 130 79 136 113
rect 182 215 198 249
rect 182 149 232 215
rect 182 115 198 149
rect 182 99 232 115
rect 268 215 354 249
rect 388 215 734 249
rect 268 149 734 215
rect 268 115 354 149
rect 388 115 734 149
rect 268 113 734 115
rect 18 73 136 79
rect 302 79 340 113
rect 374 79 412 113
rect 446 79 484 113
rect 518 79 556 113
rect 590 79 628 113
rect 662 79 700 113
rect 804 215 874 249
rect 770 149 874 215
rect 804 115 874 149
rect 770 99 874 115
rect 910 249 1028 265
rect 910 215 926 249
rect 960 215 1028 249
rect 910 149 1028 215
rect 910 115 926 149
rect 960 115 1028 149
rect 910 113 1028 115
rect 268 73 734 79
rect 910 79 916 113
rect 950 79 988 113
rect 1022 79 1028 113
rect 910 73 1028 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
<< viali >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 415 797 449 831
rect 511 797 545 831
rect 607 797 641 831
rect 703 797 737 831
rect 799 797 833 831
rect 895 797 929 831
rect 991 797 1025 831
rect 112 701 146 735
rect 184 701 218 735
rect 256 701 290 735
rect 328 701 340 735
rect 340 701 362 735
rect 400 701 434 735
rect 472 701 506 735
rect 617 701 651 735
rect 689 715 723 735
rect 689 701 698 715
rect 698 701 723 715
rect 761 701 795 735
rect 833 701 867 735
rect 905 701 939 735
rect 24 79 58 113
rect 96 79 130 113
rect 268 79 302 113
rect 340 79 374 113
rect 412 79 446 113
rect 484 79 518 113
rect 556 79 590 113
rect 628 79 662 113
rect 700 79 734 113
rect 916 79 950 113
rect 988 79 1022 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
rect 415 -17 449 17
rect 511 -17 545 17
rect 607 -17 641 17
rect 703 -17 737 17
rect 799 -17 833 17
rect 895 -17 929 17
rect 991 -17 1025 17
<< metal1 >>
rect 0 831 1056 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 415 831
rect 449 797 511 831
rect 545 797 607 831
rect 641 797 703 831
rect 737 797 799 831
rect 833 797 895 831
rect 929 797 991 831
rect 1025 797 1056 831
rect 0 791 1056 797
rect 0 735 1056 763
rect 0 701 112 735
rect 146 701 184 735
rect 218 701 256 735
rect 290 701 328 735
rect 362 701 400 735
rect 434 701 472 735
rect 506 701 617 735
rect 651 701 689 735
rect 723 701 761 735
rect 795 701 833 735
rect 867 701 905 735
rect 939 701 1056 735
rect 0 689 1056 701
rect 0 113 1056 125
rect 0 79 24 113
rect 58 79 96 113
rect 130 79 268 113
rect 302 79 340 113
rect 374 79 412 113
rect 446 79 484 113
rect 518 79 556 113
rect 590 79 628 113
rect 662 79 700 113
rect 734 79 916 113
rect 950 79 988 113
rect 1022 79 1056 113
rect 0 51 1056 79
rect 0 17 1056 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 415 17
rect 449 -17 511 17
rect 545 -17 607 17
rect 641 -17 703 17
rect 737 -17 799 17
rect 833 -17 895 17
rect 929 -17 991 17
rect 1025 -17 1056 17
rect 0 -23 1056 -17
<< labels >>
rlabel comment s 0 0 0 0 4 xor2_1
flabel metal1 s 0 51 1056 125 0 FreeSans 340 0 0 0 VGND
port 3 nsew ground bidirectional
flabel metal1 s 0 0 1056 23 0 FreeSans 340 0 0 0 VNB
port 4 nsew ground bidirectional
flabel metal1 s 0 689 1056 763 0 FreeSans 340 0 0 0 VPWR
port 6 nsew power bidirectional
flabel metal1 s 0 791 1056 814 0 FreeSans 340 0 0 0 VPB
port 5 nsew power bidirectional
flabel locali s 415 390 449 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 511 390 545 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 607 390 641 424 0 FreeSans 340 0 0 0 A
port 1 nsew signal input
flabel locali s 799 168 833 202 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 799 242 833 276 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 799 316 833 350 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 799 390 833 424 0 FreeSans 340 0 0 0 X
port 7 nsew signal output
flabel locali s 703 316 737 350 0 FreeSans 340 0 0 0 B
port 2 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 1056 814
string GDS_END 743414
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 731354
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
<< end >>
