/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/npn_05v5/sky130_fd_pr__npn_05v5_W1p00L1p00.model.spice