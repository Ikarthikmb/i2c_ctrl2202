magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1169 203
rect 29 -17 63 21
<< locali >>
rect 745 393 787 425
rect 1009 393 1059 425
rect 745 359 1059 393
rect 1009 325 1059 359
rect 158 289 620 323
rect 158 257 192 289
rect 97 215 192 257
rect 586 257 620 289
rect 251 215 541 255
rect 586 215 791 257
rect 1009 283 1179 325
rect 1101 95 1179 283
rect 917 61 1179 95
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 17 393 80 493
rect 114 427 164 527
rect 198 393 248 493
rect 282 427 332 527
rect 366 393 416 493
rect 478 425 528 493
rect 562 427 612 527
rect 646 459 871 493
rect 646 425 711 459
rect 821 427 871 459
rect 925 427 975 527
rect 17 391 416 393
rect 17 357 696 391
rect 1093 359 1179 527
rect 17 179 63 357
rect 662 325 696 357
rect 662 291 961 325
rect 927 249 961 291
rect 927 215 1059 249
rect 17 129 172 179
rect 206 145 424 181
rect 206 95 256 145
rect 21 51 256 95
rect 290 17 324 111
rect 358 51 424 145
rect 486 17 520 181
rect 554 145 1067 181
rect 554 51 620 145
rect 654 17 688 111
rect 722 51 795 145
rect 1001 129 1067 145
rect 829 17 863 111
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< obsm1 >>
rect 481 456 539 465
rect 665 456 723 465
rect 481 428 723 456
rect 481 419 539 428
rect 665 419 723 428
<< labels >>
rlabel locali s 251 215 541 255 6 A
port 1 nsew signal input
rlabel locali s 586 215 791 257 6 B
port 2 nsew signal input
rlabel locali s 586 257 620 289 6 B
port 2 nsew signal input
rlabel locali s 97 215 192 257 6 B
port 2 nsew signal input
rlabel locali s 158 257 192 289 6 B
port 2 nsew signal input
rlabel locali s 158 289 620 323 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1169 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 917 61 1179 95 6 Y
port 7 nsew signal output
rlabel locali s 1101 95 1179 283 6 Y
port 7 nsew signal output
rlabel locali s 1009 283 1179 325 6 Y
port 7 nsew signal output
rlabel locali s 1009 325 1059 359 6 Y
port 7 nsew signal output
rlabel locali s 745 359 1059 393 6 Y
port 7 nsew signal output
rlabel locali s 1009 393 1059 425 6 Y
port 7 nsew signal output
rlabel locali s 745 393 787 425 6 Y
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 500234
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 491554
<< end >>
