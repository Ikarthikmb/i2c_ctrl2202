magic
tech sky130B
timestamp 1644511149
<< pwell >>
rect -13 -13 163 1513
<< nsubdiff >>
rect 0 0 150 1500
use sky130_fd_io__gnd2gnd_strap  sky130_fd_io__gnd2gnd_strap_0
timestamp 1644511149
transform 1 0 0 0 1 0
box 0 0 150 1500
<< properties >>
string GDS_END 15525138
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 15524954
<< end >>
