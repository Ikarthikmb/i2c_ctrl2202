magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect 25 436 791 1168
<< pwell >>
rect 79 -22 751 230
<< mvnmos >>
rect 158 4 278 204
rect 362 4 482 204
rect 538 4 658 204
<< mvpmos >>
rect 158 502 278 1102
rect 362 502 482 1102
rect 538 502 658 1102
<< mvndiff >>
rect 105 192 158 204
rect 105 158 113 192
rect 147 158 158 192
rect 105 124 158 158
rect 105 90 113 124
rect 147 90 158 124
rect 105 56 158 90
rect 105 22 113 56
rect 147 22 158 56
rect 105 4 158 22
rect 278 192 362 204
rect 278 158 303 192
rect 337 158 362 192
rect 278 124 362 158
rect 278 90 303 124
rect 337 90 362 124
rect 278 56 362 90
rect 278 22 303 56
rect 337 22 362 56
rect 278 4 362 22
rect 482 192 538 204
rect 482 158 493 192
rect 527 158 538 192
rect 482 124 538 158
rect 482 90 493 124
rect 527 90 538 124
rect 482 56 538 90
rect 482 22 493 56
rect 527 22 538 56
rect 482 4 538 22
rect 658 192 725 204
rect 658 158 683 192
rect 717 158 725 192
rect 658 124 725 158
rect 658 90 683 124
rect 717 90 725 124
rect 658 56 725 90
rect 658 22 683 56
rect 717 22 725 56
rect 658 4 725 22
<< mvpdiff >>
rect 91 1090 158 1102
rect 91 1056 99 1090
rect 133 1056 158 1090
rect 91 1022 158 1056
rect 91 988 99 1022
rect 133 988 158 1022
rect 91 954 158 988
rect 91 920 99 954
rect 133 920 158 954
rect 91 886 158 920
rect 91 852 99 886
rect 133 852 158 886
rect 91 818 158 852
rect 91 784 99 818
rect 133 784 158 818
rect 91 750 158 784
rect 91 716 99 750
rect 133 716 158 750
rect 91 682 158 716
rect 91 648 99 682
rect 133 648 158 682
rect 91 614 158 648
rect 91 580 99 614
rect 133 580 158 614
rect 91 502 158 580
rect 278 1090 362 1102
rect 278 1056 303 1090
rect 337 1056 362 1090
rect 278 1022 362 1056
rect 278 988 303 1022
rect 337 988 362 1022
rect 278 954 362 988
rect 278 920 303 954
rect 337 920 362 954
rect 278 886 362 920
rect 278 852 303 886
rect 337 852 362 886
rect 278 818 362 852
rect 278 784 303 818
rect 337 784 362 818
rect 278 750 362 784
rect 278 716 303 750
rect 337 716 362 750
rect 278 682 362 716
rect 278 648 303 682
rect 337 648 362 682
rect 278 614 362 648
rect 278 580 303 614
rect 337 580 362 614
rect 278 502 362 580
rect 482 1090 538 1102
rect 482 1056 493 1090
rect 527 1056 538 1090
rect 482 1022 538 1056
rect 482 988 493 1022
rect 527 988 538 1022
rect 482 954 538 988
rect 482 920 493 954
rect 527 920 538 954
rect 482 886 538 920
rect 482 852 493 886
rect 527 852 538 886
rect 482 818 538 852
rect 482 784 493 818
rect 527 784 538 818
rect 482 750 538 784
rect 482 716 493 750
rect 527 716 538 750
rect 482 682 538 716
rect 482 648 493 682
rect 527 648 538 682
rect 482 614 538 648
rect 482 580 493 614
rect 527 580 538 614
rect 482 502 538 580
rect 658 1090 725 1102
rect 658 1056 683 1090
rect 717 1056 725 1090
rect 658 1022 725 1056
rect 658 988 683 1022
rect 717 988 725 1022
rect 658 954 725 988
rect 658 920 683 954
rect 717 920 725 954
rect 658 886 725 920
rect 658 852 683 886
rect 717 852 725 886
rect 658 818 725 852
rect 658 784 683 818
rect 717 784 725 818
rect 658 750 725 784
rect 658 716 683 750
rect 717 716 725 750
rect 658 682 725 716
rect 658 648 683 682
rect 717 648 725 682
rect 658 614 725 648
rect 658 580 683 614
rect 717 580 725 614
rect 658 502 725 580
<< mvndiffc >>
rect 113 158 147 192
rect 113 90 147 124
rect 113 22 147 56
rect 303 158 337 192
rect 303 90 337 124
rect 303 22 337 56
rect 493 158 527 192
rect 493 90 527 124
rect 493 22 527 56
rect 683 158 717 192
rect 683 90 717 124
rect 683 22 717 56
<< mvpdiffc >>
rect 99 1056 133 1090
rect 99 988 133 1022
rect 99 920 133 954
rect 99 852 133 886
rect 99 784 133 818
rect 99 716 133 750
rect 99 648 133 682
rect 99 580 133 614
rect 303 1056 337 1090
rect 303 988 337 1022
rect 303 920 337 954
rect 303 852 337 886
rect 303 784 337 818
rect 303 716 337 750
rect 303 648 337 682
rect 303 580 337 614
rect 493 1056 527 1090
rect 493 988 527 1022
rect 493 920 527 954
rect 493 852 527 886
rect 493 784 527 818
rect 493 716 527 750
rect 493 648 527 682
rect 493 580 527 614
rect 683 1056 717 1090
rect 683 988 717 1022
rect 683 920 717 954
rect 683 852 717 886
rect 683 784 717 818
rect 683 716 717 750
rect 683 648 717 682
rect 683 580 717 614
<< poly >>
rect 158 1102 278 1128
rect 362 1102 482 1128
rect 538 1102 658 1128
rect 158 454 278 502
rect 158 420 201 454
rect 235 420 278 454
rect 158 386 278 420
rect 158 352 201 386
rect 235 352 278 386
rect 158 204 278 352
rect 362 454 482 502
rect 362 420 405 454
rect 439 420 482 454
rect 362 386 482 420
rect 362 352 405 386
rect 439 352 482 386
rect 362 204 482 352
rect 538 454 658 502
rect 538 420 581 454
rect 615 420 658 454
rect 538 386 658 420
rect 538 352 581 386
rect 615 352 658 386
rect 538 204 658 352
rect 158 -22 278 4
rect 362 -22 482 4
rect 538 -22 658 4
<< polycont >>
rect 201 420 235 454
rect 201 352 235 386
rect 405 420 439 454
rect 405 352 439 386
rect 581 420 615 454
rect 581 352 615 386
<< locali >>
rect 683 1136 717 1176
rect 91 1090 140 1107
rect 91 1056 99 1090
rect 133 1056 140 1090
rect 91 1022 140 1056
rect 91 988 99 1022
rect 133 988 140 1022
rect 91 954 140 988
rect 91 920 99 954
rect 133 920 140 954
rect 91 886 140 920
rect 91 852 99 886
rect 133 852 140 886
rect 91 818 140 852
rect 91 784 99 818
rect 133 784 140 818
rect 91 750 140 784
rect 91 716 99 750
rect 133 716 140 750
rect 91 682 140 716
rect 91 648 99 682
rect 133 648 140 682
rect 91 614 140 648
rect 91 580 99 614
rect 133 580 140 614
rect 91 298 140 580
rect 303 1090 337 1106
rect 303 1022 337 1056
rect 303 954 337 988
rect 303 886 337 920
rect 303 818 337 852
rect 303 750 337 784
rect 303 682 337 716
rect 303 614 337 648
rect 303 564 337 580
rect 493 1090 527 1106
rect 493 1022 527 1056
rect 493 954 527 988
rect 493 886 527 920
rect 493 818 527 852
rect 493 750 527 784
rect 493 682 527 716
rect 493 614 527 648
rect 493 564 527 580
rect 683 1090 717 1102
rect 683 1022 717 1030
rect 683 954 717 988
rect 683 886 717 920
rect 683 818 717 852
rect 683 750 717 784
rect 683 682 717 716
rect 683 614 717 648
rect 683 564 717 580
rect 185 420 201 454
rect 235 420 251 454
rect 185 386 251 420
rect 185 352 201 386
rect 235 352 251 386
rect 389 420 405 454
rect 439 420 455 454
rect 389 386 455 420
rect 389 352 405 386
rect 439 352 455 386
rect 565 420 581 454
rect 615 420 631 454
rect 565 386 631 420
rect 565 352 581 386
rect 615 352 631 386
rect 91 242 537 298
rect 105 192 158 242
rect 105 158 113 192
rect 147 158 158 192
rect 105 124 158 158
rect 105 90 113 124
rect 147 90 158 124
rect 105 56 158 90
rect 105 22 113 56
rect 147 22 158 56
rect 105 6 158 22
rect 303 192 337 208
rect 303 124 337 158
rect 303 59 337 90
rect 303 -13 337 22
rect 482 192 537 242
rect 482 158 493 192
rect 527 158 537 192
rect 482 124 537 158
rect 482 90 493 124
rect 527 90 537 124
rect 482 56 537 90
rect 482 22 493 56
rect 527 22 537 56
rect 482 6 537 22
rect 683 192 717 208
rect 683 124 717 158
rect 683 59 717 90
rect 303 -85 337 -47
rect 683 -13 717 22
rect 683 -85 717 -47
<< viali >>
rect 683 1102 717 1136
rect 683 1056 717 1064
rect 683 1030 717 1056
rect 303 56 337 59
rect 303 25 337 56
rect 683 56 717 59
rect 683 25 717 56
rect 303 -47 337 -13
rect 303 -119 337 -85
rect 683 -47 717 -13
rect 683 -119 717 -85
<< metal1 >>
rect 260 1136 768 1276
rect 260 1102 683 1136
rect 717 1102 768 1136
rect 260 1064 768 1102
rect 260 1030 683 1064
rect 717 1030 768 1064
rect 260 1018 768 1030
rect 282 59 768 71
rect 282 25 303 59
rect 337 25 683 59
rect 717 25 768 59
rect 282 -13 768 25
rect 282 -47 303 -13
rect 337 -47 683 -13
rect 717 -47 768 -13
rect 282 -85 768 -47
rect 282 -119 303 -85
rect 337 -119 683 -85
rect 717 -119 768 -85
rect 282 -131 768 -119
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808139  sky130_fd_pr__model__nfet_highvoltage__example_55959141808139_0
timestamp 1644511149
transform -1 0 658 0 -1 204
box -42 0 338 97
use sky130_fd_pr__model__nfet_highvoltage__example_55959141808183  sky130_fd_pr__model__nfet_highvoltage__example_55959141808183_0
timestamp 1644511149
transform -1 0 278 0 -1 204
box -42 0 148 97
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_0
timestamp 1644511149
transform 1 0 158 0 -1 1102
box -42 0 145 300
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808141  sky130_fd_pr__model__pfet_highvoltage__example_55959141808141_1
timestamp 1644511149
transform 1 0 362 0 -1 1102
box -42 0 145 300
use sky130_fd_pr__model__pfet_highvoltage__example_55959141808184  sky130_fd_pr__model__pfet_highvoltage__example_55959141808184_0
timestamp 1644511149
transform -1 0 658 0 -1 1102
box -42 0 148 267
use sky130_fd_pr__via_l1m1__example_559591418084  sky130_fd_pr__via_l1m1__example_559591418084_0
timestamp 1644511149
transform 0 -1 717 -1 0 1136
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_0
timestamp 1644511149
transform 0 -1 337 -1 0 59
box 0 0 1 1
use sky130_fd_pr__via_l1m1__example_5595914180897  sky130_fd_pr__via_l1m1__example_5595914180897_1
timestamp 1644511149
transform 0 -1 717 -1 0 59
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_0
timestamp 1644511149
transform 0 -1 251 -1 0 470
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_1
timestamp 1644511149
transform 0 -1 455 -1 0 470
box 0 0 1 1
use sky130_fd_pr__via_pol1__example_559591418083  sky130_fd_pr__via_pol1__example_559591418083_2
timestamp 1644511149
transform 0 -1 631 -1 0 470
box 0 0 1 1
<< properties >>
string GDS_END 37332626
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 37331094
<< end >>
