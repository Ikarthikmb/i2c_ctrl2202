magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 1 21 367 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 259 47 289 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 259 297 289 497
<< ndiff >>
rect 27 99 79 177
rect 27 65 35 99
rect 69 65 79 99
rect 27 47 79 65
rect 109 47 163 177
rect 193 47 259 177
rect 289 161 341 177
rect 289 127 299 161
rect 333 127 341 161
rect 289 93 341 127
rect 289 59 299 93
rect 333 59 341 93
rect 289 47 341 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 349 79 383
rect 27 315 35 349
rect 69 315 79 349
rect 27 297 79 315
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 417 163 451
rect 109 383 119 417
rect 153 383 163 417
rect 109 349 163 383
rect 109 315 119 349
rect 153 315 163 349
rect 109 297 163 315
rect 193 485 259 497
rect 193 451 203 485
rect 237 451 259 485
rect 193 417 259 451
rect 193 383 203 417
rect 237 383 259 417
rect 193 297 259 383
rect 289 485 341 497
rect 289 451 299 485
rect 333 451 341 485
rect 289 417 341 451
rect 289 383 299 417
rect 333 383 341 417
rect 289 349 341 383
rect 289 315 299 349
rect 333 315 341 349
rect 289 297 341 315
<< ndiffc >>
rect 35 65 69 99
rect 299 127 333 161
rect 299 59 333 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 35 315 69 349
rect 119 451 153 485
rect 119 383 153 417
rect 119 315 153 349
rect 203 451 237 485
rect 203 383 237 417
rect 299 451 333 485
rect 299 383 333 417
rect 299 315 333 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 259 497 289 523
rect 79 265 109 297
rect 22 249 109 265
rect 22 215 32 249
rect 66 215 109 249
rect 22 199 109 215
rect 79 177 109 199
rect 163 265 193 297
rect 259 265 289 297
rect 163 249 217 265
rect 163 215 173 249
rect 207 215 217 249
rect 163 199 217 215
rect 259 249 338 265
rect 259 215 294 249
rect 328 215 338 249
rect 259 199 338 215
rect 163 177 193 199
rect 259 177 289 199
rect 79 21 109 47
rect 163 21 193 47
rect 259 21 289 47
<< polycont >>
rect 32 215 66 249
rect 173 215 207 249
rect 294 215 328 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 18 485 69 527
rect 18 451 35 485
rect 18 417 69 451
rect 18 383 35 417
rect 18 349 69 383
rect 18 315 35 349
rect 18 299 69 315
rect 103 485 169 493
rect 103 451 119 485
rect 153 451 169 485
rect 103 417 169 451
rect 103 383 119 417
rect 153 383 169 417
rect 103 349 169 383
rect 203 485 249 527
rect 237 451 249 485
rect 203 417 249 451
rect 237 383 249 417
rect 203 367 249 383
rect 283 485 349 493
rect 283 451 299 485
rect 333 451 349 485
rect 283 417 349 451
rect 283 383 299 417
rect 333 383 349 417
rect 103 315 119 349
rect 153 333 169 349
rect 283 349 349 383
rect 283 333 299 349
rect 153 315 299 333
rect 333 315 349 349
rect 103 299 349 315
rect 22 249 66 265
rect 22 215 32 249
rect 22 149 66 215
rect 103 119 139 299
rect 173 249 248 265
rect 207 215 248 249
rect 173 153 248 215
rect 289 249 351 265
rect 289 215 294 249
rect 328 215 351 249
rect 289 199 351 215
rect 283 161 349 165
rect 283 127 299 161
rect 333 127 349 161
rect 283 119 349 127
rect 18 99 69 115
rect 18 65 35 99
rect 18 17 69 65
rect 103 93 349 119
rect 103 59 299 93
rect 333 59 349 93
rect 103 51 349 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
<< metal1 >>
rect 0 561 368 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 368 561
rect 0 496 368 527
rect 0 17 368 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 368 17
rect 0 -48 368 -17
<< labels >>
flabel locali s 122 85 156 119 0 FreeSans 250 0 0 0 Y
port 8 nsew signal output
flabel locali s 306 221 340 255 0 FreeSans 250 0 0 0 A
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 250 0 0 0 C
port 3 nsew signal input
flabel locali s 214 221 248 255 0 FreeSans 250 0 0 0 B
port 2 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand3_1
rlabel metal1 s 0 -48 368 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 368 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 368 544
string GDS_END 1834052
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1829710
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 9.200 0.000 
<< end >>
