magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< pwell >>
rect 1992 3688 2144 3844
<< obsli1 >>
rect 271 4592 1996 4601
rect 2353 4592 4078 4601
rect 271 4558 1997 4592
rect 2353 4558 4079 4592
rect 271 4549 1996 4558
rect 2353 4549 4078 4558
rect 93 4308 4257 4468
rect 93 2646 235 4308
rect 290 3540 324 4274
rect 360 3574 394 4308
rect 430 3540 464 4274
rect 500 3574 534 4308
rect 570 3540 604 4274
rect 640 3574 674 4308
rect 710 3540 744 4274
rect 780 3574 814 4308
rect 850 3540 884 4274
rect 920 3574 954 4308
rect 990 3540 1024 4274
rect 1060 3577 1208 4308
rect 1060 3576 1180 3577
rect 290 3414 1052 3540
rect 290 2680 324 3414
rect 360 2646 394 3380
rect 430 2680 464 3414
rect 500 2646 534 3380
rect 570 2680 604 3414
rect 640 2646 674 3380
rect 710 2680 744 3414
rect 780 2646 814 3380
rect 850 2680 884 3414
rect 920 2646 954 3380
rect 990 2680 1024 3414
rect 1088 3378 1180 3576
rect 1244 3540 1278 4274
rect 1314 3574 1348 4308
rect 1384 3540 1418 4274
rect 1454 3574 1488 4308
rect 1524 3540 1558 4274
rect 1594 3574 1628 4308
rect 1664 3540 1698 4274
rect 1734 3574 1768 4308
rect 1804 3540 1838 4274
rect 1874 3574 1908 4308
rect 1944 3540 1978 4274
rect 1216 3414 1978 3540
rect 1060 2646 1208 3378
rect 1244 2680 1278 3414
rect 1314 2646 1348 3380
rect 1384 2680 1418 3414
rect 1454 2646 1488 3380
rect 1524 2680 1558 3414
rect 1594 2646 1628 3380
rect 1664 2680 1698 3414
rect 1734 2646 1768 3380
rect 1804 2680 1838 3414
rect 1874 2646 1908 3380
rect 1944 2680 1978 3414
rect 2033 2646 2317 4308
rect 2372 3540 2406 4274
rect 2442 3574 2476 4308
rect 2512 3540 2546 4274
rect 2582 3574 2616 4308
rect 2652 3540 2686 4274
rect 2722 3574 2756 4308
rect 2792 3540 2826 4274
rect 2862 3574 2896 4308
rect 2932 3540 2966 4274
rect 3002 3574 3036 4308
rect 3072 3540 3106 4274
rect 3142 3577 3290 4308
rect 3142 3576 3262 3577
rect 2372 3414 3134 3540
rect 2372 2680 2406 3414
rect 2442 2646 2476 3380
rect 2512 2680 2546 3414
rect 2582 2646 2616 3380
rect 2652 2680 2686 3414
rect 2722 2646 2756 3380
rect 2792 2680 2826 3414
rect 2862 2646 2896 3380
rect 2932 2680 2966 3414
rect 3002 2646 3036 3380
rect 3072 2680 3106 3414
rect 3170 3378 3262 3576
rect 3326 3540 3360 4274
rect 3396 3574 3430 4308
rect 3466 3540 3500 4274
rect 3536 3574 3570 4308
rect 3606 3540 3640 4274
rect 3676 3574 3710 4308
rect 3746 3540 3780 4274
rect 3816 3574 3850 4308
rect 3886 3540 3920 4274
rect 3956 3574 3990 4308
rect 4026 3540 4060 4274
rect 3298 3414 4060 3540
rect 3142 2646 3290 3378
rect 3326 2680 3360 3414
rect 3396 2646 3430 3380
rect 3466 2680 3500 3414
rect 3536 2646 3570 3380
rect 3606 2680 3640 3414
rect 3676 2646 3710 3380
rect 3746 2680 3780 3414
rect 3816 2646 3850 3380
rect 3886 2680 3920 3414
rect 3956 2646 3990 3380
rect 4026 2680 4060 3414
rect 4115 2646 4257 4308
rect 93 2486 4257 2646
rect 271 2422 1996 2431
rect 2353 2422 4078 2431
rect 271 2388 1997 2422
rect 2353 2388 4079 2422
rect 271 2379 1996 2388
rect 2353 2379 4078 2388
rect 271 2284 1996 2293
rect 2353 2284 4078 2293
rect 271 2250 1997 2284
rect 2353 2250 4079 2284
rect 271 2241 1996 2250
rect 2353 2241 4078 2250
rect 93 2000 4257 2160
rect 93 338 235 2000
rect 290 1232 324 1966
rect 360 1266 394 2000
rect 430 1232 464 1966
rect 500 1266 534 2000
rect 570 1232 604 1966
rect 640 1266 674 2000
rect 710 1232 744 1966
rect 780 1266 814 2000
rect 850 1232 884 1966
rect 920 1266 954 2000
rect 990 1232 1024 1966
rect 1060 1269 1208 2000
rect 1060 1268 1180 1269
rect 290 1106 1052 1232
rect 290 372 324 1106
rect 360 338 394 1072
rect 430 372 464 1106
rect 500 338 534 1072
rect 570 372 604 1106
rect 640 338 674 1072
rect 710 372 744 1106
rect 780 338 814 1072
rect 850 372 884 1106
rect 920 338 954 1072
rect 990 372 1024 1106
rect 1088 1070 1180 1268
rect 1244 1232 1278 1966
rect 1314 1266 1348 2000
rect 1384 1232 1418 1966
rect 1454 1266 1488 2000
rect 1524 1232 1558 1966
rect 1594 1266 1628 2000
rect 1664 1232 1698 1966
rect 1734 1266 1768 2000
rect 1804 1232 1838 1966
rect 1874 1266 1908 2000
rect 1944 1232 1978 1966
rect 1216 1106 1978 1232
rect 1060 338 1208 1070
rect 1244 372 1278 1106
rect 1314 338 1348 1072
rect 1384 372 1418 1106
rect 1454 338 1488 1072
rect 1524 372 1558 1106
rect 1594 338 1628 1072
rect 1664 372 1698 1106
rect 1734 338 1768 1072
rect 1804 372 1838 1106
rect 1874 338 1908 1072
rect 1944 372 1978 1106
rect 2033 338 2317 2000
rect 2372 1232 2406 1966
rect 2442 1266 2476 2000
rect 2512 1232 2546 1966
rect 2582 1266 2616 2000
rect 2652 1232 2686 1966
rect 2722 1266 2756 2000
rect 2792 1232 2826 1966
rect 2862 1266 2896 2000
rect 2932 1232 2966 1966
rect 3002 1266 3036 2000
rect 3072 1232 3106 1966
rect 3142 1269 3290 2000
rect 3142 1268 3262 1269
rect 2372 1106 3134 1232
rect 2372 372 2406 1106
rect 2442 338 2476 1072
rect 2512 372 2546 1106
rect 2582 338 2616 1072
rect 2652 372 2686 1106
rect 2722 338 2756 1072
rect 2792 372 2826 1106
rect 2862 338 2896 1072
rect 2932 372 2966 1106
rect 3002 338 3036 1072
rect 3072 372 3106 1106
rect 3170 1070 3262 1268
rect 3326 1232 3360 1966
rect 3396 1266 3430 2000
rect 3466 1232 3500 1966
rect 3536 1266 3570 2000
rect 3606 1232 3640 1966
rect 3676 1266 3710 2000
rect 3746 1232 3780 1966
rect 3816 1266 3850 2000
rect 3886 1232 3920 1966
rect 3956 1266 3990 2000
rect 4026 1232 4060 1966
rect 3298 1106 4060 1232
rect 3142 338 3290 1070
rect 3326 372 3360 1106
rect 3396 338 3430 1072
rect 3466 372 3500 1106
rect 3536 338 3570 1072
rect 3606 372 3640 1106
rect 3676 338 3710 1072
rect 3746 372 3780 1106
rect 3816 338 3850 1072
rect 3886 372 3920 1106
rect 3956 338 3990 1072
rect 4026 372 4060 1106
rect 4115 338 4257 2000
rect 93 178 4257 338
rect 271 114 1996 123
rect 2353 114 4078 123
rect 271 80 1997 114
rect 2353 80 4079 114
rect 271 71 1996 80
rect 2353 71 4078 80
<< obsm1 >>
rect 93 4629 4257 4659
rect 93 4362 243 4629
rect 271 4392 1996 4601
rect 93 4308 1024 4362
rect 93 4218 262 4308
rect 1052 4274 1216 4392
rect 2024 4362 2325 4629
rect 2353 4392 4078 4601
rect 1244 4308 3106 4362
rect 290 4246 1978 4274
rect 93 4190 1024 4218
rect 93 4106 262 4190
rect 1052 4162 1216 4246
rect 2006 4218 2344 4308
rect 3134 4274 3298 4392
rect 4106 4362 4257 4629
rect 3326 4308 4257 4362
rect 2372 4246 4060 4274
rect 1244 4190 3106 4218
rect 290 4134 1978 4162
rect 93 4078 1024 4106
rect 93 3994 262 4078
rect 1052 4050 1216 4134
rect 2006 4106 2344 4190
rect 3134 4162 3298 4246
rect 4088 4218 4257 4308
rect 3326 4190 4257 4218
rect 2372 4134 4060 4162
rect 1244 4078 3106 4106
rect 290 4022 1978 4050
rect 93 3966 1024 3994
rect 93 3882 262 3966
rect 1052 3938 1216 4022
rect 2006 3994 2344 4078
rect 3134 4050 3298 4134
rect 4088 4106 4257 4190
rect 3326 4078 4257 4106
rect 2372 4022 4060 4050
rect 1244 3966 3106 3994
rect 290 3910 1978 3938
rect 93 3854 1024 3882
rect 93 3770 262 3854
rect 1052 3826 1216 3910
rect 2006 3882 2344 3966
rect 3134 3938 3298 4022
rect 4088 3994 4257 4078
rect 3326 3966 4257 3994
rect 2372 3910 4060 3938
rect 1244 3854 3106 3882
rect 290 3798 1978 3826
rect 93 3742 1024 3770
rect 93 3658 262 3742
rect 1052 3714 1216 3798
rect 2006 3770 2344 3854
rect 3134 3826 3298 3910
rect 4088 3882 4257 3966
rect 3326 3854 4257 3882
rect 2372 3798 4060 3826
rect 1244 3742 3106 3770
rect 290 3686 1978 3714
rect 93 3630 1024 3658
rect 93 3324 262 3630
rect 1052 3602 1216 3686
rect 2006 3658 2344 3742
rect 3134 3714 3298 3798
rect 4088 3770 4257 3854
rect 3326 3742 4257 3770
rect 2372 3686 4060 3714
rect 1244 3630 3106 3658
rect 290 3574 1978 3602
rect 1052 3540 1216 3574
rect 290 3414 1978 3540
rect 1052 3380 1216 3414
rect 290 3352 1978 3380
rect 93 3296 1024 3324
rect 93 3212 262 3296
rect 1052 3268 1216 3352
rect 2006 3324 2344 3630
rect 3134 3602 3298 3686
rect 4088 3658 4257 3742
rect 3326 3630 4257 3658
rect 2372 3574 4060 3602
rect 3134 3540 3298 3574
rect 2372 3414 4060 3540
rect 3134 3380 3298 3414
rect 2372 3352 4060 3380
rect 1244 3296 3106 3324
rect 290 3240 1978 3268
rect 93 3184 1024 3212
rect 93 3100 262 3184
rect 1052 3156 1216 3240
rect 2006 3212 2344 3296
rect 3134 3268 3298 3352
rect 4088 3324 4257 3630
rect 3326 3296 4257 3324
rect 2372 3240 4060 3268
rect 1244 3184 3106 3212
rect 290 3128 1978 3156
rect 93 3072 1024 3100
rect 93 2988 262 3072
rect 1052 3044 1216 3128
rect 2006 3100 2344 3184
rect 3134 3156 3298 3240
rect 4088 3212 4257 3296
rect 3326 3184 4257 3212
rect 2372 3128 4060 3156
rect 1244 3072 3106 3100
rect 290 3016 1978 3044
rect 93 2960 1024 2988
rect 93 2876 262 2960
rect 1052 2932 1216 3016
rect 2006 2988 2344 3072
rect 3134 3044 3298 3128
rect 4088 3100 4257 3184
rect 3326 3072 4257 3100
rect 2372 3016 4060 3044
rect 1244 2960 3106 2988
rect 290 2904 1978 2932
rect 93 2848 1024 2876
rect 93 2764 262 2848
rect 1052 2820 1216 2904
rect 2006 2876 2344 2960
rect 3134 2932 3298 3016
rect 4088 2988 4257 3072
rect 3326 2960 4257 2988
rect 2372 2904 4060 2932
rect 1244 2848 3106 2876
rect 290 2792 1978 2820
rect 93 2736 1024 2764
rect 93 2646 262 2736
rect 1052 2708 1216 2792
rect 2006 2764 2344 2848
rect 3134 2820 3298 2904
rect 4088 2876 4257 2960
rect 3326 2848 4257 2876
rect 2372 2792 4060 2820
rect 1244 2736 3106 2764
rect 290 2680 1978 2708
rect 93 2592 1024 2646
rect 93 2351 243 2592
rect 1052 2562 1216 2680
rect 2006 2646 2344 2736
rect 3134 2708 3298 2792
rect 4088 2764 4257 2848
rect 3326 2736 4257 2764
rect 2372 2680 4060 2708
rect 1244 2592 3106 2646
rect 271 2379 1996 2562
rect 2024 2351 2325 2592
rect 3134 2562 3298 2680
rect 4088 2646 4257 2736
rect 3326 2592 4257 2646
rect 2353 2379 4078 2562
rect 4106 2351 4257 2592
rect 93 2321 4257 2351
rect 93 2054 243 2321
rect 271 2084 1996 2293
rect 93 2000 1024 2054
rect 93 1910 262 2000
rect 1052 1966 1216 2084
rect 2024 2054 2325 2321
rect 2353 2084 4078 2293
rect 1244 2000 3106 2054
rect 290 1938 1978 1966
rect 93 1882 1024 1910
rect 93 1798 262 1882
rect 1052 1854 1216 1938
rect 2006 1910 2344 2000
rect 3134 1966 3298 2084
rect 4106 2054 4257 2321
rect 3326 2000 4257 2054
rect 2372 1938 4060 1966
rect 1244 1882 3106 1910
rect 290 1826 1978 1854
rect 93 1770 1024 1798
rect 93 1686 262 1770
rect 1052 1742 1216 1826
rect 2006 1798 2344 1882
rect 3134 1854 3298 1938
rect 4088 1910 4257 2000
rect 3326 1882 4257 1910
rect 2372 1826 4060 1854
rect 1244 1770 3106 1798
rect 290 1714 1978 1742
rect 93 1658 1024 1686
rect 93 1574 262 1658
rect 1052 1630 1216 1714
rect 2006 1686 2344 1770
rect 3134 1742 3298 1826
rect 4088 1798 4257 1882
rect 3326 1770 4257 1798
rect 2372 1714 4060 1742
rect 1244 1658 3106 1686
rect 290 1602 1978 1630
rect 93 1546 1024 1574
rect 93 1462 262 1546
rect 1052 1518 1216 1602
rect 2006 1574 2344 1658
rect 3134 1630 3298 1714
rect 4088 1686 4257 1770
rect 3326 1658 4257 1686
rect 2372 1602 4060 1630
rect 1244 1546 3106 1574
rect 290 1490 1978 1518
rect 93 1434 1024 1462
rect 93 1350 262 1434
rect 1052 1406 1216 1490
rect 2006 1462 2344 1546
rect 3134 1518 3298 1602
rect 4088 1574 4257 1658
rect 3326 1546 4257 1574
rect 2372 1490 4060 1518
rect 1244 1434 3106 1462
rect 290 1378 1978 1406
rect 93 1322 1024 1350
rect 93 1016 262 1322
rect 1052 1294 1216 1378
rect 2006 1350 2344 1434
rect 3134 1406 3298 1490
rect 4088 1462 4257 1546
rect 3326 1434 4257 1462
rect 2372 1378 4060 1406
rect 1244 1322 3106 1350
rect 290 1266 1978 1294
rect 1052 1232 1216 1266
rect 290 1106 1978 1232
rect 1052 1072 1216 1106
rect 290 1044 1978 1072
rect 93 988 1024 1016
rect 93 904 262 988
rect 1052 960 1216 1044
rect 2006 1016 2344 1322
rect 3134 1294 3298 1378
rect 4088 1350 4257 1434
rect 3326 1322 4257 1350
rect 2372 1266 4060 1294
rect 3134 1232 3298 1266
rect 2372 1106 4060 1232
rect 3134 1072 3298 1106
rect 2372 1044 4060 1072
rect 1244 988 3106 1016
rect 290 932 1978 960
rect 93 876 1024 904
rect 93 792 262 876
rect 1052 848 1216 932
rect 2006 904 2344 988
rect 3134 960 3298 1044
rect 4088 1016 4257 1322
rect 3326 988 4257 1016
rect 2372 932 4060 960
rect 1244 876 3106 904
rect 290 820 1978 848
rect 93 764 1024 792
rect 93 680 262 764
rect 1052 736 1216 820
rect 2006 792 2344 876
rect 3134 848 3298 932
rect 4088 904 4257 988
rect 3326 876 4257 904
rect 2372 820 4060 848
rect 1244 764 3106 792
rect 290 708 1978 736
rect 93 652 1024 680
rect 93 568 262 652
rect 1052 624 1216 708
rect 2006 680 2344 764
rect 3134 736 3298 820
rect 4088 792 4257 876
rect 3326 764 4257 792
rect 2372 708 4060 736
rect 1244 652 3106 680
rect 290 596 1978 624
rect 93 540 1024 568
rect 93 456 262 540
rect 1052 512 1216 596
rect 2006 568 2344 652
rect 3134 624 3298 708
rect 4088 680 4257 764
rect 3326 652 4257 680
rect 2372 596 4060 624
rect 1244 540 3106 568
rect 290 484 1978 512
rect 93 428 1024 456
rect 93 338 262 428
rect 1052 400 1216 484
rect 2006 456 2344 540
rect 3134 512 3298 596
rect 4088 568 4257 652
rect 3326 540 4257 568
rect 2372 484 4060 512
rect 1244 428 3106 456
rect 290 372 1978 400
rect 93 284 1024 338
rect 93 43 243 284
rect 1052 254 1216 372
rect 2006 338 2344 428
rect 3134 400 3298 484
rect 4088 456 4257 540
rect 3326 428 4257 456
rect 2372 372 4060 400
rect 1244 284 3106 338
rect 271 71 1996 254
rect 2024 43 2325 284
rect 3134 254 3298 372
rect 4088 338 4257 428
rect 3326 284 4257 338
rect 2353 71 4078 254
rect 4106 43 4257 284
rect 93 13 4257 43
<< obsm2 >>
rect 65 4392 4285 4644
rect 65 2562 169 4392
rect 198 4308 1024 4362
rect 198 4274 262 4308
rect 198 4246 1024 4274
rect 198 4162 262 4246
rect 1052 4218 1216 4392
rect 1244 4308 2070 4362
rect 2006 4274 2070 4308
rect 1244 4246 2070 4274
rect 290 4190 1978 4218
rect 198 4134 1024 4162
rect 198 4050 262 4134
rect 1052 4106 1216 4190
rect 2006 4162 2070 4246
rect 1244 4134 2070 4162
rect 290 4078 1978 4106
rect 198 4022 1024 4050
rect 198 3938 262 4022
rect 1052 3994 1216 4078
rect 2006 4050 2070 4134
rect 1244 4022 2070 4050
rect 290 3966 1978 3994
rect 198 3910 1024 3938
rect 198 3826 262 3910
rect 1052 3882 1216 3966
rect 2006 3938 2070 4022
rect 1244 3910 2070 3938
rect 290 3854 1978 3882
rect 198 3798 1024 3826
rect 198 3714 262 3798
rect 1052 3770 1216 3854
rect 2006 3826 2070 3910
rect 1244 3798 2070 3826
rect 290 3742 1978 3770
rect 198 3686 1024 3714
rect 198 3602 262 3686
rect 1052 3658 1216 3742
rect 2006 3714 2070 3798
rect 1244 3686 2070 3714
rect 290 3630 1978 3658
rect 198 3574 1024 3602
rect 198 3380 262 3574
rect 1052 3540 1216 3630
rect 2006 3602 2070 3686
rect 1244 3574 2070 3602
rect 290 3414 1978 3540
rect 198 3352 1024 3380
rect 198 3268 262 3352
rect 1052 3324 1216 3414
rect 2006 3380 2070 3574
rect 1244 3352 2070 3380
rect 290 3296 1978 3324
rect 198 3240 1024 3268
rect 198 3156 262 3240
rect 1052 3212 1216 3296
rect 2006 3268 2070 3352
rect 1244 3240 2070 3268
rect 290 3184 1978 3212
rect 198 3128 1024 3156
rect 198 3044 262 3128
rect 1052 3100 1216 3184
rect 2006 3156 2070 3240
rect 1244 3128 2070 3156
rect 290 3072 1978 3100
rect 198 3016 1024 3044
rect 198 2932 262 3016
rect 1052 2988 1216 3072
rect 2006 3044 2070 3128
rect 1244 3016 2070 3044
rect 290 2960 1978 2988
rect 198 2904 1024 2932
rect 198 2820 262 2904
rect 1052 2876 1216 2960
rect 2006 2932 2070 3016
rect 1244 2904 2070 2932
rect 290 2848 1978 2876
rect 198 2792 1024 2820
rect 198 2708 262 2792
rect 1052 2764 1216 2848
rect 2006 2820 2070 2904
rect 1244 2792 2070 2820
rect 290 2736 1978 2764
rect 198 2680 1024 2708
rect 198 2646 262 2680
rect 198 2592 1024 2646
rect 1052 2562 1216 2736
rect 2006 2708 2070 2792
rect 1244 2680 2070 2708
rect 2006 2646 2070 2680
rect 1244 2592 2070 2646
rect 2098 2562 2251 4392
rect 2280 4308 3106 4362
rect 2280 4274 2344 4308
rect 2280 4246 3106 4274
rect 2280 4162 2344 4246
rect 3134 4218 3298 4392
rect 3326 4308 4152 4362
rect 4088 4274 4152 4308
rect 3326 4246 4152 4274
rect 2372 4190 4060 4218
rect 2280 4134 3106 4162
rect 2280 4050 2344 4134
rect 3134 4106 3298 4190
rect 4088 4162 4152 4246
rect 3326 4134 4152 4162
rect 2372 4078 4060 4106
rect 2280 4022 3106 4050
rect 2280 3938 2344 4022
rect 3134 3994 3298 4078
rect 4088 4050 4152 4134
rect 3326 4022 4152 4050
rect 2372 3966 4060 3994
rect 2280 3910 3106 3938
rect 2280 3826 2344 3910
rect 3134 3882 3298 3966
rect 4088 3938 4152 4022
rect 3326 3910 4152 3938
rect 2372 3854 4060 3882
rect 2280 3798 3106 3826
rect 2280 3714 2344 3798
rect 3134 3770 3298 3854
rect 4088 3826 4152 3910
rect 3326 3798 4152 3826
rect 2372 3742 4060 3770
rect 2280 3686 3106 3714
rect 2280 3602 2344 3686
rect 3134 3658 3298 3742
rect 4088 3714 4152 3798
rect 3326 3686 4152 3714
rect 2372 3630 4060 3658
rect 2280 3574 3106 3602
rect 2280 3380 2344 3574
rect 3134 3540 3298 3630
rect 4088 3602 4152 3686
rect 3326 3574 4152 3602
rect 2372 3414 4060 3540
rect 2280 3352 3106 3380
rect 2280 3268 2344 3352
rect 3134 3324 3298 3414
rect 4088 3380 4152 3574
rect 3326 3352 4152 3380
rect 2372 3296 4060 3324
rect 2280 3240 3106 3268
rect 2280 3156 2344 3240
rect 3134 3212 3298 3296
rect 4088 3268 4152 3352
rect 3326 3240 4152 3268
rect 2372 3184 4060 3212
rect 2280 3128 3106 3156
rect 2280 3044 2344 3128
rect 3134 3100 3298 3184
rect 4088 3156 4152 3240
rect 3326 3128 4152 3156
rect 2372 3072 4060 3100
rect 2280 3016 3106 3044
rect 2280 2932 2344 3016
rect 3134 2988 3298 3072
rect 4088 3044 4152 3128
rect 3326 3016 4152 3044
rect 2372 2960 4060 2988
rect 2280 2904 3106 2932
rect 2280 2820 2344 2904
rect 3134 2876 3298 2960
rect 4088 2932 4152 3016
rect 3326 2904 4152 2932
rect 2372 2848 4060 2876
rect 2280 2792 3106 2820
rect 2280 2708 2344 2792
rect 3134 2764 3298 2848
rect 4088 2820 4152 2904
rect 3326 2792 4152 2820
rect 2372 2736 4060 2764
rect 2280 2680 3106 2708
rect 2280 2646 2344 2680
rect 2280 2592 3106 2646
rect 3134 2562 3298 2736
rect 4088 2708 4152 2792
rect 3326 2680 4152 2708
rect 4088 2646 4152 2680
rect 3326 2592 4152 2646
rect 4180 2562 4285 4392
rect 65 2084 4285 2562
rect 65 254 169 2084
rect 198 2000 1024 2054
rect 198 1966 262 2000
rect 198 1938 1024 1966
rect 198 1854 262 1938
rect 1052 1910 1216 2084
rect 1244 2000 2070 2054
rect 2006 1966 2070 2000
rect 1244 1938 2070 1966
rect 290 1882 1978 1910
rect 198 1826 1024 1854
rect 198 1742 262 1826
rect 1052 1798 1216 1882
rect 2006 1854 2070 1938
rect 1244 1826 2070 1854
rect 290 1770 1978 1798
rect 198 1714 1024 1742
rect 198 1630 262 1714
rect 1052 1686 1216 1770
rect 2006 1742 2070 1826
rect 1244 1714 2070 1742
rect 290 1658 1978 1686
rect 198 1602 1024 1630
rect 198 1518 262 1602
rect 1052 1574 1216 1658
rect 2006 1630 2070 1714
rect 1244 1602 2070 1630
rect 290 1546 1978 1574
rect 198 1490 1024 1518
rect 198 1406 262 1490
rect 1052 1462 1216 1546
rect 2006 1518 2070 1602
rect 1244 1490 2070 1518
rect 290 1434 1978 1462
rect 198 1378 1024 1406
rect 198 1294 262 1378
rect 1052 1350 1216 1434
rect 2006 1406 2070 1490
rect 1244 1378 2070 1406
rect 290 1322 1978 1350
rect 198 1266 1024 1294
rect 198 1072 262 1266
rect 1052 1232 1216 1322
rect 2006 1294 2070 1378
rect 1244 1266 2070 1294
rect 290 1106 1978 1232
rect 198 1044 1024 1072
rect 198 960 262 1044
rect 1052 1016 1216 1106
rect 2006 1072 2070 1266
rect 1244 1044 2070 1072
rect 290 988 1978 1016
rect 198 932 1024 960
rect 198 848 262 932
rect 1052 904 1216 988
rect 2006 960 2070 1044
rect 1244 932 2070 960
rect 290 876 1978 904
rect 198 820 1024 848
rect 198 736 262 820
rect 1052 792 1216 876
rect 2006 848 2070 932
rect 1244 820 2070 848
rect 290 764 1978 792
rect 198 708 1024 736
rect 198 624 262 708
rect 1052 680 1216 764
rect 2006 736 2070 820
rect 1244 708 2070 736
rect 290 652 1978 680
rect 198 596 1024 624
rect 198 512 262 596
rect 1052 568 1216 652
rect 2006 624 2070 708
rect 1244 596 2070 624
rect 290 540 1978 568
rect 198 484 1024 512
rect 198 400 262 484
rect 1052 456 1216 540
rect 2006 512 2070 596
rect 1244 484 2070 512
rect 290 428 1978 456
rect 198 372 1024 400
rect 198 338 262 372
rect 198 284 1024 338
rect 1052 254 1216 428
rect 2006 400 2070 484
rect 1244 372 2070 400
rect 2006 338 2070 372
rect 1244 284 2070 338
rect 2098 254 2251 2084
rect 2280 2000 3106 2054
rect 2280 1966 2344 2000
rect 2280 1938 3106 1966
rect 2280 1854 2344 1938
rect 3134 1910 3298 2084
rect 3326 2000 4152 2054
rect 4088 1966 4152 2000
rect 3326 1938 4152 1966
rect 2372 1882 4060 1910
rect 2280 1826 3106 1854
rect 2280 1742 2344 1826
rect 3134 1798 3298 1882
rect 4088 1854 4152 1938
rect 3326 1826 4152 1854
rect 2372 1770 4060 1798
rect 2280 1714 3106 1742
rect 2280 1630 2344 1714
rect 3134 1686 3298 1770
rect 4088 1742 4152 1826
rect 3326 1714 4152 1742
rect 2372 1658 4060 1686
rect 2280 1602 3106 1630
rect 2280 1518 2344 1602
rect 3134 1574 3298 1658
rect 4088 1630 4152 1714
rect 3326 1602 4152 1630
rect 2372 1546 4060 1574
rect 2280 1490 3106 1518
rect 2280 1406 2344 1490
rect 3134 1462 3298 1546
rect 4088 1518 4152 1602
rect 3326 1490 4152 1518
rect 2372 1434 4060 1462
rect 2280 1378 3106 1406
rect 2280 1294 2344 1378
rect 3134 1350 3298 1434
rect 4088 1406 4152 1490
rect 3326 1378 4152 1406
rect 2372 1322 4060 1350
rect 2280 1266 3106 1294
rect 2280 1072 2344 1266
rect 3134 1232 3298 1322
rect 4088 1294 4152 1378
rect 3326 1266 4152 1294
rect 2372 1106 4060 1232
rect 2280 1044 3106 1072
rect 2280 960 2344 1044
rect 3134 1016 3298 1106
rect 4088 1072 4152 1266
rect 3326 1044 4152 1072
rect 2372 988 4060 1016
rect 2280 932 3106 960
rect 2280 848 2344 932
rect 3134 904 3298 988
rect 4088 960 4152 1044
rect 3326 932 4152 960
rect 2372 876 4060 904
rect 2280 820 3106 848
rect 2280 736 2344 820
rect 3134 792 3298 876
rect 4088 848 4152 932
rect 3326 820 4152 848
rect 2372 764 4060 792
rect 2280 708 3106 736
rect 2280 624 2344 708
rect 3134 680 3298 764
rect 4088 736 4152 820
rect 3326 708 4152 736
rect 2372 652 4060 680
rect 2280 596 3106 624
rect 2280 512 2344 596
rect 3134 568 3298 652
rect 4088 624 4152 708
rect 3326 596 4152 624
rect 2372 540 4060 568
rect 2280 484 3106 512
rect 2280 400 2344 484
rect 3134 456 3298 540
rect 4088 512 4152 596
rect 3326 484 4152 512
rect 2372 428 4060 456
rect 2280 372 3106 400
rect 2280 338 2344 372
rect 2280 284 3106 338
rect 3134 254 3298 428
rect 4088 400 4152 484
rect 3326 372 4152 400
rect 4088 338 4152 372
rect 3326 284 4152 338
rect 4180 254 4285 2084
rect 65 28 4285 254
<< obsm3 >>
rect 60 28 126 4644
rect 193 4527 2075 4593
rect 193 4347 259 4527
rect 319 4407 1949 4467
rect 193 4287 1041 4347
rect 193 4107 259 4287
rect 1101 4227 1167 4407
rect 2009 4347 2075 4527
rect 1227 4287 2075 4347
rect 319 4167 1949 4227
rect 193 4047 1041 4107
rect 193 3867 259 4047
rect 1101 3987 1167 4167
rect 2009 4107 2075 4287
rect 1227 4047 2075 4107
rect 319 3927 1949 3987
rect 193 3807 1041 3867
rect 193 3627 259 3807
rect 1101 3747 1167 3927
rect 2009 3867 2075 4047
rect 1227 3807 2075 3867
rect 319 3687 1949 3747
rect 193 3567 1041 3627
rect 193 3381 259 3567
rect 1101 3507 1167 3687
rect 2009 3627 2075 3807
rect 1227 3567 2075 3627
rect 319 3441 1949 3507
rect 193 3321 1041 3381
rect 193 3141 259 3321
rect 1101 3261 1167 3441
rect 2009 3381 2075 3567
rect 1227 3321 2075 3381
rect 319 3201 1949 3261
rect 193 3081 1041 3141
rect 193 2901 259 3081
rect 1101 3021 1167 3201
rect 2009 3141 2075 3321
rect 1227 3081 2075 3141
rect 319 2961 1949 3021
rect 193 2841 1041 2901
rect 193 2661 259 2841
rect 1101 2781 1167 2961
rect 2009 2901 2075 3081
rect 1227 2841 2075 2901
rect 319 2721 1949 2781
rect 193 2601 1041 2661
rect 193 2421 259 2601
rect 1101 2541 1167 2721
rect 2009 2661 2075 2841
rect 1227 2601 2075 2661
rect 319 2481 1949 2541
rect 2009 2421 2075 2601
rect 193 2355 2075 2421
rect 193 2219 2075 2285
rect 193 2039 259 2219
rect 319 2099 1949 2159
rect 193 1979 1041 2039
rect 193 1799 259 1979
rect 1101 1919 1167 2099
rect 2009 2039 2075 2219
rect 1227 1979 2075 2039
rect 319 1859 1949 1919
rect 193 1739 1041 1799
rect 193 1559 259 1739
rect 1101 1679 1167 1859
rect 2009 1799 2075 1979
rect 1227 1739 2075 1799
rect 319 1619 1949 1679
rect 193 1499 1041 1559
rect 193 1319 259 1499
rect 1101 1439 1167 1619
rect 2009 1559 2075 1739
rect 1227 1499 2075 1559
rect 319 1379 1949 1439
rect 193 1259 1041 1319
rect 193 1073 259 1259
rect 1101 1199 1167 1379
rect 2009 1319 2075 1499
rect 1227 1259 2075 1319
rect 319 1133 1949 1199
rect 193 1013 1041 1073
rect 193 833 259 1013
rect 1101 953 1167 1133
rect 2009 1073 2075 1259
rect 1227 1013 2075 1073
rect 319 893 1949 953
rect 193 773 1041 833
rect 193 593 259 773
rect 1101 713 1167 893
rect 2009 833 2075 1013
rect 1227 773 2075 833
rect 319 653 1949 713
rect 193 533 1041 593
rect 193 353 259 533
rect 1101 473 1167 653
rect 2009 593 2075 773
rect 1227 533 2075 593
rect 319 413 1949 473
rect 193 293 1041 353
rect 193 113 259 293
rect 1101 233 1167 413
rect 2009 353 2075 533
rect 1227 293 2075 353
rect 319 173 1949 233
rect 2009 113 2075 293
rect 193 47 2075 113
rect 2142 28 2208 4644
rect 2275 4527 4157 4593
rect 2275 4347 2341 4527
rect 2401 4407 4031 4467
rect 2275 4287 3123 4347
rect 2275 4107 2341 4287
rect 3183 4227 3249 4407
rect 4091 4347 4157 4527
rect 3309 4287 4157 4347
rect 2401 4167 4031 4227
rect 2275 4047 3123 4107
rect 2275 3867 2341 4047
rect 3183 3987 3249 4167
rect 4091 4107 4157 4287
rect 3309 4047 4157 4107
rect 2401 3927 4031 3987
rect 2275 3807 3123 3867
rect 2275 3627 2341 3807
rect 3183 3747 3249 3927
rect 4091 3867 4157 4047
rect 3309 3807 4157 3867
rect 2401 3687 4031 3747
rect 2275 3567 3123 3627
rect 2275 3381 2341 3567
rect 3183 3507 3249 3687
rect 4091 3627 4157 3807
rect 3309 3567 4157 3627
rect 2401 3441 4031 3507
rect 2275 3321 3123 3381
rect 2275 3141 2341 3321
rect 3183 3261 3249 3441
rect 4091 3381 4157 3567
rect 3309 3321 4157 3381
rect 2401 3201 4031 3261
rect 2275 3081 3123 3141
rect 2275 2901 2341 3081
rect 3183 3021 3249 3201
rect 4091 3141 4157 3321
rect 3309 3081 4157 3141
rect 2401 2961 4031 3021
rect 2275 2841 3123 2901
rect 2275 2661 2341 2841
rect 3183 2781 3249 2961
rect 4091 2901 4157 3081
rect 3309 2841 4157 2901
rect 2401 2721 4031 2781
rect 2275 2601 3123 2661
rect 2275 2421 2341 2601
rect 3183 2541 3249 2721
rect 4091 2661 4157 2841
rect 3309 2601 4157 2661
rect 2401 2481 4031 2541
rect 4091 2421 4157 2601
rect 2275 2355 4157 2421
rect 2275 2219 4157 2285
rect 2275 2039 2341 2219
rect 2401 2099 4031 2159
rect 2275 1979 3123 2039
rect 2275 1799 2341 1979
rect 3183 1919 3249 2099
rect 4091 2039 4157 2219
rect 3309 1979 4157 2039
rect 2401 1859 4031 1919
rect 2275 1739 3123 1799
rect 2275 1559 2341 1739
rect 3183 1679 3249 1859
rect 4091 1799 4157 1979
rect 3309 1739 4157 1799
rect 2401 1619 4031 1679
rect 2275 1499 3123 1559
rect 2275 1319 2341 1499
rect 3183 1439 3249 1619
rect 4091 1559 4157 1739
rect 3309 1499 4157 1559
rect 2401 1379 4031 1439
rect 2275 1259 3123 1319
rect 2275 1073 2341 1259
rect 3183 1199 3249 1379
rect 4091 1319 4157 1499
rect 3309 1259 4157 1319
rect 2401 1133 4031 1199
rect 2275 1013 3123 1073
rect 2275 833 2341 1013
rect 3183 953 3249 1133
rect 4091 1073 4157 1259
rect 3309 1013 4157 1073
rect 2401 893 4031 953
rect 2275 773 3123 833
rect 2275 593 2341 773
rect 3183 713 3249 893
rect 4091 833 4157 1013
rect 3309 773 4157 833
rect 2401 653 4031 713
rect 2275 533 3123 593
rect 2275 353 2341 533
rect 3183 473 3249 653
rect 4091 593 4157 773
rect 3309 533 4157 593
rect 2401 413 4031 473
rect 2275 293 3123 353
rect 2275 113 2341 293
rect 3183 233 3249 413
rect 4091 353 4157 533
rect 3309 293 4157 353
rect 2401 173 4031 233
rect 4091 113 4157 293
rect 2275 47 4157 113
rect 4224 28 4290 4644
<< metal4 >>
rect 60 28 126 4644
rect 193 4587 2009 4593
rect 193 4527 2075 4587
rect 193 2421 259 4527
rect 319 3507 379 4467
rect 439 3567 499 4527
rect 559 3507 619 4467
rect 679 3567 739 4527
rect 799 3507 859 4467
rect 919 3567 1002 4527
rect 1062 3507 1167 4467
rect 1227 3567 1349 4527
rect 1409 3507 1469 4467
rect 1529 3567 1589 4527
rect 1649 3507 1709 4467
rect 1769 3567 1829 4527
rect 1889 3507 1949 4467
rect 319 3441 1949 3507
rect 319 2481 379 3441
rect 439 2421 499 3381
rect 559 2481 619 3441
rect 679 2421 739 3381
rect 799 2481 859 3441
rect 919 2421 1002 3381
rect 1062 2481 1167 3441
rect 1227 2421 1349 3381
rect 1409 2481 1469 3441
rect 1529 2421 1589 3381
rect 1649 2481 1709 3441
rect 1769 2421 1829 3381
rect 1889 2481 1949 3441
rect 2009 2421 2075 4527
rect 193 2355 2075 2421
rect 193 2279 2009 2285
rect 193 2219 2075 2279
rect 193 113 259 2219
rect 319 1199 379 2159
rect 439 1259 499 2219
rect 559 1199 619 2159
rect 679 1259 739 2219
rect 799 1199 859 2159
rect 919 1259 1002 2219
rect 1062 1199 1167 2159
rect 1227 1259 1349 2219
rect 1409 1199 1469 2159
rect 1529 1259 1589 2219
rect 1649 1199 1709 2159
rect 1769 1259 1829 2219
rect 1889 1199 1949 2159
rect 319 1133 1949 1199
rect 319 173 379 1133
rect 439 113 499 1073
rect 559 173 619 1133
rect 679 113 739 1073
rect 799 173 859 1133
rect 919 113 1002 1073
rect 1062 173 1167 1133
rect 1227 113 1349 1073
rect 1409 173 1469 1133
rect 1529 113 1589 1073
rect 1649 173 1709 1133
rect 1769 113 1829 1073
rect 1889 173 1949 1133
rect 2009 113 2075 2219
rect 193 47 2075 113
rect 2142 28 2208 4644
rect 2275 4587 4091 4593
rect 2275 4527 4157 4587
rect 2275 2421 2341 4527
rect 2401 3507 2461 4467
rect 2521 3567 2581 4527
rect 2641 3507 2701 4467
rect 2761 3567 2821 4527
rect 2881 3507 2941 4467
rect 3001 3567 3084 4527
rect 3144 3507 3249 4467
rect 3309 3567 3431 4527
rect 3491 3507 3551 4467
rect 3611 3567 3671 4527
rect 3731 3507 3791 4467
rect 3851 3567 3911 4527
rect 3971 3507 4031 4467
rect 2401 3441 4031 3507
rect 2401 2481 2461 3441
rect 2521 2421 2581 3381
rect 2641 2481 2701 3441
rect 2761 2421 2821 3381
rect 2881 2481 2941 3441
rect 3001 2421 3084 3381
rect 3144 2481 3249 3441
rect 3309 2421 3431 3381
rect 3491 2481 3551 3441
rect 3611 2421 3671 3381
rect 3731 2481 3791 3441
rect 3851 2421 3911 3381
rect 3971 2481 4031 3441
rect 4091 2421 4157 4527
rect 2275 2355 4157 2421
rect 2275 2279 4091 2285
rect 2275 2219 4157 2279
rect 2275 113 2341 2219
rect 2401 1199 2461 2159
rect 2521 1259 2581 2219
rect 2641 1199 2701 2159
rect 2761 1259 2821 2219
rect 2881 1199 2941 2159
rect 3001 1259 3084 2219
rect 3144 1199 3249 2159
rect 3309 1259 3431 2219
rect 3491 1199 3551 2159
rect 3611 1259 3671 2219
rect 3731 1199 3791 2159
rect 3851 1259 3911 2219
rect 3971 1199 4031 2159
rect 2401 1133 4031 1199
rect 2401 173 2461 1133
rect 2521 113 2581 1073
rect 2641 173 2701 1133
rect 2761 113 2821 1073
rect 2881 173 2941 1133
rect 3001 113 3084 1073
rect 3144 173 3249 1133
rect 3309 113 3431 1073
rect 3491 173 3551 1133
rect 3611 113 3671 1073
rect 3731 173 3791 1133
rect 3851 113 3911 1073
rect 3971 173 4031 1133
rect 4091 113 4157 2219
rect 2275 47 4157 113
rect 4224 28 4290 4644
<< metal5 >>
rect 0 13 4350 4659
<< labels >>
rlabel metal4 s 4224 28 4290 4644 6 C0
port 1 nsew
rlabel metal4 s 3971 3507 4031 4467 6 C0
port 1 nsew
rlabel metal4 s 3971 2481 4031 3441 6 C0
port 1 nsew
rlabel metal4 s 3971 1199 4031 2159 6 C0
port 1 nsew
rlabel metal4 s 3971 173 4031 1133 6 C0
port 1 nsew
rlabel metal4 s 3731 3507 3791 4467 6 C0
port 1 nsew
rlabel metal4 s 3731 2481 3791 3441 6 C0
port 1 nsew
rlabel metal4 s 3731 1199 3791 2159 6 C0
port 1 nsew
rlabel metal4 s 3731 173 3791 1133 6 C0
port 1 nsew
rlabel metal4 s 3491 3507 3551 4467 6 C0
port 1 nsew
rlabel metal4 s 3491 2481 3551 3441 6 C0
port 1 nsew
rlabel metal4 s 3491 1199 3551 2159 6 C0
port 1 nsew
rlabel metal4 s 3491 173 3551 1133 6 C0
port 1 nsew
rlabel metal4 s 3144 3507 3249 4467 6 C0
port 1 nsew
rlabel metal4 s 3144 2481 3249 3441 6 C0
port 1 nsew
rlabel metal4 s 3144 1199 3249 2159 6 C0
port 1 nsew
rlabel metal4 s 3144 173 3249 1133 6 C0
port 1 nsew
rlabel metal4 s 2881 3507 2941 4467 6 C0
port 1 nsew
rlabel metal4 s 2881 2481 2941 3441 6 C0
port 1 nsew
rlabel metal4 s 2881 1199 2941 2159 6 C0
port 1 nsew
rlabel metal4 s 2881 173 2941 1133 6 C0
port 1 nsew
rlabel metal4 s 2641 3507 2701 4467 6 C0
port 1 nsew
rlabel metal4 s 2641 2481 2701 3441 6 C0
port 1 nsew
rlabel metal4 s 2641 1199 2701 2159 6 C0
port 1 nsew
rlabel metal4 s 2641 173 2701 1133 6 C0
port 1 nsew
rlabel metal4 s 2401 3507 2461 4467 6 C0
port 1 nsew
rlabel metal4 s 2401 3441 4031 3507 6 C0
port 1 nsew
rlabel metal4 s 2401 2481 2461 3441 6 C0
port 1 nsew
rlabel metal4 s 2401 1199 2461 2159 6 C0
port 1 nsew
rlabel metal4 s 2401 1133 4031 1199 6 C0
port 1 nsew
rlabel metal4 s 2401 173 2461 1133 6 C0
port 1 nsew
rlabel metal4 s 2142 28 2208 4644 6 C0
port 1 nsew
rlabel metal4 s 1889 3507 1949 4467 6 C0
port 1 nsew
rlabel metal4 s 1889 2481 1949 3441 6 C0
port 1 nsew
rlabel metal4 s 1889 1199 1949 2159 6 C0
port 1 nsew
rlabel metal4 s 1889 173 1949 1133 6 C0
port 1 nsew
rlabel metal4 s 1649 3507 1709 4467 6 C0
port 1 nsew
rlabel metal4 s 1649 2481 1709 3441 6 C0
port 1 nsew
rlabel metal4 s 1649 1199 1709 2159 6 C0
port 1 nsew
rlabel metal4 s 1649 173 1709 1133 6 C0
port 1 nsew
rlabel metal4 s 1409 3507 1469 4467 6 C0
port 1 nsew
rlabel metal4 s 1409 2481 1469 3441 6 C0
port 1 nsew
rlabel metal4 s 1409 1199 1469 2159 6 C0
port 1 nsew
rlabel metal4 s 1409 173 1469 1133 6 C0
port 1 nsew
rlabel metal4 s 1062 3507 1167 4467 6 C0
port 1 nsew
rlabel metal4 s 1062 2481 1167 3441 6 C0
port 1 nsew
rlabel metal4 s 1062 1199 1167 2159 6 C0
port 1 nsew
rlabel metal4 s 1062 173 1167 1133 6 C0
port 1 nsew
rlabel metal4 s 799 3507 859 4467 6 C0
port 1 nsew
rlabel metal4 s 799 2481 859 3441 6 C0
port 1 nsew
rlabel metal4 s 799 1199 859 2159 6 C0
port 1 nsew
rlabel metal4 s 799 173 859 1133 6 C0
port 1 nsew
rlabel metal4 s 559 3507 619 4467 6 C0
port 1 nsew
rlabel metal4 s 559 2481 619 3441 6 C0
port 1 nsew
rlabel metal4 s 559 1199 619 2159 6 C0
port 1 nsew
rlabel metal4 s 559 173 619 1133 6 C0
port 1 nsew
rlabel metal4 s 319 3507 379 4467 6 C0
port 1 nsew
rlabel metal4 s 319 3441 1949 3507 6 C0
port 1 nsew
rlabel metal4 s 319 2481 379 3441 6 C0
port 1 nsew
rlabel metal4 s 319 1199 379 2159 6 C0
port 1 nsew
rlabel metal4 s 319 1133 1949 1199 6 C0
port 1 nsew
rlabel metal4 s 319 173 379 1133 6 C0
port 1 nsew
rlabel metal4 s 60 28 126 4644 6 C0
port 1 nsew
rlabel metal5 s 0 13 4350 4659 6 M5
port 2 nsew
rlabel metal4 s 4091 2421 4157 4527 6 SUB
port 3 nsew
rlabel metal4 s 4091 113 4157 2219 6 SUB
port 3 nsew
rlabel metal4 s 3851 3567 3911 4527 6 SUB
port 3 nsew
rlabel metal4 s 3851 2421 3911 3381 6 SUB
port 3 nsew
rlabel metal4 s 3851 1259 3911 2219 6 SUB
port 3 nsew
rlabel metal4 s 3851 113 3911 1073 6 SUB
port 3 nsew
rlabel metal4 s 3611 3567 3671 4527 6 SUB
port 3 nsew
rlabel metal4 s 3611 2421 3671 3381 6 SUB
port 3 nsew
rlabel metal4 s 3611 1259 3671 2219 6 SUB
port 3 nsew
rlabel metal4 s 3611 113 3671 1073 6 SUB
port 3 nsew
rlabel metal4 s 3309 3567 3431 4527 6 SUB
port 3 nsew
rlabel metal4 s 3309 2421 3431 3381 6 SUB
port 3 nsew
rlabel metal4 s 3309 1259 3431 2219 6 SUB
port 3 nsew
rlabel metal4 s 3309 113 3431 1073 6 SUB
port 3 nsew
rlabel metal4 s 3001 3567 3084 4527 6 SUB
port 3 nsew
rlabel metal4 s 3001 2421 3084 3381 6 SUB
port 3 nsew
rlabel metal4 s 3001 1259 3084 2219 6 SUB
port 3 nsew
rlabel metal4 s 3001 113 3084 1073 6 SUB
port 3 nsew
rlabel metal4 s 2761 3567 2821 4527 6 SUB
port 3 nsew
rlabel metal4 s 2761 2421 2821 3381 6 SUB
port 3 nsew
rlabel metal4 s 2761 1259 2821 2219 6 SUB
port 3 nsew
rlabel metal4 s 2761 113 2821 1073 6 SUB
port 3 nsew
rlabel metal4 s 2521 3567 2581 4527 6 SUB
port 3 nsew
rlabel metal4 s 2521 2421 2581 3381 6 SUB
port 3 nsew
rlabel metal4 s 2521 1259 2581 2219 6 SUB
port 3 nsew
rlabel metal4 s 2521 113 2581 1073 6 SUB
port 3 nsew
rlabel metal4 s 2275 4587 4091 4593 6 SUB
port 3 nsew
rlabel metal4 s 2275 4527 4157 4587 6 SUB
port 3 nsew
rlabel metal4 s 2275 2421 2341 4527 6 SUB
port 3 nsew
rlabel metal4 s 2275 2355 4157 2421 6 SUB
port 3 nsew
rlabel metal4 s 2275 2279 4091 2285 6 SUB
port 3 nsew
rlabel metal4 s 2275 2219 4157 2279 6 SUB
port 3 nsew
rlabel metal4 s 2275 113 2341 2219 6 SUB
port 3 nsew
rlabel metal4 s 2275 47 4157 113 6 SUB
port 3 nsew
rlabel metal4 s 2009 2421 2075 4527 6 SUB
port 3 nsew
rlabel metal4 s 2009 113 2075 2219 6 SUB
port 3 nsew
rlabel metal4 s 1769 3567 1829 4527 6 SUB
port 3 nsew
rlabel metal4 s 1769 2421 1829 3381 6 SUB
port 3 nsew
rlabel metal4 s 1769 1259 1829 2219 6 SUB
port 3 nsew
rlabel metal4 s 1769 113 1829 1073 6 SUB
port 3 nsew
rlabel metal4 s 1529 3567 1589 4527 6 SUB
port 3 nsew
rlabel metal4 s 1529 2421 1589 3381 6 SUB
port 3 nsew
rlabel metal4 s 1529 1259 1589 2219 6 SUB
port 3 nsew
rlabel metal4 s 1529 113 1589 1073 6 SUB
port 3 nsew
rlabel metal4 s 1227 3567 1349 4527 6 SUB
port 3 nsew
rlabel metal4 s 1227 2421 1349 3381 6 SUB
port 3 nsew
rlabel metal4 s 1227 1259 1349 2219 6 SUB
port 3 nsew
rlabel metal4 s 1227 113 1349 1073 6 SUB
port 3 nsew
rlabel metal4 s 919 3567 1002 4527 6 SUB
port 3 nsew
rlabel metal4 s 919 2421 1002 3381 6 SUB
port 3 nsew
rlabel metal4 s 919 1259 1002 2219 6 SUB
port 3 nsew
rlabel metal4 s 919 113 1002 1073 6 SUB
port 3 nsew
rlabel metal4 s 679 3567 739 4527 6 SUB
port 3 nsew
rlabel metal4 s 679 2421 739 3381 6 SUB
port 3 nsew
rlabel metal4 s 679 1259 739 2219 6 SUB
port 3 nsew
rlabel metal4 s 679 113 739 1073 6 SUB
port 3 nsew
rlabel metal4 s 439 3567 499 4527 6 SUB
port 3 nsew
rlabel metal4 s 439 2421 499 3381 6 SUB
port 3 nsew
rlabel metal4 s 439 1259 499 2219 6 SUB
port 3 nsew
rlabel metal4 s 439 113 499 1073 6 SUB
port 3 nsew
rlabel metal4 s 193 4587 2009 4593 6 SUB
port 3 nsew
rlabel metal4 s 193 4527 2075 4587 6 SUB
port 3 nsew
rlabel metal4 s 193 2421 259 4527 6 SUB
port 3 nsew
rlabel metal4 s 193 2355 2075 2421 6 SUB
port 3 nsew
rlabel metal4 s 193 2279 2009 2285 6 SUB
port 3 nsew
rlabel metal4 s 193 2219 2075 2279 6 SUB
port 3 nsew
rlabel metal4 s 193 113 259 2219 6 SUB
port 3 nsew
rlabel metal4 s 193 47 2075 113 6 SUB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 -5 4350 4659
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 847346
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 846912
<< end >>
