magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect 4658 -327 6685 -248
rect 7568 -327 7874 -277
rect 4658 -980 7874 -327
rect 4964 -1029 6129 -980
rect 6021 -1146 6129 -1029
rect 6530 -1351 7874 -980
rect 6530 -1393 7568 -1351
<< pwell >>
rect 6413 -1509 7747 -1479
rect 6305 -2122 7747 -1509
rect 6413 -2131 7747 -2122
<< mvnmos >>
rect 6492 -2105 6612 -1505
rect 6668 -2105 6788 -1505
rect 6844 -2105 6964 -1505
rect 7020 -2105 7140 -1505
rect 7196 -2105 7316 -1505
rect 7372 -2105 7492 -1505
rect 7548 -2105 7668 -1505
<< mvpmos >>
rect 4777 -914 4877 -314
rect 4933 -914 5033 -314
rect 5089 -914 5189 -314
rect 5369 -914 5469 -314
rect 5525 -914 5625 -314
rect 5681 -914 5781 -314
rect 5837 -914 5937 -314
rect 6117 -914 6217 -314
rect 6273 -914 6373 -314
rect 6649 -477 7449 -393
rect 7724 -596 7808 -396
rect 6649 -691 7449 -607
rect 6649 -885 7449 -801
rect 7724 -852 7808 -652
rect 6649 -1111 7449 -1027
rect 7724 -1232 7808 -1032
rect 6649 -1327 7449 -1243
<< mvndiff >>
rect 6439 -1583 6492 -1505
rect 6439 -1617 6447 -1583
rect 6481 -1617 6492 -1583
rect 6439 -1651 6492 -1617
rect 6439 -1685 6447 -1651
rect 6481 -1685 6492 -1651
rect 6439 -1719 6492 -1685
rect 6439 -1753 6447 -1719
rect 6481 -1753 6492 -1719
rect 6439 -1787 6492 -1753
rect 6439 -1821 6447 -1787
rect 6481 -1821 6492 -1787
rect 6439 -1855 6492 -1821
rect 6439 -1889 6447 -1855
rect 6481 -1889 6492 -1855
rect 6439 -1923 6492 -1889
rect 6439 -1957 6447 -1923
rect 6481 -1957 6492 -1923
rect 6439 -1991 6492 -1957
rect 6439 -2025 6447 -1991
rect 6481 -2025 6492 -1991
rect 6439 -2059 6492 -2025
rect 6439 -2093 6447 -2059
rect 6481 -2093 6492 -2059
rect 6439 -2105 6492 -2093
rect 6612 -1583 6668 -1505
rect 6612 -1617 6623 -1583
rect 6657 -1617 6668 -1583
rect 6612 -1651 6668 -1617
rect 6612 -1685 6623 -1651
rect 6657 -1685 6668 -1651
rect 6612 -1719 6668 -1685
rect 6612 -1753 6623 -1719
rect 6657 -1753 6668 -1719
rect 6612 -1787 6668 -1753
rect 6612 -1821 6623 -1787
rect 6657 -1821 6668 -1787
rect 6612 -1855 6668 -1821
rect 6612 -1889 6623 -1855
rect 6657 -1889 6668 -1855
rect 6612 -1923 6668 -1889
rect 6612 -1957 6623 -1923
rect 6657 -1957 6668 -1923
rect 6612 -1991 6668 -1957
rect 6612 -2025 6623 -1991
rect 6657 -2025 6668 -1991
rect 6612 -2059 6668 -2025
rect 6612 -2093 6623 -2059
rect 6657 -2093 6668 -2059
rect 6612 -2105 6668 -2093
rect 6788 -1583 6844 -1505
rect 6788 -1617 6799 -1583
rect 6833 -1617 6844 -1583
rect 6788 -1651 6844 -1617
rect 6788 -1685 6799 -1651
rect 6833 -1685 6844 -1651
rect 6788 -1719 6844 -1685
rect 6788 -1753 6799 -1719
rect 6833 -1753 6844 -1719
rect 6788 -1787 6844 -1753
rect 6788 -1821 6799 -1787
rect 6833 -1821 6844 -1787
rect 6788 -1855 6844 -1821
rect 6788 -1889 6799 -1855
rect 6833 -1889 6844 -1855
rect 6788 -1923 6844 -1889
rect 6788 -1957 6799 -1923
rect 6833 -1957 6844 -1923
rect 6788 -1991 6844 -1957
rect 6788 -2025 6799 -1991
rect 6833 -2025 6844 -1991
rect 6788 -2059 6844 -2025
rect 6788 -2093 6799 -2059
rect 6833 -2093 6844 -2059
rect 6788 -2105 6844 -2093
rect 6964 -1583 7020 -1505
rect 6964 -1617 6975 -1583
rect 7009 -1617 7020 -1583
rect 6964 -1651 7020 -1617
rect 6964 -1685 6975 -1651
rect 7009 -1685 7020 -1651
rect 6964 -1719 7020 -1685
rect 6964 -1753 6975 -1719
rect 7009 -1753 7020 -1719
rect 6964 -1787 7020 -1753
rect 6964 -1821 6975 -1787
rect 7009 -1821 7020 -1787
rect 6964 -1855 7020 -1821
rect 6964 -1889 6975 -1855
rect 7009 -1889 7020 -1855
rect 6964 -1923 7020 -1889
rect 6964 -1957 6975 -1923
rect 7009 -1957 7020 -1923
rect 6964 -1991 7020 -1957
rect 6964 -2025 6975 -1991
rect 7009 -2025 7020 -1991
rect 6964 -2059 7020 -2025
rect 6964 -2093 6975 -2059
rect 7009 -2093 7020 -2059
rect 6964 -2105 7020 -2093
rect 7140 -1583 7196 -1505
rect 7140 -1617 7151 -1583
rect 7185 -1617 7196 -1583
rect 7140 -1651 7196 -1617
rect 7140 -1685 7151 -1651
rect 7185 -1685 7196 -1651
rect 7140 -1719 7196 -1685
rect 7140 -1753 7151 -1719
rect 7185 -1753 7196 -1719
rect 7140 -1787 7196 -1753
rect 7140 -1821 7151 -1787
rect 7185 -1821 7196 -1787
rect 7140 -1855 7196 -1821
rect 7140 -1889 7151 -1855
rect 7185 -1889 7196 -1855
rect 7140 -1923 7196 -1889
rect 7140 -1957 7151 -1923
rect 7185 -1957 7196 -1923
rect 7140 -1991 7196 -1957
rect 7140 -2025 7151 -1991
rect 7185 -2025 7196 -1991
rect 7140 -2059 7196 -2025
rect 7140 -2093 7151 -2059
rect 7185 -2093 7196 -2059
rect 7140 -2105 7196 -2093
rect 7316 -1583 7372 -1505
rect 7316 -1617 7327 -1583
rect 7361 -1617 7372 -1583
rect 7316 -1651 7372 -1617
rect 7316 -1685 7327 -1651
rect 7361 -1685 7372 -1651
rect 7316 -1719 7372 -1685
rect 7316 -1753 7327 -1719
rect 7361 -1753 7372 -1719
rect 7316 -1787 7372 -1753
rect 7316 -1821 7327 -1787
rect 7361 -1821 7372 -1787
rect 7316 -1855 7372 -1821
rect 7316 -1889 7327 -1855
rect 7361 -1889 7372 -1855
rect 7316 -1923 7372 -1889
rect 7316 -1957 7327 -1923
rect 7361 -1957 7372 -1923
rect 7316 -1991 7372 -1957
rect 7316 -2025 7327 -1991
rect 7361 -2025 7372 -1991
rect 7316 -2059 7372 -2025
rect 7316 -2093 7327 -2059
rect 7361 -2093 7372 -2059
rect 7316 -2105 7372 -2093
rect 7492 -1583 7548 -1505
rect 7492 -1617 7503 -1583
rect 7537 -1617 7548 -1583
rect 7492 -1651 7548 -1617
rect 7492 -1685 7503 -1651
rect 7537 -1685 7548 -1651
rect 7492 -1719 7548 -1685
rect 7492 -1753 7503 -1719
rect 7537 -1753 7548 -1719
rect 7492 -1787 7548 -1753
rect 7492 -1821 7503 -1787
rect 7537 -1821 7548 -1787
rect 7492 -1855 7548 -1821
rect 7492 -1889 7503 -1855
rect 7537 -1889 7548 -1855
rect 7492 -1923 7548 -1889
rect 7492 -1957 7503 -1923
rect 7537 -1957 7548 -1923
rect 7492 -1991 7548 -1957
rect 7492 -2025 7503 -1991
rect 7537 -2025 7548 -1991
rect 7492 -2059 7548 -2025
rect 7492 -2093 7503 -2059
rect 7537 -2093 7548 -2059
rect 7492 -2105 7548 -2093
rect 7668 -1583 7721 -1505
rect 7668 -1617 7679 -1583
rect 7713 -1617 7721 -1583
rect 7668 -1651 7721 -1617
rect 7668 -1685 7679 -1651
rect 7713 -1685 7721 -1651
rect 7668 -1719 7721 -1685
rect 7668 -1753 7679 -1719
rect 7713 -1753 7721 -1719
rect 7668 -1787 7721 -1753
rect 7668 -1821 7679 -1787
rect 7713 -1821 7721 -1787
rect 7668 -1855 7721 -1821
rect 7668 -1889 7679 -1855
rect 7713 -1889 7721 -1855
rect 7668 -1923 7721 -1889
rect 7668 -1957 7679 -1923
rect 7713 -1957 7721 -1923
rect 7668 -1991 7721 -1957
rect 7668 -2025 7679 -1991
rect 7713 -2025 7721 -1991
rect 7668 -2059 7721 -2025
rect 7668 -2093 7679 -2059
rect 7713 -2093 7721 -2059
rect 7668 -2105 7721 -2093
<< mvpdiff >>
rect 4724 -326 4777 -314
rect 4724 -360 4732 -326
rect 4766 -360 4777 -326
rect 4724 -394 4777 -360
rect 4724 -428 4732 -394
rect 4766 -428 4777 -394
rect 4724 -462 4777 -428
rect 4724 -496 4732 -462
rect 4766 -496 4777 -462
rect 4724 -530 4777 -496
rect 4724 -564 4732 -530
rect 4766 -564 4777 -530
rect 4724 -598 4777 -564
rect 4724 -632 4732 -598
rect 4766 -632 4777 -598
rect 4724 -666 4777 -632
rect 4724 -700 4732 -666
rect 4766 -700 4777 -666
rect 4724 -734 4777 -700
rect 4724 -768 4732 -734
rect 4766 -768 4777 -734
rect 4724 -802 4777 -768
rect 4724 -836 4732 -802
rect 4766 -836 4777 -802
rect 4724 -914 4777 -836
rect 4877 -326 4933 -314
rect 4877 -360 4888 -326
rect 4922 -360 4933 -326
rect 4877 -394 4933 -360
rect 4877 -428 4888 -394
rect 4922 -428 4933 -394
rect 4877 -462 4933 -428
rect 4877 -496 4888 -462
rect 4922 -496 4933 -462
rect 4877 -530 4933 -496
rect 4877 -564 4888 -530
rect 4922 -564 4933 -530
rect 4877 -598 4933 -564
rect 4877 -632 4888 -598
rect 4922 -632 4933 -598
rect 4877 -666 4933 -632
rect 4877 -700 4888 -666
rect 4922 -700 4933 -666
rect 4877 -734 4933 -700
rect 4877 -768 4888 -734
rect 4922 -768 4933 -734
rect 4877 -802 4933 -768
rect 4877 -836 4888 -802
rect 4922 -836 4933 -802
rect 4877 -914 4933 -836
rect 5033 -326 5089 -314
rect 5033 -360 5044 -326
rect 5078 -360 5089 -326
rect 5033 -394 5089 -360
rect 5033 -428 5044 -394
rect 5078 -428 5089 -394
rect 5033 -462 5089 -428
rect 5033 -496 5044 -462
rect 5078 -496 5089 -462
rect 5033 -530 5089 -496
rect 5033 -564 5044 -530
rect 5078 -564 5089 -530
rect 5033 -598 5089 -564
rect 5033 -632 5044 -598
rect 5078 -632 5089 -598
rect 5033 -666 5089 -632
rect 5033 -700 5044 -666
rect 5078 -700 5089 -666
rect 5033 -734 5089 -700
rect 5033 -768 5044 -734
rect 5078 -768 5089 -734
rect 5033 -802 5089 -768
rect 5033 -836 5044 -802
rect 5078 -836 5089 -802
rect 5033 -914 5089 -836
rect 5189 -326 5242 -314
rect 5189 -360 5200 -326
rect 5234 -360 5242 -326
rect 5189 -394 5242 -360
rect 5189 -428 5200 -394
rect 5234 -428 5242 -394
rect 5189 -462 5242 -428
rect 5189 -496 5200 -462
rect 5234 -496 5242 -462
rect 5189 -530 5242 -496
rect 5189 -564 5200 -530
rect 5234 -564 5242 -530
rect 5189 -598 5242 -564
rect 5189 -632 5200 -598
rect 5234 -632 5242 -598
rect 5189 -666 5242 -632
rect 5189 -700 5200 -666
rect 5234 -700 5242 -666
rect 5189 -734 5242 -700
rect 5189 -768 5200 -734
rect 5234 -768 5242 -734
rect 5189 -802 5242 -768
rect 5189 -836 5200 -802
rect 5234 -836 5242 -802
rect 5189 -914 5242 -836
rect 5316 -326 5369 -314
rect 5316 -360 5324 -326
rect 5358 -360 5369 -326
rect 5316 -394 5369 -360
rect 5316 -428 5324 -394
rect 5358 -428 5369 -394
rect 5316 -462 5369 -428
rect 5316 -496 5324 -462
rect 5358 -496 5369 -462
rect 5316 -530 5369 -496
rect 5316 -564 5324 -530
rect 5358 -564 5369 -530
rect 5316 -598 5369 -564
rect 5316 -632 5324 -598
rect 5358 -632 5369 -598
rect 5316 -666 5369 -632
rect 5316 -700 5324 -666
rect 5358 -700 5369 -666
rect 5316 -734 5369 -700
rect 5316 -768 5324 -734
rect 5358 -768 5369 -734
rect 5316 -802 5369 -768
rect 5316 -836 5324 -802
rect 5358 -836 5369 -802
rect 5316 -914 5369 -836
rect 5469 -326 5525 -314
rect 5469 -360 5480 -326
rect 5514 -360 5525 -326
rect 5469 -394 5525 -360
rect 5469 -428 5480 -394
rect 5514 -428 5525 -394
rect 5469 -462 5525 -428
rect 5469 -496 5480 -462
rect 5514 -496 5525 -462
rect 5469 -530 5525 -496
rect 5469 -564 5480 -530
rect 5514 -564 5525 -530
rect 5469 -598 5525 -564
rect 5469 -632 5480 -598
rect 5514 -632 5525 -598
rect 5469 -666 5525 -632
rect 5469 -700 5480 -666
rect 5514 -700 5525 -666
rect 5469 -734 5525 -700
rect 5469 -768 5480 -734
rect 5514 -768 5525 -734
rect 5469 -802 5525 -768
rect 5469 -836 5480 -802
rect 5514 -836 5525 -802
rect 5469 -914 5525 -836
rect 5625 -326 5681 -314
rect 5625 -360 5636 -326
rect 5670 -360 5681 -326
rect 5625 -394 5681 -360
rect 5625 -428 5636 -394
rect 5670 -428 5681 -394
rect 5625 -462 5681 -428
rect 5625 -496 5636 -462
rect 5670 -496 5681 -462
rect 5625 -530 5681 -496
rect 5625 -564 5636 -530
rect 5670 -564 5681 -530
rect 5625 -598 5681 -564
rect 5625 -632 5636 -598
rect 5670 -632 5681 -598
rect 5625 -666 5681 -632
rect 5625 -700 5636 -666
rect 5670 -700 5681 -666
rect 5625 -734 5681 -700
rect 5625 -768 5636 -734
rect 5670 -768 5681 -734
rect 5625 -802 5681 -768
rect 5625 -836 5636 -802
rect 5670 -836 5681 -802
rect 5625 -914 5681 -836
rect 5781 -326 5837 -314
rect 5781 -360 5792 -326
rect 5826 -360 5837 -326
rect 5781 -394 5837 -360
rect 5781 -428 5792 -394
rect 5826 -428 5837 -394
rect 5781 -462 5837 -428
rect 5781 -496 5792 -462
rect 5826 -496 5837 -462
rect 5781 -530 5837 -496
rect 5781 -564 5792 -530
rect 5826 -564 5837 -530
rect 5781 -598 5837 -564
rect 5781 -632 5792 -598
rect 5826 -632 5837 -598
rect 5781 -666 5837 -632
rect 5781 -700 5792 -666
rect 5826 -700 5837 -666
rect 5781 -734 5837 -700
rect 5781 -768 5792 -734
rect 5826 -768 5837 -734
rect 5781 -802 5837 -768
rect 5781 -836 5792 -802
rect 5826 -836 5837 -802
rect 5781 -914 5837 -836
rect 5937 -326 5990 -314
rect 5937 -360 5948 -326
rect 5982 -360 5990 -326
rect 5937 -394 5990 -360
rect 5937 -428 5948 -394
rect 5982 -428 5990 -394
rect 5937 -462 5990 -428
rect 5937 -496 5948 -462
rect 5982 -496 5990 -462
rect 5937 -530 5990 -496
rect 5937 -564 5948 -530
rect 5982 -564 5990 -530
rect 5937 -598 5990 -564
rect 5937 -632 5948 -598
rect 5982 -632 5990 -598
rect 5937 -666 5990 -632
rect 5937 -700 5948 -666
rect 5982 -700 5990 -666
rect 5937 -734 5990 -700
rect 5937 -768 5948 -734
rect 5982 -768 5990 -734
rect 5937 -802 5990 -768
rect 5937 -836 5948 -802
rect 5982 -836 5990 -802
rect 5937 -914 5990 -836
rect 6064 -326 6117 -314
rect 6064 -360 6072 -326
rect 6106 -360 6117 -326
rect 6064 -394 6117 -360
rect 6064 -428 6072 -394
rect 6106 -428 6117 -394
rect 6064 -462 6117 -428
rect 6064 -496 6072 -462
rect 6106 -496 6117 -462
rect 6064 -530 6117 -496
rect 6064 -564 6072 -530
rect 6106 -564 6117 -530
rect 6064 -598 6117 -564
rect 6064 -632 6072 -598
rect 6106 -632 6117 -598
rect 6064 -666 6117 -632
rect 6064 -700 6072 -666
rect 6106 -700 6117 -666
rect 6064 -734 6117 -700
rect 6064 -768 6072 -734
rect 6106 -768 6117 -734
rect 6064 -802 6117 -768
rect 6064 -836 6072 -802
rect 6106 -836 6117 -802
rect 6064 -914 6117 -836
rect 6217 -326 6273 -314
rect 6217 -360 6228 -326
rect 6262 -360 6273 -326
rect 6217 -394 6273 -360
rect 6217 -428 6228 -394
rect 6262 -428 6273 -394
rect 6217 -462 6273 -428
rect 6217 -496 6228 -462
rect 6262 -496 6273 -462
rect 6217 -530 6273 -496
rect 6217 -564 6228 -530
rect 6262 -564 6273 -530
rect 6217 -598 6273 -564
rect 6217 -632 6228 -598
rect 6262 -632 6273 -598
rect 6217 -666 6273 -632
rect 6217 -700 6228 -666
rect 6262 -700 6273 -666
rect 6217 -734 6273 -700
rect 6217 -768 6228 -734
rect 6262 -768 6273 -734
rect 6217 -802 6273 -768
rect 6217 -836 6228 -802
rect 6262 -836 6273 -802
rect 6217 -914 6273 -836
rect 6373 -326 6426 -314
rect 6373 -360 6384 -326
rect 6418 -360 6426 -326
rect 6373 -394 6426 -360
rect 7724 -351 7808 -343
rect 7724 -385 7736 -351
rect 7770 -385 7808 -351
rect 6373 -428 6384 -394
rect 6418 -428 6426 -394
rect 6373 -462 6426 -428
rect 6373 -496 6384 -462
rect 6418 -496 6426 -462
rect 6596 -431 6649 -393
rect 6596 -465 6604 -431
rect 6638 -465 6649 -431
rect 6596 -477 6649 -465
rect 7449 -431 7502 -393
rect 7724 -396 7808 -385
rect 7449 -465 7460 -431
rect 7494 -465 7502 -431
rect 7449 -477 7502 -465
rect 6373 -530 6426 -496
rect 6373 -564 6384 -530
rect 6418 -564 6426 -530
rect 6373 -598 6426 -564
rect 6373 -632 6384 -598
rect 6418 -632 6426 -598
rect 6373 -666 6426 -632
rect 6373 -700 6384 -666
rect 6418 -700 6426 -666
rect 6596 -645 6649 -607
rect 6596 -679 6604 -645
rect 6638 -679 6649 -645
rect 6596 -691 6649 -679
rect 7449 -645 7502 -607
rect 7449 -679 7460 -645
rect 7494 -679 7502 -645
rect 7449 -691 7502 -679
rect 7724 -607 7808 -596
rect 7724 -641 7736 -607
rect 7770 -641 7808 -607
rect 7724 -652 7808 -641
rect 6373 -734 6426 -700
rect 6373 -768 6384 -734
rect 6418 -768 6426 -734
rect 6373 -802 6426 -768
rect 6373 -836 6384 -802
rect 6418 -836 6426 -802
rect 6373 -914 6426 -836
rect 6596 -813 6649 -801
rect 6596 -847 6604 -813
rect 6638 -847 6649 -813
rect 6596 -885 6649 -847
rect 7449 -813 7502 -801
rect 7449 -847 7460 -813
rect 7494 -847 7502 -813
rect 7449 -885 7502 -847
rect 7724 -863 7808 -852
rect 7724 -897 7736 -863
rect 7770 -897 7808 -863
rect 7724 -905 7808 -897
rect 7724 -987 7808 -979
rect 7724 -1021 7736 -987
rect 7770 -1021 7808 -987
rect 6596 -1065 6649 -1027
rect 6596 -1099 6604 -1065
rect 6638 -1099 6649 -1065
rect 6596 -1111 6649 -1099
rect 7449 -1065 7502 -1027
rect 7724 -1032 7808 -1021
rect 7449 -1099 7460 -1065
rect 7494 -1099 7502 -1065
rect 7449 -1111 7502 -1099
rect 7724 -1243 7808 -1232
rect 6596 -1281 6649 -1243
rect 6596 -1315 6604 -1281
rect 6638 -1315 6649 -1281
rect 6596 -1327 6649 -1315
rect 7449 -1281 7502 -1243
rect 7449 -1315 7460 -1281
rect 7494 -1315 7502 -1281
rect 7724 -1277 7736 -1243
rect 7770 -1277 7808 -1243
rect 7724 -1285 7808 -1277
rect 7449 -1327 7502 -1315
<< mvndiffc >>
rect 6447 -1617 6481 -1583
rect 6447 -1685 6481 -1651
rect 6447 -1753 6481 -1719
rect 6447 -1821 6481 -1787
rect 6447 -1889 6481 -1855
rect 6447 -1957 6481 -1923
rect 6447 -2025 6481 -1991
rect 6447 -2093 6481 -2059
rect 6623 -1617 6657 -1583
rect 6623 -1685 6657 -1651
rect 6623 -1753 6657 -1719
rect 6623 -1821 6657 -1787
rect 6623 -1889 6657 -1855
rect 6623 -1957 6657 -1923
rect 6623 -2025 6657 -1991
rect 6623 -2093 6657 -2059
rect 6799 -1617 6833 -1583
rect 6799 -1685 6833 -1651
rect 6799 -1753 6833 -1719
rect 6799 -1821 6833 -1787
rect 6799 -1889 6833 -1855
rect 6799 -1957 6833 -1923
rect 6799 -2025 6833 -1991
rect 6799 -2093 6833 -2059
rect 6975 -1617 7009 -1583
rect 6975 -1685 7009 -1651
rect 6975 -1753 7009 -1719
rect 6975 -1821 7009 -1787
rect 6975 -1889 7009 -1855
rect 6975 -1957 7009 -1923
rect 6975 -2025 7009 -1991
rect 6975 -2093 7009 -2059
rect 7151 -1617 7185 -1583
rect 7151 -1685 7185 -1651
rect 7151 -1753 7185 -1719
rect 7151 -1821 7185 -1787
rect 7151 -1889 7185 -1855
rect 7151 -1957 7185 -1923
rect 7151 -2025 7185 -1991
rect 7151 -2093 7185 -2059
rect 7327 -1617 7361 -1583
rect 7327 -1685 7361 -1651
rect 7327 -1753 7361 -1719
rect 7327 -1821 7361 -1787
rect 7327 -1889 7361 -1855
rect 7327 -1957 7361 -1923
rect 7327 -2025 7361 -1991
rect 7327 -2093 7361 -2059
rect 7503 -1617 7537 -1583
rect 7503 -1685 7537 -1651
rect 7503 -1753 7537 -1719
rect 7503 -1821 7537 -1787
rect 7503 -1889 7537 -1855
rect 7503 -1957 7537 -1923
rect 7503 -2025 7537 -1991
rect 7503 -2093 7537 -2059
rect 7679 -1617 7713 -1583
rect 7679 -1685 7713 -1651
rect 7679 -1753 7713 -1719
rect 7679 -1821 7713 -1787
rect 7679 -1889 7713 -1855
rect 7679 -1957 7713 -1923
rect 7679 -2025 7713 -1991
rect 7679 -2093 7713 -2059
<< mvpdiffc >>
rect 4732 -360 4766 -326
rect 4732 -428 4766 -394
rect 4732 -496 4766 -462
rect 4732 -564 4766 -530
rect 4732 -632 4766 -598
rect 4732 -700 4766 -666
rect 4732 -768 4766 -734
rect 4732 -836 4766 -802
rect 4888 -360 4922 -326
rect 4888 -428 4922 -394
rect 4888 -496 4922 -462
rect 4888 -564 4922 -530
rect 4888 -632 4922 -598
rect 4888 -700 4922 -666
rect 4888 -768 4922 -734
rect 4888 -836 4922 -802
rect 5044 -360 5078 -326
rect 5044 -428 5078 -394
rect 5044 -496 5078 -462
rect 5044 -564 5078 -530
rect 5044 -632 5078 -598
rect 5044 -700 5078 -666
rect 5044 -768 5078 -734
rect 5044 -836 5078 -802
rect 5200 -360 5234 -326
rect 5200 -428 5234 -394
rect 5200 -496 5234 -462
rect 5200 -564 5234 -530
rect 5200 -632 5234 -598
rect 5200 -700 5234 -666
rect 5200 -768 5234 -734
rect 5200 -836 5234 -802
rect 5324 -360 5358 -326
rect 5324 -428 5358 -394
rect 5324 -496 5358 -462
rect 5324 -564 5358 -530
rect 5324 -632 5358 -598
rect 5324 -700 5358 -666
rect 5324 -768 5358 -734
rect 5324 -836 5358 -802
rect 5480 -360 5514 -326
rect 5480 -428 5514 -394
rect 5480 -496 5514 -462
rect 5480 -564 5514 -530
rect 5480 -632 5514 -598
rect 5480 -700 5514 -666
rect 5480 -768 5514 -734
rect 5480 -836 5514 -802
rect 5636 -360 5670 -326
rect 5636 -428 5670 -394
rect 5636 -496 5670 -462
rect 5636 -564 5670 -530
rect 5636 -632 5670 -598
rect 5636 -700 5670 -666
rect 5636 -768 5670 -734
rect 5636 -836 5670 -802
rect 5792 -360 5826 -326
rect 5792 -428 5826 -394
rect 5792 -496 5826 -462
rect 5792 -564 5826 -530
rect 5792 -632 5826 -598
rect 5792 -700 5826 -666
rect 5792 -768 5826 -734
rect 5792 -836 5826 -802
rect 5948 -360 5982 -326
rect 5948 -428 5982 -394
rect 5948 -496 5982 -462
rect 5948 -564 5982 -530
rect 5948 -632 5982 -598
rect 5948 -700 5982 -666
rect 5948 -768 5982 -734
rect 5948 -836 5982 -802
rect 6072 -360 6106 -326
rect 6072 -428 6106 -394
rect 6072 -496 6106 -462
rect 6072 -564 6106 -530
rect 6072 -632 6106 -598
rect 6072 -700 6106 -666
rect 6072 -768 6106 -734
rect 6072 -836 6106 -802
rect 6228 -360 6262 -326
rect 6228 -428 6262 -394
rect 6228 -496 6262 -462
rect 6228 -564 6262 -530
rect 6228 -632 6262 -598
rect 6228 -700 6262 -666
rect 6228 -768 6262 -734
rect 6228 -836 6262 -802
rect 6384 -360 6418 -326
rect 7736 -385 7770 -351
rect 6384 -428 6418 -394
rect 6384 -496 6418 -462
rect 6604 -465 6638 -431
rect 7460 -465 7494 -431
rect 6384 -564 6418 -530
rect 6384 -632 6418 -598
rect 6384 -700 6418 -666
rect 6604 -679 6638 -645
rect 7460 -679 7494 -645
rect 7736 -641 7770 -607
rect 6384 -768 6418 -734
rect 6384 -836 6418 -802
rect 6604 -847 6638 -813
rect 7460 -847 7494 -813
rect 7736 -897 7770 -863
rect 7736 -1021 7770 -987
rect 6604 -1099 6638 -1065
rect 7460 -1099 7494 -1065
rect 6604 -1315 6638 -1281
rect 7460 -1315 7494 -1281
rect 7736 -1277 7770 -1243
<< psubdiff >>
rect 6331 -1559 6365 -1535
rect 6331 -1627 6365 -1593
rect 6331 -1695 6365 -1661
rect 6331 -1763 6365 -1729
rect 6331 -1831 6365 -1797
rect 6331 -1900 6365 -1865
rect 6331 -1969 6365 -1934
rect 6331 -2038 6365 -2003
rect 6331 -2096 6365 -2072
<< psubdiffcont >>
rect 6331 -1593 6365 -1559
rect 6331 -1661 6365 -1627
rect 6331 -1729 6365 -1695
rect 6331 -1797 6365 -1763
rect 6331 -1865 6365 -1831
rect 6331 -1934 6365 -1900
rect 6331 -2003 6365 -1969
rect 6331 -2072 6365 -2038
<< poly >>
rect 4777 -314 4877 -282
rect 4933 -314 5033 -282
rect 5089 -314 5189 -282
rect 5369 -314 5469 -282
rect 5525 -314 5625 -282
rect 5681 -314 5781 -282
rect 5837 -314 5937 -282
rect 6117 -314 6217 -282
rect 6273 -314 6373 -282
rect 6649 -393 7449 -361
rect 7626 -412 7724 -396
rect 7626 -446 7642 -412
rect 7676 -446 7724 -412
rect 6649 -525 7449 -477
rect 6649 -559 6665 -525
rect 6699 -559 6739 -525
rect 6773 -559 6813 -525
rect 6847 -559 6887 -525
rect 6921 -559 6961 -525
rect 6995 -559 7034 -525
rect 7068 -559 7107 -525
rect 7141 -559 7180 -525
rect 7214 -559 7253 -525
rect 7287 -559 7326 -525
rect 7360 -559 7399 -525
rect 7433 -559 7449 -525
rect 6649 -607 7449 -559
rect 7626 -484 7724 -446
rect 7626 -518 7642 -484
rect 7676 -518 7724 -484
rect 7626 -556 7724 -518
rect 7626 -590 7642 -556
rect 7676 -590 7724 -556
rect 7626 -596 7724 -590
rect 7808 -596 7840 -396
rect 7626 -629 7692 -596
rect 7626 -663 7642 -629
rect 7676 -652 7692 -629
rect 7676 -663 7724 -652
rect 6649 -723 7449 -691
rect 7626 -702 7724 -663
rect 7626 -736 7642 -702
rect 7676 -736 7724 -702
rect 6649 -801 7449 -769
rect 7626 -775 7724 -736
rect 7626 -809 7642 -775
rect 7676 -809 7724 -775
rect 7626 -852 7724 -809
rect 7808 -852 7840 -652
rect 4777 -946 4877 -914
rect 4933 -946 5033 -914
rect 5089 -946 5189 -914
rect 4777 -962 5189 -946
rect 4777 -996 4793 -962
rect 4827 -996 4863 -962
rect 4897 -996 4932 -962
rect 4966 -996 5001 -962
rect 5035 -996 5070 -962
rect 5104 -996 5139 -962
rect 5173 -996 5189 -962
rect 4777 -1012 5189 -996
rect 5369 -946 5469 -914
rect 5525 -946 5625 -914
rect 5681 -946 5781 -914
rect 5837 -946 5937 -914
rect 5369 -962 5937 -946
rect 5369 -996 5385 -962
rect 5419 -996 5456 -962
rect 5490 -996 5527 -962
rect 5561 -996 5599 -962
rect 5633 -996 5671 -962
rect 5705 -996 5743 -962
rect 5777 -996 5815 -962
rect 5849 -996 5887 -962
rect 5921 -996 5937 -962
rect 5369 -1012 5937 -996
rect 6117 -963 6217 -914
rect 6117 -997 6167 -963
rect 6201 -997 6217 -963
rect 6117 -1031 6217 -997
rect 6117 -1065 6167 -1031
rect 6201 -1065 6217 -1031
rect 6117 -1081 6217 -1065
rect 6273 -963 6373 -914
rect 6273 -997 6306 -963
rect 6340 -997 6373 -963
rect 6273 -1031 6373 -997
rect 6649 -939 7449 -885
rect 6649 -973 6665 -939
rect 6699 -973 6738 -939
rect 6772 -973 6811 -939
rect 6845 -973 6884 -939
rect 6918 -973 6957 -939
rect 6991 -973 7030 -939
rect 7064 -973 7103 -939
rect 7137 -973 7177 -939
rect 7211 -973 7251 -939
rect 7285 -973 7325 -939
rect 7359 -973 7399 -939
rect 7433 -973 7449 -939
rect 6649 -1027 7449 -973
rect 6273 -1065 6306 -1031
rect 6340 -1065 6373 -1031
rect 6273 -1081 6373 -1065
rect 7626 -1093 7724 -1032
rect 6649 -1160 7449 -1111
rect 6649 -1194 6675 -1160
rect 6709 -1194 6744 -1160
rect 6778 -1194 6813 -1160
rect 6847 -1194 6881 -1160
rect 6915 -1194 6949 -1160
rect 6983 -1194 7017 -1160
rect 7051 -1194 7085 -1160
rect 7119 -1194 7153 -1160
rect 7187 -1194 7221 -1160
rect 7255 -1194 7289 -1160
rect 7323 -1194 7357 -1160
rect 7391 -1194 7449 -1160
rect 6649 -1243 7449 -1194
rect 7626 -1127 7642 -1093
rect 7676 -1127 7724 -1093
rect 7626 -1178 7724 -1127
rect 7626 -1212 7642 -1178
rect 7676 -1212 7724 -1178
rect 7626 -1232 7724 -1212
rect 7808 -1232 7840 -1032
rect 6649 -1359 7449 -1327
rect 6468 -1423 6612 -1407
rect 6468 -1457 6484 -1423
rect 6518 -1457 6562 -1423
rect 6596 -1457 6612 -1423
rect 6468 -1473 6612 -1457
rect 6492 -1505 6612 -1473
rect 6668 -1423 6964 -1407
rect 6668 -1457 6684 -1423
rect 6718 -1457 6761 -1423
rect 6795 -1457 6838 -1423
rect 6872 -1457 6914 -1423
rect 6948 -1457 6964 -1423
rect 6668 -1473 6964 -1457
rect 6668 -1505 6788 -1473
rect 6844 -1505 6964 -1473
rect 7020 -1423 7316 -1359
rect 7020 -1457 7036 -1423
rect 7070 -1457 7113 -1423
rect 7147 -1457 7190 -1423
rect 7224 -1457 7266 -1423
rect 7300 -1457 7316 -1423
rect 7020 -1473 7316 -1457
rect 7020 -1505 7140 -1473
rect 7196 -1505 7316 -1473
rect 7372 -1423 7668 -1407
rect 7372 -1457 7388 -1423
rect 7422 -1457 7464 -1423
rect 7498 -1457 7541 -1423
rect 7575 -1457 7618 -1423
rect 7652 -1457 7668 -1423
rect 7372 -1473 7668 -1457
rect 7372 -1505 7492 -1473
rect 7548 -1505 7668 -1473
rect 6492 -2137 6612 -2105
rect 6668 -2137 6788 -2105
rect 6844 -2137 6964 -2105
rect 7020 -2137 7140 -2105
rect 7196 -2137 7316 -2105
rect 7372 -2137 7492 -2105
rect 7548 -2137 7668 -2105
<< polycont >>
rect 7642 -446 7676 -412
rect 6665 -559 6699 -525
rect 6739 -559 6773 -525
rect 6813 -559 6847 -525
rect 6887 -559 6921 -525
rect 6961 -559 6995 -525
rect 7034 -559 7068 -525
rect 7107 -559 7141 -525
rect 7180 -559 7214 -525
rect 7253 -559 7287 -525
rect 7326 -559 7360 -525
rect 7399 -559 7433 -525
rect 7642 -518 7676 -484
rect 7642 -590 7676 -556
rect 7642 -663 7676 -629
rect 7642 -736 7676 -702
rect 7642 -809 7676 -775
rect 4793 -996 4827 -962
rect 4863 -996 4897 -962
rect 4932 -996 4966 -962
rect 5001 -996 5035 -962
rect 5070 -996 5104 -962
rect 5139 -996 5173 -962
rect 5385 -996 5419 -962
rect 5456 -996 5490 -962
rect 5527 -996 5561 -962
rect 5599 -996 5633 -962
rect 5671 -996 5705 -962
rect 5743 -996 5777 -962
rect 5815 -996 5849 -962
rect 5887 -996 5921 -962
rect 6167 -997 6201 -963
rect 6167 -1065 6201 -1031
rect 6306 -997 6340 -963
rect 6665 -973 6699 -939
rect 6738 -973 6772 -939
rect 6811 -973 6845 -939
rect 6884 -973 6918 -939
rect 6957 -973 6991 -939
rect 7030 -973 7064 -939
rect 7103 -973 7137 -939
rect 7177 -973 7211 -939
rect 7251 -973 7285 -939
rect 7325 -973 7359 -939
rect 7399 -973 7433 -939
rect 6306 -1065 6340 -1031
rect 6675 -1194 6709 -1160
rect 6744 -1194 6778 -1160
rect 6813 -1194 6847 -1160
rect 6881 -1194 6915 -1160
rect 6949 -1194 6983 -1160
rect 7017 -1194 7051 -1160
rect 7085 -1194 7119 -1160
rect 7153 -1194 7187 -1160
rect 7221 -1194 7255 -1160
rect 7289 -1194 7323 -1160
rect 7357 -1194 7391 -1160
rect 7642 -1127 7676 -1093
rect 7642 -1212 7676 -1178
rect 6484 -1457 6518 -1423
rect 6562 -1457 6596 -1423
rect 6684 -1457 6718 -1423
rect 6761 -1457 6795 -1423
rect 6838 -1457 6872 -1423
rect 6914 -1457 6948 -1423
rect 7036 -1457 7070 -1423
rect 7113 -1457 7147 -1423
rect 7190 -1457 7224 -1423
rect 7266 -1457 7300 -1423
rect 7388 -1457 7422 -1423
rect 7464 -1457 7498 -1423
rect 7541 -1457 7575 -1423
rect 7618 -1457 7652 -1423
<< locali >>
rect 4732 -326 4766 -310
rect 4732 -394 4766 -360
rect 4888 -326 4922 -310
rect 4888 -379 4922 -360
rect 5044 -326 5078 -310
rect 4886 -394 4924 -379
rect 4886 -413 4888 -394
rect 4732 -462 4766 -428
rect 4732 -530 4766 -524
rect 4732 -586 4766 -564
rect 4732 -666 4766 -632
rect 4732 -734 4766 -700
rect 4732 -802 4766 -768
rect 4732 -852 4766 -836
rect 4922 -413 4924 -394
rect 5044 -394 5078 -360
rect 5200 -326 5234 -310
rect 5200 -379 5234 -360
rect 5324 -326 5358 -310
rect 4888 -462 4922 -428
rect 4888 -530 4922 -496
rect 4888 -598 4922 -564
rect 4888 -666 4922 -632
rect 4888 -734 4922 -700
rect 4888 -802 4922 -768
rect 4888 -852 4922 -836
rect 5191 -394 5229 -379
rect 5191 -413 5200 -394
rect 5324 -394 5358 -360
rect 5044 -462 5078 -428
rect 5044 -530 5078 -524
rect 5044 -586 5078 -564
rect 5044 -666 5078 -632
rect 5044 -734 5078 -700
rect 5044 -802 5078 -768
rect 5044 -852 5078 -836
rect 5200 -462 5234 -428
rect 5324 -462 5358 -428
rect 5480 -326 5514 -310
rect 5480 -394 5514 -360
rect 5480 -462 5514 -428
rect 5200 -530 5234 -496
rect 5358 -496 5367 -465
rect 5329 -499 5367 -496
rect 5636 -326 5670 -310
rect 5636 -394 5670 -360
rect 5636 -462 5670 -428
rect 5200 -598 5234 -564
rect 5200 -666 5234 -632
rect 5200 -734 5234 -700
rect 5200 -802 5234 -768
rect 5200 -852 5234 -836
rect 5324 -530 5358 -499
rect 5480 -530 5514 -496
rect 5632 -496 5636 -465
rect 5792 -326 5826 -310
rect 5792 -394 5826 -360
rect 5792 -462 5826 -428
rect 5632 -499 5670 -496
rect 5948 -326 5982 -310
rect 5948 -394 5982 -360
rect 5948 -462 5982 -428
rect 5324 -598 5358 -564
rect 5478 -564 5480 -542
rect 5636 -530 5670 -499
rect 5514 -564 5516 -542
rect 5478 -576 5516 -564
rect 5324 -666 5358 -632
rect 5324 -734 5358 -700
rect 5324 -802 5358 -768
rect 5324 -852 5358 -836
rect 5480 -598 5514 -576
rect 5480 -666 5514 -632
rect 5480 -734 5514 -700
rect 5480 -802 5514 -768
rect 5480 -852 5514 -836
rect 5636 -598 5670 -564
rect 5792 -530 5826 -496
rect 5945 -496 5948 -465
rect 6072 -326 6106 -310
rect 6072 -394 6106 -360
rect 6228 -326 6262 -310
rect 6228 -379 6262 -360
rect 6384 -326 6418 -310
rect 6072 -462 6106 -428
rect 5982 -496 5983 -465
rect 5945 -499 5983 -496
rect 5792 -598 5826 -564
rect 5636 -666 5670 -632
rect 5791 -632 5792 -620
rect 5948 -530 5982 -499
rect 6072 -530 6106 -496
rect 5948 -598 5982 -564
rect 6071 -564 6072 -542
rect 6228 -394 6266 -379
rect 6194 -428 6228 -413
rect 6262 -413 6266 -394
rect 6262 -428 6300 -413
rect 6194 -462 6300 -428
rect 6194 -496 6228 -462
rect 6262 -496 6300 -462
rect 6194 -530 6300 -496
rect 6106 -564 6109 -542
rect 6071 -576 6109 -564
rect 6194 -564 6228 -530
rect 6262 -564 6300 -530
rect 5826 -632 5829 -620
rect 5791 -654 5829 -632
rect 5636 -734 5670 -700
rect 5792 -666 5826 -654
rect 5792 -734 5826 -700
rect 5636 -802 5670 -768
rect 5636 -852 5670 -836
rect 5712 -815 5746 -777
rect 4777 -909 5309 -886
rect 4777 -943 5186 -909
rect 5220 -943 5258 -909
rect 5292 -943 5309 -909
rect 4777 -962 5309 -943
rect 5712 -962 5746 -849
rect 5948 -666 5982 -632
rect 5948 -734 5982 -700
rect 5792 -802 5826 -768
rect 5792 -852 5826 -836
rect 5872 -815 5906 -777
rect 5872 -962 5906 -849
rect 5948 -802 5982 -768
rect 5948 -852 5982 -836
rect 6072 -598 6106 -576
rect 6072 -666 6106 -632
rect 6072 -734 6106 -700
rect 6072 -802 6106 -768
rect 6072 -852 6106 -836
rect 6194 -598 6300 -564
rect 6194 -632 6228 -598
rect 6262 -632 6300 -598
rect 6384 -394 6418 -360
rect 7460 -353 7461 -319
rect 7495 -353 7533 -319
rect 6557 -413 6595 -379
rect 6629 -413 6638 -379
rect 6384 -462 6418 -428
rect 6604 -431 6638 -413
rect 6604 -481 6638 -465
rect 7460 -431 7567 -353
rect 7720 -385 7736 -351
rect 7770 -385 7786 -351
rect 7494 -465 7567 -431
rect 7460 -481 7567 -465
rect 7642 -412 7676 -396
rect 6384 -530 6418 -496
rect 7642 -484 7676 -446
rect 6384 -598 6418 -564
rect 6531 -518 7642 -515
rect 7720 -412 7786 -385
rect 7720 -446 7732 -412
rect 7766 -446 7786 -412
rect 7720 -484 7786 -446
rect 7720 -518 7732 -484
rect 7766 -518 7786 -484
rect 6531 -523 7676 -518
rect 6531 -557 6543 -523
rect 6577 -557 6615 -523
rect 6649 -525 7676 -523
rect 6649 -557 6665 -525
rect 6531 -559 6665 -557
rect 6699 -559 6739 -525
rect 6773 -559 6813 -525
rect 6847 -559 6887 -525
rect 6921 -559 6961 -525
rect 6995 -559 7034 -525
rect 7068 -559 7107 -525
rect 7141 -559 7180 -525
rect 7214 -559 7253 -525
rect 7287 -559 7326 -525
rect 7360 -559 7399 -525
rect 7433 -556 7676 -525
rect 7433 -559 7642 -556
rect 6531 -575 7642 -559
rect 6194 -666 6300 -632
rect 6418 -632 6422 -620
rect 6384 -654 6422 -632
rect 7642 -629 7676 -590
rect 6604 -645 6638 -629
rect 6194 -700 6228 -666
rect 6262 -700 6300 -666
rect 6194 -734 6300 -700
rect 6194 -768 6228 -734
rect 6262 -768 6300 -734
rect 6194 -802 6300 -768
rect 6194 -833 6228 -802
rect 6262 -833 6300 -802
rect 6262 -836 6266 -833
rect 6228 -867 6266 -836
rect 6384 -666 6418 -654
rect 6384 -734 6418 -700
rect 6384 -802 6418 -768
rect 6604 -813 6638 -679
rect 7460 -645 7608 -629
rect 7494 -649 7608 -645
rect 7460 -683 7466 -679
rect 7500 -683 7538 -649
rect 7572 -683 7608 -649
rect 7460 -695 7608 -683
rect 6384 -852 6418 -836
rect 6495 -867 6533 -833
rect 6567 -867 6569 -833
rect 6604 -863 6638 -847
rect 7460 -798 7494 -797
rect 7460 -813 7532 -798
rect 7494 -847 7532 -813
rect 6137 -943 6175 -909
rect 4777 -996 4793 -962
rect 4827 -996 4863 -962
rect 4897 -996 4932 -962
rect 4966 -996 5001 -962
rect 5035 -996 5070 -962
rect 5104 -996 5139 -962
rect 5173 -996 5309 -962
rect 5369 -996 5385 -962
rect 5419 -996 5456 -962
rect 5490 -996 5527 -962
rect 5561 -996 5599 -962
rect 5633 -996 5671 -962
rect 5705 -996 5743 -962
rect 5777 -996 5815 -962
rect 5849 -996 5887 -962
rect 5921 -996 5937 -962
rect 6167 -963 6201 -943
rect 4777 -1000 5309 -996
rect 6167 -1031 6201 -997
rect 6167 -1081 6201 -1065
rect 6266 -963 6373 -914
rect 6266 -997 6306 -963
rect 6340 -997 6373 -963
rect 6266 -1031 6373 -997
rect 6266 -1065 6306 -1031
rect 6340 -1065 6373 -1031
rect 6266 -1306 6373 -1065
rect 6461 -1016 6569 -867
rect 7460 -895 7532 -847
rect 6649 -939 7449 -933
rect 6649 -973 6665 -939
rect 6699 -973 6738 -939
rect 6772 -973 6811 -939
rect 6845 -973 6884 -939
rect 6918 -973 6957 -939
rect 6991 -973 7030 -939
rect 7064 -973 7103 -939
rect 7137 -973 7177 -939
rect 7211 -973 7251 -939
rect 7285 -973 7325 -939
rect 7359 -973 7399 -939
rect 7433 -973 7449 -939
rect 6649 -979 7449 -973
rect 7491 -959 7532 -895
rect 7566 -863 7608 -695
rect 7642 -702 7676 -663
rect 7719 -607 7919 -562
rect 7719 -641 7736 -607
rect 7770 -641 7919 -607
rect 7719 -674 7919 -641
rect 7642 -775 7676 -736
rect 7642 -825 7676 -809
rect 7721 -740 7787 -735
rect 7721 -774 7732 -740
rect 7766 -774 7787 -740
rect 7721 -812 7787 -774
rect 7721 -846 7732 -812
rect 7766 -846 7787 -812
rect 7721 -863 7787 -846
rect 7566 -897 7736 -863
rect 7770 -897 7787 -863
rect 7566 -925 7787 -897
rect 6461 -1065 6638 -1016
rect 6461 -1099 6604 -1065
rect 6461 -1116 6638 -1099
rect 7020 -1159 7315 -979
rect 7491 -987 7786 -959
rect 7491 -991 7736 -987
rect 7770 -991 7786 -987
rect 7491 -1015 7524 -991
rect 7558 -1025 7598 -991
rect 7632 -1025 7671 -991
rect 7705 -1021 7736 -991
rect 7705 -1025 7744 -1021
rect 7778 -1025 7786 -991
rect 7460 -1065 7498 -1049
rect 7494 -1099 7536 -1065
rect 6659 -1160 7407 -1159
rect 6659 -1194 6675 -1160
rect 6709 -1194 6744 -1160
rect 6778 -1194 6813 -1160
rect 6847 -1194 6881 -1160
rect 6915 -1194 6949 -1160
rect 6983 -1194 7017 -1160
rect 7051 -1194 7085 -1160
rect 7119 -1194 7153 -1160
rect 7187 -1194 7221 -1160
rect 7255 -1194 7289 -1160
rect 7323 -1194 7357 -1160
rect 7391 -1194 7407 -1160
rect 6659 -1195 7407 -1194
rect 6266 -1340 6267 -1306
rect 6301 -1340 6339 -1306
rect 6266 -1346 6373 -1340
rect 6479 -1253 6517 -1219
rect 6551 -1253 6570 -1219
rect 6445 -1423 6570 -1253
rect 6604 -1281 6638 -1265
rect 6638 -1315 6843 -1289
rect 6604 -1316 6843 -1315
rect 6604 -1350 6736 -1316
rect 6770 -1350 6808 -1316
rect 6842 -1350 6843 -1316
rect 6604 -1355 6843 -1350
rect 6725 -1423 6767 -1407
rect 6801 -1423 6843 -1407
rect 6877 -1423 6918 -1407
rect 7020 -1423 7315 -1195
rect 7460 -1281 7536 -1099
rect 7570 -1093 7676 -1059
rect 7570 -1127 7642 -1093
rect 7570 -1178 7676 -1127
rect 7570 -1212 7642 -1178
rect 7570 -1213 7676 -1212
rect 7604 -1247 7642 -1213
rect 7822 -1243 7919 -674
rect 7494 -1315 7536 -1281
rect 7460 -1331 7536 -1315
rect 7720 -1277 7736 -1243
rect 7770 -1277 7919 -1243
rect 7720 -1339 7919 -1277
rect 7429 -1423 7471 -1407
rect 7505 -1423 7547 -1407
rect 7581 -1423 7622 -1407
rect 6445 -1457 6484 -1423
rect 6518 -1457 6562 -1423
rect 6596 -1457 6612 -1423
rect 6668 -1457 6684 -1423
rect 6725 -1441 6761 -1423
rect 6801 -1441 6838 -1423
rect 6877 -1441 6914 -1423
rect 6952 -1441 6964 -1423
rect 6718 -1457 6761 -1441
rect 6795 -1457 6838 -1441
rect 6872 -1457 6914 -1441
rect 6948 -1457 6964 -1441
rect 7020 -1457 7036 -1423
rect 7070 -1457 7113 -1423
rect 7147 -1457 7190 -1423
rect 7224 -1457 7266 -1423
rect 7300 -1457 7316 -1423
rect 7372 -1457 7388 -1423
rect 7429 -1441 7464 -1423
rect 7505 -1441 7541 -1423
rect 7581 -1441 7618 -1423
rect 7656 -1441 7668 -1423
rect 7422 -1457 7464 -1441
rect 7498 -1457 7541 -1441
rect 7575 -1457 7618 -1441
rect 7652 -1457 7668 -1441
rect 7020 -1487 7315 -1457
rect 7020 -1521 7080 -1487
rect 7114 -1521 7152 -1487
rect 7186 -1521 7315 -1487
rect 7020 -1523 7315 -1521
rect 6331 -1559 6481 -1535
rect 6365 -1583 6481 -1559
rect 6365 -1620 6447 -1583
rect 6331 -1627 6481 -1620
rect 6365 -1651 6481 -1627
rect 6365 -1692 6447 -1651
rect 6331 -1695 6481 -1692
rect 6365 -1719 6481 -1695
rect 6365 -1729 6447 -1719
rect 6331 -1753 6447 -1729
rect 6331 -1763 6481 -1753
rect 6365 -1787 6481 -1763
rect 6365 -1797 6447 -1787
rect 6331 -1821 6447 -1797
rect 6331 -1831 6481 -1821
rect 6365 -1855 6481 -1831
rect 6365 -1865 6447 -1855
rect 6331 -1889 6447 -1865
rect 6331 -1900 6481 -1889
rect 6365 -1923 6481 -1900
rect 6365 -1934 6447 -1923
rect 6331 -1957 6447 -1934
rect 6331 -1969 6481 -1957
rect 6365 -1991 6481 -1969
rect 6365 -2003 6447 -1991
rect 6331 -2025 6447 -2003
rect 6331 -2038 6481 -2025
rect 6365 -2059 6481 -2038
rect 6365 -2072 6447 -2059
rect 6331 -2093 6447 -2072
rect 6331 -2096 6481 -2093
rect 6447 -2109 6481 -2096
rect 6623 -1583 6657 -1567
rect 6623 -1651 6657 -1617
rect 6623 -1719 6657 -1685
rect 6623 -1787 6657 -1753
rect 6623 -1855 6657 -1821
rect 6623 -1923 6657 -1889
rect 6623 -1991 6657 -1957
rect 6623 -2059 6657 -2025
rect 6623 -2122 6657 -2093
rect 6799 -1583 6833 -1567
rect 6799 -1651 6833 -1620
rect 6799 -1719 6833 -1692
rect 6799 -1787 6833 -1753
rect 6799 -1855 6833 -1821
rect 6799 -1923 6833 -1889
rect 6799 -1991 6833 -1957
rect 6799 -2059 6833 -2025
rect 6799 -2109 6833 -2093
rect 6975 -1583 7009 -1567
rect 6975 -1651 7009 -1617
rect 6975 -1719 7009 -1685
rect 6975 -1787 7009 -1753
rect 6975 -1855 7009 -1821
rect 6975 -1923 7009 -1889
rect 6975 -1991 7009 -1957
rect 6975 -2059 7009 -2025
rect 6975 -2122 7009 -2093
rect 7151 -1583 7185 -1567
rect 7151 -1651 7185 -1620
rect 7151 -1719 7185 -1692
rect 7151 -1787 7185 -1753
rect 7151 -1855 7185 -1821
rect 7151 -1923 7185 -1889
rect 7151 -1991 7185 -1957
rect 7151 -2059 7185 -2025
rect 7151 -2109 7185 -2093
rect 7327 -1583 7361 -1567
rect 7327 -1651 7361 -1617
rect 7327 -1719 7361 -1685
rect 7327 -1787 7361 -1753
rect 7327 -1855 7361 -1821
rect 7327 -1923 7361 -1889
rect 7327 -1991 7361 -1957
rect 7327 -2059 7361 -2025
rect 7327 -2122 7361 -2093
rect 7503 -1583 7537 -1567
rect 7503 -1651 7537 -1620
rect 7503 -1719 7537 -1692
rect 7503 -1787 7537 -1753
rect 7503 -1855 7537 -1821
rect 7503 -1923 7537 -1889
rect 7503 -1991 7537 -1957
rect 7503 -2059 7537 -2025
rect 7503 -2109 7537 -2093
rect 7679 -1583 7713 -1567
rect 7679 -1651 7713 -1617
rect 7679 -1719 7713 -1685
rect 7679 -1787 7713 -1753
rect 7679 -1855 7713 -1821
rect 7679 -1923 7713 -1889
rect 7679 -1991 7713 -1957
rect 7679 -2059 7713 -2025
rect 7679 -2122 7713 -2093
rect 6632 -2156 6670 -2122
rect 6976 -2156 7014 -2122
rect 7330 -2156 7368 -2122
rect 7674 -2156 7712 -2122
<< viali >>
rect 4852 -413 4886 -379
rect 4732 -496 4766 -490
rect 4732 -524 4766 -496
rect 4732 -598 4766 -586
rect 4732 -620 4766 -598
rect 4924 -413 4958 -379
rect 5157 -413 5191 -379
rect 5229 -394 5263 -379
rect 5229 -413 5234 -394
rect 5234 -413 5263 -394
rect 5044 -496 5078 -490
rect 5044 -524 5078 -496
rect 5044 -598 5078 -586
rect 5044 -620 5078 -598
rect 5295 -496 5324 -465
rect 5324 -496 5329 -465
rect 5295 -499 5329 -496
rect 5367 -499 5401 -465
rect 5598 -499 5632 -465
rect 5670 -499 5704 -465
rect 5444 -576 5478 -542
rect 5516 -576 5550 -542
rect 5911 -499 5945 -465
rect 5983 -499 6017 -465
rect 5757 -654 5791 -620
rect 6037 -576 6071 -542
rect 6194 -413 6228 -379
rect 6266 -413 6300 -379
rect 6109 -576 6143 -542
rect 5829 -654 5863 -620
rect 5712 -777 5746 -743
rect 5712 -849 5746 -815
rect 5186 -943 5220 -909
rect 5258 -943 5292 -909
rect 5872 -777 5906 -743
rect 5872 -849 5906 -815
rect 7461 -353 7495 -319
rect 7533 -353 7567 -319
rect 6523 -413 6557 -379
rect 6595 -413 6629 -379
rect 7732 -446 7766 -412
rect 7732 -518 7766 -484
rect 6543 -557 6577 -523
rect 6615 -557 6649 -523
rect 6350 -654 6384 -620
rect 6422 -654 6456 -620
rect 6194 -867 6228 -833
rect 6266 -867 6300 -833
rect 7466 -679 7494 -649
rect 7494 -679 7500 -649
rect 7466 -683 7500 -679
rect 7538 -683 7572 -649
rect 6461 -867 6495 -833
rect 6533 -867 6567 -833
rect 6103 -943 6137 -909
rect 6175 -943 6209 -909
rect 7732 -774 7766 -740
rect 7732 -846 7766 -812
rect 7524 -1025 7558 -991
rect 7598 -1025 7632 -991
rect 7671 -1025 7705 -991
rect 7744 -1021 7770 -991
rect 7770 -1021 7778 -991
rect 7744 -1025 7778 -1021
rect 6267 -1340 6301 -1306
rect 6339 -1340 6373 -1306
rect 6445 -1253 6479 -1219
rect 6517 -1253 6551 -1219
rect 6736 -1350 6770 -1316
rect 6808 -1350 6842 -1316
rect 6691 -1423 6725 -1407
rect 6767 -1423 6801 -1407
rect 6843 -1423 6877 -1407
rect 6918 -1423 6952 -1407
rect 7570 -1247 7604 -1213
rect 7642 -1247 7676 -1213
rect 7395 -1423 7429 -1407
rect 7471 -1423 7505 -1407
rect 7547 -1423 7581 -1407
rect 7622 -1423 7656 -1407
rect 6691 -1441 6718 -1423
rect 6718 -1441 6725 -1423
rect 6767 -1441 6795 -1423
rect 6795 -1441 6801 -1423
rect 6843 -1441 6872 -1423
rect 6872 -1441 6877 -1423
rect 6918 -1441 6948 -1423
rect 6948 -1441 6952 -1423
rect 7395 -1441 7422 -1423
rect 7422 -1441 7429 -1423
rect 7471 -1441 7498 -1423
rect 7498 -1441 7505 -1423
rect 7547 -1441 7575 -1423
rect 7575 -1441 7581 -1423
rect 7622 -1441 7652 -1423
rect 7652 -1441 7656 -1423
rect 7080 -1521 7114 -1487
rect 7152 -1521 7186 -1487
rect 6331 -1593 6365 -1586
rect 6331 -1620 6365 -1593
rect 6447 -1617 6481 -1586
rect 6447 -1620 6481 -1617
rect 6331 -1661 6365 -1658
rect 6331 -1692 6365 -1661
rect 6447 -1685 6481 -1658
rect 6447 -1692 6481 -1685
rect 6799 -1617 6833 -1586
rect 6799 -1620 6833 -1617
rect 6799 -1685 6833 -1658
rect 6799 -1692 6833 -1685
rect 7151 -1617 7185 -1586
rect 7151 -1620 7185 -1617
rect 7151 -1685 7185 -1658
rect 7151 -1692 7185 -1685
rect 7503 -1617 7537 -1586
rect 7503 -1620 7537 -1617
rect 7503 -1685 7537 -1658
rect 7503 -1692 7537 -1685
rect 6598 -2156 6632 -2122
rect 6670 -2156 6704 -2122
rect 6942 -2156 6976 -2122
rect 7014 -2156 7048 -2122
rect 7296 -2156 7330 -2122
rect 7368 -2156 7402 -2122
rect 7640 -2156 7674 -2122
rect 7712 -2156 7746 -2122
<< metal1 >>
rect 7449 -319 7872 -313
rect 7449 -353 7461 -319
rect 7495 -353 7533 -319
rect 7567 -353 7820 -319
rect 7449 -359 7820 -353
tri 7773 -373 7787 -359 ne
rect 7787 -371 7820 -359
rect 7787 -373 7872 -371
rect 4840 -379 6313 -373
rect 6424 -379 6641 -373
rect 4840 -413 4852 -379
rect 4886 -413 4924 -379
rect 4958 -413 5157 -379
rect 5191 -413 5229 -379
rect 5263 -413 6194 -379
rect 6228 -413 6266 -379
rect 6300 -413 6313 -379
tri 6390 -413 6424 -379 se
rect 4840 -419 6313 -413
tri 6384 -419 6390 -413 se
rect 6390 -419 6424 -413
tri 6364 -439 6384 -419 se
rect 6384 -431 6424 -419
rect 6476 -413 6523 -379
rect 6557 -413 6595 -379
rect 6629 -413 6641 -379
tri 7787 -400 7814 -373 ne
rect 7814 -383 7872 -373
rect 7814 -400 7820 -383
rect 6476 -419 6641 -413
rect 7726 -412 7772 -400
tri 7814 -406 7820 -400 ne
rect 6476 -431 6489 -419
rect 6384 -439 6489 -431
tri 6489 -439 6509 -419 nw
tri 6357 -446 6364 -439 se
rect 6364 -441 6487 -439
tri 6487 -441 6489 -439 nw
rect 6364 -443 6482 -441
rect 6364 -446 6424 -443
tri 6344 -459 6357 -446 se
rect 6357 -459 6424 -446
rect 5283 -465 6424 -459
rect 4726 -490 5084 -478
rect 4726 -524 4732 -490
rect 4766 -524 5044 -490
rect 5078 -524 5084 -490
rect 5283 -499 5295 -465
rect 5329 -499 5367 -465
rect 5401 -499 5598 -465
rect 5632 -499 5670 -465
rect 5704 -499 5911 -465
rect 5945 -499 5983 -465
rect 6017 -495 6424 -465
rect 6476 -446 6482 -443
tri 6482 -446 6487 -441 nw
rect 7726 -446 7732 -412
rect 7766 -446 7772 -412
rect 7820 -441 7872 -435
tri 6476 -452 6482 -446 nw
rect 6017 -499 6476 -495
rect 5283 -501 6476 -499
rect 7726 -484 7772 -446
rect 5283 -505 6364 -501
tri 6364 -505 6368 -501 nw
rect 4726 -586 5084 -524
rect 6529 -523 6661 -517
rect 5432 -542 6155 -536
rect 5432 -576 5444 -542
rect 5478 -576 5516 -542
rect 5550 -576 6037 -542
rect 6071 -576 6109 -542
rect 6143 -576 6155 -542
rect 5432 -582 6155 -576
rect 6529 -557 6543 -523
rect 6577 -557 6587 -523
rect 6649 -557 6661 -523
rect 6529 -575 6587 -557
rect 6639 -575 6661 -557
rect 4726 -620 4732 -586
rect 4766 -620 5044 -586
rect 5078 -620 5084 -586
rect 6529 -587 6661 -575
rect 4726 -632 5084 -620
rect 5745 -620 6468 -614
rect 5745 -654 5757 -620
rect 5791 -654 5829 -620
rect 5863 -654 6350 -620
rect 6384 -654 6422 -620
rect 6456 -654 6468 -620
rect 5745 -660 6468 -654
rect 6529 -639 6587 -587
rect 6639 -623 6661 -587
rect 6529 -645 6639 -639
tri 6639 -645 6661 -623 nw
rect 7726 -518 7732 -484
rect 7766 -518 7772 -484
rect 6529 -649 6635 -645
tri 6635 -649 6639 -645 nw
rect 7454 -646 7584 -640
rect 7454 -649 7473 -646
rect 7525 -649 7584 -646
rect 6529 -660 6624 -649
tri 6624 -660 6635 -649 nw
rect 6529 -683 6601 -660
tri 6601 -683 6624 -660 nw
rect 7454 -683 7466 -649
rect 7525 -683 7538 -649
rect 7572 -683 7584 -649
rect 6529 -689 6595 -683
tri 6595 -689 6601 -683 nw
tri 6487 -731 6529 -689 se
rect 6529 -731 6553 -689
tri 6553 -731 6595 -689 nw
rect 7454 -698 7473 -683
rect 7525 -698 7584 -683
rect 7454 -710 7584 -698
rect 5706 -740 6544 -731
tri 6544 -740 6553 -731 nw
rect 5706 -743 6510 -740
rect 5706 -777 5712 -743
rect 5746 -777 5872 -743
rect 5906 -774 6510 -743
tri 6510 -774 6544 -740 nw
rect 7454 -762 7473 -710
rect 7525 -762 7584 -710
rect 7454 -768 7584 -762
rect 7726 -740 7772 -518
rect 7726 -774 7732 -740
rect 7766 -774 7772 -740
rect 5906 -777 6507 -774
tri 6507 -777 6510 -774 nw
rect 5706 -812 6061 -777
tri 6061 -812 6096 -777 nw
rect 7726 -812 7772 -774
rect 5706 -815 6040 -812
rect 5706 -849 5712 -815
rect 5746 -849 5872 -815
rect 5906 -833 6040 -815
tri 6040 -833 6061 -812 nw
rect 6182 -833 6579 -827
rect 5906 -849 6012 -833
rect 5706 -861 6012 -849
tri 6012 -861 6040 -833 nw
rect 6182 -867 6194 -833
rect 6228 -867 6266 -833
rect 6300 -867 6461 -833
rect 6495 -867 6533 -833
rect 6567 -867 6579 -833
rect 7726 -846 7732 -812
rect 7766 -846 7772 -812
rect 7726 -858 7772 -846
rect 6182 -873 6579 -867
rect 5174 -949 5180 -897
rect 5232 -949 5246 -897
rect 5298 -949 5304 -897
rect 6091 -909 6221 -903
rect 6091 -943 6103 -909
rect 6137 -943 6175 -909
rect 6209 -943 6221 -909
rect 6091 -949 6221 -943
rect 7512 -991 7790 -985
rect 7512 -1025 7524 -991
rect 7558 -1025 7598 -991
rect 7632 -1025 7671 -991
rect 7705 -1025 7744 -991
rect 7778 -1025 7790 -991
rect 7512 -1031 7790 -1025
tri 6695 -1211 6699 -1207 se
rect 6699 -1211 7688 -1207
rect 5399 -1263 5405 -1211
rect 5457 -1263 5469 -1211
rect 5521 -1219 6563 -1211
tri 6693 -1213 6695 -1211 se
rect 6695 -1213 7688 -1211
rect 5521 -1253 6445 -1219
rect 6479 -1253 6517 -1219
rect 6551 -1253 6563 -1219
tri 6659 -1247 6693 -1213 se
rect 6693 -1247 7570 -1213
rect 7604 -1247 7642 -1213
rect 7676 -1247 7688 -1213
rect 5521 -1263 6563 -1253
tri 6643 -1263 6659 -1247 se
rect 6659 -1253 7688 -1247
tri 7795 -1253 7820 -1228 se
rect 7820 -1234 7872 -1228
rect 6659 -1263 6699 -1253
tri 6633 -1273 6643 -1263 se
rect 6643 -1273 6699 -1263
tri 6699 -1273 6719 -1253 nw
tri 7775 -1273 7795 -1253 se
rect 7795 -1273 7820 -1253
tri 6606 -1300 6633 -1273 se
rect 6633 -1300 6672 -1273
tri 6672 -1300 6699 -1273 nw
tri 7748 -1300 7775 -1273 se
rect 7775 -1286 7820 -1273
rect 7775 -1298 7872 -1286
rect 7775 -1300 7820 -1298
rect 6255 -1306 6656 -1300
rect 6255 -1340 6267 -1306
rect 6301 -1340 6339 -1306
rect 6373 -1316 6656 -1306
tri 6656 -1316 6672 -1300 nw
tri 7738 -1310 7748 -1300 se
rect 7748 -1310 7820 -1300
rect 6724 -1316 7820 -1310
rect 6373 -1340 6626 -1316
rect 6255 -1346 6626 -1340
tri 6626 -1346 6656 -1316 nw
rect 6724 -1350 6736 -1316
rect 6770 -1350 6808 -1316
rect 6842 -1350 7820 -1316
rect 6724 -1356 7872 -1350
rect 6587 -1447 6593 -1395
rect 6645 -1447 6657 -1395
rect 6709 -1401 6715 -1395
tri 6715 -1401 6721 -1395 sw
rect 6709 -1407 7668 -1401
rect 6725 -1441 6767 -1407
rect 6801 -1441 6843 -1407
rect 6877 -1441 6918 -1407
rect 6952 -1441 7395 -1407
rect 7429 -1441 7471 -1407
rect 7505 -1441 7547 -1407
rect 7581 -1441 7622 -1407
rect 7656 -1441 7668 -1407
rect 6709 -1447 7668 -1441
rect 7068 -1487 7198 -1481
rect 7068 -1521 7080 -1487
rect 7114 -1521 7152 -1487
rect 7186 -1521 7198 -1487
rect 7068 -1527 7198 -1521
rect 6325 -1586 6371 -1574
rect 6325 -1620 6331 -1586
rect 6365 -1620 6371 -1586
rect 6325 -1658 6371 -1620
rect 6325 -1692 6331 -1658
rect 6365 -1692 6371 -1658
rect 6325 -1704 6371 -1692
rect 6441 -1586 7543 -1574
rect 6441 -1620 6447 -1586
rect 6481 -1620 6799 -1586
rect 6833 -1620 7151 -1586
rect 7185 -1620 7503 -1586
rect 7537 -1620 7543 -1586
rect 6441 -1658 7543 -1620
rect 6441 -1692 6447 -1658
rect 6481 -1692 6799 -1658
rect 6833 -1692 7151 -1658
rect 7185 -1692 7503 -1658
rect 7537 -1692 7543 -1658
rect 6441 -1704 7543 -1692
rect 6476 -2162 6482 -2110
rect 6534 -2162 6546 -2110
rect 6598 -2116 6604 -2110
tri 7410 -2116 7416 -2110 se
rect 7416 -2116 7422 -2110
rect 6598 -2122 7060 -2116
rect 6632 -2156 6670 -2122
rect 6704 -2156 6942 -2122
rect 6976 -2156 7014 -2122
rect 7048 -2156 7060 -2122
rect 6598 -2162 7060 -2156
rect 7284 -2122 7422 -2116
rect 7284 -2156 7296 -2122
rect 7330 -2156 7368 -2122
rect 7402 -2156 7422 -2122
rect 7284 -2162 7422 -2156
rect 7474 -2162 7486 -2110
rect 7538 -2116 7544 -2110
tri 7544 -2116 7550 -2110 sw
rect 7538 -2122 7758 -2116
rect 7538 -2156 7640 -2122
rect 7674 -2156 7712 -2122
rect 7746 -2156 7758 -2122
rect 7538 -2162 7758 -2156
<< via1 >>
rect 7820 -371 7872 -319
rect 6424 -431 6476 -379
rect 6424 -495 6476 -443
rect 7820 -435 7872 -383
rect 6587 -557 6615 -523
rect 6615 -557 6639 -523
rect 6587 -575 6639 -557
rect 6587 -639 6639 -587
rect 7473 -649 7525 -646
rect 7473 -683 7500 -649
rect 7500 -683 7525 -649
rect 7473 -698 7525 -683
rect 7473 -762 7525 -710
rect 5180 -909 5232 -897
rect 5180 -943 5186 -909
rect 5186 -943 5220 -909
rect 5220 -943 5232 -909
rect 5180 -949 5232 -943
rect 5246 -909 5298 -897
rect 5246 -943 5258 -909
rect 5258 -943 5292 -909
rect 5292 -943 5298 -909
rect 5246 -949 5298 -943
rect 5405 -1263 5457 -1211
rect 5469 -1263 5521 -1211
rect 7820 -1286 7872 -1234
rect 7820 -1350 7872 -1298
rect 6593 -1447 6645 -1395
rect 6657 -1407 6709 -1395
rect 6657 -1441 6691 -1407
rect 6691 -1441 6709 -1407
rect 6657 -1447 6709 -1441
rect 6482 -2162 6534 -2110
rect 6546 -2162 6598 -2110
rect 7422 -2162 7474 -2110
rect 7486 -2162 7538 -2110
<< metal2 >>
rect 7820 -319 7872 -313
rect 6424 -379 6476 -373
rect 6424 -443 6476 -431
rect 6424 -501 6476 -495
tri 6424 -507 6430 -501 ne
rect 5174 -949 5180 -897
rect 5232 -949 5246 -897
rect 5298 -949 5349 -897
tri 5349 -949 5401 -897 sw
tri 5327 -952 5330 -949 ne
rect 5330 -952 5401 -949
tri 5401 -952 5404 -949 sw
tri 5330 -971 5349 -952 ne
rect 5349 -971 5404 -952
tri 5349 -1026 5404 -971 ne
tri 5404 -1026 5478 -952 sw
tri 5404 -1048 5426 -1026 ne
tri 5399 -1211 5426 -1184 se
rect 5426 -1211 5478 -1026
tri 5478 -1211 5505 -1184 sw
rect 5399 -1263 5405 -1211
rect 5457 -1263 5469 -1211
rect 5521 -1263 5527 -1211
rect 6430 -2070 6476 -501
rect 7820 -383 7872 -371
rect 6587 -523 6639 -517
rect 6587 -587 6639 -575
rect 6587 -645 6639 -639
rect 6587 -646 6638 -645
tri 6638 -646 6639 -645 nw
rect 7473 -646 7525 -640
rect 6587 -1350 6633 -646
tri 6633 -651 6638 -646 nw
rect 7473 -710 7525 -698
rect 7473 -768 7525 -762
tri 7473 -787 7492 -768 ne
tri 6633 -1350 6670 -1313 sw
rect 6587 -1395 6670 -1350
tri 6670 -1395 6715 -1350 sw
rect 6587 -1447 6593 -1395
rect 6645 -1447 6657 -1395
rect 6709 -1447 6715 -1395
tri 6476 -2070 6485 -2061 sw
rect 6430 -2081 6485 -2070
tri 6430 -2110 6459 -2081 ne
rect 6459 -2110 6485 -2081
tri 6485 -2110 6525 -2070 sw
tri 7452 -2110 7492 -2070 se
rect 7492 -2110 7525 -768
rect 7820 -1234 7872 -435
rect 7820 -1298 7872 -1286
rect 7820 -1356 7872 -1350
tri 7525 -2110 7544 -2091 sw
tri 6459 -2127 6476 -2110 ne
rect 6476 -2162 6482 -2110
rect 6534 -2162 6546 -2110
rect 6598 -2162 6604 -2110
rect 7416 -2162 7422 -2110
rect 7474 -2162 7486 -2110
rect 7538 -2162 7544 -2110
use sky130_fd_pr__nfet_01v8__example_55959141808116  sky130_fd_pr__nfet_01v8__example_55959141808116_0
timestamp 1644511149
transform -1 0 7140 0 1 -2105
box -28 0 148 267
use sky130_fd_pr__nfet_01v8__example_55959141808116  sky130_fd_pr__nfet_01v8__example_55959141808116_1
timestamp 1644511149
transform 1 0 7196 0 1 -2105
box -28 0 148 267
use sky130_fd_pr__nfet_01v8__example_55959141808116  sky130_fd_pr__nfet_01v8__example_55959141808116_2
timestamp 1644511149
transform 1 0 6492 0 1 -2105
box -28 0 148 267
use sky130_fd_pr__nfet_01v8__example_55959141808631  sky130_fd_pr__nfet_01v8__example_55959141808631_0
timestamp 1644511149
transform 1 0 7372 0 1 -2105
box -28 0 324 267
use sky130_fd_pr__nfet_01v8__example_55959141808631  sky130_fd_pr__nfet_01v8__example_55959141808631_1
timestamp 1644511149
transform -1 0 6964 0 1 -2105
box -28 0 324 267
use sky130_fd_pr__pfet_01v8__example_55959141808354  sky130_fd_pr__pfet_01v8__example_55959141808354_0
timestamp 1644511149
transform 1 0 6649 0 1 -1111
box -28 0 828 29
use sky130_fd_pr__pfet_01v8__example_55959141808354  sky130_fd_pr__pfet_01v8__example_55959141808354_1
timestamp 1644511149
transform -1 0 7449 0 1 -477
box -28 0 828 29
use sky130_fd_pr__pfet_01v8__example_55959141808354  sky130_fd_pr__pfet_01v8__example_55959141808354_2
timestamp 1644511149
transform 1 0 6649 0 1 -1327
box -28 0 828 29
use sky130_fd_pr__pfet_01v8__example_55959141808626  sky130_fd_pr__pfet_01v8__example_55959141808626_0
timestamp 1644511149
transform 1 0 5369 0 -1 -314
box -28 0 284 267
use sky130_fd_pr__pfet_01v8__example_55959141808626  sky130_fd_pr__pfet_01v8__example_55959141808626_1
timestamp 1644511149
transform 1 0 5681 0 -1 -314
box -28 0 284 267
use sky130_fd_pr__pfet_01v8__example_55959141808627  sky130_fd_pr__pfet_01v8__example_55959141808627_0
timestamp 1644511149
transform 1 0 4777 0 -1 -314
box -28 0 440 267
use sky130_fd_pr__pfet_01v8__example_55959141808628  sky130_fd_pr__pfet_01v8__example_55959141808628_0
timestamp 1644511149
transform -1 0 6217 0 -1 -314
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808628  sky130_fd_pr__pfet_01v8__example_55959141808628_1
timestamp 1644511149
transform 1 0 6273 0 -1 -314
box -28 0 128 267
use sky130_fd_pr__pfet_01v8__example_55959141808629  sky130_fd_pr__pfet_01v8__example_55959141808629_0
timestamp 1644511149
transform 0 1 7724 -1 0 -652
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808629  sky130_fd_pr__pfet_01v8__example_55959141808629_1
timestamp 1644511149
transform 0 1 7724 1 0 -596
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808629  sky130_fd_pr__pfet_01v8__example_55959141808629_2
timestamp 1644511149
transform 0 1 7724 -1 0 -1032
box -28 0 228 29
use sky130_fd_pr__pfet_01v8__example_55959141808630  sky130_fd_pr__pfet_01v8__example_55959141808630_0
timestamp 1644511149
transform -1 0 7449 0 -1 -801
box -28 0 828 29
use sky130_fd_pr__pfet_01v8__example_55959141808630  sky130_fd_pr__pfet_01v8__example_55959141808630_1
timestamp 1644511149
transform 1 0 6649 0 1 -691
box -28 0 828 29
<< labels >>
flabel metal1 s 6890 -1437 6918 -1409 3 FreeSans 280 0 0 0 DRVLO_H_N
port 1 nsew
flabel metal1 s 7330 -2152 7358 -2124 3 FreeSans 280 0 0 0 PD_I2C_H
port 2 nsew
flabel metal1 s 7108 -1514 7136 -1486 3 FreeSans 280 0 0 0 PDEN_H_N
port 3 nsew
flabel metal1 s 6978 -2151 7006 -2123 3 FreeSans 280 0 0 0 PD_H
port 4 nsew
flabel metal1 s 7576 -1019 7604 -991 3 FreeSans 280 0 0 0 VCC_IO
port 5 nsew
flabel metal1 s 6488 -1253 6516 -1225 3 FreeSans 280 180 0 0 I2C_MODE_H
port 6 nsew
flabel metal1 s 7066 -1651 7094 -1623 3 FreeSans 280 0 0 0 VGND_IO
port 7 nsew
flabel metal1 s 6169 -941 6197 -913 3 FreeSans 280 0 0 0 EN_FAST_N[0]
port 8 nsew
flabel metal1 s 7590 -1243 7618 -1215 3 FreeSans 280 0 0 0 EN_FAST_N[1]
port 9 nsew
flabel metal1 s 4869 -554 4897 -526 3 FreeSans 280 0 0 0 VCC_IO
port 5 nsew
flabel comment s 6823 -2142 6823 -2142 0 FreeSans 440 0 0 0 PD_H
flabel comment s 7498 -2142 7498 -2142 0 FreeSans 440 0 0 0 PD_I2C_H
<< properties >>
string GDS_END 7485436
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7455964
<< end >>
