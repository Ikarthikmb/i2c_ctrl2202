/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/sky130A/libs.tech/ngspice/capacitors/sky130_fd_pr__model__cap_mim.model.spice