/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/rf_pfet_01v8/sky130_fd_pr__rf_pfet_01v8_bM02W5p00L0p25.spice