magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< dnwell >>
rect 88 579 15088 5356
<< nwell >>
rect -36 5150 15191 5489
rect -36 785 469 5150
rect 14753 785 15191 5150
rect -36 423 15191 785
<< pwell >>
rect 529 4760 14693 4982
rect 529 4084 751 4760
rect 14471 4084 14693 4760
rect 529 3032 14693 4084
rect 529 2483 751 3032
rect 1552 2483 1840 3032
rect 2544 2483 2832 3032
rect 3536 2483 3824 3032
rect 4528 2483 4816 3032
rect 5520 2483 5808 3032
rect 6512 2483 6800 3032
rect 7504 2483 7792 3032
rect 8496 2483 8784 3032
rect 9488 2483 9776 3032
rect 10480 2483 10768 3032
rect 11472 2483 11760 3032
rect 12464 2483 12752 3032
rect 13456 2483 13744 3032
rect 14471 2483 14693 3032
rect 529 1431 14693 2483
rect 529 1174 751 1431
rect 14471 1174 14693 1431
rect 529 952 14693 1174
<< mvnmos >>
rect 924 3058 1044 4058
rect 1354 3058 1474 4058
rect 1916 3058 2036 4058
rect 2346 3058 2466 4058
rect 2908 3058 3028 4058
rect 3338 3058 3458 4058
rect 3900 3058 4020 4058
rect 4330 3058 4450 4058
rect 4892 3058 5012 4058
rect 5322 3058 5442 4058
rect 5884 3058 6004 4058
rect 6314 3058 6434 4058
rect 6876 3058 6996 4058
rect 7306 3058 7426 4058
rect 7868 3058 7988 4058
rect 8298 3058 8418 4058
rect 8860 3058 8980 4058
rect 9290 3058 9410 4058
rect 9852 3058 9972 4058
rect 10282 3058 10402 4058
rect 10844 3058 10964 4058
rect 11274 3058 11394 4058
rect 11836 3058 11956 4058
rect 12266 3058 12386 4058
rect 12828 3058 12948 4058
rect 13258 3058 13378 4058
rect 13820 3058 13940 4058
rect 14178 3058 14298 4058
rect 924 1457 1044 2457
rect 1354 1457 1474 2457
rect 1916 1457 2036 2457
rect 2346 1457 2466 2457
rect 2908 1457 3028 2457
rect 3338 1457 3458 2457
rect 3900 1457 4020 2457
rect 4330 1457 4450 2457
rect 4892 1457 5012 2457
rect 5322 1457 5442 2457
rect 5884 1457 6004 2457
rect 6314 1457 6434 2457
rect 6876 1457 6996 2457
rect 7306 1457 7426 2457
rect 7868 1457 7988 2457
rect 8298 1457 8418 2457
rect 8860 1457 8980 2457
rect 9290 1457 9410 2457
rect 9852 1457 9972 2457
rect 10282 1457 10402 2457
rect 10844 1457 10964 2457
rect 11274 1457 11394 2457
rect 11836 1457 11956 2457
rect 12266 1457 12386 2457
rect 12828 1457 12948 2457
rect 13258 1457 13378 2457
rect 13820 1457 13940 2457
rect 14178 1457 14298 2457
<< mvndiff >>
rect 787 4046 924 4058
rect 787 4012 802 4046
rect 836 4012 924 4046
rect 787 3978 924 4012
rect 787 3944 802 3978
rect 836 3944 924 3978
rect 787 3910 924 3944
rect 787 3876 802 3910
rect 836 3876 924 3910
rect 787 3842 924 3876
rect 787 3808 802 3842
rect 836 3808 924 3842
rect 787 3774 924 3808
rect 787 3740 802 3774
rect 836 3740 924 3774
rect 787 3706 924 3740
rect 787 3672 802 3706
rect 836 3672 924 3706
rect 787 3638 924 3672
rect 787 3604 802 3638
rect 836 3604 924 3638
rect 787 3570 924 3604
rect 787 3536 802 3570
rect 836 3536 924 3570
rect 787 3502 924 3536
rect 787 3468 802 3502
rect 836 3468 924 3502
rect 787 3434 924 3468
rect 787 3400 802 3434
rect 836 3400 924 3434
rect 787 3366 924 3400
rect 787 3332 802 3366
rect 836 3332 924 3366
rect 787 3298 924 3332
rect 787 3264 802 3298
rect 836 3264 924 3298
rect 787 3230 924 3264
rect 787 3196 802 3230
rect 836 3196 924 3230
rect 787 3162 924 3196
rect 787 3128 802 3162
rect 836 3128 924 3162
rect 787 3058 924 3128
rect 1044 4046 1354 4058
rect 1044 4012 1146 4046
rect 1180 4012 1218 4046
rect 1252 4012 1354 4046
rect 1044 3978 1354 4012
rect 1044 3944 1146 3978
rect 1180 3944 1218 3978
rect 1252 3944 1354 3978
rect 1044 3910 1354 3944
rect 1044 3876 1146 3910
rect 1180 3876 1218 3910
rect 1252 3876 1354 3910
rect 1044 3842 1354 3876
rect 1044 3808 1146 3842
rect 1180 3808 1218 3842
rect 1252 3808 1354 3842
rect 1044 3774 1354 3808
rect 1044 3740 1146 3774
rect 1180 3740 1218 3774
rect 1252 3740 1354 3774
rect 1044 3706 1354 3740
rect 1044 3672 1146 3706
rect 1180 3672 1218 3706
rect 1252 3672 1354 3706
rect 1044 3638 1354 3672
rect 1044 3604 1146 3638
rect 1180 3604 1218 3638
rect 1252 3604 1354 3638
rect 1044 3570 1354 3604
rect 1044 3536 1146 3570
rect 1180 3536 1218 3570
rect 1252 3536 1354 3570
rect 1044 3502 1354 3536
rect 1044 3468 1146 3502
rect 1180 3468 1218 3502
rect 1252 3468 1354 3502
rect 1044 3434 1354 3468
rect 1044 3400 1146 3434
rect 1180 3400 1218 3434
rect 1252 3400 1354 3434
rect 1044 3366 1354 3400
rect 1044 3332 1146 3366
rect 1180 3332 1218 3366
rect 1252 3332 1354 3366
rect 1044 3298 1354 3332
rect 1044 3264 1146 3298
rect 1180 3264 1218 3298
rect 1252 3264 1354 3298
rect 1044 3230 1354 3264
rect 1044 3196 1146 3230
rect 1180 3196 1218 3230
rect 1252 3196 1354 3230
rect 1044 3162 1354 3196
rect 1044 3128 1146 3162
rect 1180 3128 1218 3162
rect 1252 3128 1354 3162
rect 1044 3058 1354 3128
rect 1474 4046 1625 4058
rect 1765 4046 1916 4058
rect 1474 4012 1576 4046
rect 1610 4012 1625 4046
rect 1765 4012 1780 4046
rect 1814 4012 1916 4046
rect 1474 3978 1625 4012
rect 1765 3978 1916 4012
rect 1474 3944 1576 3978
rect 1610 3944 1625 3978
rect 1765 3944 1780 3978
rect 1814 3944 1916 3978
rect 1474 3910 1625 3944
rect 1765 3910 1916 3944
rect 1474 3876 1576 3910
rect 1610 3876 1625 3910
rect 1765 3876 1780 3910
rect 1814 3876 1916 3910
rect 1474 3842 1625 3876
rect 1765 3842 1916 3876
rect 1474 3808 1576 3842
rect 1610 3808 1625 3842
rect 1765 3808 1780 3842
rect 1814 3808 1916 3842
rect 1474 3774 1625 3808
rect 1765 3774 1916 3808
rect 1474 3740 1576 3774
rect 1610 3740 1625 3774
rect 1765 3740 1780 3774
rect 1814 3740 1916 3774
rect 1474 3706 1625 3740
rect 1765 3706 1916 3740
rect 1474 3672 1576 3706
rect 1610 3672 1625 3706
rect 1765 3672 1780 3706
rect 1814 3672 1916 3706
rect 1474 3638 1625 3672
rect 1765 3638 1916 3672
rect 1474 3604 1576 3638
rect 1610 3604 1625 3638
rect 1765 3604 1780 3638
rect 1814 3604 1916 3638
rect 1474 3570 1625 3604
rect 1765 3570 1916 3604
rect 1474 3536 1576 3570
rect 1610 3536 1625 3570
rect 1765 3536 1780 3570
rect 1814 3536 1916 3570
rect 1474 3502 1625 3536
rect 1765 3502 1916 3536
rect 1474 3468 1576 3502
rect 1610 3468 1625 3502
rect 1765 3468 1780 3502
rect 1814 3468 1916 3502
rect 1474 3434 1625 3468
rect 1765 3434 1916 3468
rect 1474 3400 1576 3434
rect 1610 3400 1625 3434
rect 1765 3400 1780 3434
rect 1814 3400 1916 3434
rect 1474 3366 1625 3400
rect 1765 3366 1916 3400
rect 1474 3332 1576 3366
rect 1610 3332 1625 3366
rect 1765 3332 1780 3366
rect 1814 3332 1916 3366
rect 1474 3298 1625 3332
rect 1765 3298 1916 3332
rect 1474 3264 1576 3298
rect 1610 3264 1625 3298
rect 1765 3264 1780 3298
rect 1814 3264 1916 3298
rect 1474 3230 1625 3264
rect 1765 3230 1916 3264
rect 1474 3196 1576 3230
rect 1610 3196 1625 3230
rect 1765 3196 1780 3230
rect 1814 3196 1916 3230
rect 1474 3162 1625 3196
rect 1765 3162 1916 3196
rect 1474 3128 1576 3162
rect 1610 3128 1625 3162
rect 1765 3128 1780 3162
rect 1814 3128 1916 3162
rect 1474 3058 1625 3128
rect 1765 3058 1916 3128
rect 2036 4046 2346 4058
rect 2036 4012 2138 4046
rect 2172 4012 2210 4046
rect 2244 4012 2346 4046
rect 2036 3978 2346 4012
rect 2036 3944 2138 3978
rect 2172 3944 2210 3978
rect 2244 3944 2346 3978
rect 2036 3910 2346 3944
rect 2036 3876 2138 3910
rect 2172 3876 2210 3910
rect 2244 3876 2346 3910
rect 2036 3842 2346 3876
rect 2036 3808 2138 3842
rect 2172 3808 2210 3842
rect 2244 3808 2346 3842
rect 2036 3774 2346 3808
rect 2036 3740 2138 3774
rect 2172 3740 2210 3774
rect 2244 3740 2346 3774
rect 2036 3706 2346 3740
rect 2036 3672 2138 3706
rect 2172 3672 2210 3706
rect 2244 3672 2346 3706
rect 2036 3638 2346 3672
rect 2036 3604 2138 3638
rect 2172 3604 2210 3638
rect 2244 3604 2346 3638
rect 2036 3570 2346 3604
rect 2036 3536 2138 3570
rect 2172 3536 2210 3570
rect 2244 3536 2346 3570
rect 2036 3502 2346 3536
rect 2036 3468 2138 3502
rect 2172 3468 2210 3502
rect 2244 3468 2346 3502
rect 2036 3434 2346 3468
rect 2036 3400 2138 3434
rect 2172 3400 2210 3434
rect 2244 3400 2346 3434
rect 2036 3366 2346 3400
rect 2036 3332 2138 3366
rect 2172 3332 2210 3366
rect 2244 3332 2346 3366
rect 2036 3298 2346 3332
rect 2036 3264 2138 3298
rect 2172 3264 2210 3298
rect 2244 3264 2346 3298
rect 2036 3230 2346 3264
rect 2036 3196 2138 3230
rect 2172 3196 2210 3230
rect 2244 3196 2346 3230
rect 2036 3162 2346 3196
rect 2036 3128 2138 3162
rect 2172 3128 2210 3162
rect 2244 3128 2346 3162
rect 2036 3058 2346 3128
rect 2466 4046 2617 4058
rect 2757 4046 2908 4058
rect 2466 4012 2568 4046
rect 2602 4012 2617 4046
rect 2757 4012 2772 4046
rect 2806 4012 2908 4046
rect 2466 3978 2617 4012
rect 2757 3978 2908 4012
rect 2466 3944 2568 3978
rect 2602 3944 2617 3978
rect 2757 3944 2772 3978
rect 2806 3944 2908 3978
rect 2466 3910 2617 3944
rect 2757 3910 2908 3944
rect 2466 3876 2568 3910
rect 2602 3876 2617 3910
rect 2757 3876 2772 3910
rect 2806 3876 2908 3910
rect 2466 3842 2617 3876
rect 2757 3842 2908 3876
rect 2466 3808 2568 3842
rect 2602 3808 2617 3842
rect 2757 3808 2772 3842
rect 2806 3808 2908 3842
rect 2466 3774 2617 3808
rect 2757 3774 2908 3808
rect 2466 3740 2568 3774
rect 2602 3740 2617 3774
rect 2757 3740 2772 3774
rect 2806 3740 2908 3774
rect 2466 3706 2617 3740
rect 2757 3706 2908 3740
rect 2466 3672 2568 3706
rect 2602 3672 2617 3706
rect 2757 3672 2772 3706
rect 2806 3672 2908 3706
rect 2466 3638 2617 3672
rect 2757 3638 2908 3672
rect 2466 3604 2568 3638
rect 2602 3604 2617 3638
rect 2757 3604 2772 3638
rect 2806 3604 2908 3638
rect 2466 3570 2617 3604
rect 2757 3570 2908 3604
rect 2466 3536 2568 3570
rect 2602 3536 2617 3570
rect 2757 3536 2772 3570
rect 2806 3536 2908 3570
rect 2466 3502 2617 3536
rect 2757 3502 2908 3536
rect 2466 3468 2568 3502
rect 2602 3468 2617 3502
rect 2757 3468 2772 3502
rect 2806 3468 2908 3502
rect 2466 3434 2617 3468
rect 2757 3434 2908 3468
rect 2466 3400 2568 3434
rect 2602 3400 2617 3434
rect 2757 3400 2772 3434
rect 2806 3400 2908 3434
rect 2466 3366 2617 3400
rect 2757 3366 2908 3400
rect 2466 3332 2568 3366
rect 2602 3332 2617 3366
rect 2757 3332 2772 3366
rect 2806 3332 2908 3366
rect 2466 3298 2617 3332
rect 2757 3298 2908 3332
rect 2466 3264 2568 3298
rect 2602 3264 2617 3298
rect 2757 3264 2772 3298
rect 2806 3264 2908 3298
rect 2466 3230 2617 3264
rect 2757 3230 2908 3264
rect 2466 3196 2568 3230
rect 2602 3196 2617 3230
rect 2757 3196 2772 3230
rect 2806 3196 2908 3230
rect 2466 3162 2617 3196
rect 2757 3162 2908 3196
rect 2466 3128 2568 3162
rect 2602 3128 2617 3162
rect 2757 3128 2772 3162
rect 2806 3128 2908 3162
rect 2466 3058 2617 3128
rect 2757 3058 2908 3128
rect 3028 4046 3338 4058
rect 3028 4012 3130 4046
rect 3164 4012 3202 4046
rect 3236 4012 3338 4046
rect 3028 3978 3338 4012
rect 3028 3944 3130 3978
rect 3164 3944 3202 3978
rect 3236 3944 3338 3978
rect 3028 3910 3338 3944
rect 3028 3876 3130 3910
rect 3164 3876 3202 3910
rect 3236 3876 3338 3910
rect 3028 3842 3338 3876
rect 3028 3808 3130 3842
rect 3164 3808 3202 3842
rect 3236 3808 3338 3842
rect 3028 3774 3338 3808
rect 3028 3740 3130 3774
rect 3164 3740 3202 3774
rect 3236 3740 3338 3774
rect 3028 3706 3338 3740
rect 3028 3672 3130 3706
rect 3164 3672 3202 3706
rect 3236 3672 3338 3706
rect 3028 3638 3338 3672
rect 3028 3604 3130 3638
rect 3164 3604 3202 3638
rect 3236 3604 3338 3638
rect 3028 3570 3338 3604
rect 3028 3536 3130 3570
rect 3164 3536 3202 3570
rect 3236 3536 3338 3570
rect 3028 3502 3338 3536
rect 3028 3468 3130 3502
rect 3164 3468 3202 3502
rect 3236 3468 3338 3502
rect 3028 3434 3338 3468
rect 3028 3400 3130 3434
rect 3164 3400 3202 3434
rect 3236 3400 3338 3434
rect 3028 3366 3338 3400
rect 3028 3332 3130 3366
rect 3164 3332 3202 3366
rect 3236 3332 3338 3366
rect 3028 3298 3338 3332
rect 3028 3264 3130 3298
rect 3164 3264 3202 3298
rect 3236 3264 3338 3298
rect 3028 3230 3338 3264
rect 3028 3196 3130 3230
rect 3164 3196 3202 3230
rect 3236 3196 3338 3230
rect 3028 3162 3338 3196
rect 3028 3128 3130 3162
rect 3164 3128 3202 3162
rect 3236 3128 3338 3162
rect 3028 3058 3338 3128
rect 3458 4046 3609 4058
rect 3749 4046 3900 4058
rect 3458 4012 3560 4046
rect 3594 4012 3609 4046
rect 3749 4012 3764 4046
rect 3798 4012 3900 4046
rect 3458 3978 3609 4012
rect 3749 3978 3900 4012
rect 3458 3944 3560 3978
rect 3594 3944 3609 3978
rect 3749 3944 3764 3978
rect 3798 3944 3900 3978
rect 3458 3910 3609 3944
rect 3749 3910 3900 3944
rect 3458 3876 3560 3910
rect 3594 3876 3609 3910
rect 3749 3876 3764 3910
rect 3798 3876 3900 3910
rect 3458 3842 3609 3876
rect 3749 3842 3900 3876
rect 3458 3808 3560 3842
rect 3594 3808 3609 3842
rect 3749 3808 3764 3842
rect 3798 3808 3900 3842
rect 3458 3774 3609 3808
rect 3749 3774 3900 3808
rect 3458 3740 3560 3774
rect 3594 3740 3609 3774
rect 3749 3740 3764 3774
rect 3798 3740 3900 3774
rect 3458 3706 3609 3740
rect 3749 3706 3900 3740
rect 3458 3672 3560 3706
rect 3594 3672 3609 3706
rect 3749 3672 3764 3706
rect 3798 3672 3900 3706
rect 3458 3638 3609 3672
rect 3749 3638 3900 3672
rect 3458 3604 3560 3638
rect 3594 3604 3609 3638
rect 3749 3604 3764 3638
rect 3798 3604 3900 3638
rect 3458 3570 3609 3604
rect 3749 3570 3900 3604
rect 3458 3536 3560 3570
rect 3594 3536 3609 3570
rect 3749 3536 3764 3570
rect 3798 3536 3900 3570
rect 3458 3502 3609 3536
rect 3749 3502 3900 3536
rect 3458 3468 3560 3502
rect 3594 3468 3609 3502
rect 3749 3468 3764 3502
rect 3798 3468 3900 3502
rect 3458 3434 3609 3468
rect 3749 3434 3900 3468
rect 3458 3400 3560 3434
rect 3594 3400 3609 3434
rect 3749 3400 3764 3434
rect 3798 3400 3900 3434
rect 3458 3366 3609 3400
rect 3749 3366 3900 3400
rect 3458 3332 3560 3366
rect 3594 3332 3609 3366
rect 3749 3332 3764 3366
rect 3798 3332 3900 3366
rect 3458 3298 3609 3332
rect 3749 3298 3900 3332
rect 3458 3264 3560 3298
rect 3594 3264 3609 3298
rect 3749 3264 3764 3298
rect 3798 3264 3900 3298
rect 3458 3230 3609 3264
rect 3749 3230 3900 3264
rect 3458 3196 3560 3230
rect 3594 3196 3609 3230
rect 3749 3196 3764 3230
rect 3798 3196 3900 3230
rect 3458 3162 3609 3196
rect 3749 3162 3900 3196
rect 3458 3128 3560 3162
rect 3594 3128 3609 3162
rect 3749 3128 3764 3162
rect 3798 3128 3900 3162
rect 3458 3058 3609 3128
rect 3749 3058 3900 3128
rect 4020 4046 4330 4058
rect 4020 4012 4122 4046
rect 4156 4012 4194 4046
rect 4228 4012 4330 4046
rect 4020 3978 4330 4012
rect 4020 3944 4122 3978
rect 4156 3944 4194 3978
rect 4228 3944 4330 3978
rect 4020 3910 4330 3944
rect 4020 3876 4122 3910
rect 4156 3876 4194 3910
rect 4228 3876 4330 3910
rect 4020 3842 4330 3876
rect 4020 3808 4122 3842
rect 4156 3808 4194 3842
rect 4228 3808 4330 3842
rect 4020 3774 4330 3808
rect 4020 3740 4122 3774
rect 4156 3740 4194 3774
rect 4228 3740 4330 3774
rect 4020 3706 4330 3740
rect 4020 3672 4122 3706
rect 4156 3672 4194 3706
rect 4228 3672 4330 3706
rect 4020 3638 4330 3672
rect 4020 3604 4122 3638
rect 4156 3604 4194 3638
rect 4228 3604 4330 3638
rect 4020 3570 4330 3604
rect 4020 3536 4122 3570
rect 4156 3536 4194 3570
rect 4228 3536 4330 3570
rect 4020 3502 4330 3536
rect 4020 3468 4122 3502
rect 4156 3468 4194 3502
rect 4228 3468 4330 3502
rect 4020 3434 4330 3468
rect 4020 3400 4122 3434
rect 4156 3400 4194 3434
rect 4228 3400 4330 3434
rect 4020 3366 4330 3400
rect 4020 3332 4122 3366
rect 4156 3332 4194 3366
rect 4228 3332 4330 3366
rect 4020 3298 4330 3332
rect 4020 3264 4122 3298
rect 4156 3264 4194 3298
rect 4228 3264 4330 3298
rect 4020 3230 4330 3264
rect 4020 3196 4122 3230
rect 4156 3196 4194 3230
rect 4228 3196 4330 3230
rect 4020 3162 4330 3196
rect 4020 3128 4122 3162
rect 4156 3128 4194 3162
rect 4228 3128 4330 3162
rect 4020 3058 4330 3128
rect 4450 4046 4601 4058
rect 4741 4046 4892 4058
rect 4450 4012 4552 4046
rect 4586 4012 4601 4046
rect 4741 4012 4756 4046
rect 4790 4012 4892 4046
rect 4450 3978 4601 4012
rect 4741 3978 4892 4012
rect 4450 3944 4552 3978
rect 4586 3944 4601 3978
rect 4741 3944 4756 3978
rect 4790 3944 4892 3978
rect 4450 3910 4601 3944
rect 4741 3910 4892 3944
rect 4450 3876 4552 3910
rect 4586 3876 4601 3910
rect 4741 3876 4756 3910
rect 4790 3876 4892 3910
rect 4450 3842 4601 3876
rect 4741 3842 4892 3876
rect 4450 3808 4552 3842
rect 4586 3808 4601 3842
rect 4741 3808 4756 3842
rect 4790 3808 4892 3842
rect 4450 3774 4601 3808
rect 4741 3774 4892 3808
rect 4450 3740 4552 3774
rect 4586 3740 4601 3774
rect 4741 3740 4756 3774
rect 4790 3740 4892 3774
rect 4450 3706 4601 3740
rect 4741 3706 4892 3740
rect 4450 3672 4552 3706
rect 4586 3672 4601 3706
rect 4741 3672 4756 3706
rect 4790 3672 4892 3706
rect 4450 3638 4601 3672
rect 4741 3638 4892 3672
rect 4450 3604 4552 3638
rect 4586 3604 4601 3638
rect 4741 3604 4756 3638
rect 4790 3604 4892 3638
rect 4450 3570 4601 3604
rect 4741 3570 4892 3604
rect 4450 3536 4552 3570
rect 4586 3536 4601 3570
rect 4741 3536 4756 3570
rect 4790 3536 4892 3570
rect 4450 3502 4601 3536
rect 4741 3502 4892 3536
rect 4450 3468 4552 3502
rect 4586 3468 4601 3502
rect 4741 3468 4756 3502
rect 4790 3468 4892 3502
rect 4450 3434 4601 3468
rect 4741 3434 4892 3468
rect 4450 3400 4552 3434
rect 4586 3400 4601 3434
rect 4741 3400 4756 3434
rect 4790 3400 4892 3434
rect 4450 3366 4601 3400
rect 4741 3366 4892 3400
rect 4450 3332 4552 3366
rect 4586 3332 4601 3366
rect 4741 3332 4756 3366
rect 4790 3332 4892 3366
rect 4450 3298 4601 3332
rect 4741 3298 4892 3332
rect 4450 3264 4552 3298
rect 4586 3264 4601 3298
rect 4741 3264 4756 3298
rect 4790 3264 4892 3298
rect 4450 3230 4601 3264
rect 4741 3230 4892 3264
rect 4450 3196 4552 3230
rect 4586 3196 4601 3230
rect 4741 3196 4756 3230
rect 4790 3196 4892 3230
rect 4450 3162 4601 3196
rect 4741 3162 4892 3196
rect 4450 3128 4552 3162
rect 4586 3128 4601 3162
rect 4741 3128 4756 3162
rect 4790 3128 4892 3162
rect 4450 3058 4601 3128
rect 4741 3058 4892 3128
rect 5012 4046 5322 4058
rect 5012 4012 5114 4046
rect 5148 4012 5186 4046
rect 5220 4012 5322 4046
rect 5012 3978 5322 4012
rect 5012 3944 5114 3978
rect 5148 3944 5186 3978
rect 5220 3944 5322 3978
rect 5012 3910 5322 3944
rect 5012 3876 5114 3910
rect 5148 3876 5186 3910
rect 5220 3876 5322 3910
rect 5012 3842 5322 3876
rect 5012 3808 5114 3842
rect 5148 3808 5186 3842
rect 5220 3808 5322 3842
rect 5012 3774 5322 3808
rect 5012 3740 5114 3774
rect 5148 3740 5186 3774
rect 5220 3740 5322 3774
rect 5012 3706 5322 3740
rect 5012 3672 5114 3706
rect 5148 3672 5186 3706
rect 5220 3672 5322 3706
rect 5012 3638 5322 3672
rect 5012 3604 5114 3638
rect 5148 3604 5186 3638
rect 5220 3604 5322 3638
rect 5012 3570 5322 3604
rect 5012 3536 5114 3570
rect 5148 3536 5186 3570
rect 5220 3536 5322 3570
rect 5012 3502 5322 3536
rect 5012 3468 5114 3502
rect 5148 3468 5186 3502
rect 5220 3468 5322 3502
rect 5012 3434 5322 3468
rect 5012 3400 5114 3434
rect 5148 3400 5186 3434
rect 5220 3400 5322 3434
rect 5012 3366 5322 3400
rect 5012 3332 5114 3366
rect 5148 3332 5186 3366
rect 5220 3332 5322 3366
rect 5012 3298 5322 3332
rect 5012 3264 5114 3298
rect 5148 3264 5186 3298
rect 5220 3264 5322 3298
rect 5012 3230 5322 3264
rect 5012 3196 5114 3230
rect 5148 3196 5186 3230
rect 5220 3196 5322 3230
rect 5012 3162 5322 3196
rect 5012 3128 5114 3162
rect 5148 3128 5186 3162
rect 5220 3128 5322 3162
rect 5012 3058 5322 3128
rect 5442 4046 5593 4058
rect 5733 4046 5884 4058
rect 5442 4012 5544 4046
rect 5578 4012 5593 4046
rect 5733 4012 5748 4046
rect 5782 4012 5884 4046
rect 5442 3978 5593 4012
rect 5733 3978 5884 4012
rect 5442 3944 5544 3978
rect 5578 3944 5593 3978
rect 5733 3944 5748 3978
rect 5782 3944 5884 3978
rect 5442 3910 5593 3944
rect 5733 3910 5884 3944
rect 5442 3876 5544 3910
rect 5578 3876 5593 3910
rect 5733 3876 5748 3910
rect 5782 3876 5884 3910
rect 5442 3842 5593 3876
rect 5733 3842 5884 3876
rect 5442 3808 5544 3842
rect 5578 3808 5593 3842
rect 5733 3808 5748 3842
rect 5782 3808 5884 3842
rect 5442 3774 5593 3808
rect 5733 3774 5884 3808
rect 5442 3740 5544 3774
rect 5578 3740 5593 3774
rect 5733 3740 5748 3774
rect 5782 3740 5884 3774
rect 5442 3706 5593 3740
rect 5733 3706 5884 3740
rect 5442 3672 5544 3706
rect 5578 3672 5593 3706
rect 5733 3672 5748 3706
rect 5782 3672 5884 3706
rect 5442 3638 5593 3672
rect 5733 3638 5884 3672
rect 5442 3604 5544 3638
rect 5578 3604 5593 3638
rect 5733 3604 5748 3638
rect 5782 3604 5884 3638
rect 5442 3570 5593 3604
rect 5733 3570 5884 3604
rect 5442 3536 5544 3570
rect 5578 3536 5593 3570
rect 5733 3536 5748 3570
rect 5782 3536 5884 3570
rect 5442 3502 5593 3536
rect 5733 3502 5884 3536
rect 5442 3468 5544 3502
rect 5578 3468 5593 3502
rect 5733 3468 5748 3502
rect 5782 3468 5884 3502
rect 5442 3434 5593 3468
rect 5733 3434 5884 3468
rect 5442 3400 5544 3434
rect 5578 3400 5593 3434
rect 5733 3400 5748 3434
rect 5782 3400 5884 3434
rect 5442 3366 5593 3400
rect 5733 3366 5884 3400
rect 5442 3332 5544 3366
rect 5578 3332 5593 3366
rect 5733 3332 5748 3366
rect 5782 3332 5884 3366
rect 5442 3298 5593 3332
rect 5733 3298 5884 3332
rect 5442 3264 5544 3298
rect 5578 3264 5593 3298
rect 5733 3264 5748 3298
rect 5782 3264 5884 3298
rect 5442 3230 5593 3264
rect 5733 3230 5884 3264
rect 5442 3196 5544 3230
rect 5578 3196 5593 3230
rect 5733 3196 5748 3230
rect 5782 3196 5884 3230
rect 5442 3162 5593 3196
rect 5733 3162 5884 3196
rect 5442 3128 5544 3162
rect 5578 3128 5593 3162
rect 5733 3128 5748 3162
rect 5782 3128 5884 3162
rect 5442 3058 5593 3128
rect 5733 3058 5884 3128
rect 6004 4046 6314 4058
rect 6004 4012 6106 4046
rect 6140 4012 6178 4046
rect 6212 4012 6314 4046
rect 6004 3978 6314 4012
rect 6004 3944 6106 3978
rect 6140 3944 6178 3978
rect 6212 3944 6314 3978
rect 6004 3910 6314 3944
rect 6004 3876 6106 3910
rect 6140 3876 6178 3910
rect 6212 3876 6314 3910
rect 6004 3842 6314 3876
rect 6004 3808 6106 3842
rect 6140 3808 6178 3842
rect 6212 3808 6314 3842
rect 6004 3774 6314 3808
rect 6004 3740 6106 3774
rect 6140 3740 6178 3774
rect 6212 3740 6314 3774
rect 6004 3706 6314 3740
rect 6004 3672 6106 3706
rect 6140 3672 6178 3706
rect 6212 3672 6314 3706
rect 6004 3638 6314 3672
rect 6004 3604 6106 3638
rect 6140 3604 6178 3638
rect 6212 3604 6314 3638
rect 6004 3570 6314 3604
rect 6004 3536 6106 3570
rect 6140 3536 6178 3570
rect 6212 3536 6314 3570
rect 6004 3502 6314 3536
rect 6004 3468 6106 3502
rect 6140 3468 6178 3502
rect 6212 3468 6314 3502
rect 6004 3434 6314 3468
rect 6004 3400 6106 3434
rect 6140 3400 6178 3434
rect 6212 3400 6314 3434
rect 6004 3366 6314 3400
rect 6004 3332 6106 3366
rect 6140 3332 6178 3366
rect 6212 3332 6314 3366
rect 6004 3298 6314 3332
rect 6004 3264 6106 3298
rect 6140 3264 6178 3298
rect 6212 3264 6314 3298
rect 6004 3230 6314 3264
rect 6004 3196 6106 3230
rect 6140 3196 6178 3230
rect 6212 3196 6314 3230
rect 6004 3162 6314 3196
rect 6004 3128 6106 3162
rect 6140 3128 6178 3162
rect 6212 3128 6314 3162
rect 6004 3058 6314 3128
rect 6434 4046 6585 4058
rect 6725 4046 6876 4058
rect 6434 4012 6536 4046
rect 6570 4012 6585 4046
rect 6725 4012 6740 4046
rect 6774 4012 6876 4046
rect 6434 3978 6585 4012
rect 6725 3978 6876 4012
rect 6434 3944 6536 3978
rect 6570 3944 6585 3978
rect 6725 3944 6740 3978
rect 6774 3944 6876 3978
rect 6434 3910 6585 3944
rect 6725 3910 6876 3944
rect 6434 3876 6536 3910
rect 6570 3876 6585 3910
rect 6725 3876 6740 3910
rect 6774 3876 6876 3910
rect 6434 3842 6585 3876
rect 6725 3842 6876 3876
rect 6434 3808 6536 3842
rect 6570 3808 6585 3842
rect 6725 3808 6740 3842
rect 6774 3808 6876 3842
rect 6434 3774 6585 3808
rect 6725 3774 6876 3808
rect 6434 3740 6536 3774
rect 6570 3740 6585 3774
rect 6725 3740 6740 3774
rect 6774 3740 6876 3774
rect 6434 3706 6585 3740
rect 6725 3706 6876 3740
rect 6434 3672 6536 3706
rect 6570 3672 6585 3706
rect 6725 3672 6740 3706
rect 6774 3672 6876 3706
rect 6434 3638 6585 3672
rect 6725 3638 6876 3672
rect 6434 3604 6536 3638
rect 6570 3604 6585 3638
rect 6725 3604 6740 3638
rect 6774 3604 6876 3638
rect 6434 3570 6585 3604
rect 6725 3570 6876 3604
rect 6434 3536 6536 3570
rect 6570 3536 6585 3570
rect 6725 3536 6740 3570
rect 6774 3536 6876 3570
rect 6434 3502 6585 3536
rect 6725 3502 6876 3536
rect 6434 3468 6536 3502
rect 6570 3468 6585 3502
rect 6725 3468 6740 3502
rect 6774 3468 6876 3502
rect 6434 3434 6585 3468
rect 6725 3434 6876 3468
rect 6434 3400 6536 3434
rect 6570 3400 6585 3434
rect 6725 3400 6740 3434
rect 6774 3400 6876 3434
rect 6434 3366 6585 3400
rect 6725 3366 6876 3400
rect 6434 3332 6536 3366
rect 6570 3332 6585 3366
rect 6725 3332 6740 3366
rect 6774 3332 6876 3366
rect 6434 3298 6585 3332
rect 6725 3298 6876 3332
rect 6434 3264 6536 3298
rect 6570 3264 6585 3298
rect 6725 3264 6740 3298
rect 6774 3264 6876 3298
rect 6434 3230 6585 3264
rect 6725 3230 6876 3264
rect 6434 3196 6536 3230
rect 6570 3196 6585 3230
rect 6725 3196 6740 3230
rect 6774 3196 6876 3230
rect 6434 3162 6585 3196
rect 6725 3162 6876 3196
rect 6434 3128 6536 3162
rect 6570 3128 6585 3162
rect 6725 3128 6740 3162
rect 6774 3128 6876 3162
rect 6434 3058 6585 3128
rect 6725 3058 6876 3128
rect 6996 4046 7306 4058
rect 6996 4012 7098 4046
rect 7132 4012 7170 4046
rect 7204 4012 7306 4046
rect 6996 3978 7306 4012
rect 6996 3944 7098 3978
rect 7132 3944 7170 3978
rect 7204 3944 7306 3978
rect 6996 3910 7306 3944
rect 6996 3876 7098 3910
rect 7132 3876 7170 3910
rect 7204 3876 7306 3910
rect 6996 3842 7306 3876
rect 6996 3808 7098 3842
rect 7132 3808 7170 3842
rect 7204 3808 7306 3842
rect 6996 3774 7306 3808
rect 6996 3740 7098 3774
rect 7132 3740 7170 3774
rect 7204 3740 7306 3774
rect 6996 3706 7306 3740
rect 6996 3672 7098 3706
rect 7132 3672 7170 3706
rect 7204 3672 7306 3706
rect 6996 3638 7306 3672
rect 6996 3604 7098 3638
rect 7132 3604 7170 3638
rect 7204 3604 7306 3638
rect 6996 3570 7306 3604
rect 6996 3536 7098 3570
rect 7132 3536 7170 3570
rect 7204 3536 7306 3570
rect 6996 3502 7306 3536
rect 6996 3468 7098 3502
rect 7132 3468 7170 3502
rect 7204 3468 7306 3502
rect 6996 3434 7306 3468
rect 6996 3400 7098 3434
rect 7132 3400 7170 3434
rect 7204 3400 7306 3434
rect 6996 3366 7306 3400
rect 6996 3332 7098 3366
rect 7132 3332 7170 3366
rect 7204 3332 7306 3366
rect 6996 3298 7306 3332
rect 6996 3264 7098 3298
rect 7132 3264 7170 3298
rect 7204 3264 7306 3298
rect 6996 3230 7306 3264
rect 6996 3196 7098 3230
rect 7132 3196 7170 3230
rect 7204 3196 7306 3230
rect 6996 3162 7306 3196
rect 6996 3128 7098 3162
rect 7132 3128 7170 3162
rect 7204 3128 7306 3162
rect 6996 3058 7306 3128
rect 7426 4046 7577 4058
rect 7717 4046 7868 4058
rect 7426 4012 7528 4046
rect 7562 4012 7577 4046
rect 7717 4012 7732 4046
rect 7766 4012 7868 4046
rect 7426 3978 7577 4012
rect 7717 3978 7868 4012
rect 7426 3944 7528 3978
rect 7562 3944 7577 3978
rect 7717 3944 7732 3978
rect 7766 3944 7868 3978
rect 7426 3910 7577 3944
rect 7717 3910 7868 3944
rect 7426 3876 7528 3910
rect 7562 3876 7577 3910
rect 7717 3876 7732 3910
rect 7766 3876 7868 3910
rect 7426 3842 7577 3876
rect 7717 3842 7868 3876
rect 7426 3808 7528 3842
rect 7562 3808 7577 3842
rect 7717 3808 7732 3842
rect 7766 3808 7868 3842
rect 7426 3774 7577 3808
rect 7717 3774 7868 3808
rect 7426 3740 7528 3774
rect 7562 3740 7577 3774
rect 7717 3740 7732 3774
rect 7766 3740 7868 3774
rect 7426 3706 7577 3740
rect 7717 3706 7868 3740
rect 7426 3672 7528 3706
rect 7562 3672 7577 3706
rect 7717 3672 7732 3706
rect 7766 3672 7868 3706
rect 7426 3638 7577 3672
rect 7717 3638 7868 3672
rect 7426 3604 7528 3638
rect 7562 3604 7577 3638
rect 7717 3604 7732 3638
rect 7766 3604 7868 3638
rect 7426 3570 7577 3604
rect 7717 3570 7868 3604
rect 7426 3536 7528 3570
rect 7562 3536 7577 3570
rect 7717 3536 7732 3570
rect 7766 3536 7868 3570
rect 7426 3502 7577 3536
rect 7717 3502 7868 3536
rect 7426 3468 7528 3502
rect 7562 3468 7577 3502
rect 7717 3468 7732 3502
rect 7766 3468 7868 3502
rect 7426 3434 7577 3468
rect 7717 3434 7868 3468
rect 7426 3400 7528 3434
rect 7562 3400 7577 3434
rect 7717 3400 7732 3434
rect 7766 3400 7868 3434
rect 7426 3366 7577 3400
rect 7717 3366 7868 3400
rect 7426 3332 7528 3366
rect 7562 3332 7577 3366
rect 7717 3332 7732 3366
rect 7766 3332 7868 3366
rect 7426 3298 7577 3332
rect 7717 3298 7868 3332
rect 7426 3264 7528 3298
rect 7562 3264 7577 3298
rect 7717 3264 7732 3298
rect 7766 3264 7868 3298
rect 7426 3230 7577 3264
rect 7717 3230 7868 3264
rect 7426 3196 7528 3230
rect 7562 3196 7577 3230
rect 7717 3196 7732 3230
rect 7766 3196 7868 3230
rect 7426 3162 7577 3196
rect 7717 3162 7868 3196
rect 7426 3128 7528 3162
rect 7562 3128 7577 3162
rect 7717 3128 7732 3162
rect 7766 3128 7868 3162
rect 7426 3058 7577 3128
rect 7717 3058 7868 3128
rect 7988 4046 8298 4058
rect 7988 4012 8090 4046
rect 8124 4012 8162 4046
rect 8196 4012 8298 4046
rect 7988 3978 8298 4012
rect 7988 3944 8090 3978
rect 8124 3944 8162 3978
rect 8196 3944 8298 3978
rect 7988 3910 8298 3944
rect 7988 3876 8090 3910
rect 8124 3876 8162 3910
rect 8196 3876 8298 3910
rect 7988 3842 8298 3876
rect 7988 3808 8090 3842
rect 8124 3808 8162 3842
rect 8196 3808 8298 3842
rect 7988 3774 8298 3808
rect 7988 3740 8090 3774
rect 8124 3740 8162 3774
rect 8196 3740 8298 3774
rect 7988 3706 8298 3740
rect 7988 3672 8090 3706
rect 8124 3672 8162 3706
rect 8196 3672 8298 3706
rect 7988 3638 8298 3672
rect 7988 3604 8090 3638
rect 8124 3604 8162 3638
rect 8196 3604 8298 3638
rect 7988 3570 8298 3604
rect 7988 3536 8090 3570
rect 8124 3536 8162 3570
rect 8196 3536 8298 3570
rect 7988 3502 8298 3536
rect 7988 3468 8090 3502
rect 8124 3468 8162 3502
rect 8196 3468 8298 3502
rect 7988 3434 8298 3468
rect 7988 3400 8090 3434
rect 8124 3400 8162 3434
rect 8196 3400 8298 3434
rect 7988 3366 8298 3400
rect 7988 3332 8090 3366
rect 8124 3332 8162 3366
rect 8196 3332 8298 3366
rect 7988 3298 8298 3332
rect 7988 3264 8090 3298
rect 8124 3264 8162 3298
rect 8196 3264 8298 3298
rect 7988 3230 8298 3264
rect 7988 3196 8090 3230
rect 8124 3196 8162 3230
rect 8196 3196 8298 3230
rect 7988 3162 8298 3196
rect 7988 3128 8090 3162
rect 8124 3128 8162 3162
rect 8196 3128 8298 3162
rect 7988 3058 8298 3128
rect 8418 4046 8569 4058
rect 8709 4046 8860 4058
rect 8418 4012 8520 4046
rect 8554 4012 8569 4046
rect 8709 4012 8724 4046
rect 8758 4012 8860 4046
rect 8418 3978 8569 4012
rect 8709 3978 8860 4012
rect 8418 3944 8520 3978
rect 8554 3944 8569 3978
rect 8709 3944 8724 3978
rect 8758 3944 8860 3978
rect 8418 3910 8569 3944
rect 8709 3910 8860 3944
rect 8418 3876 8520 3910
rect 8554 3876 8569 3910
rect 8709 3876 8724 3910
rect 8758 3876 8860 3910
rect 8418 3842 8569 3876
rect 8709 3842 8860 3876
rect 8418 3808 8520 3842
rect 8554 3808 8569 3842
rect 8709 3808 8724 3842
rect 8758 3808 8860 3842
rect 8418 3774 8569 3808
rect 8709 3774 8860 3808
rect 8418 3740 8520 3774
rect 8554 3740 8569 3774
rect 8709 3740 8724 3774
rect 8758 3740 8860 3774
rect 8418 3706 8569 3740
rect 8709 3706 8860 3740
rect 8418 3672 8520 3706
rect 8554 3672 8569 3706
rect 8709 3672 8724 3706
rect 8758 3672 8860 3706
rect 8418 3638 8569 3672
rect 8709 3638 8860 3672
rect 8418 3604 8520 3638
rect 8554 3604 8569 3638
rect 8709 3604 8724 3638
rect 8758 3604 8860 3638
rect 8418 3570 8569 3604
rect 8709 3570 8860 3604
rect 8418 3536 8520 3570
rect 8554 3536 8569 3570
rect 8709 3536 8724 3570
rect 8758 3536 8860 3570
rect 8418 3502 8569 3536
rect 8709 3502 8860 3536
rect 8418 3468 8520 3502
rect 8554 3468 8569 3502
rect 8709 3468 8724 3502
rect 8758 3468 8860 3502
rect 8418 3434 8569 3468
rect 8709 3434 8860 3468
rect 8418 3400 8520 3434
rect 8554 3400 8569 3434
rect 8709 3400 8724 3434
rect 8758 3400 8860 3434
rect 8418 3366 8569 3400
rect 8709 3366 8860 3400
rect 8418 3332 8520 3366
rect 8554 3332 8569 3366
rect 8709 3332 8724 3366
rect 8758 3332 8860 3366
rect 8418 3298 8569 3332
rect 8709 3298 8860 3332
rect 8418 3264 8520 3298
rect 8554 3264 8569 3298
rect 8709 3264 8724 3298
rect 8758 3264 8860 3298
rect 8418 3230 8569 3264
rect 8709 3230 8860 3264
rect 8418 3196 8520 3230
rect 8554 3196 8569 3230
rect 8709 3196 8724 3230
rect 8758 3196 8860 3230
rect 8418 3162 8569 3196
rect 8709 3162 8860 3196
rect 8418 3128 8520 3162
rect 8554 3128 8569 3162
rect 8709 3128 8724 3162
rect 8758 3128 8860 3162
rect 8418 3058 8569 3128
rect 8709 3058 8860 3128
rect 8980 4046 9290 4058
rect 8980 4012 9082 4046
rect 9116 4012 9154 4046
rect 9188 4012 9290 4046
rect 8980 3978 9290 4012
rect 8980 3944 9082 3978
rect 9116 3944 9154 3978
rect 9188 3944 9290 3978
rect 8980 3910 9290 3944
rect 8980 3876 9082 3910
rect 9116 3876 9154 3910
rect 9188 3876 9290 3910
rect 8980 3842 9290 3876
rect 8980 3808 9082 3842
rect 9116 3808 9154 3842
rect 9188 3808 9290 3842
rect 8980 3774 9290 3808
rect 8980 3740 9082 3774
rect 9116 3740 9154 3774
rect 9188 3740 9290 3774
rect 8980 3706 9290 3740
rect 8980 3672 9082 3706
rect 9116 3672 9154 3706
rect 9188 3672 9290 3706
rect 8980 3638 9290 3672
rect 8980 3604 9082 3638
rect 9116 3604 9154 3638
rect 9188 3604 9290 3638
rect 8980 3570 9290 3604
rect 8980 3536 9082 3570
rect 9116 3536 9154 3570
rect 9188 3536 9290 3570
rect 8980 3502 9290 3536
rect 8980 3468 9082 3502
rect 9116 3468 9154 3502
rect 9188 3468 9290 3502
rect 8980 3434 9290 3468
rect 8980 3400 9082 3434
rect 9116 3400 9154 3434
rect 9188 3400 9290 3434
rect 8980 3366 9290 3400
rect 8980 3332 9082 3366
rect 9116 3332 9154 3366
rect 9188 3332 9290 3366
rect 8980 3298 9290 3332
rect 8980 3264 9082 3298
rect 9116 3264 9154 3298
rect 9188 3264 9290 3298
rect 8980 3230 9290 3264
rect 8980 3196 9082 3230
rect 9116 3196 9154 3230
rect 9188 3196 9290 3230
rect 8980 3162 9290 3196
rect 8980 3128 9082 3162
rect 9116 3128 9154 3162
rect 9188 3128 9290 3162
rect 8980 3058 9290 3128
rect 9410 4046 9561 4058
rect 9701 4046 9852 4058
rect 9410 4012 9512 4046
rect 9546 4012 9561 4046
rect 9701 4012 9716 4046
rect 9750 4012 9852 4046
rect 9410 3978 9561 4012
rect 9701 3978 9852 4012
rect 9410 3944 9512 3978
rect 9546 3944 9561 3978
rect 9701 3944 9716 3978
rect 9750 3944 9852 3978
rect 9410 3910 9561 3944
rect 9701 3910 9852 3944
rect 9410 3876 9512 3910
rect 9546 3876 9561 3910
rect 9701 3876 9716 3910
rect 9750 3876 9852 3910
rect 9410 3842 9561 3876
rect 9701 3842 9852 3876
rect 9410 3808 9512 3842
rect 9546 3808 9561 3842
rect 9701 3808 9716 3842
rect 9750 3808 9852 3842
rect 9410 3774 9561 3808
rect 9701 3774 9852 3808
rect 9410 3740 9512 3774
rect 9546 3740 9561 3774
rect 9701 3740 9716 3774
rect 9750 3740 9852 3774
rect 9410 3706 9561 3740
rect 9701 3706 9852 3740
rect 9410 3672 9512 3706
rect 9546 3672 9561 3706
rect 9701 3672 9716 3706
rect 9750 3672 9852 3706
rect 9410 3638 9561 3672
rect 9701 3638 9852 3672
rect 9410 3604 9512 3638
rect 9546 3604 9561 3638
rect 9701 3604 9716 3638
rect 9750 3604 9852 3638
rect 9410 3570 9561 3604
rect 9701 3570 9852 3604
rect 9410 3536 9512 3570
rect 9546 3536 9561 3570
rect 9701 3536 9716 3570
rect 9750 3536 9852 3570
rect 9410 3502 9561 3536
rect 9701 3502 9852 3536
rect 9410 3468 9512 3502
rect 9546 3468 9561 3502
rect 9701 3468 9716 3502
rect 9750 3468 9852 3502
rect 9410 3434 9561 3468
rect 9701 3434 9852 3468
rect 9410 3400 9512 3434
rect 9546 3400 9561 3434
rect 9701 3400 9716 3434
rect 9750 3400 9852 3434
rect 9410 3366 9561 3400
rect 9701 3366 9852 3400
rect 9410 3332 9512 3366
rect 9546 3332 9561 3366
rect 9701 3332 9716 3366
rect 9750 3332 9852 3366
rect 9410 3298 9561 3332
rect 9701 3298 9852 3332
rect 9410 3264 9512 3298
rect 9546 3264 9561 3298
rect 9701 3264 9716 3298
rect 9750 3264 9852 3298
rect 9410 3230 9561 3264
rect 9701 3230 9852 3264
rect 9410 3196 9512 3230
rect 9546 3196 9561 3230
rect 9701 3196 9716 3230
rect 9750 3196 9852 3230
rect 9410 3162 9561 3196
rect 9701 3162 9852 3196
rect 9410 3128 9512 3162
rect 9546 3128 9561 3162
rect 9701 3128 9716 3162
rect 9750 3128 9852 3162
rect 9410 3058 9561 3128
rect 9701 3058 9852 3128
rect 9972 4046 10282 4058
rect 9972 4012 10074 4046
rect 10108 4012 10146 4046
rect 10180 4012 10282 4046
rect 9972 3978 10282 4012
rect 9972 3944 10074 3978
rect 10108 3944 10146 3978
rect 10180 3944 10282 3978
rect 9972 3910 10282 3944
rect 9972 3876 10074 3910
rect 10108 3876 10146 3910
rect 10180 3876 10282 3910
rect 9972 3842 10282 3876
rect 9972 3808 10074 3842
rect 10108 3808 10146 3842
rect 10180 3808 10282 3842
rect 9972 3774 10282 3808
rect 9972 3740 10074 3774
rect 10108 3740 10146 3774
rect 10180 3740 10282 3774
rect 9972 3706 10282 3740
rect 9972 3672 10074 3706
rect 10108 3672 10146 3706
rect 10180 3672 10282 3706
rect 9972 3638 10282 3672
rect 9972 3604 10074 3638
rect 10108 3604 10146 3638
rect 10180 3604 10282 3638
rect 9972 3570 10282 3604
rect 9972 3536 10074 3570
rect 10108 3536 10146 3570
rect 10180 3536 10282 3570
rect 9972 3502 10282 3536
rect 9972 3468 10074 3502
rect 10108 3468 10146 3502
rect 10180 3468 10282 3502
rect 9972 3434 10282 3468
rect 9972 3400 10074 3434
rect 10108 3400 10146 3434
rect 10180 3400 10282 3434
rect 9972 3366 10282 3400
rect 9972 3332 10074 3366
rect 10108 3332 10146 3366
rect 10180 3332 10282 3366
rect 9972 3298 10282 3332
rect 9972 3264 10074 3298
rect 10108 3264 10146 3298
rect 10180 3264 10282 3298
rect 9972 3230 10282 3264
rect 9972 3196 10074 3230
rect 10108 3196 10146 3230
rect 10180 3196 10282 3230
rect 9972 3162 10282 3196
rect 9972 3128 10074 3162
rect 10108 3128 10146 3162
rect 10180 3128 10282 3162
rect 9972 3058 10282 3128
rect 10402 4046 10553 4058
rect 10693 4046 10844 4058
rect 10402 4012 10504 4046
rect 10538 4012 10553 4046
rect 10693 4012 10708 4046
rect 10742 4012 10844 4046
rect 10402 3978 10553 4012
rect 10693 3978 10844 4012
rect 10402 3944 10504 3978
rect 10538 3944 10553 3978
rect 10693 3944 10708 3978
rect 10742 3944 10844 3978
rect 10402 3910 10553 3944
rect 10693 3910 10844 3944
rect 10402 3876 10504 3910
rect 10538 3876 10553 3910
rect 10693 3876 10708 3910
rect 10742 3876 10844 3910
rect 10402 3842 10553 3876
rect 10693 3842 10844 3876
rect 10402 3808 10504 3842
rect 10538 3808 10553 3842
rect 10693 3808 10708 3842
rect 10742 3808 10844 3842
rect 10402 3774 10553 3808
rect 10693 3774 10844 3808
rect 10402 3740 10504 3774
rect 10538 3740 10553 3774
rect 10693 3740 10708 3774
rect 10742 3740 10844 3774
rect 10402 3706 10553 3740
rect 10693 3706 10844 3740
rect 10402 3672 10504 3706
rect 10538 3672 10553 3706
rect 10693 3672 10708 3706
rect 10742 3672 10844 3706
rect 10402 3638 10553 3672
rect 10693 3638 10844 3672
rect 10402 3604 10504 3638
rect 10538 3604 10553 3638
rect 10693 3604 10708 3638
rect 10742 3604 10844 3638
rect 10402 3570 10553 3604
rect 10693 3570 10844 3604
rect 10402 3536 10504 3570
rect 10538 3536 10553 3570
rect 10693 3536 10708 3570
rect 10742 3536 10844 3570
rect 10402 3502 10553 3536
rect 10693 3502 10844 3536
rect 10402 3468 10504 3502
rect 10538 3468 10553 3502
rect 10693 3468 10708 3502
rect 10742 3468 10844 3502
rect 10402 3434 10553 3468
rect 10693 3434 10844 3468
rect 10402 3400 10504 3434
rect 10538 3400 10553 3434
rect 10693 3400 10708 3434
rect 10742 3400 10844 3434
rect 10402 3366 10553 3400
rect 10693 3366 10844 3400
rect 10402 3332 10504 3366
rect 10538 3332 10553 3366
rect 10693 3332 10708 3366
rect 10742 3332 10844 3366
rect 10402 3298 10553 3332
rect 10693 3298 10844 3332
rect 10402 3264 10504 3298
rect 10538 3264 10553 3298
rect 10693 3264 10708 3298
rect 10742 3264 10844 3298
rect 10402 3230 10553 3264
rect 10693 3230 10844 3264
rect 10402 3196 10504 3230
rect 10538 3196 10553 3230
rect 10693 3196 10708 3230
rect 10742 3196 10844 3230
rect 10402 3162 10553 3196
rect 10693 3162 10844 3196
rect 10402 3128 10504 3162
rect 10538 3128 10553 3162
rect 10693 3128 10708 3162
rect 10742 3128 10844 3162
rect 10402 3058 10553 3128
rect 10693 3058 10844 3128
rect 10964 4046 11274 4058
rect 10964 4012 11066 4046
rect 11100 4012 11138 4046
rect 11172 4012 11274 4046
rect 10964 3978 11274 4012
rect 10964 3944 11066 3978
rect 11100 3944 11138 3978
rect 11172 3944 11274 3978
rect 10964 3910 11274 3944
rect 10964 3876 11066 3910
rect 11100 3876 11138 3910
rect 11172 3876 11274 3910
rect 10964 3842 11274 3876
rect 10964 3808 11066 3842
rect 11100 3808 11138 3842
rect 11172 3808 11274 3842
rect 10964 3774 11274 3808
rect 10964 3740 11066 3774
rect 11100 3740 11138 3774
rect 11172 3740 11274 3774
rect 10964 3706 11274 3740
rect 10964 3672 11066 3706
rect 11100 3672 11138 3706
rect 11172 3672 11274 3706
rect 10964 3638 11274 3672
rect 10964 3604 11066 3638
rect 11100 3604 11138 3638
rect 11172 3604 11274 3638
rect 10964 3570 11274 3604
rect 10964 3536 11066 3570
rect 11100 3536 11138 3570
rect 11172 3536 11274 3570
rect 10964 3502 11274 3536
rect 10964 3468 11066 3502
rect 11100 3468 11138 3502
rect 11172 3468 11274 3502
rect 10964 3434 11274 3468
rect 10964 3400 11066 3434
rect 11100 3400 11138 3434
rect 11172 3400 11274 3434
rect 10964 3366 11274 3400
rect 10964 3332 11066 3366
rect 11100 3332 11138 3366
rect 11172 3332 11274 3366
rect 10964 3298 11274 3332
rect 10964 3264 11066 3298
rect 11100 3264 11138 3298
rect 11172 3264 11274 3298
rect 10964 3230 11274 3264
rect 10964 3196 11066 3230
rect 11100 3196 11138 3230
rect 11172 3196 11274 3230
rect 10964 3162 11274 3196
rect 10964 3128 11066 3162
rect 11100 3128 11138 3162
rect 11172 3128 11274 3162
rect 10964 3058 11274 3128
rect 11394 4046 11545 4058
rect 11685 4046 11836 4058
rect 11394 4012 11496 4046
rect 11530 4012 11545 4046
rect 11685 4012 11700 4046
rect 11734 4012 11836 4046
rect 11394 3978 11545 4012
rect 11685 3978 11836 4012
rect 11394 3944 11496 3978
rect 11530 3944 11545 3978
rect 11685 3944 11700 3978
rect 11734 3944 11836 3978
rect 11394 3910 11545 3944
rect 11685 3910 11836 3944
rect 11394 3876 11496 3910
rect 11530 3876 11545 3910
rect 11685 3876 11700 3910
rect 11734 3876 11836 3910
rect 11394 3842 11545 3876
rect 11685 3842 11836 3876
rect 11394 3808 11496 3842
rect 11530 3808 11545 3842
rect 11685 3808 11700 3842
rect 11734 3808 11836 3842
rect 11394 3774 11545 3808
rect 11685 3774 11836 3808
rect 11394 3740 11496 3774
rect 11530 3740 11545 3774
rect 11685 3740 11700 3774
rect 11734 3740 11836 3774
rect 11394 3706 11545 3740
rect 11685 3706 11836 3740
rect 11394 3672 11496 3706
rect 11530 3672 11545 3706
rect 11685 3672 11700 3706
rect 11734 3672 11836 3706
rect 11394 3638 11545 3672
rect 11685 3638 11836 3672
rect 11394 3604 11496 3638
rect 11530 3604 11545 3638
rect 11685 3604 11700 3638
rect 11734 3604 11836 3638
rect 11394 3570 11545 3604
rect 11685 3570 11836 3604
rect 11394 3536 11496 3570
rect 11530 3536 11545 3570
rect 11685 3536 11700 3570
rect 11734 3536 11836 3570
rect 11394 3502 11545 3536
rect 11685 3502 11836 3536
rect 11394 3468 11496 3502
rect 11530 3468 11545 3502
rect 11685 3468 11700 3502
rect 11734 3468 11836 3502
rect 11394 3434 11545 3468
rect 11685 3434 11836 3468
rect 11394 3400 11496 3434
rect 11530 3400 11545 3434
rect 11685 3400 11700 3434
rect 11734 3400 11836 3434
rect 11394 3366 11545 3400
rect 11685 3366 11836 3400
rect 11394 3332 11496 3366
rect 11530 3332 11545 3366
rect 11685 3332 11700 3366
rect 11734 3332 11836 3366
rect 11394 3298 11545 3332
rect 11685 3298 11836 3332
rect 11394 3264 11496 3298
rect 11530 3264 11545 3298
rect 11685 3264 11700 3298
rect 11734 3264 11836 3298
rect 11394 3230 11545 3264
rect 11685 3230 11836 3264
rect 11394 3196 11496 3230
rect 11530 3196 11545 3230
rect 11685 3196 11700 3230
rect 11734 3196 11836 3230
rect 11394 3162 11545 3196
rect 11685 3162 11836 3196
rect 11394 3128 11496 3162
rect 11530 3128 11545 3162
rect 11685 3128 11700 3162
rect 11734 3128 11836 3162
rect 11394 3058 11545 3128
rect 11685 3058 11836 3128
rect 11956 4046 12266 4058
rect 11956 4012 12058 4046
rect 12092 4012 12130 4046
rect 12164 4012 12266 4046
rect 11956 3978 12266 4012
rect 11956 3944 12058 3978
rect 12092 3944 12130 3978
rect 12164 3944 12266 3978
rect 11956 3910 12266 3944
rect 11956 3876 12058 3910
rect 12092 3876 12130 3910
rect 12164 3876 12266 3910
rect 11956 3842 12266 3876
rect 11956 3808 12058 3842
rect 12092 3808 12130 3842
rect 12164 3808 12266 3842
rect 11956 3774 12266 3808
rect 11956 3740 12058 3774
rect 12092 3740 12130 3774
rect 12164 3740 12266 3774
rect 11956 3706 12266 3740
rect 11956 3672 12058 3706
rect 12092 3672 12130 3706
rect 12164 3672 12266 3706
rect 11956 3638 12266 3672
rect 11956 3604 12058 3638
rect 12092 3604 12130 3638
rect 12164 3604 12266 3638
rect 11956 3570 12266 3604
rect 11956 3536 12058 3570
rect 12092 3536 12130 3570
rect 12164 3536 12266 3570
rect 11956 3502 12266 3536
rect 11956 3468 12058 3502
rect 12092 3468 12130 3502
rect 12164 3468 12266 3502
rect 11956 3434 12266 3468
rect 11956 3400 12058 3434
rect 12092 3400 12130 3434
rect 12164 3400 12266 3434
rect 11956 3366 12266 3400
rect 11956 3332 12058 3366
rect 12092 3332 12130 3366
rect 12164 3332 12266 3366
rect 11956 3298 12266 3332
rect 11956 3264 12058 3298
rect 12092 3264 12130 3298
rect 12164 3264 12266 3298
rect 11956 3230 12266 3264
rect 11956 3196 12058 3230
rect 12092 3196 12130 3230
rect 12164 3196 12266 3230
rect 11956 3162 12266 3196
rect 11956 3128 12058 3162
rect 12092 3128 12130 3162
rect 12164 3128 12266 3162
rect 11956 3058 12266 3128
rect 12386 4046 12537 4058
rect 12677 4046 12828 4058
rect 12386 4012 12488 4046
rect 12522 4012 12537 4046
rect 12677 4012 12692 4046
rect 12726 4012 12828 4046
rect 12386 3978 12537 4012
rect 12677 3978 12828 4012
rect 12386 3944 12488 3978
rect 12522 3944 12537 3978
rect 12677 3944 12692 3978
rect 12726 3944 12828 3978
rect 12386 3910 12537 3944
rect 12677 3910 12828 3944
rect 12386 3876 12488 3910
rect 12522 3876 12537 3910
rect 12677 3876 12692 3910
rect 12726 3876 12828 3910
rect 12386 3842 12537 3876
rect 12677 3842 12828 3876
rect 12386 3808 12488 3842
rect 12522 3808 12537 3842
rect 12677 3808 12692 3842
rect 12726 3808 12828 3842
rect 12386 3774 12537 3808
rect 12677 3774 12828 3808
rect 12386 3740 12488 3774
rect 12522 3740 12537 3774
rect 12677 3740 12692 3774
rect 12726 3740 12828 3774
rect 12386 3706 12537 3740
rect 12677 3706 12828 3740
rect 12386 3672 12488 3706
rect 12522 3672 12537 3706
rect 12677 3672 12692 3706
rect 12726 3672 12828 3706
rect 12386 3638 12537 3672
rect 12677 3638 12828 3672
rect 12386 3604 12488 3638
rect 12522 3604 12537 3638
rect 12677 3604 12692 3638
rect 12726 3604 12828 3638
rect 12386 3570 12537 3604
rect 12677 3570 12828 3604
rect 12386 3536 12488 3570
rect 12522 3536 12537 3570
rect 12677 3536 12692 3570
rect 12726 3536 12828 3570
rect 12386 3502 12537 3536
rect 12677 3502 12828 3536
rect 12386 3468 12488 3502
rect 12522 3468 12537 3502
rect 12677 3468 12692 3502
rect 12726 3468 12828 3502
rect 12386 3434 12537 3468
rect 12677 3434 12828 3468
rect 12386 3400 12488 3434
rect 12522 3400 12537 3434
rect 12677 3400 12692 3434
rect 12726 3400 12828 3434
rect 12386 3366 12537 3400
rect 12677 3366 12828 3400
rect 12386 3332 12488 3366
rect 12522 3332 12537 3366
rect 12677 3332 12692 3366
rect 12726 3332 12828 3366
rect 12386 3298 12537 3332
rect 12677 3298 12828 3332
rect 12386 3264 12488 3298
rect 12522 3264 12537 3298
rect 12677 3264 12692 3298
rect 12726 3264 12828 3298
rect 12386 3230 12537 3264
rect 12677 3230 12828 3264
rect 12386 3196 12488 3230
rect 12522 3196 12537 3230
rect 12677 3196 12692 3230
rect 12726 3196 12828 3230
rect 12386 3162 12537 3196
rect 12677 3162 12828 3196
rect 12386 3128 12488 3162
rect 12522 3128 12537 3162
rect 12677 3128 12692 3162
rect 12726 3128 12828 3162
rect 12386 3058 12537 3128
rect 12677 3058 12828 3128
rect 12948 4046 13258 4058
rect 12948 4012 13050 4046
rect 13084 4012 13122 4046
rect 13156 4012 13258 4046
rect 12948 3978 13258 4012
rect 12948 3944 13050 3978
rect 13084 3944 13122 3978
rect 13156 3944 13258 3978
rect 12948 3910 13258 3944
rect 12948 3876 13050 3910
rect 13084 3876 13122 3910
rect 13156 3876 13258 3910
rect 12948 3842 13258 3876
rect 12948 3808 13050 3842
rect 13084 3808 13122 3842
rect 13156 3808 13258 3842
rect 12948 3774 13258 3808
rect 12948 3740 13050 3774
rect 13084 3740 13122 3774
rect 13156 3740 13258 3774
rect 12948 3706 13258 3740
rect 12948 3672 13050 3706
rect 13084 3672 13122 3706
rect 13156 3672 13258 3706
rect 12948 3638 13258 3672
rect 12948 3604 13050 3638
rect 13084 3604 13122 3638
rect 13156 3604 13258 3638
rect 12948 3570 13258 3604
rect 12948 3536 13050 3570
rect 13084 3536 13122 3570
rect 13156 3536 13258 3570
rect 12948 3502 13258 3536
rect 12948 3468 13050 3502
rect 13084 3468 13122 3502
rect 13156 3468 13258 3502
rect 12948 3434 13258 3468
rect 12948 3400 13050 3434
rect 13084 3400 13122 3434
rect 13156 3400 13258 3434
rect 12948 3366 13258 3400
rect 12948 3332 13050 3366
rect 13084 3332 13122 3366
rect 13156 3332 13258 3366
rect 12948 3298 13258 3332
rect 12948 3264 13050 3298
rect 13084 3264 13122 3298
rect 13156 3264 13258 3298
rect 12948 3230 13258 3264
rect 12948 3196 13050 3230
rect 13084 3196 13122 3230
rect 13156 3196 13258 3230
rect 12948 3162 13258 3196
rect 12948 3128 13050 3162
rect 13084 3128 13122 3162
rect 13156 3128 13258 3162
rect 12948 3058 13258 3128
rect 13378 4046 13529 4058
rect 13669 4046 13820 4058
rect 13378 4012 13480 4046
rect 13514 4012 13529 4046
rect 13669 4012 13684 4046
rect 13718 4012 13820 4046
rect 13378 3978 13529 4012
rect 13669 3978 13820 4012
rect 13378 3944 13480 3978
rect 13514 3944 13529 3978
rect 13669 3944 13684 3978
rect 13718 3944 13820 3978
rect 13378 3910 13529 3944
rect 13669 3910 13820 3944
rect 13378 3876 13480 3910
rect 13514 3876 13529 3910
rect 13669 3876 13684 3910
rect 13718 3876 13820 3910
rect 13378 3842 13529 3876
rect 13669 3842 13820 3876
rect 13378 3808 13480 3842
rect 13514 3808 13529 3842
rect 13669 3808 13684 3842
rect 13718 3808 13820 3842
rect 13378 3774 13529 3808
rect 13669 3774 13820 3808
rect 13378 3740 13480 3774
rect 13514 3740 13529 3774
rect 13669 3740 13684 3774
rect 13718 3740 13820 3774
rect 13378 3706 13529 3740
rect 13669 3706 13820 3740
rect 13378 3672 13480 3706
rect 13514 3672 13529 3706
rect 13669 3672 13684 3706
rect 13718 3672 13820 3706
rect 13378 3638 13529 3672
rect 13669 3638 13820 3672
rect 13378 3604 13480 3638
rect 13514 3604 13529 3638
rect 13669 3604 13684 3638
rect 13718 3604 13820 3638
rect 13378 3570 13529 3604
rect 13669 3570 13820 3604
rect 13378 3536 13480 3570
rect 13514 3536 13529 3570
rect 13669 3536 13684 3570
rect 13718 3536 13820 3570
rect 13378 3502 13529 3536
rect 13669 3502 13820 3536
rect 13378 3468 13480 3502
rect 13514 3468 13529 3502
rect 13669 3468 13684 3502
rect 13718 3468 13820 3502
rect 13378 3434 13529 3468
rect 13669 3434 13820 3468
rect 13378 3400 13480 3434
rect 13514 3400 13529 3434
rect 13669 3400 13684 3434
rect 13718 3400 13820 3434
rect 13378 3366 13529 3400
rect 13669 3366 13820 3400
rect 13378 3332 13480 3366
rect 13514 3332 13529 3366
rect 13669 3332 13684 3366
rect 13718 3332 13820 3366
rect 13378 3298 13529 3332
rect 13669 3298 13820 3332
rect 13378 3264 13480 3298
rect 13514 3264 13529 3298
rect 13669 3264 13684 3298
rect 13718 3264 13820 3298
rect 13378 3230 13529 3264
rect 13669 3230 13820 3264
rect 13378 3196 13480 3230
rect 13514 3196 13529 3230
rect 13669 3196 13684 3230
rect 13718 3196 13820 3230
rect 13378 3162 13529 3196
rect 13669 3162 13820 3196
rect 13378 3128 13480 3162
rect 13514 3128 13529 3162
rect 13669 3128 13684 3162
rect 13718 3128 13820 3162
rect 13378 3058 13529 3128
rect 13669 3058 13820 3128
rect 13940 4046 14178 4058
rect 13940 4012 14042 4046
rect 14076 4012 14178 4046
rect 13940 3978 14178 4012
rect 13940 3944 14042 3978
rect 14076 3944 14178 3978
rect 13940 3910 14178 3944
rect 13940 3876 14042 3910
rect 14076 3876 14178 3910
rect 13940 3842 14178 3876
rect 13940 3808 14042 3842
rect 14076 3808 14178 3842
rect 13940 3774 14178 3808
rect 13940 3740 14042 3774
rect 14076 3740 14178 3774
rect 13940 3706 14178 3740
rect 13940 3672 14042 3706
rect 14076 3672 14178 3706
rect 13940 3638 14178 3672
rect 13940 3604 14042 3638
rect 14076 3604 14178 3638
rect 13940 3570 14178 3604
rect 13940 3536 14042 3570
rect 14076 3536 14178 3570
rect 13940 3502 14178 3536
rect 13940 3468 14042 3502
rect 14076 3468 14178 3502
rect 13940 3434 14178 3468
rect 13940 3400 14042 3434
rect 14076 3400 14178 3434
rect 13940 3366 14178 3400
rect 13940 3332 14042 3366
rect 14076 3332 14178 3366
rect 13940 3298 14178 3332
rect 13940 3264 14042 3298
rect 14076 3264 14178 3298
rect 13940 3230 14178 3264
rect 13940 3196 14042 3230
rect 14076 3196 14178 3230
rect 13940 3162 14178 3196
rect 13940 3128 14042 3162
rect 14076 3128 14178 3162
rect 13940 3058 14178 3128
rect 14298 4046 14435 4058
rect 14298 4012 14386 4046
rect 14420 4012 14435 4046
rect 14298 3978 14435 4012
rect 14298 3944 14386 3978
rect 14420 3944 14435 3978
rect 14298 3910 14435 3944
rect 14298 3876 14386 3910
rect 14420 3876 14435 3910
rect 14298 3842 14435 3876
rect 14298 3808 14386 3842
rect 14420 3808 14435 3842
rect 14298 3774 14435 3808
rect 14298 3740 14386 3774
rect 14420 3740 14435 3774
rect 14298 3706 14435 3740
rect 14298 3672 14386 3706
rect 14420 3672 14435 3706
rect 14298 3638 14435 3672
rect 14298 3604 14386 3638
rect 14420 3604 14435 3638
rect 14298 3570 14435 3604
rect 14298 3536 14386 3570
rect 14420 3536 14435 3570
rect 14298 3502 14435 3536
rect 14298 3468 14386 3502
rect 14420 3468 14435 3502
rect 14298 3434 14435 3468
rect 14298 3400 14386 3434
rect 14420 3400 14435 3434
rect 14298 3366 14435 3400
rect 14298 3332 14386 3366
rect 14420 3332 14435 3366
rect 14298 3298 14435 3332
rect 14298 3264 14386 3298
rect 14420 3264 14435 3298
rect 14298 3230 14435 3264
rect 14298 3196 14386 3230
rect 14420 3196 14435 3230
rect 14298 3162 14435 3196
rect 14298 3128 14386 3162
rect 14420 3128 14435 3162
rect 14298 3058 14435 3128
rect 787 2445 924 2457
rect 787 2411 802 2445
rect 836 2411 924 2445
rect 787 2377 924 2411
rect 787 2343 802 2377
rect 836 2343 924 2377
rect 787 2309 924 2343
rect 787 2275 802 2309
rect 836 2275 924 2309
rect 787 2241 924 2275
rect 787 2207 802 2241
rect 836 2207 924 2241
rect 787 2173 924 2207
rect 787 2139 802 2173
rect 836 2139 924 2173
rect 787 2105 924 2139
rect 787 2071 802 2105
rect 836 2071 924 2105
rect 787 2037 924 2071
rect 787 2003 802 2037
rect 836 2003 924 2037
rect 787 1969 924 2003
rect 787 1935 802 1969
rect 836 1935 924 1969
rect 787 1901 924 1935
rect 787 1867 802 1901
rect 836 1867 924 1901
rect 787 1833 924 1867
rect 787 1799 802 1833
rect 836 1799 924 1833
rect 787 1765 924 1799
rect 787 1731 802 1765
rect 836 1731 924 1765
rect 787 1697 924 1731
rect 787 1663 802 1697
rect 836 1663 924 1697
rect 787 1629 924 1663
rect 787 1595 802 1629
rect 836 1595 924 1629
rect 787 1561 924 1595
rect 787 1527 802 1561
rect 836 1527 924 1561
rect 787 1457 924 1527
rect 1044 2445 1354 2457
rect 1044 2411 1146 2445
rect 1180 2411 1218 2445
rect 1252 2411 1354 2445
rect 1044 2377 1354 2411
rect 1044 2343 1146 2377
rect 1180 2343 1218 2377
rect 1252 2343 1354 2377
rect 1044 2309 1354 2343
rect 1044 2275 1146 2309
rect 1180 2275 1218 2309
rect 1252 2275 1354 2309
rect 1044 2241 1354 2275
rect 1044 2207 1146 2241
rect 1180 2207 1218 2241
rect 1252 2207 1354 2241
rect 1044 2173 1354 2207
rect 1044 2139 1146 2173
rect 1180 2139 1218 2173
rect 1252 2139 1354 2173
rect 1044 2105 1354 2139
rect 1044 2071 1146 2105
rect 1180 2071 1218 2105
rect 1252 2071 1354 2105
rect 1044 2037 1354 2071
rect 1044 2003 1146 2037
rect 1180 2003 1218 2037
rect 1252 2003 1354 2037
rect 1044 1969 1354 2003
rect 1044 1935 1146 1969
rect 1180 1935 1218 1969
rect 1252 1935 1354 1969
rect 1044 1901 1354 1935
rect 1044 1867 1146 1901
rect 1180 1867 1218 1901
rect 1252 1867 1354 1901
rect 1044 1833 1354 1867
rect 1044 1799 1146 1833
rect 1180 1799 1218 1833
rect 1252 1799 1354 1833
rect 1044 1765 1354 1799
rect 1044 1731 1146 1765
rect 1180 1731 1218 1765
rect 1252 1731 1354 1765
rect 1044 1697 1354 1731
rect 1044 1663 1146 1697
rect 1180 1663 1218 1697
rect 1252 1663 1354 1697
rect 1044 1629 1354 1663
rect 1044 1595 1146 1629
rect 1180 1595 1218 1629
rect 1252 1595 1354 1629
rect 1044 1561 1354 1595
rect 1044 1527 1146 1561
rect 1180 1527 1218 1561
rect 1252 1527 1354 1561
rect 1044 1457 1354 1527
rect 1474 2445 1625 2457
rect 1765 2445 1916 2457
rect 1474 2411 1576 2445
rect 1610 2411 1625 2445
rect 1765 2411 1780 2445
rect 1814 2411 1916 2445
rect 1474 2377 1625 2411
rect 1765 2377 1916 2411
rect 1474 2343 1576 2377
rect 1610 2343 1625 2377
rect 1765 2343 1780 2377
rect 1814 2343 1916 2377
rect 1474 2309 1625 2343
rect 1765 2309 1916 2343
rect 1474 2275 1576 2309
rect 1610 2275 1625 2309
rect 1765 2275 1780 2309
rect 1814 2275 1916 2309
rect 1474 2241 1625 2275
rect 1765 2241 1916 2275
rect 1474 2207 1576 2241
rect 1610 2207 1625 2241
rect 1765 2207 1780 2241
rect 1814 2207 1916 2241
rect 1474 2173 1625 2207
rect 1765 2173 1916 2207
rect 1474 2139 1576 2173
rect 1610 2139 1625 2173
rect 1765 2139 1780 2173
rect 1814 2139 1916 2173
rect 1474 2105 1625 2139
rect 1765 2105 1916 2139
rect 1474 2071 1576 2105
rect 1610 2071 1625 2105
rect 1765 2071 1780 2105
rect 1814 2071 1916 2105
rect 1474 2037 1625 2071
rect 1765 2037 1916 2071
rect 1474 2003 1576 2037
rect 1610 2003 1625 2037
rect 1765 2003 1780 2037
rect 1814 2003 1916 2037
rect 1474 1969 1625 2003
rect 1765 1969 1916 2003
rect 1474 1935 1576 1969
rect 1610 1935 1625 1969
rect 1765 1935 1780 1969
rect 1814 1935 1916 1969
rect 1474 1901 1625 1935
rect 1765 1901 1916 1935
rect 1474 1867 1576 1901
rect 1610 1867 1625 1901
rect 1765 1867 1780 1901
rect 1814 1867 1916 1901
rect 1474 1833 1625 1867
rect 1765 1833 1916 1867
rect 1474 1799 1576 1833
rect 1610 1799 1625 1833
rect 1765 1799 1780 1833
rect 1814 1799 1916 1833
rect 1474 1765 1625 1799
rect 1765 1765 1916 1799
rect 1474 1731 1576 1765
rect 1610 1731 1625 1765
rect 1765 1731 1780 1765
rect 1814 1731 1916 1765
rect 1474 1697 1625 1731
rect 1765 1697 1916 1731
rect 1474 1663 1576 1697
rect 1610 1663 1625 1697
rect 1765 1663 1780 1697
rect 1814 1663 1916 1697
rect 1474 1629 1625 1663
rect 1765 1629 1916 1663
rect 1474 1595 1576 1629
rect 1610 1595 1625 1629
rect 1765 1595 1780 1629
rect 1814 1595 1916 1629
rect 1474 1561 1625 1595
rect 1765 1561 1916 1595
rect 1474 1527 1576 1561
rect 1610 1527 1625 1561
rect 1765 1527 1780 1561
rect 1814 1527 1916 1561
rect 1474 1457 1625 1527
rect 1765 1457 1916 1527
rect 2036 2445 2346 2457
rect 2036 2411 2138 2445
rect 2172 2411 2210 2445
rect 2244 2411 2346 2445
rect 2036 2377 2346 2411
rect 2036 2343 2138 2377
rect 2172 2343 2210 2377
rect 2244 2343 2346 2377
rect 2036 2309 2346 2343
rect 2036 2275 2138 2309
rect 2172 2275 2210 2309
rect 2244 2275 2346 2309
rect 2036 2241 2346 2275
rect 2036 2207 2138 2241
rect 2172 2207 2210 2241
rect 2244 2207 2346 2241
rect 2036 2173 2346 2207
rect 2036 2139 2138 2173
rect 2172 2139 2210 2173
rect 2244 2139 2346 2173
rect 2036 2105 2346 2139
rect 2036 2071 2138 2105
rect 2172 2071 2210 2105
rect 2244 2071 2346 2105
rect 2036 2037 2346 2071
rect 2036 2003 2138 2037
rect 2172 2003 2210 2037
rect 2244 2003 2346 2037
rect 2036 1969 2346 2003
rect 2036 1935 2138 1969
rect 2172 1935 2210 1969
rect 2244 1935 2346 1969
rect 2036 1901 2346 1935
rect 2036 1867 2138 1901
rect 2172 1867 2210 1901
rect 2244 1867 2346 1901
rect 2036 1833 2346 1867
rect 2036 1799 2138 1833
rect 2172 1799 2210 1833
rect 2244 1799 2346 1833
rect 2036 1765 2346 1799
rect 2036 1731 2138 1765
rect 2172 1731 2210 1765
rect 2244 1731 2346 1765
rect 2036 1697 2346 1731
rect 2036 1663 2138 1697
rect 2172 1663 2210 1697
rect 2244 1663 2346 1697
rect 2036 1629 2346 1663
rect 2036 1595 2138 1629
rect 2172 1595 2210 1629
rect 2244 1595 2346 1629
rect 2036 1561 2346 1595
rect 2036 1527 2138 1561
rect 2172 1527 2210 1561
rect 2244 1527 2346 1561
rect 2036 1457 2346 1527
rect 2466 2445 2617 2457
rect 2757 2445 2908 2457
rect 2466 2411 2568 2445
rect 2602 2411 2617 2445
rect 2757 2411 2772 2445
rect 2806 2411 2908 2445
rect 2466 2377 2617 2411
rect 2757 2377 2908 2411
rect 2466 2343 2568 2377
rect 2602 2343 2617 2377
rect 2757 2343 2772 2377
rect 2806 2343 2908 2377
rect 2466 2309 2617 2343
rect 2757 2309 2908 2343
rect 2466 2275 2568 2309
rect 2602 2275 2617 2309
rect 2757 2275 2772 2309
rect 2806 2275 2908 2309
rect 2466 2241 2617 2275
rect 2757 2241 2908 2275
rect 2466 2207 2568 2241
rect 2602 2207 2617 2241
rect 2757 2207 2772 2241
rect 2806 2207 2908 2241
rect 2466 2173 2617 2207
rect 2757 2173 2908 2207
rect 2466 2139 2568 2173
rect 2602 2139 2617 2173
rect 2757 2139 2772 2173
rect 2806 2139 2908 2173
rect 2466 2105 2617 2139
rect 2757 2105 2908 2139
rect 2466 2071 2568 2105
rect 2602 2071 2617 2105
rect 2757 2071 2772 2105
rect 2806 2071 2908 2105
rect 2466 2037 2617 2071
rect 2757 2037 2908 2071
rect 2466 2003 2568 2037
rect 2602 2003 2617 2037
rect 2757 2003 2772 2037
rect 2806 2003 2908 2037
rect 2466 1969 2617 2003
rect 2757 1969 2908 2003
rect 2466 1935 2568 1969
rect 2602 1935 2617 1969
rect 2757 1935 2772 1969
rect 2806 1935 2908 1969
rect 2466 1901 2617 1935
rect 2757 1901 2908 1935
rect 2466 1867 2568 1901
rect 2602 1867 2617 1901
rect 2757 1867 2772 1901
rect 2806 1867 2908 1901
rect 2466 1833 2617 1867
rect 2757 1833 2908 1867
rect 2466 1799 2568 1833
rect 2602 1799 2617 1833
rect 2757 1799 2772 1833
rect 2806 1799 2908 1833
rect 2466 1765 2617 1799
rect 2757 1765 2908 1799
rect 2466 1731 2568 1765
rect 2602 1731 2617 1765
rect 2757 1731 2772 1765
rect 2806 1731 2908 1765
rect 2466 1697 2617 1731
rect 2757 1697 2908 1731
rect 2466 1663 2568 1697
rect 2602 1663 2617 1697
rect 2757 1663 2772 1697
rect 2806 1663 2908 1697
rect 2466 1629 2617 1663
rect 2757 1629 2908 1663
rect 2466 1595 2568 1629
rect 2602 1595 2617 1629
rect 2757 1595 2772 1629
rect 2806 1595 2908 1629
rect 2466 1561 2617 1595
rect 2757 1561 2908 1595
rect 2466 1527 2568 1561
rect 2602 1527 2617 1561
rect 2757 1527 2772 1561
rect 2806 1527 2908 1561
rect 2466 1457 2617 1527
rect 2757 1457 2908 1527
rect 3028 2445 3338 2457
rect 3028 2411 3130 2445
rect 3164 2411 3202 2445
rect 3236 2411 3338 2445
rect 3028 2377 3338 2411
rect 3028 2343 3130 2377
rect 3164 2343 3202 2377
rect 3236 2343 3338 2377
rect 3028 2309 3338 2343
rect 3028 2275 3130 2309
rect 3164 2275 3202 2309
rect 3236 2275 3338 2309
rect 3028 2241 3338 2275
rect 3028 2207 3130 2241
rect 3164 2207 3202 2241
rect 3236 2207 3338 2241
rect 3028 2173 3338 2207
rect 3028 2139 3130 2173
rect 3164 2139 3202 2173
rect 3236 2139 3338 2173
rect 3028 2105 3338 2139
rect 3028 2071 3130 2105
rect 3164 2071 3202 2105
rect 3236 2071 3338 2105
rect 3028 2037 3338 2071
rect 3028 2003 3130 2037
rect 3164 2003 3202 2037
rect 3236 2003 3338 2037
rect 3028 1969 3338 2003
rect 3028 1935 3130 1969
rect 3164 1935 3202 1969
rect 3236 1935 3338 1969
rect 3028 1901 3338 1935
rect 3028 1867 3130 1901
rect 3164 1867 3202 1901
rect 3236 1867 3338 1901
rect 3028 1833 3338 1867
rect 3028 1799 3130 1833
rect 3164 1799 3202 1833
rect 3236 1799 3338 1833
rect 3028 1765 3338 1799
rect 3028 1731 3130 1765
rect 3164 1731 3202 1765
rect 3236 1731 3338 1765
rect 3028 1697 3338 1731
rect 3028 1663 3130 1697
rect 3164 1663 3202 1697
rect 3236 1663 3338 1697
rect 3028 1629 3338 1663
rect 3028 1595 3130 1629
rect 3164 1595 3202 1629
rect 3236 1595 3338 1629
rect 3028 1561 3338 1595
rect 3028 1527 3130 1561
rect 3164 1527 3202 1561
rect 3236 1527 3338 1561
rect 3028 1457 3338 1527
rect 3458 2445 3609 2457
rect 3749 2445 3900 2457
rect 3458 2411 3560 2445
rect 3594 2411 3609 2445
rect 3749 2411 3764 2445
rect 3798 2411 3900 2445
rect 3458 2377 3609 2411
rect 3749 2377 3900 2411
rect 3458 2343 3560 2377
rect 3594 2343 3609 2377
rect 3749 2343 3764 2377
rect 3798 2343 3900 2377
rect 3458 2309 3609 2343
rect 3749 2309 3900 2343
rect 3458 2275 3560 2309
rect 3594 2275 3609 2309
rect 3749 2275 3764 2309
rect 3798 2275 3900 2309
rect 3458 2241 3609 2275
rect 3749 2241 3900 2275
rect 3458 2207 3560 2241
rect 3594 2207 3609 2241
rect 3749 2207 3764 2241
rect 3798 2207 3900 2241
rect 3458 2173 3609 2207
rect 3749 2173 3900 2207
rect 3458 2139 3560 2173
rect 3594 2139 3609 2173
rect 3749 2139 3764 2173
rect 3798 2139 3900 2173
rect 3458 2105 3609 2139
rect 3749 2105 3900 2139
rect 3458 2071 3560 2105
rect 3594 2071 3609 2105
rect 3749 2071 3764 2105
rect 3798 2071 3900 2105
rect 3458 2037 3609 2071
rect 3749 2037 3900 2071
rect 3458 2003 3560 2037
rect 3594 2003 3609 2037
rect 3749 2003 3764 2037
rect 3798 2003 3900 2037
rect 3458 1969 3609 2003
rect 3749 1969 3900 2003
rect 3458 1935 3560 1969
rect 3594 1935 3609 1969
rect 3749 1935 3764 1969
rect 3798 1935 3900 1969
rect 3458 1901 3609 1935
rect 3749 1901 3900 1935
rect 3458 1867 3560 1901
rect 3594 1867 3609 1901
rect 3749 1867 3764 1901
rect 3798 1867 3900 1901
rect 3458 1833 3609 1867
rect 3749 1833 3900 1867
rect 3458 1799 3560 1833
rect 3594 1799 3609 1833
rect 3749 1799 3764 1833
rect 3798 1799 3900 1833
rect 3458 1765 3609 1799
rect 3749 1765 3900 1799
rect 3458 1731 3560 1765
rect 3594 1731 3609 1765
rect 3749 1731 3764 1765
rect 3798 1731 3900 1765
rect 3458 1697 3609 1731
rect 3749 1697 3900 1731
rect 3458 1663 3560 1697
rect 3594 1663 3609 1697
rect 3749 1663 3764 1697
rect 3798 1663 3900 1697
rect 3458 1629 3609 1663
rect 3749 1629 3900 1663
rect 3458 1595 3560 1629
rect 3594 1595 3609 1629
rect 3749 1595 3764 1629
rect 3798 1595 3900 1629
rect 3458 1561 3609 1595
rect 3749 1561 3900 1595
rect 3458 1527 3560 1561
rect 3594 1527 3609 1561
rect 3749 1527 3764 1561
rect 3798 1527 3900 1561
rect 3458 1457 3609 1527
rect 3749 1457 3900 1527
rect 4020 2445 4330 2457
rect 4020 2411 4122 2445
rect 4156 2411 4194 2445
rect 4228 2411 4330 2445
rect 4020 2377 4330 2411
rect 4020 2343 4122 2377
rect 4156 2343 4194 2377
rect 4228 2343 4330 2377
rect 4020 2309 4330 2343
rect 4020 2275 4122 2309
rect 4156 2275 4194 2309
rect 4228 2275 4330 2309
rect 4020 2241 4330 2275
rect 4020 2207 4122 2241
rect 4156 2207 4194 2241
rect 4228 2207 4330 2241
rect 4020 2173 4330 2207
rect 4020 2139 4122 2173
rect 4156 2139 4194 2173
rect 4228 2139 4330 2173
rect 4020 2105 4330 2139
rect 4020 2071 4122 2105
rect 4156 2071 4194 2105
rect 4228 2071 4330 2105
rect 4020 2037 4330 2071
rect 4020 2003 4122 2037
rect 4156 2003 4194 2037
rect 4228 2003 4330 2037
rect 4020 1969 4330 2003
rect 4020 1935 4122 1969
rect 4156 1935 4194 1969
rect 4228 1935 4330 1969
rect 4020 1901 4330 1935
rect 4020 1867 4122 1901
rect 4156 1867 4194 1901
rect 4228 1867 4330 1901
rect 4020 1833 4330 1867
rect 4020 1799 4122 1833
rect 4156 1799 4194 1833
rect 4228 1799 4330 1833
rect 4020 1765 4330 1799
rect 4020 1731 4122 1765
rect 4156 1731 4194 1765
rect 4228 1731 4330 1765
rect 4020 1697 4330 1731
rect 4020 1663 4122 1697
rect 4156 1663 4194 1697
rect 4228 1663 4330 1697
rect 4020 1629 4330 1663
rect 4020 1595 4122 1629
rect 4156 1595 4194 1629
rect 4228 1595 4330 1629
rect 4020 1561 4330 1595
rect 4020 1527 4122 1561
rect 4156 1527 4194 1561
rect 4228 1527 4330 1561
rect 4020 1457 4330 1527
rect 4450 2445 4601 2457
rect 4741 2445 4892 2457
rect 4450 2411 4552 2445
rect 4586 2411 4601 2445
rect 4741 2411 4756 2445
rect 4790 2411 4892 2445
rect 4450 2377 4601 2411
rect 4741 2377 4892 2411
rect 4450 2343 4552 2377
rect 4586 2343 4601 2377
rect 4741 2343 4756 2377
rect 4790 2343 4892 2377
rect 4450 2309 4601 2343
rect 4741 2309 4892 2343
rect 4450 2275 4552 2309
rect 4586 2275 4601 2309
rect 4741 2275 4756 2309
rect 4790 2275 4892 2309
rect 4450 2241 4601 2275
rect 4741 2241 4892 2275
rect 4450 2207 4552 2241
rect 4586 2207 4601 2241
rect 4741 2207 4756 2241
rect 4790 2207 4892 2241
rect 4450 2173 4601 2207
rect 4741 2173 4892 2207
rect 4450 2139 4552 2173
rect 4586 2139 4601 2173
rect 4741 2139 4756 2173
rect 4790 2139 4892 2173
rect 4450 2105 4601 2139
rect 4741 2105 4892 2139
rect 4450 2071 4552 2105
rect 4586 2071 4601 2105
rect 4741 2071 4756 2105
rect 4790 2071 4892 2105
rect 4450 2037 4601 2071
rect 4741 2037 4892 2071
rect 4450 2003 4552 2037
rect 4586 2003 4601 2037
rect 4741 2003 4756 2037
rect 4790 2003 4892 2037
rect 4450 1969 4601 2003
rect 4741 1969 4892 2003
rect 4450 1935 4552 1969
rect 4586 1935 4601 1969
rect 4741 1935 4756 1969
rect 4790 1935 4892 1969
rect 4450 1901 4601 1935
rect 4741 1901 4892 1935
rect 4450 1867 4552 1901
rect 4586 1867 4601 1901
rect 4741 1867 4756 1901
rect 4790 1867 4892 1901
rect 4450 1833 4601 1867
rect 4741 1833 4892 1867
rect 4450 1799 4552 1833
rect 4586 1799 4601 1833
rect 4741 1799 4756 1833
rect 4790 1799 4892 1833
rect 4450 1765 4601 1799
rect 4741 1765 4892 1799
rect 4450 1731 4552 1765
rect 4586 1731 4601 1765
rect 4741 1731 4756 1765
rect 4790 1731 4892 1765
rect 4450 1697 4601 1731
rect 4741 1697 4892 1731
rect 4450 1663 4552 1697
rect 4586 1663 4601 1697
rect 4741 1663 4756 1697
rect 4790 1663 4892 1697
rect 4450 1629 4601 1663
rect 4741 1629 4892 1663
rect 4450 1595 4552 1629
rect 4586 1595 4601 1629
rect 4741 1595 4756 1629
rect 4790 1595 4892 1629
rect 4450 1561 4601 1595
rect 4741 1561 4892 1595
rect 4450 1527 4552 1561
rect 4586 1527 4601 1561
rect 4741 1527 4756 1561
rect 4790 1527 4892 1561
rect 4450 1457 4601 1527
rect 4741 1457 4892 1527
rect 5012 2445 5322 2457
rect 5012 2411 5114 2445
rect 5148 2411 5186 2445
rect 5220 2411 5322 2445
rect 5012 2377 5322 2411
rect 5012 2343 5114 2377
rect 5148 2343 5186 2377
rect 5220 2343 5322 2377
rect 5012 2309 5322 2343
rect 5012 2275 5114 2309
rect 5148 2275 5186 2309
rect 5220 2275 5322 2309
rect 5012 2241 5322 2275
rect 5012 2207 5114 2241
rect 5148 2207 5186 2241
rect 5220 2207 5322 2241
rect 5012 2173 5322 2207
rect 5012 2139 5114 2173
rect 5148 2139 5186 2173
rect 5220 2139 5322 2173
rect 5012 2105 5322 2139
rect 5012 2071 5114 2105
rect 5148 2071 5186 2105
rect 5220 2071 5322 2105
rect 5012 2037 5322 2071
rect 5012 2003 5114 2037
rect 5148 2003 5186 2037
rect 5220 2003 5322 2037
rect 5012 1969 5322 2003
rect 5012 1935 5114 1969
rect 5148 1935 5186 1969
rect 5220 1935 5322 1969
rect 5012 1901 5322 1935
rect 5012 1867 5114 1901
rect 5148 1867 5186 1901
rect 5220 1867 5322 1901
rect 5012 1833 5322 1867
rect 5012 1799 5114 1833
rect 5148 1799 5186 1833
rect 5220 1799 5322 1833
rect 5012 1765 5322 1799
rect 5012 1731 5114 1765
rect 5148 1731 5186 1765
rect 5220 1731 5322 1765
rect 5012 1697 5322 1731
rect 5012 1663 5114 1697
rect 5148 1663 5186 1697
rect 5220 1663 5322 1697
rect 5012 1629 5322 1663
rect 5012 1595 5114 1629
rect 5148 1595 5186 1629
rect 5220 1595 5322 1629
rect 5012 1561 5322 1595
rect 5012 1527 5114 1561
rect 5148 1527 5186 1561
rect 5220 1527 5322 1561
rect 5012 1457 5322 1527
rect 5442 2445 5593 2457
rect 5733 2445 5884 2457
rect 5442 2411 5544 2445
rect 5578 2411 5593 2445
rect 5733 2411 5748 2445
rect 5782 2411 5884 2445
rect 5442 2377 5593 2411
rect 5733 2377 5884 2411
rect 5442 2343 5544 2377
rect 5578 2343 5593 2377
rect 5733 2343 5748 2377
rect 5782 2343 5884 2377
rect 5442 2309 5593 2343
rect 5733 2309 5884 2343
rect 5442 2275 5544 2309
rect 5578 2275 5593 2309
rect 5733 2275 5748 2309
rect 5782 2275 5884 2309
rect 5442 2241 5593 2275
rect 5733 2241 5884 2275
rect 5442 2207 5544 2241
rect 5578 2207 5593 2241
rect 5733 2207 5748 2241
rect 5782 2207 5884 2241
rect 5442 2173 5593 2207
rect 5733 2173 5884 2207
rect 5442 2139 5544 2173
rect 5578 2139 5593 2173
rect 5733 2139 5748 2173
rect 5782 2139 5884 2173
rect 5442 2105 5593 2139
rect 5733 2105 5884 2139
rect 5442 2071 5544 2105
rect 5578 2071 5593 2105
rect 5733 2071 5748 2105
rect 5782 2071 5884 2105
rect 5442 2037 5593 2071
rect 5733 2037 5884 2071
rect 5442 2003 5544 2037
rect 5578 2003 5593 2037
rect 5733 2003 5748 2037
rect 5782 2003 5884 2037
rect 5442 1969 5593 2003
rect 5733 1969 5884 2003
rect 5442 1935 5544 1969
rect 5578 1935 5593 1969
rect 5733 1935 5748 1969
rect 5782 1935 5884 1969
rect 5442 1901 5593 1935
rect 5733 1901 5884 1935
rect 5442 1867 5544 1901
rect 5578 1867 5593 1901
rect 5733 1867 5748 1901
rect 5782 1867 5884 1901
rect 5442 1833 5593 1867
rect 5733 1833 5884 1867
rect 5442 1799 5544 1833
rect 5578 1799 5593 1833
rect 5733 1799 5748 1833
rect 5782 1799 5884 1833
rect 5442 1765 5593 1799
rect 5733 1765 5884 1799
rect 5442 1731 5544 1765
rect 5578 1731 5593 1765
rect 5733 1731 5748 1765
rect 5782 1731 5884 1765
rect 5442 1697 5593 1731
rect 5733 1697 5884 1731
rect 5442 1663 5544 1697
rect 5578 1663 5593 1697
rect 5733 1663 5748 1697
rect 5782 1663 5884 1697
rect 5442 1629 5593 1663
rect 5733 1629 5884 1663
rect 5442 1595 5544 1629
rect 5578 1595 5593 1629
rect 5733 1595 5748 1629
rect 5782 1595 5884 1629
rect 5442 1561 5593 1595
rect 5733 1561 5884 1595
rect 5442 1527 5544 1561
rect 5578 1527 5593 1561
rect 5733 1527 5748 1561
rect 5782 1527 5884 1561
rect 5442 1457 5593 1527
rect 5733 1457 5884 1527
rect 6004 2445 6314 2457
rect 6004 2411 6106 2445
rect 6140 2411 6178 2445
rect 6212 2411 6314 2445
rect 6004 2377 6314 2411
rect 6004 2343 6106 2377
rect 6140 2343 6178 2377
rect 6212 2343 6314 2377
rect 6004 2309 6314 2343
rect 6004 2275 6106 2309
rect 6140 2275 6178 2309
rect 6212 2275 6314 2309
rect 6004 2241 6314 2275
rect 6004 2207 6106 2241
rect 6140 2207 6178 2241
rect 6212 2207 6314 2241
rect 6004 2173 6314 2207
rect 6004 2139 6106 2173
rect 6140 2139 6178 2173
rect 6212 2139 6314 2173
rect 6004 2105 6314 2139
rect 6004 2071 6106 2105
rect 6140 2071 6178 2105
rect 6212 2071 6314 2105
rect 6004 2037 6314 2071
rect 6004 2003 6106 2037
rect 6140 2003 6178 2037
rect 6212 2003 6314 2037
rect 6004 1969 6314 2003
rect 6004 1935 6106 1969
rect 6140 1935 6178 1969
rect 6212 1935 6314 1969
rect 6004 1901 6314 1935
rect 6004 1867 6106 1901
rect 6140 1867 6178 1901
rect 6212 1867 6314 1901
rect 6004 1833 6314 1867
rect 6004 1799 6106 1833
rect 6140 1799 6178 1833
rect 6212 1799 6314 1833
rect 6004 1765 6314 1799
rect 6004 1731 6106 1765
rect 6140 1731 6178 1765
rect 6212 1731 6314 1765
rect 6004 1697 6314 1731
rect 6004 1663 6106 1697
rect 6140 1663 6178 1697
rect 6212 1663 6314 1697
rect 6004 1629 6314 1663
rect 6004 1595 6106 1629
rect 6140 1595 6178 1629
rect 6212 1595 6314 1629
rect 6004 1561 6314 1595
rect 6004 1527 6106 1561
rect 6140 1527 6178 1561
rect 6212 1527 6314 1561
rect 6004 1457 6314 1527
rect 6434 2445 6585 2457
rect 6725 2445 6876 2457
rect 6434 2411 6536 2445
rect 6570 2411 6585 2445
rect 6725 2411 6740 2445
rect 6774 2411 6876 2445
rect 6434 2377 6585 2411
rect 6725 2377 6876 2411
rect 6434 2343 6536 2377
rect 6570 2343 6585 2377
rect 6725 2343 6740 2377
rect 6774 2343 6876 2377
rect 6434 2309 6585 2343
rect 6725 2309 6876 2343
rect 6434 2275 6536 2309
rect 6570 2275 6585 2309
rect 6725 2275 6740 2309
rect 6774 2275 6876 2309
rect 6434 2241 6585 2275
rect 6725 2241 6876 2275
rect 6434 2207 6536 2241
rect 6570 2207 6585 2241
rect 6725 2207 6740 2241
rect 6774 2207 6876 2241
rect 6434 2173 6585 2207
rect 6725 2173 6876 2207
rect 6434 2139 6536 2173
rect 6570 2139 6585 2173
rect 6725 2139 6740 2173
rect 6774 2139 6876 2173
rect 6434 2105 6585 2139
rect 6725 2105 6876 2139
rect 6434 2071 6536 2105
rect 6570 2071 6585 2105
rect 6725 2071 6740 2105
rect 6774 2071 6876 2105
rect 6434 2037 6585 2071
rect 6725 2037 6876 2071
rect 6434 2003 6536 2037
rect 6570 2003 6585 2037
rect 6725 2003 6740 2037
rect 6774 2003 6876 2037
rect 6434 1969 6585 2003
rect 6725 1969 6876 2003
rect 6434 1935 6536 1969
rect 6570 1935 6585 1969
rect 6725 1935 6740 1969
rect 6774 1935 6876 1969
rect 6434 1901 6585 1935
rect 6725 1901 6876 1935
rect 6434 1867 6536 1901
rect 6570 1867 6585 1901
rect 6725 1867 6740 1901
rect 6774 1867 6876 1901
rect 6434 1833 6585 1867
rect 6725 1833 6876 1867
rect 6434 1799 6536 1833
rect 6570 1799 6585 1833
rect 6725 1799 6740 1833
rect 6774 1799 6876 1833
rect 6434 1765 6585 1799
rect 6725 1765 6876 1799
rect 6434 1731 6536 1765
rect 6570 1731 6585 1765
rect 6725 1731 6740 1765
rect 6774 1731 6876 1765
rect 6434 1697 6585 1731
rect 6725 1697 6876 1731
rect 6434 1663 6536 1697
rect 6570 1663 6585 1697
rect 6725 1663 6740 1697
rect 6774 1663 6876 1697
rect 6434 1629 6585 1663
rect 6725 1629 6876 1663
rect 6434 1595 6536 1629
rect 6570 1595 6585 1629
rect 6725 1595 6740 1629
rect 6774 1595 6876 1629
rect 6434 1561 6585 1595
rect 6725 1561 6876 1595
rect 6434 1527 6536 1561
rect 6570 1527 6585 1561
rect 6725 1527 6740 1561
rect 6774 1527 6876 1561
rect 6434 1457 6585 1527
rect 6725 1457 6876 1527
rect 6996 2445 7306 2457
rect 6996 2411 7098 2445
rect 7132 2411 7170 2445
rect 7204 2411 7306 2445
rect 6996 2377 7306 2411
rect 6996 2343 7098 2377
rect 7132 2343 7170 2377
rect 7204 2343 7306 2377
rect 6996 2309 7306 2343
rect 6996 2275 7098 2309
rect 7132 2275 7170 2309
rect 7204 2275 7306 2309
rect 6996 2241 7306 2275
rect 6996 2207 7098 2241
rect 7132 2207 7170 2241
rect 7204 2207 7306 2241
rect 6996 2173 7306 2207
rect 6996 2139 7098 2173
rect 7132 2139 7170 2173
rect 7204 2139 7306 2173
rect 6996 2105 7306 2139
rect 6996 2071 7098 2105
rect 7132 2071 7170 2105
rect 7204 2071 7306 2105
rect 6996 2037 7306 2071
rect 6996 2003 7098 2037
rect 7132 2003 7170 2037
rect 7204 2003 7306 2037
rect 6996 1969 7306 2003
rect 6996 1935 7098 1969
rect 7132 1935 7170 1969
rect 7204 1935 7306 1969
rect 6996 1901 7306 1935
rect 6996 1867 7098 1901
rect 7132 1867 7170 1901
rect 7204 1867 7306 1901
rect 6996 1833 7306 1867
rect 6996 1799 7098 1833
rect 7132 1799 7170 1833
rect 7204 1799 7306 1833
rect 6996 1765 7306 1799
rect 6996 1731 7098 1765
rect 7132 1731 7170 1765
rect 7204 1731 7306 1765
rect 6996 1697 7306 1731
rect 6996 1663 7098 1697
rect 7132 1663 7170 1697
rect 7204 1663 7306 1697
rect 6996 1629 7306 1663
rect 6996 1595 7098 1629
rect 7132 1595 7170 1629
rect 7204 1595 7306 1629
rect 6996 1561 7306 1595
rect 6996 1527 7098 1561
rect 7132 1527 7170 1561
rect 7204 1527 7306 1561
rect 6996 1457 7306 1527
rect 7426 2445 7577 2457
rect 7717 2445 7868 2457
rect 7426 2411 7528 2445
rect 7562 2411 7577 2445
rect 7717 2411 7732 2445
rect 7766 2411 7868 2445
rect 7426 2377 7577 2411
rect 7717 2377 7868 2411
rect 7426 2343 7528 2377
rect 7562 2343 7577 2377
rect 7717 2343 7732 2377
rect 7766 2343 7868 2377
rect 7426 2309 7577 2343
rect 7717 2309 7868 2343
rect 7426 2275 7528 2309
rect 7562 2275 7577 2309
rect 7717 2275 7732 2309
rect 7766 2275 7868 2309
rect 7426 2241 7577 2275
rect 7717 2241 7868 2275
rect 7426 2207 7528 2241
rect 7562 2207 7577 2241
rect 7717 2207 7732 2241
rect 7766 2207 7868 2241
rect 7426 2173 7577 2207
rect 7717 2173 7868 2207
rect 7426 2139 7528 2173
rect 7562 2139 7577 2173
rect 7717 2139 7732 2173
rect 7766 2139 7868 2173
rect 7426 2105 7577 2139
rect 7717 2105 7868 2139
rect 7426 2071 7528 2105
rect 7562 2071 7577 2105
rect 7717 2071 7732 2105
rect 7766 2071 7868 2105
rect 7426 2037 7577 2071
rect 7717 2037 7868 2071
rect 7426 2003 7528 2037
rect 7562 2003 7577 2037
rect 7717 2003 7732 2037
rect 7766 2003 7868 2037
rect 7426 1969 7577 2003
rect 7717 1969 7868 2003
rect 7426 1935 7528 1969
rect 7562 1935 7577 1969
rect 7717 1935 7732 1969
rect 7766 1935 7868 1969
rect 7426 1901 7577 1935
rect 7717 1901 7868 1935
rect 7426 1867 7528 1901
rect 7562 1867 7577 1901
rect 7717 1867 7732 1901
rect 7766 1867 7868 1901
rect 7426 1833 7577 1867
rect 7717 1833 7868 1867
rect 7426 1799 7528 1833
rect 7562 1799 7577 1833
rect 7717 1799 7732 1833
rect 7766 1799 7868 1833
rect 7426 1765 7577 1799
rect 7717 1765 7868 1799
rect 7426 1731 7528 1765
rect 7562 1731 7577 1765
rect 7717 1731 7732 1765
rect 7766 1731 7868 1765
rect 7426 1697 7577 1731
rect 7717 1697 7868 1731
rect 7426 1663 7528 1697
rect 7562 1663 7577 1697
rect 7717 1663 7732 1697
rect 7766 1663 7868 1697
rect 7426 1629 7577 1663
rect 7717 1629 7868 1663
rect 7426 1595 7528 1629
rect 7562 1595 7577 1629
rect 7717 1595 7732 1629
rect 7766 1595 7868 1629
rect 7426 1561 7577 1595
rect 7717 1561 7868 1595
rect 7426 1527 7528 1561
rect 7562 1527 7577 1561
rect 7717 1527 7732 1561
rect 7766 1527 7868 1561
rect 7426 1457 7577 1527
rect 7717 1457 7868 1527
rect 7988 2445 8298 2457
rect 7988 2411 8090 2445
rect 8124 2411 8162 2445
rect 8196 2411 8298 2445
rect 7988 2377 8298 2411
rect 7988 2343 8090 2377
rect 8124 2343 8162 2377
rect 8196 2343 8298 2377
rect 7988 2309 8298 2343
rect 7988 2275 8090 2309
rect 8124 2275 8162 2309
rect 8196 2275 8298 2309
rect 7988 2241 8298 2275
rect 7988 2207 8090 2241
rect 8124 2207 8162 2241
rect 8196 2207 8298 2241
rect 7988 2173 8298 2207
rect 7988 2139 8090 2173
rect 8124 2139 8162 2173
rect 8196 2139 8298 2173
rect 7988 2105 8298 2139
rect 7988 2071 8090 2105
rect 8124 2071 8162 2105
rect 8196 2071 8298 2105
rect 7988 2037 8298 2071
rect 7988 2003 8090 2037
rect 8124 2003 8162 2037
rect 8196 2003 8298 2037
rect 7988 1969 8298 2003
rect 7988 1935 8090 1969
rect 8124 1935 8162 1969
rect 8196 1935 8298 1969
rect 7988 1901 8298 1935
rect 7988 1867 8090 1901
rect 8124 1867 8162 1901
rect 8196 1867 8298 1901
rect 7988 1833 8298 1867
rect 7988 1799 8090 1833
rect 8124 1799 8162 1833
rect 8196 1799 8298 1833
rect 7988 1765 8298 1799
rect 7988 1731 8090 1765
rect 8124 1731 8162 1765
rect 8196 1731 8298 1765
rect 7988 1697 8298 1731
rect 7988 1663 8090 1697
rect 8124 1663 8162 1697
rect 8196 1663 8298 1697
rect 7988 1629 8298 1663
rect 7988 1595 8090 1629
rect 8124 1595 8162 1629
rect 8196 1595 8298 1629
rect 7988 1561 8298 1595
rect 7988 1527 8090 1561
rect 8124 1527 8162 1561
rect 8196 1527 8298 1561
rect 7988 1457 8298 1527
rect 8418 2445 8569 2457
rect 8709 2445 8860 2457
rect 8418 2411 8520 2445
rect 8554 2411 8569 2445
rect 8709 2411 8724 2445
rect 8758 2411 8860 2445
rect 8418 2377 8569 2411
rect 8709 2377 8860 2411
rect 8418 2343 8520 2377
rect 8554 2343 8569 2377
rect 8709 2343 8724 2377
rect 8758 2343 8860 2377
rect 8418 2309 8569 2343
rect 8709 2309 8860 2343
rect 8418 2275 8520 2309
rect 8554 2275 8569 2309
rect 8709 2275 8724 2309
rect 8758 2275 8860 2309
rect 8418 2241 8569 2275
rect 8709 2241 8860 2275
rect 8418 2207 8520 2241
rect 8554 2207 8569 2241
rect 8709 2207 8724 2241
rect 8758 2207 8860 2241
rect 8418 2173 8569 2207
rect 8709 2173 8860 2207
rect 8418 2139 8520 2173
rect 8554 2139 8569 2173
rect 8709 2139 8724 2173
rect 8758 2139 8860 2173
rect 8418 2105 8569 2139
rect 8709 2105 8860 2139
rect 8418 2071 8520 2105
rect 8554 2071 8569 2105
rect 8709 2071 8724 2105
rect 8758 2071 8860 2105
rect 8418 2037 8569 2071
rect 8709 2037 8860 2071
rect 8418 2003 8520 2037
rect 8554 2003 8569 2037
rect 8709 2003 8724 2037
rect 8758 2003 8860 2037
rect 8418 1969 8569 2003
rect 8709 1969 8860 2003
rect 8418 1935 8520 1969
rect 8554 1935 8569 1969
rect 8709 1935 8724 1969
rect 8758 1935 8860 1969
rect 8418 1901 8569 1935
rect 8709 1901 8860 1935
rect 8418 1867 8520 1901
rect 8554 1867 8569 1901
rect 8709 1867 8724 1901
rect 8758 1867 8860 1901
rect 8418 1833 8569 1867
rect 8709 1833 8860 1867
rect 8418 1799 8520 1833
rect 8554 1799 8569 1833
rect 8709 1799 8724 1833
rect 8758 1799 8860 1833
rect 8418 1765 8569 1799
rect 8709 1765 8860 1799
rect 8418 1731 8520 1765
rect 8554 1731 8569 1765
rect 8709 1731 8724 1765
rect 8758 1731 8860 1765
rect 8418 1697 8569 1731
rect 8709 1697 8860 1731
rect 8418 1663 8520 1697
rect 8554 1663 8569 1697
rect 8709 1663 8724 1697
rect 8758 1663 8860 1697
rect 8418 1629 8569 1663
rect 8709 1629 8860 1663
rect 8418 1595 8520 1629
rect 8554 1595 8569 1629
rect 8709 1595 8724 1629
rect 8758 1595 8860 1629
rect 8418 1561 8569 1595
rect 8709 1561 8860 1595
rect 8418 1527 8520 1561
rect 8554 1527 8569 1561
rect 8709 1527 8724 1561
rect 8758 1527 8860 1561
rect 8418 1457 8569 1527
rect 8709 1457 8860 1527
rect 8980 2445 9290 2457
rect 8980 2411 9082 2445
rect 9116 2411 9154 2445
rect 9188 2411 9290 2445
rect 8980 2377 9290 2411
rect 8980 2343 9082 2377
rect 9116 2343 9154 2377
rect 9188 2343 9290 2377
rect 8980 2309 9290 2343
rect 8980 2275 9082 2309
rect 9116 2275 9154 2309
rect 9188 2275 9290 2309
rect 8980 2241 9290 2275
rect 8980 2207 9082 2241
rect 9116 2207 9154 2241
rect 9188 2207 9290 2241
rect 8980 2173 9290 2207
rect 8980 2139 9082 2173
rect 9116 2139 9154 2173
rect 9188 2139 9290 2173
rect 8980 2105 9290 2139
rect 8980 2071 9082 2105
rect 9116 2071 9154 2105
rect 9188 2071 9290 2105
rect 8980 2037 9290 2071
rect 8980 2003 9082 2037
rect 9116 2003 9154 2037
rect 9188 2003 9290 2037
rect 8980 1969 9290 2003
rect 8980 1935 9082 1969
rect 9116 1935 9154 1969
rect 9188 1935 9290 1969
rect 8980 1901 9290 1935
rect 8980 1867 9082 1901
rect 9116 1867 9154 1901
rect 9188 1867 9290 1901
rect 8980 1833 9290 1867
rect 8980 1799 9082 1833
rect 9116 1799 9154 1833
rect 9188 1799 9290 1833
rect 8980 1765 9290 1799
rect 8980 1731 9082 1765
rect 9116 1731 9154 1765
rect 9188 1731 9290 1765
rect 8980 1697 9290 1731
rect 8980 1663 9082 1697
rect 9116 1663 9154 1697
rect 9188 1663 9290 1697
rect 8980 1629 9290 1663
rect 8980 1595 9082 1629
rect 9116 1595 9154 1629
rect 9188 1595 9290 1629
rect 8980 1561 9290 1595
rect 8980 1527 9082 1561
rect 9116 1527 9154 1561
rect 9188 1527 9290 1561
rect 8980 1457 9290 1527
rect 9410 2445 9561 2457
rect 9701 2445 9852 2457
rect 9410 2411 9512 2445
rect 9546 2411 9561 2445
rect 9701 2411 9716 2445
rect 9750 2411 9852 2445
rect 9410 2377 9561 2411
rect 9701 2377 9852 2411
rect 9410 2343 9512 2377
rect 9546 2343 9561 2377
rect 9701 2343 9716 2377
rect 9750 2343 9852 2377
rect 9410 2309 9561 2343
rect 9701 2309 9852 2343
rect 9410 2275 9512 2309
rect 9546 2275 9561 2309
rect 9701 2275 9716 2309
rect 9750 2275 9852 2309
rect 9410 2241 9561 2275
rect 9701 2241 9852 2275
rect 9410 2207 9512 2241
rect 9546 2207 9561 2241
rect 9701 2207 9716 2241
rect 9750 2207 9852 2241
rect 9410 2173 9561 2207
rect 9701 2173 9852 2207
rect 9410 2139 9512 2173
rect 9546 2139 9561 2173
rect 9701 2139 9716 2173
rect 9750 2139 9852 2173
rect 9410 2105 9561 2139
rect 9701 2105 9852 2139
rect 9410 2071 9512 2105
rect 9546 2071 9561 2105
rect 9701 2071 9716 2105
rect 9750 2071 9852 2105
rect 9410 2037 9561 2071
rect 9701 2037 9852 2071
rect 9410 2003 9512 2037
rect 9546 2003 9561 2037
rect 9701 2003 9716 2037
rect 9750 2003 9852 2037
rect 9410 1969 9561 2003
rect 9701 1969 9852 2003
rect 9410 1935 9512 1969
rect 9546 1935 9561 1969
rect 9701 1935 9716 1969
rect 9750 1935 9852 1969
rect 9410 1901 9561 1935
rect 9701 1901 9852 1935
rect 9410 1867 9512 1901
rect 9546 1867 9561 1901
rect 9701 1867 9716 1901
rect 9750 1867 9852 1901
rect 9410 1833 9561 1867
rect 9701 1833 9852 1867
rect 9410 1799 9512 1833
rect 9546 1799 9561 1833
rect 9701 1799 9716 1833
rect 9750 1799 9852 1833
rect 9410 1765 9561 1799
rect 9701 1765 9852 1799
rect 9410 1731 9512 1765
rect 9546 1731 9561 1765
rect 9701 1731 9716 1765
rect 9750 1731 9852 1765
rect 9410 1697 9561 1731
rect 9701 1697 9852 1731
rect 9410 1663 9512 1697
rect 9546 1663 9561 1697
rect 9701 1663 9716 1697
rect 9750 1663 9852 1697
rect 9410 1629 9561 1663
rect 9701 1629 9852 1663
rect 9410 1595 9512 1629
rect 9546 1595 9561 1629
rect 9701 1595 9716 1629
rect 9750 1595 9852 1629
rect 9410 1561 9561 1595
rect 9701 1561 9852 1595
rect 9410 1527 9512 1561
rect 9546 1527 9561 1561
rect 9701 1527 9716 1561
rect 9750 1527 9852 1561
rect 9410 1457 9561 1527
rect 9701 1457 9852 1527
rect 9972 2445 10282 2457
rect 9972 2411 10074 2445
rect 10108 2411 10146 2445
rect 10180 2411 10282 2445
rect 9972 2377 10282 2411
rect 9972 2343 10074 2377
rect 10108 2343 10146 2377
rect 10180 2343 10282 2377
rect 9972 2309 10282 2343
rect 9972 2275 10074 2309
rect 10108 2275 10146 2309
rect 10180 2275 10282 2309
rect 9972 2241 10282 2275
rect 9972 2207 10074 2241
rect 10108 2207 10146 2241
rect 10180 2207 10282 2241
rect 9972 2173 10282 2207
rect 9972 2139 10074 2173
rect 10108 2139 10146 2173
rect 10180 2139 10282 2173
rect 9972 2105 10282 2139
rect 9972 2071 10074 2105
rect 10108 2071 10146 2105
rect 10180 2071 10282 2105
rect 9972 2037 10282 2071
rect 9972 2003 10074 2037
rect 10108 2003 10146 2037
rect 10180 2003 10282 2037
rect 9972 1969 10282 2003
rect 9972 1935 10074 1969
rect 10108 1935 10146 1969
rect 10180 1935 10282 1969
rect 9972 1901 10282 1935
rect 9972 1867 10074 1901
rect 10108 1867 10146 1901
rect 10180 1867 10282 1901
rect 9972 1833 10282 1867
rect 9972 1799 10074 1833
rect 10108 1799 10146 1833
rect 10180 1799 10282 1833
rect 9972 1765 10282 1799
rect 9972 1731 10074 1765
rect 10108 1731 10146 1765
rect 10180 1731 10282 1765
rect 9972 1697 10282 1731
rect 9972 1663 10074 1697
rect 10108 1663 10146 1697
rect 10180 1663 10282 1697
rect 9972 1629 10282 1663
rect 9972 1595 10074 1629
rect 10108 1595 10146 1629
rect 10180 1595 10282 1629
rect 9972 1561 10282 1595
rect 9972 1527 10074 1561
rect 10108 1527 10146 1561
rect 10180 1527 10282 1561
rect 9972 1457 10282 1527
rect 10402 2445 10553 2457
rect 10693 2445 10844 2457
rect 10402 2411 10504 2445
rect 10538 2411 10553 2445
rect 10693 2411 10708 2445
rect 10742 2411 10844 2445
rect 10402 2377 10553 2411
rect 10693 2377 10844 2411
rect 10402 2343 10504 2377
rect 10538 2343 10553 2377
rect 10693 2343 10708 2377
rect 10742 2343 10844 2377
rect 10402 2309 10553 2343
rect 10693 2309 10844 2343
rect 10402 2275 10504 2309
rect 10538 2275 10553 2309
rect 10693 2275 10708 2309
rect 10742 2275 10844 2309
rect 10402 2241 10553 2275
rect 10693 2241 10844 2275
rect 10402 2207 10504 2241
rect 10538 2207 10553 2241
rect 10693 2207 10708 2241
rect 10742 2207 10844 2241
rect 10402 2173 10553 2207
rect 10693 2173 10844 2207
rect 10402 2139 10504 2173
rect 10538 2139 10553 2173
rect 10693 2139 10708 2173
rect 10742 2139 10844 2173
rect 10402 2105 10553 2139
rect 10693 2105 10844 2139
rect 10402 2071 10504 2105
rect 10538 2071 10553 2105
rect 10693 2071 10708 2105
rect 10742 2071 10844 2105
rect 10402 2037 10553 2071
rect 10693 2037 10844 2071
rect 10402 2003 10504 2037
rect 10538 2003 10553 2037
rect 10693 2003 10708 2037
rect 10742 2003 10844 2037
rect 10402 1969 10553 2003
rect 10693 1969 10844 2003
rect 10402 1935 10504 1969
rect 10538 1935 10553 1969
rect 10693 1935 10708 1969
rect 10742 1935 10844 1969
rect 10402 1901 10553 1935
rect 10693 1901 10844 1935
rect 10402 1867 10504 1901
rect 10538 1867 10553 1901
rect 10693 1867 10708 1901
rect 10742 1867 10844 1901
rect 10402 1833 10553 1867
rect 10693 1833 10844 1867
rect 10402 1799 10504 1833
rect 10538 1799 10553 1833
rect 10693 1799 10708 1833
rect 10742 1799 10844 1833
rect 10402 1765 10553 1799
rect 10693 1765 10844 1799
rect 10402 1731 10504 1765
rect 10538 1731 10553 1765
rect 10693 1731 10708 1765
rect 10742 1731 10844 1765
rect 10402 1697 10553 1731
rect 10693 1697 10844 1731
rect 10402 1663 10504 1697
rect 10538 1663 10553 1697
rect 10693 1663 10708 1697
rect 10742 1663 10844 1697
rect 10402 1629 10553 1663
rect 10693 1629 10844 1663
rect 10402 1595 10504 1629
rect 10538 1595 10553 1629
rect 10693 1595 10708 1629
rect 10742 1595 10844 1629
rect 10402 1561 10553 1595
rect 10693 1561 10844 1595
rect 10402 1527 10504 1561
rect 10538 1527 10553 1561
rect 10693 1527 10708 1561
rect 10742 1527 10844 1561
rect 10402 1457 10553 1527
rect 10693 1457 10844 1527
rect 10964 2445 11274 2457
rect 10964 2411 11066 2445
rect 11100 2411 11138 2445
rect 11172 2411 11274 2445
rect 10964 2377 11274 2411
rect 10964 2343 11066 2377
rect 11100 2343 11138 2377
rect 11172 2343 11274 2377
rect 10964 2309 11274 2343
rect 10964 2275 11066 2309
rect 11100 2275 11138 2309
rect 11172 2275 11274 2309
rect 10964 2241 11274 2275
rect 10964 2207 11066 2241
rect 11100 2207 11138 2241
rect 11172 2207 11274 2241
rect 10964 2173 11274 2207
rect 10964 2139 11066 2173
rect 11100 2139 11138 2173
rect 11172 2139 11274 2173
rect 10964 2105 11274 2139
rect 10964 2071 11066 2105
rect 11100 2071 11138 2105
rect 11172 2071 11274 2105
rect 10964 2037 11274 2071
rect 10964 2003 11066 2037
rect 11100 2003 11138 2037
rect 11172 2003 11274 2037
rect 10964 1969 11274 2003
rect 10964 1935 11066 1969
rect 11100 1935 11138 1969
rect 11172 1935 11274 1969
rect 10964 1901 11274 1935
rect 10964 1867 11066 1901
rect 11100 1867 11138 1901
rect 11172 1867 11274 1901
rect 10964 1833 11274 1867
rect 10964 1799 11066 1833
rect 11100 1799 11138 1833
rect 11172 1799 11274 1833
rect 10964 1765 11274 1799
rect 10964 1731 11066 1765
rect 11100 1731 11138 1765
rect 11172 1731 11274 1765
rect 10964 1697 11274 1731
rect 10964 1663 11066 1697
rect 11100 1663 11138 1697
rect 11172 1663 11274 1697
rect 10964 1629 11274 1663
rect 10964 1595 11066 1629
rect 11100 1595 11138 1629
rect 11172 1595 11274 1629
rect 10964 1561 11274 1595
rect 10964 1527 11066 1561
rect 11100 1527 11138 1561
rect 11172 1527 11274 1561
rect 10964 1457 11274 1527
rect 11394 2445 11545 2457
rect 11685 2445 11836 2457
rect 11394 2411 11496 2445
rect 11530 2411 11545 2445
rect 11685 2411 11700 2445
rect 11734 2411 11836 2445
rect 11394 2377 11545 2411
rect 11685 2377 11836 2411
rect 11394 2343 11496 2377
rect 11530 2343 11545 2377
rect 11685 2343 11700 2377
rect 11734 2343 11836 2377
rect 11394 2309 11545 2343
rect 11685 2309 11836 2343
rect 11394 2275 11496 2309
rect 11530 2275 11545 2309
rect 11685 2275 11700 2309
rect 11734 2275 11836 2309
rect 11394 2241 11545 2275
rect 11685 2241 11836 2275
rect 11394 2207 11496 2241
rect 11530 2207 11545 2241
rect 11685 2207 11700 2241
rect 11734 2207 11836 2241
rect 11394 2173 11545 2207
rect 11685 2173 11836 2207
rect 11394 2139 11496 2173
rect 11530 2139 11545 2173
rect 11685 2139 11700 2173
rect 11734 2139 11836 2173
rect 11394 2105 11545 2139
rect 11685 2105 11836 2139
rect 11394 2071 11496 2105
rect 11530 2071 11545 2105
rect 11685 2071 11700 2105
rect 11734 2071 11836 2105
rect 11394 2037 11545 2071
rect 11685 2037 11836 2071
rect 11394 2003 11496 2037
rect 11530 2003 11545 2037
rect 11685 2003 11700 2037
rect 11734 2003 11836 2037
rect 11394 1969 11545 2003
rect 11685 1969 11836 2003
rect 11394 1935 11496 1969
rect 11530 1935 11545 1969
rect 11685 1935 11700 1969
rect 11734 1935 11836 1969
rect 11394 1901 11545 1935
rect 11685 1901 11836 1935
rect 11394 1867 11496 1901
rect 11530 1867 11545 1901
rect 11685 1867 11700 1901
rect 11734 1867 11836 1901
rect 11394 1833 11545 1867
rect 11685 1833 11836 1867
rect 11394 1799 11496 1833
rect 11530 1799 11545 1833
rect 11685 1799 11700 1833
rect 11734 1799 11836 1833
rect 11394 1765 11545 1799
rect 11685 1765 11836 1799
rect 11394 1731 11496 1765
rect 11530 1731 11545 1765
rect 11685 1731 11700 1765
rect 11734 1731 11836 1765
rect 11394 1697 11545 1731
rect 11685 1697 11836 1731
rect 11394 1663 11496 1697
rect 11530 1663 11545 1697
rect 11685 1663 11700 1697
rect 11734 1663 11836 1697
rect 11394 1629 11545 1663
rect 11685 1629 11836 1663
rect 11394 1595 11496 1629
rect 11530 1595 11545 1629
rect 11685 1595 11700 1629
rect 11734 1595 11836 1629
rect 11394 1561 11545 1595
rect 11685 1561 11836 1595
rect 11394 1527 11496 1561
rect 11530 1527 11545 1561
rect 11685 1527 11700 1561
rect 11734 1527 11836 1561
rect 11394 1457 11545 1527
rect 11685 1457 11836 1527
rect 11956 2445 12266 2457
rect 11956 2411 12058 2445
rect 12092 2411 12130 2445
rect 12164 2411 12266 2445
rect 11956 2377 12266 2411
rect 11956 2343 12058 2377
rect 12092 2343 12130 2377
rect 12164 2343 12266 2377
rect 11956 2309 12266 2343
rect 11956 2275 12058 2309
rect 12092 2275 12130 2309
rect 12164 2275 12266 2309
rect 11956 2241 12266 2275
rect 11956 2207 12058 2241
rect 12092 2207 12130 2241
rect 12164 2207 12266 2241
rect 11956 2173 12266 2207
rect 11956 2139 12058 2173
rect 12092 2139 12130 2173
rect 12164 2139 12266 2173
rect 11956 2105 12266 2139
rect 11956 2071 12058 2105
rect 12092 2071 12130 2105
rect 12164 2071 12266 2105
rect 11956 2037 12266 2071
rect 11956 2003 12058 2037
rect 12092 2003 12130 2037
rect 12164 2003 12266 2037
rect 11956 1969 12266 2003
rect 11956 1935 12058 1969
rect 12092 1935 12130 1969
rect 12164 1935 12266 1969
rect 11956 1901 12266 1935
rect 11956 1867 12058 1901
rect 12092 1867 12130 1901
rect 12164 1867 12266 1901
rect 11956 1833 12266 1867
rect 11956 1799 12058 1833
rect 12092 1799 12130 1833
rect 12164 1799 12266 1833
rect 11956 1765 12266 1799
rect 11956 1731 12058 1765
rect 12092 1731 12130 1765
rect 12164 1731 12266 1765
rect 11956 1697 12266 1731
rect 11956 1663 12058 1697
rect 12092 1663 12130 1697
rect 12164 1663 12266 1697
rect 11956 1629 12266 1663
rect 11956 1595 12058 1629
rect 12092 1595 12130 1629
rect 12164 1595 12266 1629
rect 11956 1561 12266 1595
rect 11956 1527 12058 1561
rect 12092 1527 12130 1561
rect 12164 1527 12266 1561
rect 11956 1457 12266 1527
rect 12386 2445 12537 2457
rect 12677 2445 12828 2457
rect 12386 2411 12488 2445
rect 12522 2411 12537 2445
rect 12677 2411 12692 2445
rect 12726 2411 12828 2445
rect 12386 2377 12537 2411
rect 12677 2377 12828 2411
rect 12386 2343 12488 2377
rect 12522 2343 12537 2377
rect 12677 2343 12692 2377
rect 12726 2343 12828 2377
rect 12386 2309 12537 2343
rect 12677 2309 12828 2343
rect 12386 2275 12488 2309
rect 12522 2275 12537 2309
rect 12677 2275 12692 2309
rect 12726 2275 12828 2309
rect 12386 2241 12537 2275
rect 12677 2241 12828 2275
rect 12386 2207 12488 2241
rect 12522 2207 12537 2241
rect 12677 2207 12692 2241
rect 12726 2207 12828 2241
rect 12386 2173 12537 2207
rect 12677 2173 12828 2207
rect 12386 2139 12488 2173
rect 12522 2139 12537 2173
rect 12677 2139 12692 2173
rect 12726 2139 12828 2173
rect 12386 2105 12537 2139
rect 12677 2105 12828 2139
rect 12386 2071 12488 2105
rect 12522 2071 12537 2105
rect 12677 2071 12692 2105
rect 12726 2071 12828 2105
rect 12386 2037 12537 2071
rect 12677 2037 12828 2071
rect 12386 2003 12488 2037
rect 12522 2003 12537 2037
rect 12677 2003 12692 2037
rect 12726 2003 12828 2037
rect 12386 1969 12537 2003
rect 12677 1969 12828 2003
rect 12386 1935 12488 1969
rect 12522 1935 12537 1969
rect 12677 1935 12692 1969
rect 12726 1935 12828 1969
rect 12386 1901 12537 1935
rect 12677 1901 12828 1935
rect 12386 1867 12488 1901
rect 12522 1867 12537 1901
rect 12677 1867 12692 1901
rect 12726 1867 12828 1901
rect 12386 1833 12537 1867
rect 12677 1833 12828 1867
rect 12386 1799 12488 1833
rect 12522 1799 12537 1833
rect 12677 1799 12692 1833
rect 12726 1799 12828 1833
rect 12386 1765 12537 1799
rect 12677 1765 12828 1799
rect 12386 1731 12488 1765
rect 12522 1731 12537 1765
rect 12677 1731 12692 1765
rect 12726 1731 12828 1765
rect 12386 1697 12537 1731
rect 12677 1697 12828 1731
rect 12386 1663 12488 1697
rect 12522 1663 12537 1697
rect 12677 1663 12692 1697
rect 12726 1663 12828 1697
rect 12386 1629 12537 1663
rect 12677 1629 12828 1663
rect 12386 1595 12488 1629
rect 12522 1595 12537 1629
rect 12677 1595 12692 1629
rect 12726 1595 12828 1629
rect 12386 1561 12537 1595
rect 12677 1561 12828 1595
rect 12386 1527 12488 1561
rect 12522 1527 12537 1561
rect 12677 1527 12692 1561
rect 12726 1527 12828 1561
rect 12386 1457 12537 1527
rect 12677 1457 12828 1527
rect 12948 2445 13258 2457
rect 12948 2411 13050 2445
rect 13084 2411 13122 2445
rect 13156 2411 13258 2445
rect 12948 2377 13258 2411
rect 12948 2343 13050 2377
rect 13084 2343 13122 2377
rect 13156 2343 13258 2377
rect 12948 2309 13258 2343
rect 12948 2275 13050 2309
rect 13084 2275 13122 2309
rect 13156 2275 13258 2309
rect 12948 2241 13258 2275
rect 12948 2207 13050 2241
rect 13084 2207 13122 2241
rect 13156 2207 13258 2241
rect 12948 2173 13258 2207
rect 12948 2139 13050 2173
rect 13084 2139 13122 2173
rect 13156 2139 13258 2173
rect 12948 2105 13258 2139
rect 12948 2071 13050 2105
rect 13084 2071 13122 2105
rect 13156 2071 13258 2105
rect 12948 2037 13258 2071
rect 12948 2003 13050 2037
rect 13084 2003 13122 2037
rect 13156 2003 13258 2037
rect 12948 1969 13258 2003
rect 12948 1935 13050 1969
rect 13084 1935 13122 1969
rect 13156 1935 13258 1969
rect 12948 1901 13258 1935
rect 12948 1867 13050 1901
rect 13084 1867 13122 1901
rect 13156 1867 13258 1901
rect 12948 1833 13258 1867
rect 12948 1799 13050 1833
rect 13084 1799 13122 1833
rect 13156 1799 13258 1833
rect 12948 1765 13258 1799
rect 12948 1731 13050 1765
rect 13084 1731 13122 1765
rect 13156 1731 13258 1765
rect 12948 1697 13258 1731
rect 12948 1663 13050 1697
rect 13084 1663 13122 1697
rect 13156 1663 13258 1697
rect 12948 1629 13258 1663
rect 12948 1595 13050 1629
rect 13084 1595 13122 1629
rect 13156 1595 13258 1629
rect 12948 1561 13258 1595
rect 12948 1527 13050 1561
rect 13084 1527 13122 1561
rect 13156 1527 13258 1561
rect 12948 1457 13258 1527
rect 13378 2445 13529 2457
rect 13669 2445 13820 2457
rect 13378 2411 13480 2445
rect 13514 2411 13529 2445
rect 13669 2411 13684 2445
rect 13718 2411 13820 2445
rect 13378 2377 13529 2411
rect 13669 2377 13820 2411
rect 13378 2343 13480 2377
rect 13514 2343 13529 2377
rect 13669 2343 13684 2377
rect 13718 2343 13820 2377
rect 13378 2309 13529 2343
rect 13669 2309 13820 2343
rect 13378 2275 13480 2309
rect 13514 2275 13529 2309
rect 13669 2275 13684 2309
rect 13718 2275 13820 2309
rect 13378 2241 13529 2275
rect 13669 2241 13820 2275
rect 13378 2207 13480 2241
rect 13514 2207 13529 2241
rect 13669 2207 13684 2241
rect 13718 2207 13820 2241
rect 13378 2173 13529 2207
rect 13669 2173 13820 2207
rect 13378 2139 13480 2173
rect 13514 2139 13529 2173
rect 13669 2139 13684 2173
rect 13718 2139 13820 2173
rect 13378 2105 13529 2139
rect 13669 2105 13820 2139
rect 13378 2071 13480 2105
rect 13514 2071 13529 2105
rect 13669 2071 13684 2105
rect 13718 2071 13820 2105
rect 13378 2037 13529 2071
rect 13669 2037 13820 2071
rect 13378 2003 13480 2037
rect 13514 2003 13529 2037
rect 13669 2003 13684 2037
rect 13718 2003 13820 2037
rect 13378 1969 13529 2003
rect 13669 1969 13820 2003
rect 13378 1935 13480 1969
rect 13514 1935 13529 1969
rect 13669 1935 13684 1969
rect 13718 1935 13820 1969
rect 13378 1901 13529 1935
rect 13669 1901 13820 1935
rect 13378 1867 13480 1901
rect 13514 1867 13529 1901
rect 13669 1867 13684 1901
rect 13718 1867 13820 1901
rect 13378 1833 13529 1867
rect 13669 1833 13820 1867
rect 13378 1799 13480 1833
rect 13514 1799 13529 1833
rect 13669 1799 13684 1833
rect 13718 1799 13820 1833
rect 13378 1765 13529 1799
rect 13669 1765 13820 1799
rect 13378 1731 13480 1765
rect 13514 1731 13529 1765
rect 13669 1731 13684 1765
rect 13718 1731 13820 1765
rect 13378 1697 13529 1731
rect 13669 1697 13820 1731
rect 13378 1663 13480 1697
rect 13514 1663 13529 1697
rect 13669 1663 13684 1697
rect 13718 1663 13820 1697
rect 13378 1629 13529 1663
rect 13669 1629 13820 1663
rect 13378 1595 13480 1629
rect 13514 1595 13529 1629
rect 13669 1595 13684 1629
rect 13718 1595 13820 1629
rect 13378 1561 13529 1595
rect 13669 1561 13820 1595
rect 13378 1527 13480 1561
rect 13514 1527 13529 1561
rect 13669 1527 13684 1561
rect 13718 1527 13820 1561
rect 13378 1457 13529 1527
rect 13669 1457 13820 1527
rect 13940 2445 14178 2457
rect 13940 2411 14042 2445
rect 14076 2411 14178 2445
rect 13940 2377 14178 2411
rect 13940 2343 14042 2377
rect 14076 2343 14178 2377
rect 13940 2309 14178 2343
rect 13940 2275 14042 2309
rect 14076 2275 14178 2309
rect 13940 2241 14178 2275
rect 13940 2207 14042 2241
rect 14076 2207 14178 2241
rect 13940 2173 14178 2207
rect 13940 2139 14042 2173
rect 14076 2139 14178 2173
rect 13940 2105 14178 2139
rect 13940 2071 14042 2105
rect 14076 2071 14178 2105
rect 13940 2037 14178 2071
rect 13940 2003 14042 2037
rect 14076 2003 14178 2037
rect 13940 1969 14178 2003
rect 13940 1935 14042 1969
rect 14076 1935 14178 1969
rect 13940 1901 14178 1935
rect 13940 1867 14042 1901
rect 14076 1867 14178 1901
rect 13940 1833 14178 1867
rect 13940 1799 14042 1833
rect 14076 1799 14178 1833
rect 13940 1765 14178 1799
rect 13940 1731 14042 1765
rect 14076 1731 14178 1765
rect 13940 1697 14178 1731
rect 13940 1663 14042 1697
rect 14076 1663 14178 1697
rect 13940 1629 14178 1663
rect 13940 1595 14042 1629
rect 14076 1595 14178 1629
rect 13940 1561 14178 1595
rect 13940 1527 14042 1561
rect 14076 1527 14178 1561
rect 13940 1457 14178 1527
rect 14298 2445 14435 2457
rect 14298 2411 14386 2445
rect 14420 2411 14435 2445
rect 14298 2377 14435 2411
rect 14298 2343 14386 2377
rect 14420 2343 14435 2377
rect 14298 2309 14435 2343
rect 14298 2275 14386 2309
rect 14420 2275 14435 2309
rect 14298 2241 14435 2275
rect 14298 2207 14386 2241
rect 14420 2207 14435 2241
rect 14298 2173 14435 2207
rect 14298 2139 14386 2173
rect 14420 2139 14435 2173
rect 14298 2105 14435 2139
rect 14298 2071 14386 2105
rect 14420 2071 14435 2105
rect 14298 2037 14435 2071
rect 14298 2003 14386 2037
rect 14420 2003 14435 2037
rect 14298 1969 14435 2003
rect 14298 1935 14386 1969
rect 14420 1935 14435 1969
rect 14298 1901 14435 1935
rect 14298 1867 14386 1901
rect 14420 1867 14435 1901
rect 14298 1833 14435 1867
rect 14298 1799 14386 1833
rect 14420 1799 14435 1833
rect 14298 1765 14435 1799
rect 14298 1731 14386 1765
rect 14420 1731 14435 1765
rect 14298 1697 14435 1731
rect 14298 1663 14386 1697
rect 14420 1663 14435 1697
rect 14298 1629 14435 1663
rect 14298 1595 14386 1629
rect 14420 1595 14435 1629
rect 14298 1561 14435 1595
rect 14298 1527 14386 1561
rect 14420 1527 14435 1561
rect 14298 1457 14435 1527
<< mvndiffc >>
rect 802 4012 836 4046
rect 802 3944 836 3978
rect 802 3876 836 3910
rect 802 3808 836 3842
rect 802 3740 836 3774
rect 802 3672 836 3706
rect 802 3604 836 3638
rect 802 3536 836 3570
rect 802 3468 836 3502
rect 802 3400 836 3434
rect 802 3332 836 3366
rect 802 3264 836 3298
rect 802 3196 836 3230
rect 802 3128 836 3162
rect 1146 4012 1180 4046
rect 1218 4012 1252 4046
rect 1146 3944 1180 3978
rect 1218 3944 1252 3978
rect 1146 3876 1180 3910
rect 1218 3876 1252 3910
rect 1146 3808 1180 3842
rect 1218 3808 1252 3842
rect 1146 3740 1180 3774
rect 1218 3740 1252 3774
rect 1146 3672 1180 3706
rect 1218 3672 1252 3706
rect 1146 3604 1180 3638
rect 1218 3604 1252 3638
rect 1146 3536 1180 3570
rect 1218 3536 1252 3570
rect 1146 3468 1180 3502
rect 1218 3468 1252 3502
rect 1146 3400 1180 3434
rect 1218 3400 1252 3434
rect 1146 3332 1180 3366
rect 1218 3332 1252 3366
rect 1146 3264 1180 3298
rect 1218 3264 1252 3298
rect 1146 3196 1180 3230
rect 1218 3196 1252 3230
rect 1146 3128 1180 3162
rect 1218 3128 1252 3162
rect 1576 4012 1610 4046
rect 1780 4012 1814 4046
rect 1576 3944 1610 3978
rect 1780 3944 1814 3978
rect 1576 3876 1610 3910
rect 1780 3876 1814 3910
rect 1576 3808 1610 3842
rect 1780 3808 1814 3842
rect 1576 3740 1610 3774
rect 1780 3740 1814 3774
rect 1576 3672 1610 3706
rect 1780 3672 1814 3706
rect 1576 3604 1610 3638
rect 1780 3604 1814 3638
rect 1576 3536 1610 3570
rect 1780 3536 1814 3570
rect 1576 3468 1610 3502
rect 1780 3468 1814 3502
rect 1576 3400 1610 3434
rect 1780 3400 1814 3434
rect 1576 3332 1610 3366
rect 1780 3332 1814 3366
rect 1576 3264 1610 3298
rect 1780 3264 1814 3298
rect 1576 3196 1610 3230
rect 1780 3196 1814 3230
rect 1576 3128 1610 3162
rect 1780 3128 1814 3162
rect 2138 4012 2172 4046
rect 2210 4012 2244 4046
rect 2138 3944 2172 3978
rect 2210 3944 2244 3978
rect 2138 3876 2172 3910
rect 2210 3876 2244 3910
rect 2138 3808 2172 3842
rect 2210 3808 2244 3842
rect 2138 3740 2172 3774
rect 2210 3740 2244 3774
rect 2138 3672 2172 3706
rect 2210 3672 2244 3706
rect 2138 3604 2172 3638
rect 2210 3604 2244 3638
rect 2138 3536 2172 3570
rect 2210 3536 2244 3570
rect 2138 3468 2172 3502
rect 2210 3468 2244 3502
rect 2138 3400 2172 3434
rect 2210 3400 2244 3434
rect 2138 3332 2172 3366
rect 2210 3332 2244 3366
rect 2138 3264 2172 3298
rect 2210 3264 2244 3298
rect 2138 3196 2172 3230
rect 2210 3196 2244 3230
rect 2138 3128 2172 3162
rect 2210 3128 2244 3162
rect 2568 4012 2602 4046
rect 2772 4012 2806 4046
rect 2568 3944 2602 3978
rect 2772 3944 2806 3978
rect 2568 3876 2602 3910
rect 2772 3876 2806 3910
rect 2568 3808 2602 3842
rect 2772 3808 2806 3842
rect 2568 3740 2602 3774
rect 2772 3740 2806 3774
rect 2568 3672 2602 3706
rect 2772 3672 2806 3706
rect 2568 3604 2602 3638
rect 2772 3604 2806 3638
rect 2568 3536 2602 3570
rect 2772 3536 2806 3570
rect 2568 3468 2602 3502
rect 2772 3468 2806 3502
rect 2568 3400 2602 3434
rect 2772 3400 2806 3434
rect 2568 3332 2602 3366
rect 2772 3332 2806 3366
rect 2568 3264 2602 3298
rect 2772 3264 2806 3298
rect 2568 3196 2602 3230
rect 2772 3196 2806 3230
rect 2568 3128 2602 3162
rect 2772 3128 2806 3162
rect 3130 4012 3164 4046
rect 3202 4012 3236 4046
rect 3130 3944 3164 3978
rect 3202 3944 3236 3978
rect 3130 3876 3164 3910
rect 3202 3876 3236 3910
rect 3130 3808 3164 3842
rect 3202 3808 3236 3842
rect 3130 3740 3164 3774
rect 3202 3740 3236 3774
rect 3130 3672 3164 3706
rect 3202 3672 3236 3706
rect 3130 3604 3164 3638
rect 3202 3604 3236 3638
rect 3130 3536 3164 3570
rect 3202 3536 3236 3570
rect 3130 3468 3164 3502
rect 3202 3468 3236 3502
rect 3130 3400 3164 3434
rect 3202 3400 3236 3434
rect 3130 3332 3164 3366
rect 3202 3332 3236 3366
rect 3130 3264 3164 3298
rect 3202 3264 3236 3298
rect 3130 3196 3164 3230
rect 3202 3196 3236 3230
rect 3130 3128 3164 3162
rect 3202 3128 3236 3162
rect 3560 4012 3594 4046
rect 3764 4012 3798 4046
rect 3560 3944 3594 3978
rect 3764 3944 3798 3978
rect 3560 3876 3594 3910
rect 3764 3876 3798 3910
rect 3560 3808 3594 3842
rect 3764 3808 3798 3842
rect 3560 3740 3594 3774
rect 3764 3740 3798 3774
rect 3560 3672 3594 3706
rect 3764 3672 3798 3706
rect 3560 3604 3594 3638
rect 3764 3604 3798 3638
rect 3560 3536 3594 3570
rect 3764 3536 3798 3570
rect 3560 3468 3594 3502
rect 3764 3468 3798 3502
rect 3560 3400 3594 3434
rect 3764 3400 3798 3434
rect 3560 3332 3594 3366
rect 3764 3332 3798 3366
rect 3560 3264 3594 3298
rect 3764 3264 3798 3298
rect 3560 3196 3594 3230
rect 3764 3196 3798 3230
rect 3560 3128 3594 3162
rect 3764 3128 3798 3162
rect 4122 4012 4156 4046
rect 4194 4012 4228 4046
rect 4122 3944 4156 3978
rect 4194 3944 4228 3978
rect 4122 3876 4156 3910
rect 4194 3876 4228 3910
rect 4122 3808 4156 3842
rect 4194 3808 4228 3842
rect 4122 3740 4156 3774
rect 4194 3740 4228 3774
rect 4122 3672 4156 3706
rect 4194 3672 4228 3706
rect 4122 3604 4156 3638
rect 4194 3604 4228 3638
rect 4122 3536 4156 3570
rect 4194 3536 4228 3570
rect 4122 3468 4156 3502
rect 4194 3468 4228 3502
rect 4122 3400 4156 3434
rect 4194 3400 4228 3434
rect 4122 3332 4156 3366
rect 4194 3332 4228 3366
rect 4122 3264 4156 3298
rect 4194 3264 4228 3298
rect 4122 3196 4156 3230
rect 4194 3196 4228 3230
rect 4122 3128 4156 3162
rect 4194 3128 4228 3162
rect 4552 4012 4586 4046
rect 4756 4012 4790 4046
rect 4552 3944 4586 3978
rect 4756 3944 4790 3978
rect 4552 3876 4586 3910
rect 4756 3876 4790 3910
rect 4552 3808 4586 3842
rect 4756 3808 4790 3842
rect 4552 3740 4586 3774
rect 4756 3740 4790 3774
rect 4552 3672 4586 3706
rect 4756 3672 4790 3706
rect 4552 3604 4586 3638
rect 4756 3604 4790 3638
rect 4552 3536 4586 3570
rect 4756 3536 4790 3570
rect 4552 3468 4586 3502
rect 4756 3468 4790 3502
rect 4552 3400 4586 3434
rect 4756 3400 4790 3434
rect 4552 3332 4586 3366
rect 4756 3332 4790 3366
rect 4552 3264 4586 3298
rect 4756 3264 4790 3298
rect 4552 3196 4586 3230
rect 4756 3196 4790 3230
rect 4552 3128 4586 3162
rect 4756 3128 4790 3162
rect 5114 4012 5148 4046
rect 5186 4012 5220 4046
rect 5114 3944 5148 3978
rect 5186 3944 5220 3978
rect 5114 3876 5148 3910
rect 5186 3876 5220 3910
rect 5114 3808 5148 3842
rect 5186 3808 5220 3842
rect 5114 3740 5148 3774
rect 5186 3740 5220 3774
rect 5114 3672 5148 3706
rect 5186 3672 5220 3706
rect 5114 3604 5148 3638
rect 5186 3604 5220 3638
rect 5114 3536 5148 3570
rect 5186 3536 5220 3570
rect 5114 3468 5148 3502
rect 5186 3468 5220 3502
rect 5114 3400 5148 3434
rect 5186 3400 5220 3434
rect 5114 3332 5148 3366
rect 5186 3332 5220 3366
rect 5114 3264 5148 3298
rect 5186 3264 5220 3298
rect 5114 3196 5148 3230
rect 5186 3196 5220 3230
rect 5114 3128 5148 3162
rect 5186 3128 5220 3162
rect 5544 4012 5578 4046
rect 5748 4012 5782 4046
rect 5544 3944 5578 3978
rect 5748 3944 5782 3978
rect 5544 3876 5578 3910
rect 5748 3876 5782 3910
rect 5544 3808 5578 3842
rect 5748 3808 5782 3842
rect 5544 3740 5578 3774
rect 5748 3740 5782 3774
rect 5544 3672 5578 3706
rect 5748 3672 5782 3706
rect 5544 3604 5578 3638
rect 5748 3604 5782 3638
rect 5544 3536 5578 3570
rect 5748 3536 5782 3570
rect 5544 3468 5578 3502
rect 5748 3468 5782 3502
rect 5544 3400 5578 3434
rect 5748 3400 5782 3434
rect 5544 3332 5578 3366
rect 5748 3332 5782 3366
rect 5544 3264 5578 3298
rect 5748 3264 5782 3298
rect 5544 3196 5578 3230
rect 5748 3196 5782 3230
rect 5544 3128 5578 3162
rect 5748 3128 5782 3162
rect 6106 4012 6140 4046
rect 6178 4012 6212 4046
rect 6106 3944 6140 3978
rect 6178 3944 6212 3978
rect 6106 3876 6140 3910
rect 6178 3876 6212 3910
rect 6106 3808 6140 3842
rect 6178 3808 6212 3842
rect 6106 3740 6140 3774
rect 6178 3740 6212 3774
rect 6106 3672 6140 3706
rect 6178 3672 6212 3706
rect 6106 3604 6140 3638
rect 6178 3604 6212 3638
rect 6106 3536 6140 3570
rect 6178 3536 6212 3570
rect 6106 3468 6140 3502
rect 6178 3468 6212 3502
rect 6106 3400 6140 3434
rect 6178 3400 6212 3434
rect 6106 3332 6140 3366
rect 6178 3332 6212 3366
rect 6106 3264 6140 3298
rect 6178 3264 6212 3298
rect 6106 3196 6140 3230
rect 6178 3196 6212 3230
rect 6106 3128 6140 3162
rect 6178 3128 6212 3162
rect 6536 4012 6570 4046
rect 6740 4012 6774 4046
rect 6536 3944 6570 3978
rect 6740 3944 6774 3978
rect 6536 3876 6570 3910
rect 6740 3876 6774 3910
rect 6536 3808 6570 3842
rect 6740 3808 6774 3842
rect 6536 3740 6570 3774
rect 6740 3740 6774 3774
rect 6536 3672 6570 3706
rect 6740 3672 6774 3706
rect 6536 3604 6570 3638
rect 6740 3604 6774 3638
rect 6536 3536 6570 3570
rect 6740 3536 6774 3570
rect 6536 3468 6570 3502
rect 6740 3468 6774 3502
rect 6536 3400 6570 3434
rect 6740 3400 6774 3434
rect 6536 3332 6570 3366
rect 6740 3332 6774 3366
rect 6536 3264 6570 3298
rect 6740 3264 6774 3298
rect 6536 3196 6570 3230
rect 6740 3196 6774 3230
rect 6536 3128 6570 3162
rect 6740 3128 6774 3162
rect 7098 4012 7132 4046
rect 7170 4012 7204 4046
rect 7098 3944 7132 3978
rect 7170 3944 7204 3978
rect 7098 3876 7132 3910
rect 7170 3876 7204 3910
rect 7098 3808 7132 3842
rect 7170 3808 7204 3842
rect 7098 3740 7132 3774
rect 7170 3740 7204 3774
rect 7098 3672 7132 3706
rect 7170 3672 7204 3706
rect 7098 3604 7132 3638
rect 7170 3604 7204 3638
rect 7098 3536 7132 3570
rect 7170 3536 7204 3570
rect 7098 3468 7132 3502
rect 7170 3468 7204 3502
rect 7098 3400 7132 3434
rect 7170 3400 7204 3434
rect 7098 3332 7132 3366
rect 7170 3332 7204 3366
rect 7098 3264 7132 3298
rect 7170 3264 7204 3298
rect 7098 3196 7132 3230
rect 7170 3196 7204 3230
rect 7098 3128 7132 3162
rect 7170 3128 7204 3162
rect 7528 4012 7562 4046
rect 7732 4012 7766 4046
rect 7528 3944 7562 3978
rect 7732 3944 7766 3978
rect 7528 3876 7562 3910
rect 7732 3876 7766 3910
rect 7528 3808 7562 3842
rect 7732 3808 7766 3842
rect 7528 3740 7562 3774
rect 7732 3740 7766 3774
rect 7528 3672 7562 3706
rect 7732 3672 7766 3706
rect 7528 3604 7562 3638
rect 7732 3604 7766 3638
rect 7528 3536 7562 3570
rect 7732 3536 7766 3570
rect 7528 3468 7562 3502
rect 7732 3468 7766 3502
rect 7528 3400 7562 3434
rect 7732 3400 7766 3434
rect 7528 3332 7562 3366
rect 7732 3332 7766 3366
rect 7528 3264 7562 3298
rect 7732 3264 7766 3298
rect 7528 3196 7562 3230
rect 7732 3196 7766 3230
rect 7528 3128 7562 3162
rect 7732 3128 7766 3162
rect 8090 4012 8124 4046
rect 8162 4012 8196 4046
rect 8090 3944 8124 3978
rect 8162 3944 8196 3978
rect 8090 3876 8124 3910
rect 8162 3876 8196 3910
rect 8090 3808 8124 3842
rect 8162 3808 8196 3842
rect 8090 3740 8124 3774
rect 8162 3740 8196 3774
rect 8090 3672 8124 3706
rect 8162 3672 8196 3706
rect 8090 3604 8124 3638
rect 8162 3604 8196 3638
rect 8090 3536 8124 3570
rect 8162 3536 8196 3570
rect 8090 3468 8124 3502
rect 8162 3468 8196 3502
rect 8090 3400 8124 3434
rect 8162 3400 8196 3434
rect 8090 3332 8124 3366
rect 8162 3332 8196 3366
rect 8090 3264 8124 3298
rect 8162 3264 8196 3298
rect 8090 3196 8124 3230
rect 8162 3196 8196 3230
rect 8090 3128 8124 3162
rect 8162 3128 8196 3162
rect 8520 4012 8554 4046
rect 8724 4012 8758 4046
rect 8520 3944 8554 3978
rect 8724 3944 8758 3978
rect 8520 3876 8554 3910
rect 8724 3876 8758 3910
rect 8520 3808 8554 3842
rect 8724 3808 8758 3842
rect 8520 3740 8554 3774
rect 8724 3740 8758 3774
rect 8520 3672 8554 3706
rect 8724 3672 8758 3706
rect 8520 3604 8554 3638
rect 8724 3604 8758 3638
rect 8520 3536 8554 3570
rect 8724 3536 8758 3570
rect 8520 3468 8554 3502
rect 8724 3468 8758 3502
rect 8520 3400 8554 3434
rect 8724 3400 8758 3434
rect 8520 3332 8554 3366
rect 8724 3332 8758 3366
rect 8520 3264 8554 3298
rect 8724 3264 8758 3298
rect 8520 3196 8554 3230
rect 8724 3196 8758 3230
rect 8520 3128 8554 3162
rect 8724 3128 8758 3162
rect 9082 4012 9116 4046
rect 9154 4012 9188 4046
rect 9082 3944 9116 3978
rect 9154 3944 9188 3978
rect 9082 3876 9116 3910
rect 9154 3876 9188 3910
rect 9082 3808 9116 3842
rect 9154 3808 9188 3842
rect 9082 3740 9116 3774
rect 9154 3740 9188 3774
rect 9082 3672 9116 3706
rect 9154 3672 9188 3706
rect 9082 3604 9116 3638
rect 9154 3604 9188 3638
rect 9082 3536 9116 3570
rect 9154 3536 9188 3570
rect 9082 3468 9116 3502
rect 9154 3468 9188 3502
rect 9082 3400 9116 3434
rect 9154 3400 9188 3434
rect 9082 3332 9116 3366
rect 9154 3332 9188 3366
rect 9082 3264 9116 3298
rect 9154 3264 9188 3298
rect 9082 3196 9116 3230
rect 9154 3196 9188 3230
rect 9082 3128 9116 3162
rect 9154 3128 9188 3162
rect 9512 4012 9546 4046
rect 9716 4012 9750 4046
rect 9512 3944 9546 3978
rect 9716 3944 9750 3978
rect 9512 3876 9546 3910
rect 9716 3876 9750 3910
rect 9512 3808 9546 3842
rect 9716 3808 9750 3842
rect 9512 3740 9546 3774
rect 9716 3740 9750 3774
rect 9512 3672 9546 3706
rect 9716 3672 9750 3706
rect 9512 3604 9546 3638
rect 9716 3604 9750 3638
rect 9512 3536 9546 3570
rect 9716 3536 9750 3570
rect 9512 3468 9546 3502
rect 9716 3468 9750 3502
rect 9512 3400 9546 3434
rect 9716 3400 9750 3434
rect 9512 3332 9546 3366
rect 9716 3332 9750 3366
rect 9512 3264 9546 3298
rect 9716 3264 9750 3298
rect 9512 3196 9546 3230
rect 9716 3196 9750 3230
rect 9512 3128 9546 3162
rect 9716 3128 9750 3162
rect 10074 4012 10108 4046
rect 10146 4012 10180 4046
rect 10074 3944 10108 3978
rect 10146 3944 10180 3978
rect 10074 3876 10108 3910
rect 10146 3876 10180 3910
rect 10074 3808 10108 3842
rect 10146 3808 10180 3842
rect 10074 3740 10108 3774
rect 10146 3740 10180 3774
rect 10074 3672 10108 3706
rect 10146 3672 10180 3706
rect 10074 3604 10108 3638
rect 10146 3604 10180 3638
rect 10074 3536 10108 3570
rect 10146 3536 10180 3570
rect 10074 3468 10108 3502
rect 10146 3468 10180 3502
rect 10074 3400 10108 3434
rect 10146 3400 10180 3434
rect 10074 3332 10108 3366
rect 10146 3332 10180 3366
rect 10074 3264 10108 3298
rect 10146 3264 10180 3298
rect 10074 3196 10108 3230
rect 10146 3196 10180 3230
rect 10074 3128 10108 3162
rect 10146 3128 10180 3162
rect 10504 4012 10538 4046
rect 10708 4012 10742 4046
rect 10504 3944 10538 3978
rect 10708 3944 10742 3978
rect 10504 3876 10538 3910
rect 10708 3876 10742 3910
rect 10504 3808 10538 3842
rect 10708 3808 10742 3842
rect 10504 3740 10538 3774
rect 10708 3740 10742 3774
rect 10504 3672 10538 3706
rect 10708 3672 10742 3706
rect 10504 3604 10538 3638
rect 10708 3604 10742 3638
rect 10504 3536 10538 3570
rect 10708 3536 10742 3570
rect 10504 3468 10538 3502
rect 10708 3468 10742 3502
rect 10504 3400 10538 3434
rect 10708 3400 10742 3434
rect 10504 3332 10538 3366
rect 10708 3332 10742 3366
rect 10504 3264 10538 3298
rect 10708 3264 10742 3298
rect 10504 3196 10538 3230
rect 10708 3196 10742 3230
rect 10504 3128 10538 3162
rect 10708 3128 10742 3162
rect 11066 4012 11100 4046
rect 11138 4012 11172 4046
rect 11066 3944 11100 3978
rect 11138 3944 11172 3978
rect 11066 3876 11100 3910
rect 11138 3876 11172 3910
rect 11066 3808 11100 3842
rect 11138 3808 11172 3842
rect 11066 3740 11100 3774
rect 11138 3740 11172 3774
rect 11066 3672 11100 3706
rect 11138 3672 11172 3706
rect 11066 3604 11100 3638
rect 11138 3604 11172 3638
rect 11066 3536 11100 3570
rect 11138 3536 11172 3570
rect 11066 3468 11100 3502
rect 11138 3468 11172 3502
rect 11066 3400 11100 3434
rect 11138 3400 11172 3434
rect 11066 3332 11100 3366
rect 11138 3332 11172 3366
rect 11066 3264 11100 3298
rect 11138 3264 11172 3298
rect 11066 3196 11100 3230
rect 11138 3196 11172 3230
rect 11066 3128 11100 3162
rect 11138 3128 11172 3162
rect 11496 4012 11530 4046
rect 11700 4012 11734 4046
rect 11496 3944 11530 3978
rect 11700 3944 11734 3978
rect 11496 3876 11530 3910
rect 11700 3876 11734 3910
rect 11496 3808 11530 3842
rect 11700 3808 11734 3842
rect 11496 3740 11530 3774
rect 11700 3740 11734 3774
rect 11496 3672 11530 3706
rect 11700 3672 11734 3706
rect 11496 3604 11530 3638
rect 11700 3604 11734 3638
rect 11496 3536 11530 3570
rect 11700 3536 11734 3570
rect 11496 3468 11530 3502
rect 11700 3468 11734 3502
rect 11496 3400 11530 3434
rect 11700 3400 11734 3434
rect 11496 3332 11530 3366
rect 11700 3332 11734 3366
rect 11496 3264 11530 3298
rect 11700 3264 11734 3298
rect 11496 3196 11530 3230
rect 11700 3196 11734 3230
rect 11496 3128 11530 3162
rect 11700 3128 11734 3162
rect 12058 4012 12092 4046
rect 12130 4012 12164 4046
rect 12058 3944 12092 3978
rect 12130 3944 12164 3978
rect 12058 3876 12092 3910
rect 12130 3876 12164 3910
rect 12058 3808 12092 3842
rect 12130 3808 12164 3842
rect 12058 3740 12092 3774
rect 12130 3740 12164 3774
rect 12058 3672 12092 3706
rect 12130 3672 12164 3706
rect 12058 3604 12092 3638
rect 12130 3604 12164 3638
rect 12058 3536 12092 3570
rect 12130 3536 12164 3570
rect 12058 3468 12092 3502
rect 12130 3468 12164 3502
rect 12058 3400 12092 3434
rect 12130 3400 12164 3434
rect 12058 3332 12092 3366
rect 12130 3332 12164 3366
rect 12058 3264 12092 3298
rect 12130 3264 12164 3298
rect 12058 3196 12092 3230
rect 12130 3196 12164 3230
rect 12058 3128 12092 3162
rect 12130 3128 12164 3162
rect 12488 4012 12522 4046
rect 12692 4012 12726 4046
rect 12488 3944 12522 3978
rect 12692 3944 12726 3978
rect 12488 3876 12522 3910
rect 12692 3876 12726 3910
rect 12488 3808 12522 3842
rect 12692 3808 12726 3842
rect 12488 3740 12522 3774
rect 12692 3740 12726 3774
rect 12488 3672 12522 3706
rect 12692 3672 12726 3706
rect 12488 3604 12522 3638
rect 12692 3604 12726 3638
rect 12488 3536 12522 3570
rect 12692 3536 12726 3570
rect 12488 3468 12522 3502
rect 12692 3468 12726 3502
rect 12488 3400 12522 3434
rect 12692 3400 12726 3434
rect 12488 3332 12522 3366
rect 12692 3332 12726 3366
rect 12488 3264 12522 3298
rect 12692 3264 12726 3298
rect 12488 3196 12522 3230
rect 12692 3196 12726 3230
rect 12488 3128 12522 3162
rect 12692 3128 12726 3162
rect 13050 4012 13084 4046
rect 13122 4012 13156 4046
rect 13050 3944 13084 3978
rect 13122 3944 13156 3978
rect 13050 3876 13084 3910
rect 13122 3876 13156 3910
rect 13050 3808 13084 3842
rect 13122 3808 13156 3842
rect 13050 3740 13084 3774
rect 13122 3740 13156 3774
rect 13050 3672 13084 3706
rect 13122 3672 13156 3706
rect 13050 3604 13084 3638
rect 13122 3604 13156 3638
rect 13050 3536 13084 3570
rect 13122 3536 13156 3570
rect 13050 3468 13084 3502
rect 13122 3468 13156 3502
rect 13050 3400 13084 3434
rect 13122 3400 13156 3434
rect 13050 3332 13084 3366
rect 13122 3332 13156 3366
rect 13050 3264 13084 3298
rect 13122 3264 13156 3298
rect 13050 3196 13084 3230
rect 13122 3196 13156 3230
rect 13050 3128 13084 3162
rect 13122 3128 13156 3162
rect 13480 4012 13514 4046
rect 13684 4012 13718 4046
rect 13480 3944 13514 3978
rect 13684 3944 13718 3978
rect 13480 3876 13514 3910
rect 13684 3876 13718 3910
rect 13480 3808 13514 3842
rect 13684 3808 13718 3842
rect 13480 3740 13514 3774
rect 13684 3740 13718 3774
rect 13480 3672 13514 3706
rect 13684 3672 13718 3706
rect 13480 3604 13514 3638
rect 13684 3604 13718 3638
rect 13480 3536 13514 3570
rect 13684 3536 13718 3570
rect 13480 3468 13514 3502
rect 13684 3468 13718 3502
rect 13480 3400 13514 3434
rect 13684 3400 13718 3434
rect 13480 3332 13514 3366
rect 13684 3332 13718 3366
rect 13480 3264 13514 3298
rect 13684 3264 13718 3298
rect 13480 3196 13514 3230
rect 13684 3196 13718 3230
rect 13480 3128 13514 3162
rect 13684 3128 13718 3162
rect 14042 4012 14076 4046
rect 14042 3944 14076 3978
rect 14042 3876 14076 3910
rect 14042 3808 14076 3842
rect 14042 3740 14076 3774
rect 14042 3672 14076 3706
rect 14042 3604 14076 3638
rect 14042 3536 14076 3570
rect 14042 3468 14076 3502
rect 14042 3400 14076 3434
rect 14042 3332 14076 3366
rect 14042 3264 14076 3298
rect 14042 3196 14076 3230
rect 14042 3128 14076 3162
rect 14386 4012 14420 4046
rect 14386 3944 14420 3978
rect 14386 3876 14420 3910
rect 14386 3808 14420 3842
rect 14386 3740 14420 3774
rect 14386 3672 14420 3706
rect 14386 3604 14420 3638
rect 14386 3536 14420 3570
rect 14386 3468 14420 3502
rect 14386 3400 14420 3434
rect 14386 3332 14420 3366
rect 14386 3264 14420 3298
rect 14386 3196 14420 3230
rect 14386 3128 14420 3162
rect 802 2411 836 2445
rect 802 2343 836 2377
rect 802 2275 836 2309
rect 802 2207 836 2241
rect 802 2139 836 2173
rect 802 2071 836 2105
rect 802 2003 836 2037
rect 802 1935 836 1969
rect 802 1867 836 1901
rect 802 1799 836 1833
rect 802 1731 836 1765
rect 802 1663 836 1697
rect 802 1595 836 1629
rect 802 1527 836 1561
rect 1146 2411 1180 2445
rect 1218 2411 1252 2445
rect 1146 2343 1180 2377
rect 1218 2343 1252 2377
rect 1146 2275 1180 2309
rect 1218 2275 1252 2309
rect 1146 2207 1180 2241
rect 1218 2207 1252 2241
rect 1146 2139 1180 2173
rect 1218 2139 1252 2173
rect 1146 2071 1180 2105
rect 1218 2071 1252 2105
rect 1146 2003 1180 2037
rect 1218 2003 1252 2037
rect 1146 1935 1180 1969
rect 1218 1935 1252 1969
rect 1146 1867 1180 1901
rect 1218 1867 1252 1901
rect 1146 1799 1180 1833
rect 1218 1799 1252 1833
rect 1146 1731 1180 1765
rect 1218 1731 1252 1765
rect 1146 1663 1180 1697
rect 1218 1663 1252 1697
rect 1146 1595 1180 1629
rect 1218 1595 1252 1629
rect 1146 1527 1180 1561
rect 1218 1527 1252 1561
rect 1576 2411 1610 2445
rect 1780 2411 1814 2445
rect 1576 2343 1610 2377
rect 1780 2343 1814 2377
rect 1576 2275 1610 2309
rect 1780 2275 1814 2309
rect 1576 2207 1610 2241
rect 1780 2207 1814 2241
rect 1576 2139 1610 2173
rect 1780 2139 1814 2173
rect 1576 2071 1610 2105
rect 1780 2071 1814 2105
rect 1576 2003 1610 2037
rect 1780 2003 1814 2037
rect 1576 1935 1610 1969
rect 1780 1935 1814 1969
rect 1576 1867 1610 1901
rect 1780 1867 1814 1901
rect 1576 1799 1610 1833
rect 1780 1799 1814 1833
rect 1576 1731 1610 1765
rect 1780 1731 1814 1765
rect 1576 1663 1610 1697
rect 1780 1663 1814 1697
rect 1576 1595 1610 1629
rect 1780 1595 1814 1629
rect 1576 1527 1610 1561
rect 1780 1527 1814 1561
rect 2138 2411 2172 2445
rect 2210 2411 2244 2445
rect 2138 2343 2172 2377
rect 2210 2343 2244 2377
rect 2138 2275 2172 2309
rect 2210 2275 2244 2309
rect 2138 2207 2172 2241
rect 2210 2207 2244 2241
rect 2138 2139 2172 2173
rect 2210 2139 2244 2173
rect 2138 2071 2172 2105
rect 2210 2071 2244 2105
rect 2138 2003 2172 2037
rect 2210 2003 2244 2037
rect 2138 1935 2172 1969
rect 2210 1935 2244 1969
rect 2138 1867 2172 1901
rect 2210 1867 2244 1901
rect 2138 1799 2172 1833
rect 2210 1799 2244 1833
rect 2138 1731 2172 1765
rect 2210 1731 2244 1765
rect 2138 1663 2172 1697
rect 2210 1663 2244 1697
rect 2138 1595 2172 1629
rect 2210 1595 2244 1629
rect 2138 1527 2172 1561
rect 2210 1527 2244 1561
rect 2568 2411 2602 2445
rect 2772 2411 2806 2445
rect 2568 2343 2602 2377
rect 2772 2343 2806 2377
rect 2568 2275 2602 2309
rect 2772 2275 2806 2309
rect 2568 2207 2602 2241
rect 2772 2207 2806 2241
rect 2568 2139 2602 2173
rect 2772 2139 2806 2173
rect 2568 2071 2602 2105
rect 2772 2071 2806 2105
rect 2568 2003 2602 2037
rect 2772 2003 2806 2037
rect 2568 1935 2602 1969
rect 2772 1935 2806 1969
rect 2568 1867 2602 1901
rect 2772 1867 2806 1901
rect 2568 1799 2602 1833
rect 2772 1799 2806 1833
rect 2568 1731 2602 1765
rect 2772 1731 2806 1765
rect 2568 1663 2602 1697
rect 2772 1663 2806 1697
rect 2568 1595 2602 1629
rect 2772 1595 2806 1629
rect 2568 1527 2602 1561
rect 2772 1527 2806 1561
rect 3130 2411 3164 2445
rect 3202 2411 3236 2445
rect 3130 2343 3164 2377
rect 3202 2343 3236 2377
rect 3130 2275 3164 2309
rect 3202 2275 3236 2309
rect 3130 2207 3164 2241
rect 3202 2207 3236 2241
rect 3130 2139 3164 2173
rect 3202 2139 3236 2173
rect 3130 2071 3164 2105
rect 3202 2071 3236 2105
rect 3130 2003 3164 2037
rect 3202 2003 3236 2037
rect 3130 1935 3164 1969
rect 3202 1935 3236 1969
rect 3130 1867 3164 1901
rect 3202 1867 3236 1901
rect 3130 1799 3164 1833
rect 3202 1799 3236 1833
rect 3130 1731 3164 1765
rect 3202 1731 3236 1765
rect 3130 1663 3164 1697
rect 3202 1663 3236 1697
rect 3130 1595 3164 1629
rect 3202 1595 3236 1629
rect 3130 1527 3164 1561
rect 3202 1527 3236 1561
rect 3560 2411 3594 2445
rect 3764 2411 3798 2445
rect 3560 2343 3594 2377
rect 3764 2343 3798 2377
rect 3560 2275 3594 2309
rect 3764 2275 3798 2309
rect 3560 2207 3594 2241
rect 3764 2207 3798 2241
rect 3560 2139 3594 2173
rect 3764 2139 3798 2173
rect 3560 2071 3594 2105
rect 3764 2071 3798 2105
rect 3560 2003 3594 2037
rect 3764 2003 3798 2037
rect 3560 1935 3594 1969
rect 3764 1935 3798 1969
rect 3560 1867 3594 1901
rect 3764 1867 3798 1901
rect 3560 1799 3594 1833
rect 3764 1799 3798 1833
rect 3560 1731 3594 1765
rect 3764 1731 3798 1765
rect 3560 1663 3594 1697
rect 3764 1663 3798 1697
rect 3560 1595 3594 1629
rect 3764 1595 3798 1629
rect 3560 1527 3594 1561
rect 3764 1527 3798 1561
rect 4122 2411 4156 2445
rect 4194 2411 4228 2445
rect 4122 2343 4156 2377
rect 4194 2343 4228 2377
rect 4122 2275 4156 2309
rect 4194 2275 4228 2309
rect 4122 2207 4156 2241
rect 4194 2207 4228 2241
rect 4122 2139 4156 2173
rect 4194 2139 4228 2173
rect 4122 2071 4156 2105
rect 4194 2071 4228 2105
rect 4122 2003 4156 2037
rect 4194 2003 4228 2037
rect 4122 1935 4156 1969
rect 4194 1935 4228 1969
rect 4122 1867 4156 1901
rect 4194 1867 4228 1901
rect 4122 1799 4156 1833
rect 4194 1799 4228 1833
rect 4122 1731 4156 1765
rect 4194 1731 4228 1765
rect 4122 1663 4156 1697
rect 4194 1663 4228 1697
rect 4122 1595 4156 1629
rect 4194 1595 4228 1629
rect 4122 1527 4156 1561
rect 4194 1527 4228 1561
rect 4552 2411 4586 2445
rect 4756 2411 4790 2445
rect 4552 2343 4586 2377
rect 4756 2343 4790 2377
rect 4552 2275 4586 2309
rect 4756 2275 4790 2309
rect 4552 2207 4586 2241
rect 4756 2207 4790 2241
rect 4552 2139 4586 2173
rect 4756 2139 4790 2173
rect 4552 2071 4586 2105
rect 4756 2071 4790 2105
rect 4552 2003 4586 2037
rect 4756 2003 4790 2037
rect 4552 1935 4586 1969
rect 4756 1935 4790 1969
rect 4552 1867 4586 1901
rect 4756 1867 4790 1901
rect 4552 1799 4586 1833
rect 4756 1799 4790 1833
rect 4552 1731 4586 1765
rect 4756 1731 4790 1765
rect 4552 1663 4586 1697
rect 4756 1663 4790 1697
rect 4552 1595 4586 1629
rect 4756 1595 4790 1629
rect 4552 1527 4586 1561
rect 4756 1527 4790 1561
rect 5114 2411 5148 2445
rect 5186 2411 5220 2445
rect 5114 2343 5148 2377
rect 5186 2343 5220 2377
rect 5114 2275 5148 2309
rect 5186 2275 5220 2309
rect 5114 2207 5148 2241
rect 5186 2207 5220 2241
rect 5114 2139 5148 2173
rect 5186 2139 5220 2173
rect 5114 2071 5148 2105
rect 5186 2071 5220 2105
rect 5114 2003 5148 2037
rect 5186 2003 5220 2037
rect 5114 1935 5148 1969
rect 5186 1935 5220 1969
rect 5114 1867 5148 1901
rect 5186 1867 5220 1901
rect 5114 1799 5148 1833
rect 5186 1799 5220 1833
rect 5114 1731 5148 1765
rect 5186 1731 5220 1765
rect 5114 1663 5148 1697
rect 5186 1663 5220 1697
rect 5114 1595 5148 1629
rect 5186 1595 5220 1629
rect 5114 1527 5148 1561
rect 5186 1527 5220 1561
rect 5544 2411 5578 2445
rect 5748 2411 5782 2445
rect 5544 2343 5578 2377
rect 5748 2343 5782 2377
rect 5544 2275 5578 2309
rect 5748 2275 5782 2309
rect 5544 2207 5578 2241
rect 5748 2207 5782 2241
rect 5544 2139 5578 2173
rect 5748 2139 5782 2173
rect 5544 2071 5578 2105
rect 5748 2071 5782 2105
rect 5544 2003 5578 2037
rect 5748 2003 5782 2037
rect 5544 1935 5578 1969
rect 5748 1935 5782 1969
rect 5544 1867 5578 1901
rect 5748 1867 5782 1901
rect 5544 1799 5578 1833
rect 5748 1799 5782 1833
rect 5544 1731 5578 1765
rect 5748 1731 5782 1765
rect 5544 1663 5578 1697
rect 5748 1663 5782 1697
rect 5544 1595 5578 1629
rect 5748 1595 5782 1629
rect 5544 1527 5578 1561
rect 5748 1527 5782 1561
rect 6106 2411 6140 2445
rect 6178 2411 6212 2445
rect 6106 2343 6140 2377
rect 6178 2343 6212 2377
rect 6106 2275 6140 2309
rect 6178 2275 6212 2309
rect 6106 2207 6140 2241
rect 6178 2207 6212 2241
rect 6106 2139 6140 2173
rect 6178 2139 6212 2173
rect 6106 2071 6140 2105
rect 6178 2071 6212 2105
rect 6106 2003 6140 2037
rect 6178 2003 6212 2037
rect 6106 1935 6140 1969
rect 6178 1935 6212 1969
rect 6106 1867 6140 1901
rect 6178 1867 6212 1901
rect 6106 1799 6140 1833
rect 6178 1799 6212 1833
rect 6106 1731 6140 1765
rect 6178 1731 6212 1765
rect 6106 1663 6140 1697
rect 6178 1663 6212 1697
rect 6106 1595 6140 1629
rect 6178 1595 6212 1629
rect 6106 1527 6140 1561
rect 6178 1527 6212 1561
rect 6536 2411 6570 2445
rect 6740 2411 6774 2445
rect 6536 2343 6570 2377
rect 6740 2343 6774 2377
rect 6536 2275 6570 2309
rect 6740 2275 6774 2309
rect 6536 2207 6570 2241
rect 6740 2207 6774 2241
rect 6536 2139 6570 2173
rect 6740 2139 6774 2173
rect 6536 2071 6570 2105
rect 6740 2071 6774 2105
rect 6536 2003 6570 2037
rect 6740 2003 6774 2037
rect 6536 1935 6570 1969
rect 6740 1935 6774 1969
rect 6536 1867 6570 1901
rect 6740 1867 6774 1901
rect 6536 1799 6570 1833
rect 6740 1799 6774 1833
rect 6536 1731 6570 1765
rect 6740 1731 6774 1765
rect 6536 1663 6570 1697
rect 6740 1663 6774 1697
rect 6536 1595 6570 1629
rect 6740 1595 6774 1629
rect 6536 1527 6570 1561
rect 6740 1527 6774 1561
rect 7098 2411 7132 2445
rect 7170 2411 7204 2445
rect 7098 2343 7132 2377
rect 7170 2343 7204 2377
rect 7098 2275 7132 2309
rect 7170 2275 7204 2309
rect 7098 2207 7132 2241
rect 7170 2207 7204 2241
rect 7098 2139 7132 2173
rect 7170 2139 7204 2173
rect 7098 2071 7132 2105
rect 7170 2071 7204 2105
rect 7098 2003 7132 2037
rect 7170 2003 7204 2037
rect 7098 1935 7132 1969
rect 7170 1935 7204 1969
rect 7098 1867 7132 1901
rect 7170 1867 7204 1901
rect 7098 1799 7132 1833
rect 7170 1799 7204 1833
rect 7098 1731 7132 1765
rect 7170 1731 7204 1765
rect 7098 1663 7132 1697
rect 7170 1663 7204 1697
rect 7098 1595 7132 1629
rect 7170 1595 7204 1629
rect 7098 1527 7132 1561
rect 7170 1527 7204 1561
rect 7528 2411 7562 2445
rect 7732 2411 7766 2445
rect 7528 2343 7562 2377
rect 7732 2343 7766 2377
rect 7528 2275 7562 2309
rect 7732 2275 7766 2309
rect 7528 2207 7562 2241
rect 7732 2207 7766 2241
rect 7528 2139 7562 2173
rect 7732 2139 7766 2173
rect 7528 2071 7562 2105
rect 7732 2071 7766 2105
rect 7528 2003 7562 2037
rect 7732 2003 7766 2037
rect 7528 1935 7562 1969
rect 7732 1935 7766 1969
rect 7528 1867 7562 1901
rect 7732 1867 7766 1901
rect 7528 1799 7562 1833
rect 7732 1799 7766 1833
rect 7528 1731 7562 1765
rect 7732 1731 7766 1765
rect 7528 1663 7562 1697
rect 7732 1663 7766 1697
rect 7528 1595 7562 1629
rect 7732 1595 7766 1629
rect 7528 1527 7562 1561
rect 7732 1527 7766 1561
rect 8090 2411 8124 2445
rect 8162 2411 8196 2445
rect 8090 2343 8124 2377
rect 8162 2343 8196 2377
rect 8090 2275 8124 2309
rect 8162 2275 8196 2309
rect 8090 2207 8124 2241
rect 8162 2207 8196 2241
rect 8090 2139 8124 2173
rect 8162 2139 8196 2173
rect 8090 2071 8124 2105
rect 8162 2071 8196 2105
rect 8090 2003 8124 2037
rect 8162 2003 8196 2037
rect 8090 1935 8124 1969
rect 8162 1935 8196 1969
rect 8090 1867 8124 1901
rect 8162 1867 8196 1901
rect 8090 1799 8124 1833
rect 8162 1799 8196 1833
rect 8090 1731 8124 1765
rect 8162 1731 8196 1765
rect 8090 1663 8124 1697
rect 8162 1663 8196 1697
rect 8090 1595 8124 1629
rect 8162 1595 8196 1629
rect 8090 1527 8124 1561
rect 8162 1527 8196 1561
rect 8520 2411 8554 2445
rect 8724 2411 8758 2445
rect 8520 2343 8554 2377
rect 8724 2343 8758 2377
rect 8520 2275 8554 2309
rect 8724 2275 8758 2309
rect 8520 2207 8554 2241
rect 8724 2207 8758 2241
rect 8520 2139 8554 2173
rect 8724 2139 8758 2173
rect 8520 2071 8554 2105
rect 8724 2071 8758 2105
rect 8520 2003 8554 2037
rect 8724 2003 8758 2037
rect 8520 1935 8554 1969
rect 8724 1935 8758 1969
rect 8520 1867 8554 1901
rect 8724 1867 8758 1901
rect 8520 1799 8554 1833
rect 8724 1799 8758 1833
rect 8520 1731 8554 1765
rect 8724 1731 8758 1765
rect 8520 1663 8554 1697
rect 8724 1663 8758 1697
rect 8520 1595 8554 1629
rect 8724 1595 8758 1629
rect 8520 1527 8554 1561
rect 8724 1527 8758 1561
rect 9082 2411 9116 2445
rect 9154 2411 9188 2445
rect 9082 2343 9116 2377
rect 9154 2343 9188 2377
rect 9082 2275 9116 2309
rect 9154 2275 9188 2309
rect 9082 2207 9116 2241
rect 9154 2207 9188 2241
rect 9082 2139 9116 2173
rect 9154 2139 9188 2173
rect 9082 2071 9116 2105
rect 9154 2071 9188 2105
rect 9082 2003 9116 2037
rect 9154 2003 9188 2037
rect 9082 1935 9116 1969
rect 9154 1935 9188 1969
rect 9082 1867 9116 1901
rect 9154 1867 9188 1901
rect 9082 1799 9116 1833
rect 9154 1799 9188 1833
rect 9082 1731 9116 1765
rect 9154 1731 9188 1765
rect 9082 1663 9116 1697
rect 9154 1663 9188 1697
rect 9082 1595 9116 1629
rect 9154 1595 9188 1629
rect 9082 1527 9116 1561
rect 9154 1527 9188 1561
rect 9512 2411 9546 2445
rect 9716 2411 9750 2445
rect 9512 2343 9546 2377
rect 9716 2343 9750 2377
rect 9512 2275 9546 2309
rect 9716 2275 9750 2309
rect 9512 2207 9546 2241
rect 9716 2207 9750 2241
rect 9512 2139 9546 2173
rect 9716 2139 9750 2173
rect 9512 2071 9546 2105
rect 9716 2071 9750 2105
rect 9512 2003 9546 2037
rect 9716 2003 9750 2037
rect 9512 1935 9546 1969
rect 9716 1935 9750 1969
rect 9512 1867 9546 1901
rect 9716 1867 9750 1901
rect 9512 1799 9546 1833
rect 9716 1799 9750 1833
rect 9512 1731 9546 1765
rect 9716 1731 9750 1765
rect 9512 1663 9546 1697
rect 9716 1663 9750 1697
rect 9512 1595 9546 1629
rect 9716 1595 9750 1629
rect 9512 1527 9546 1561
rect 9716 1527 9750 1561
rect 10074 2411 10108 2445
rect 10146 2411 10180 2445
rect 10074 2343 10108 2377
rect 10146 2343 10180 2377
rect 10074 2275 10108 2309
rect 10146 2275 10180 2309
rect 10074 2207 10108 2241
rect 10146 2207 10180 2241
rect 10074 2139 10108 2173
rect 10146 2139 10180 2173
rect 10074 2071 10108 2105
rect 10146 2071 10180 2105
rect 10074 2003 10108 2037
rect 10146 2003 10180 2037
rect 10074 1935 10108 1969
rect 10146 1935 10180 1969
rect 10074 1867 10108 1901
rect 10146 1867 10180 1901
rect 10074 1799 10108 1833
rect 10146 1799 10180 1833
rect 10074 1731 10108 1765
rect 10146 1731 10180 1765
rect 10074 1663 10108 1697
rect 10146 1663 10180 1697
rect 10074 1595 10108 1629
rect 10146 1595 10180 1629
rect 10074 1527 10108 1561
rect 10146 1527 10180 1561
rect 10504 2411 10538 2445
rect 10708 2411 10742 2445
rect 10504 2343 10538 2377
rect 10708 2343 10742 2377
rect 10504 2275 10538 2309
rect 10708 2275 10742 2309
rect 10504 2207 10538 2241
rect 10708 2207 10742 2241
rect 10504 2139 10538 2173
rect 10708 2139 10742 2173
rect 10504 2071 10538 2105
rect 10708 2071 10742 2105
rect 10504 2003 10538 2037
rect 10708 2003 10742 2037
rect 10504 1935 10538 1969
rect 10708 1935 10742 1969
rect 10504 1867 10538 1901
rect 10708 1867 10742 1901
rect 10504 1799 10538 1833
rect 10708 1799 10742 1833
rect 10504 1731 10538 1765
rect 10708 1731 10742 1765
rect 10504 1663 10538 1697
rect 10708 1663 10742 1697
rect 10504 1595 10538 1629
rect 10708 1595 10742 1629
rect 10504 1527 10538 1561
rect 10708 1527 10742 1561
rect 11066 2411 11100 2445
rect 11138 2411 11172 2445
rect 11066 2343 11100 2377
rect 11138 2343 11172 2377
rect 11066 2275 11100 2309
rect 11138 2275 11172 2309
rect 11066 2207 11100 2241
rect 11138 2207 11172 2241
rect 11066 2139 11100 2173
rect 11138 2139 11172 2173
rect 11066 2071 11100 2105
rect 11138 2071 11172 2105
rect 11066 2003 11100 2037
rect 11138 2003 11172 2037
rect 11066 1935 11100 1969
rect 11138 1935 11172 1969
rect 11066 1867 11100 1901
rect 11138 1867 11172 1901
rect 11066 1799 11100 1833
rect 11138 1799 11172 1833
rect 11066 1731 11100 1765
rect 11138 1731 11172 1765
rect 11066 1663 11100 1697
rect 11138 1663 11172 1697
rect 11066 1595 11100 1629
rect 11138 1595 11172 1629
rect 11066 1527 11100 1561
rect 11138 1527 11172 1561
rect 11496 2411 11530 2445
rect 11700 2411 11734 2445
rect 11496 2343 11530 2377
rect 11700 2343 11734 2377
rect 11496 2275 11530 2309
rect 11700 2275 11734 2309
rect 11496 2207 11530 2241
rect 11700 2207 11734 2241
rect 11496 2139 11530 2173
rect 11700 2139 11734 2173
rect 11496 2071 11530 2105
rect 11700 2071 11734 2105
rect 11496 2003 11530 2037
rect 11700 2003 11734 2037
rect 11496 1935 11530 1969
rect 11700 1935 11734 1969
rect 11496 1867 11530 1901
rect 11700 1867 11734 1901
rect 11496 1799 11530 1833
rect 11700 1799 11734 1833
rect 11496 1731 11530 1765
rect 11700 1731 11734 1765
rect 11496 1663 11530 1697
rect 11700 1663 11734 1697
rect 11496 1595 11530 1629
rect 11700 1595 11734 1629
rect 11496 1527 11530 1561
rect 11700 1527 11734 1561
rect 12058 2411 12092 2445
rect 12130 2411 12164 2445
rect 12058 2343 12092 2377
rect 12130 2343 12164 2377
rect 12058 2275 12092 2309
rect 12130 2275 12164 2309
rect 12058 2207 12092 2241
rect 12130 2207 12164 2241
rect 12058 2139 12092 2173
rect 12130 2139 12164 2173
rect 12058 2071 12092 2105
rect 12130 2071 12164 2105
rect 12058 2003 12092 2037
rect 12130 2003 12164 2037
rect 12058 1935 12092 1969
rect 12130 1935 12164 1969
rect 12058 1867 12092 1901
rect 12130 1867 12164 1901
rect 12058 1799 12092 1833
rect 12130 1799 12164 1833
rect 12058 1731 12092 1765
rect 12130 1731 12164 1765
rect 12058 1663 12092 1697
rect 12130 1663 12164 1697
rect 12058 1595 12092 1629
rect 12130 1595 12164 1629
rect 12058 1527 12092 1561
rect 12130 1527 12164 1561
rect 12488 2411 12522 2445
rect 12692 2411 12726 2445
rect 12488 2343 12522 2377
rect 12692 2343 12726 2377
rect 12488 2275 12522 2309
rect 12692 2275 12726 2309
rect 12488 2207 12522 2241
rect 12692 2207 12726 2241
rect 12488 2139 12522 2173
rect 12692 2139 12726 2173
rect 12488 2071 12522 2105
rect 12692 2071 12726 2105
rect 12488 2003 12522 2037
rect 12692 2003 12726 2037
rect 12488 1935 12522 1969
rect 12692 1935 12726 1969
rect 12488 1867 12522 1901
rect 12692 1867 12726 1901
rect 12488 1799 12522 1833
rect 12692 1799 12726 1833
rect 12488 1731 12522 1765
rect 12692 1731 12726 1765
rect 12488 1663 12522 1697
rect 12692 1663 12726 1697
rect 12488 1595 12522 1629
rect 12692 1595 12726 1629
rect 12488 1527 12522 1561
rect 12692 1527 12726 1561
rect 13050 2411 13084 2445
rect 13122 2411 13156 2445
rect 13050 2343 13084 2377
rect 13122 2343 13156 2377
rect 13050 2275 13084 2309
rect 13122 2275 13156 2309
rect 13050 2207 13084 2241
rect 13122 2207 13156 2241
rect 13050 2139 13084 2173
rect 13122 2139 13156 2173
rect 13050 2071 13084 2105
rect 13122 2071 13156 2105
rect 13050 2003 13084 2037
rect 13122 2003 13156 2037
rect 13050 1935 13084 1969
rect 13122 1935 13156 1969
rect 13050 1867 13084 1901
rect 13122 1867 13156 1901
rect 13050 1799 13084 1833
rect 13122 1799 13156 1833
rect 13050 1731 13084 1765
rect 13122 1731 13156 1765
rect 13050 1663 13084 1697
rect 13122 1663 13156 1697
rect 13050 1595 13084 1629
rect 13122 1595 13156 1629
rect 13050 1527 13084 1561
rect 13122 1527 13156 1561
rect 13480 2411 13514 2445
rect 13684 2411 13718 2445
rect 13480 2343 13514 2377
rect 13684 2343 13718 2377
rect 13480 2275 13514 2309
rect 13684 2275 13718 2309
rect 13480 2207 13514 2241
rect 13684 2207 13718 2241
rect 13480 2139 13514 2173
rect 13684 2139 13718 2173
rect 13480 2071 13514 2105
rect 13684 2071 13718 2105
rect 13480 2003 13514 2037
rect 13684 2003 13718 2037
rect 13480 1935 13514 1969
rect 13684 1935 13718 1969
rect 13480 1867 13514 1901
rect 13684 1867 13718 1901
rect 13480 1799 13514 1833
rect 13684 1799 13718 1833
rect 13480 1731 13514 1765
rect 13684 1731 13718 1765
rect 13480 1663 13514 1697
rect 13684 1663 13718 1697
rect 13480 1595 13514 1629
rect 13684 1595 13718 1629
rect 13480 1527 13514 1561
rect 13684 1527 13718 1561
rect 14042 2411 14076 2445
rect 14042 2343 14076 2377
rect 14042 2275 14076 2309
rect 14042 2207 14076 2241
rect 14042 2139 14076 2173
rect 14042 2071 14076 2105
rect 14042 2003 14076 2037
rect 14042 1935 14076 1969
rect 14042 1867 14076 1901
rect 14042 1799 14076 1833
rect 14042 1731 14076 1765
rect 14042 1663 14076 1697
rect 14042 1595 14076 1629
rect 14042 1527 14076 1561
rect 14386 2411 14420 2445
rect 14386 2343 14420 2377
rect 14386 2275 14420 2309
rect 14386 2207 14420 2241
rect 14386 2139 14420 2173
rect 14386 2071 14420 2105
rect 14386 2003 14420 2037
rect 14386 1935 14420 1969
rect 14386 1867 14420 1901
rect 14386 1799 14420 1833
rect 14386 1731 14420 1765
rect 14386 1663 14420 1697
rect 14386 1595 14420 1629
rect 14386 1527 14420 1561
<< nsubdiff >>
rect 14948 490 14990 579
<< mvpsubdiff >>
rect 555 4922 657 4956
rect 14495 4922 14530 4956
rect 14564 4922 14599 4956
rect 14633 4922 14667 4956
rect 589 4888 657 4922
rect 14461 4888 14667 4922
rect 555 4854 623 4888
rect 14461 4854 14496 4888
rect 14530 4854 14565 4888
rect 14599 4854 14667 4888
rect 555 4850 691 4854
rect 589 4819 691 4850
rect 589 4816 623 4819
rect 555 4785 623 4816
rect 657 4786 691 4819
rect 14393 4844 14667 4854
rect 14393 4820 14633 4844
rect 14393 4786 14428 4820
rect 14462 4786 14497 4820
rect 14531 4818 14633 4820
rect 14531 4786 14565 4818
rect 657 4785 725 4786
rect 555 4778 725 4785
rect 589 4751 725 4778
rect 589 4750 691 4751
rect 589 4744 623 4750
rect 555 4716 623 4744
rect 657 4717 691 4750
rect 657 4716 725 4717
rect 555 4706 725 4716
rect 589 4682 725 4706
rect 589 4681 691 4682
rect 589 4672 623 4681
rect 555 4647 623 4672
rect 657 4648 691 4681
rect 657 4647 725 4648
rect 555 4634 725 4647
rect 589 4613 725 4634
rect 589 4600 623 4613
rect 555 4563 623 4600
rect 589 4529 623 4563
rect 555 4492 623 4529
rect 589 4458 623 4492
rect 555 4421 623 4458
rect 589 4387 623 4421
rect 555 4350 623 4387
rect 589 4316 623 4350
rect 555 4279 623 4316
rect 589 4245 623 4279
rect 555 4208 623 4245
rect 589 4174 623 4208
rect 555 4137 623 4174
rect 589 4103 623 4137
rect 14497 4784 14565 4786
rect 14599 4810 14633 4818
rect 14599 4784 14667 4810
rect 14497 4771 14667 4784
rect 14497 4750 14633 4771
rect 14531 4748 14633 4750
rect 14531 4716 14565 4748
rect 14497 4714 14565 4716
rect 14599 4737 14633 4748
rect 14599 4714 14667 4737
rect 14497 4698 14667 4714
rect 14497 4680 14633 4698
rect 14531 4678 14633 4680
rect 14531 4646 14565 4678
rect 14497 4644 14565 4646
rect 14599 4664 14633 4678
rect 14599 4644 14667 4664
rect 14497 4625 14667 4644
rect 14497 4610 14633 4625
rect 14531 4608 14633 4610
rect 14531 4576 14565 4608
rect 14497 4574 14565 4576
rect 14599 4591 14633 4608
rect 14599 4574 14667 4591
rect 14497 4552 14667 4574
rect 14497 4540 14633 4552
rect 14531 4538 14633 4540
rect 14531 4506 14565 4538
rect 14497 4504 14565 4506
rect 14599 4518 14633 4538
rect 14599 4504 14667 4518
rect 14497 4479 14667 4504
rect 14497 4470 14633 4479
rect 14531 4468 14633 4470
rect 14531 4436 14565 4468
rect 14497 4434 14565 4436
rect 14599 4445 14633 4468
rect 14599 4434 14667 4445
rect 14497 4406 14667 4434
rect 14497 4399 14633 4406
rect 14531 4398 14633 4399
rect 14531 4365 14565 4398
rect 14497 4364 14565 4365
rect 14599 4372 14633 4398
rect 14599 4364 14667 4372
rect 14497 4333 14667 4364
rect 14497 4328 14633 4333
rect 14531 4294 14565 4328
rect 14599 4299 14633 4328
rect 14599 4294 14667 4299
rect 14497 4260 14667 4294
rect 14497 4257 14633 4260
rect 555 4058 725 4103
rect 14531 4223 14565 4257
rect 14599 4226 14633 4257
rect 14599 4223 14667 4226
rect 14497 4186 14667 4223
rect 14531 4152 14565 4186
rect 14599 4152 14633 4186
rect 14497 4115 14667 4152
rect 14497 4081 14565 4115
rect 14599 4081 14633 4115
rect 14497 4058 14667 4081
rect 555 4041 787 4058
rect 589 4007 623 4041
rect 657 4034 787 4041
rect 657 4007 734 4034
rect 555 4000 734 4007
rect 768 4000 787 4034
rect 555 3970 787 4000
rect 589 3936 623 3970
rect 657 3966 787 3970
rect 657 3936 734 3966
rect 555 3932 734 3936
rect 768 3932 787 3966
rect 555 3898 787 3932
rect 555 3896 734 3898
rect 589 3862 623 3896
rect 657 3864 734 3896
rect 768 3864 787 3898
rect 657 3862 787 3864
rect 555 3830 787 3862
rect 555 3825 734 3830
rect 589 3791 623 3825
rect 657 3796 734 3825
rect 768 3796 787 3830
rect 657 3791 787 3796
rect 555 3762 787 3791
rect 555 3751 734 3762
rect 589 3717 623 3751
rect 657 3728 734 3751
rect 768 3728 787 3762
rect 657 3717 787 3728
rect 555 3694 787 3717
rect 555 3680 734 3694
rect 589 3646 623 3680
rect 657 3660 734 3680
rect 768 3660 787 3694
rect 657 3646 787 3660
rect 555 3626 787 3646
rect 555 3606 734 3626
rect 589 3572 623 3606
rect 657 3592 734 3606
rect 768 3592 787 3626
rect 657 3572 787 3592
rect 555 3558 787 3572
rect 555 3535 734 3558
rect 589 3501 623 3535
rect 657 3524 734 3535
rect 768 3524 787 3558
rect 657 3501 787 3524
rect 555 3490 787 3501
rect 555 3461 734 3490
rect 589 3427 623 3461
rect 657 3456 734 3461
rect 768 3456 787 3490
rect 657 3427 787 3456
rect 555 3422 787 3427
rect 555 3390 734 3422
rect 589 3356 623 3390
rect 657 3388 734 3390
rect 768 3388 787 3422
rect 657 3356 787 3388
rect 555 3354 787 3356
rect 555 3320 734 3354
rect 768 3320 787 3354
rect 555 3316 787 3320
rect 589 3282 623 3316
rect 657 3286 787 3316
rect 657 3282 734 3286
rect 555 3252 734 3282
rect 768 3252 787 3286
rect 555 3245 787 3252
rect 589 3211 623 3245
rect 657 3218 787 3245
rect 657 3211 734 3218
rect 555 3184 734 3211
rect 768 3184 787 3218
rect 555 3151 787 3184
rect 589 3117 623 3151
rect 657 3150 787 3151
rect 657 3117 734 3150
rect 555 3116 734 3117
rect 768 3116 787 3150
rect 555 3081 787 3116
rect 657 3058 787 3081
rect 1625 4046 1765 4058
rect 1625 4012 1678 4046
rect 1712 4012 1765 4046
rect 1625 3978 1765 4012
rect 1625 3944 1678 3978
rect 1712 3944 1765 3978
rect 1625 3910 1765 3944
rect 1625 3876 1678 3910
rect 1712 3876 1765 3910
rect 1625 3842 1765 3876
rect 1625 3808 1678 3842
rect 1712 3808 1765 3842
rect 1625 3774 1765 3808
rect 1625 3740 1678 3774
rect 1712 3740 1765 3774
rect 1625 3706 1765 3740
rect 1625 3672 1678 3706
rect 1712 3672 1765 3706
rect 1625 3638 1765 3672
rect 1625 3604 1678 3638
rect 1712 3604 1765 3638
rect 1625 3570 1765 3604
rect 1625 3536 1678 3570
rect 1712 3536 1765 3570
rect 1625 3502 1765 3536
rect 1625 3468 1678 3502
rect 1712 3468 1765 3502
rect 1625 3434 1765 3468
rect 1625 3400 1678 3434
rect 1712 3400 1765 3434
rect 1625 3366 1765 3400
rect 1625 3332 1678 3366
rect 1712 3332 1765 3366
rect 1625 3298 1765 3332
rect 1625 3264 1678 3298
rect 1712 3264 1765 3298
rect 1625 3230 1765 3264
rect 1625 3196 1678 3230
rect 1712 3196 1765 3230
rect 1625 3162 1765 3196
rect 1625 3128 1678 3162
rect 1712 3128 1765 3162
rect 1625 3058 1765 3128
rect 2617 4046 2757 4058
rect 2617 4012 2670 4046
rect 2704 4012 2757 4046
rect 2617 3978 2757 4012
rect 2617 3944 2670 3978
rect 2704 3944 2757 3978
rect 2617 3910 2757 3944
rect 2617 3876 2670 3910
rect 2704 3876 2757 3910
rect 2617 3842 2757 3876
rect 2617 3808 2670 3842
rect 2704 3808 2757 3842
rect 2617 3774 2757 3808
rect 2617 3740 2670 3774
rect 2704 3740 2757 3774
rect 2617 3706 2757 3740
rect 2617 3672 2670 3706
rect 2704 3672 2757 3706
rect 2617 3638 2757 3672
rect 2617 3604 2670 3638
rect 2704 3604 2757 3638
rect 2617 3570 2757 3604
rect 2617 3536 2670 3570
rect 2704 3536 2757 3570
rect 2617 3502 2757 3536
rect 2617 3468 2670 3502
rect 2704 3468 2757 3502
rect 2617 3434 2757 3468
rect 2617 3400 2670 3434
rect 2704 3400 2757 3434
rect 2617 3366 2757 3400
rect 2617 3332 2670 3366
rect 2704 3332 2757 3366
rect 2617 3298 2757 3332
rect 2617 3264 2670 3298
rect 2704 3264 2757 3298
rect 2617 3230 2757 3264
rect 2617 3196 2670 3230
rect 2704 3196 2757 3230
rect 2617 3162 2757 3196
rect 2617 3128 2670 3162
rect 2704 3128 2757 3162
rect 2617 3058 2757 3128
rect 3609 4046 3749 4058
rect 3609 4012 3662 4046
rect 3696 4012 3749 4046
rect 3609 3978 3749 4012
rect 3609 3944 3662 3978
rect 3696 3944 3749 3978
rect 3609 3910 3749 3944
rect 3609 3876 3662 3910
rect 3696 3876 3749 3910
rect 3609 3842 3749 3876
rect 3609 3808 3662 3842
rect 3696 3808 3749 3842
rect 3609 3774 3749 3808
rect 3609 3740 3662 3774
rect 3696 3740 3749 3774
rect 3609 3706 3749 3740
rect 3609 3672 3662 3706
rect 3696 3672 3749 3706
rect 3609 3638 3749 3672
rect 3609 3604 3662 3638
rect 3696 3604 3749 3638
rect 3609 3570 3749 3604
rect 3609 3536 3662 3570
rect 3696 3536 3749 3570
rect 3609 3502 3749 3536
rect 3609 3468 3662 3502
rect 3696 3468 3749 3502
rect 3609 3434 3749 3468
rect 3609 3400 3662 3434
rect 3696 3400 3749 3434
rect 3609 3366 3749 3400
rect 3609 3332 3662 3366
rect 3696 3332 3749 3366
rect 3609 3298 3749 3332
rect 3609 3264 3662 3298
rect 3696 3264 3749 3298
rect 3609 3230 3749 3264
rect 3609 3196 3662 3230
rect 3696 3196 3749 3230
rect 3609 3162 3749 3196
rect 3609 3128 3662 3162
rect 3696 3128 3749 3162
rect 3609 3058 3749 3128
rect 4601 4046 4741 4058
rect 4601 4012 4654 4046
rect 4688 4012 4741 4046
rect 4601 3978 4741 4012
rect 4601 3944 4654 3978
rect 4688 3944 4741 3978
rect 4601 3910 4741 3944
rect 4601 3876 4654 3910
rect 4688 3876 4741 3910
rect 4601 3842 4741 3876
rect 4601 3808 4654 3842
rect 4688 3808 4741 3842
rect 4601 3774 4741 3808
rect 4601 3740 4654 3774
rect 4688 3740 4741 3774
rect 4601 3706 4741 3740
rect 4601 3672 4654 3706
rect 4688 3672 4741 3706
rect 4601 3638 4741 3672
rect 4601 3604 4654 3638
rect 4688 3604 4741 3638
rect 4601 3570 4741 3604
rect 4601 3536 4654 3570
rect 4688 3536 4741 3570
rect 4601 3502 4741 3536
rect 4601 3468 4654 3502
rect 4688 3468 4741 3502
rect 4601 3434 4741 3468
rect 4601 3400 4654 3434
rect 4688 3400 4741 3434
rect 4601 3366 4741 3400
rect 4601 3332 4654 3366
rect 4688 3332 4741 3366
rect 4601 3298 4741 3332
rect 4601 3264 4654 3298
rect 4688 3264 4741 3298
rect 4601 3230 4741 3264
rect 4601 3196 4654 3230
rect 4688 3196 4741 3230
rect 4601 3162 4741 3196
rect 4601 3128 4654 3162
rect 4688 3128 4741 3162
rect 4601 3058 4741 3128
rect 5593 4046 5733 4058
rect 5593 4012 5646 4046
rect 5680 4012 5733 4046
rect 5593 3978 5733 4012
rect 5593 3944 5646 3978
rect 5680 3944 5733 3978
rect 5593 3910 5733 3944
rect 5593 3876 5646 3910
rect 5680 3876 5733 3910
rect 5593 3842 5733 3876
rect 5593 3808 5646 3842
rect 5680 3808 5733 3842
rect 5593 3774 5733 3808
rect 5593 3740 5646 3774
rect 5680 3740 5733 3774
rect 5593 3706 5733 3740
rect 5593 3672 5646 3706
rect 5680 3672 5733 3706
rect 5593 3638 5733 3672
rect 5593 3604 5646 3638
rect 5680 3604 5733 3638
rect 5593 3570 5733 3604
rect 5593 3536 5646 3570
rect 5680 3536 5733 3570
rect 5593 3502 5733 3536
rect 5593 3468 5646 3502
rect 5680 3468 5733 3502
rect 5593 3434 5733 3468
rect 5593 3400 5646 3434
rect 5680 3400 5733 3434
rect 5593 3366 5733 3400
rect 5593 3332 5646 3366
rect 5680 3332 5733 3366
rect 5593 3298 5733 3332
rect 5593 3264 5646 3298
rect 5680 3264 5733 3298
rect 5593 3230 5733 3264
rect 5593 3196 5646 3230
rect 5680 3196 5733 3230
rect 5593 3162 5733 3196
rect 5593 3128 5646 3162
rect 5680 3128 5733 3162
rect 5593 3058 5733 3128
rect 6585 4046 6725 4058
rect 6585 4012 6638 4046
rect 6672 4012 6725 4046
rect 6585 3978 6725 4012
rect 6585 3944 6638 3978
rect 6672 3944 6725 3978
rect 6585 3910 6725 3944
rect 6585 3876 6638 3910
rect 6672 3876 6725 3910
rect 6585 3842 6725 3876
rect 6585 3808 6638 3842
rect 6672 3808 6725 3842
rect 6585 3774 6725 3808
rect 6585 3740 6638 3774
rect 6672 3740 6725 3774
rect 6585 3706 6725 3740
rect 6585 3672 6638 3706
rect 6672 3672 6725 3706
rect 6585 3638 6725 3672
rect 6585 3604 6638 3638
rect 6672 3604 6725 3638
rect 6585 3570 6725 3604
rect 6585 3536 6638 3570
rect 6672 3536 6725 3570
rect 6585 3502 6725 3536
rect 6585 3468 6638 3502
rect 6672 3468 6725 3502
rect 6585 3434 6725 3468
rect 6585 3400 6638 3434
rect 6672 3400 6725 3434
rect 6585 3366 6725 3400
rect 6585 3332 6638 3366
rect 6672 3332 6725 3366
rect 6585 3298 6725 3332
rect 6585 3264 6638 3298
rect 6672 3264 6725 3298
rect 6585 3230 6725 3264
rect 6585 3196 6638 3230
rect 6672 3196 6725 3230
rect 6585 3162 6725 3196
rect 6585 3128 6638 3162
rect 6672 3128 6725 3162
rect 6585 3058 6725 3128
rect 7577 4046 7717 4058
rect 7577 4012 7630 4046
rect 7664 4012 7717 4046
rect 7577 3978 7717 4012
rect 7577 3944 7630 3978
rect 7664 3944 7717 3978
rect 7577 3910 7717 3944
rect 7577 3876 7630 3910
rect 7664 3876 7717 3910
rect 7577 3842 7717 3876
rect 7577 3808 7630 3842
rect 7664 3808 7717 3842
rect 7577 3774 7717 3808
rect 7577 3740 7630 3774
rect 7664 3740 7717 3774
rect 7577 3706 7717 3740
rect 7577 3672 7630 3706
rect 7664 3672 7717 3706
rect 7577 3638 7717 3672
rect 7577 3604 7630 3638
rect 7664 3604 7717 3638
rect 7577 3570 7717 3604
rect 7577 3536 7630 3570
rect 7664 3536 7717 3570
rect 7577 3502 7717 3536
rect 7577 3468 7630 3502
rect 7664 3468 7717 3502
rect 7577 3434 7717 3468
rect 7577 3400 7630 3434
rect 7664 3400 7717 3434
rect 7577 3366 7717 3400
rect 7577 3332 7630 3366
rect 7664 3332 7717 3366
rect 7577 3298 7717 3332
rect 7577 3264 7630 3298
rect 7664 3264 7717 3298
rect 7577 3230 7717 3264
rect 7577 3196 7630 3230
rect 7664 3196 7717 3230
rect 7577 3162 7717 3196
rect 7577 3128 7630 3162
rect 7664 3128 7717 3162
rect 7577 3058 7717 3128
rect 8569 4046 8709 4058
rect 8569 4012 8622 4046
rect 8656 4012 8709 4046
rect 8569 3978 8709 4012
rect 8569 3944 8622 3978
rect 8656 3944 8709 3978
rect 8569 3910 8709 3944
rect 8569 3876 8622 3910
rect 8656 3876 8709 3910
rect 8569 3842 8709 3876
rect 8569 3808 8622 3842
rect 8656 3808 8709 3842
rect 8569 3774 8709 3808
rect 8569 3740 8622 3774
rect 8656 3740 8709 3774
rect 8569 3706 8709 3740
rect 8569 3672 8622 3706
rect 8656 3672 8709 3706
rect 8569 3638 8709 3672
rect 8569 3604 8622 3638
rect 8656 3604 8709 3638
rect 8569 3570 8709 3604
rect 8569 3536 8622 3570
rect 8656 3536 8709 3570
rect 8569 3502 8709 3536
rect 8569 3468 8622 3502
rect 8656 3468 8709 3502
rect 8569 3434 8709 3468
rect 8569 3400 8622 3434
rect 8656 3400 8709 3434
rect 8569 3366 8709 3400
rect 8569 3332 8622 3366
rect 8656 3332 8709 3366
rect 8569 3298 8709 3332
rect 8569 3264 8622 3298
rect 8656 3264 8709 3298
rect 8569 3230 8709 3264
rect 8569 3196 8622 3230
rect 8656 3196 8709 3230
rect 8569 3162 8709 3196
rect 8569 3128 8622 3162
rect 8656 3128 8709 3162
rect 8569 3058 8709 3128
rect 9561 4046 9701 4058
rect 9561 4012 9614 4046
rect 9648 4012 9701 4046
rect 9561 3978 9701 4012
rect 9561 3944 9614 3978
rect 9648 3944 9701 3978
rect 9561 3910 9701 3944
rect 9561 3876 9614 3910
rect 9648 3876 9701 3910
rect 9561 3842 9701 3876
rect 9561 3808 9614 3842
rect 9648 3808 9701 3842
rect 9561 3774 9701 3808
rect 9561 3740 9614 3774
rect 9648 3740 9701 3774
rect 9561 3706 9701 3740
rect 9561 3672 9614 3706
rect 9648 3672 9701 3706
rect 9561 3638 9701 3672
rect 9561 3604 9614 3638
rect 9648 3604 9701 3638
rect 9561 3570 9701 3604
rect 9561 3536 9614 3570
rect 9648 3536 9701 3570
rect 9561 3502 9701 3536
rect 9561 3468 9614 3502
rect 9648 3468 9701 3502
rect 9561 3434 9701 3468
rect 9561 3400 9614 3434
rect 9648 3400 9701 3434
rect 9561 3366 9701 3400
rect 9561 3332 9614 3366
rect 9648 3332 9701 3366
rect 9561 3298 9701 3332
rect 9561 3264 9614 3298
rect 9648 3264 9701 3298
rect 9561 3230 9701 3264
rect 9561 3196 9614 3230
rect 9648 3196 9701 3230
rect 9561 3162 9701 3196
rect 9561 3128 9614 3162
rect 9648 3128 9701 3162
rect 9561 3058 9701 3128
rect 10553 4046 10693 4058
rect 10553 4012 10606 4046
rect 10640 4012 10693 4046
rect 10553 3978 10693 4012
rect 10553 3944 10606 3978
rect 10640 3944 10693 3978
rect 10553 3910 10693 3944
rect 10553 3876 10606 3910
rect 10640 3876 10693 3910
rect 10553 3842 10693 3876
rect 10553 3808 10606 3842
rect 10640 3808 10693 3842
rect 10553 3774 10693 3808
rect 10553 3740 10606 3774
rect 10640 3740 10693 3774
rect 10553 3706 10693 3740
rect 10553 3672 10606 3706
rect 10640 3672 10693 3706
rect 10553 3638 10693 3672
rect 10553 3604 10606 3638
rect 10640 3604 10693 3638
rect 10553 3570 10693 3604
rect 10553 3536 10606 3570
rect 10640 3536 10693 3570
rect 10553 3502 10693 3536
rect 10553 3468 10606 3502
rect 10640 3468 10693 3502
rect 10553 3434 10693 3468
rect 10553 3400 10606 3434
rect 10640 3400 10693 3434
rect 10553 3366 10693 3400
rect 10553 3332 10606 3366
rect 10640 3332 10693 3366
rect 10553 3298 10693 3332
rect 10553 3264 10606 3298
rect 10640 3264 10693 3298
rect 10553 3230 10693 3264
rect 10553 3196 10606 3230
rect 10640 3196 10693 3230
rect 10553 3162 10693 3196
rect 10553 3128 10606 3162
rect 10640 3128 10693 3162
rect 10553 3058 10693 3128
rect 11545 4046 11685 4058
rect 11545 4012 11598 4046
rect 11632 4012 11685 4046
rect 11545 3978 11685 4012
rect 11545 3944 11598 3978
rect 11632 3944 11685 3978
rect 11545 3910 11685 3944
rect 11545 3876 11598 3910
rect 11632 3876 11685 3910
rect 11545 3842 11685 3876
rect 11545 3808 11598 3842
rect 11632 3808 11685 3842
rect 11545 3774 11685 3808
rect 11545 3740 11598 3774
rect 11632 3740 11685 3774
rect 11545 3706 11685 3740
rect 11545 3672 11598 3706
rect 11632 3672 11685 3706
rect 11545 3638 11685 3672
rect 11545 3604 11598 3638
rect 11632 3604 11685 3638
rect 11545 3570 11685 3604
rect 11545 3536 11598 3570
rect 11632 3536 11685 3570
rect 11545 3502 11685 3536
rect 11545 3468 11598 3502
rect 11632 3468 11685 3502
rect 11545 3434 11685 3468
rect 11545 3400 11598 3434
rect 11632 3400 11685 3434
rect 11545 3366 11685 3400
rect 11545 3332 11598 3366
rect 11632 3332 11685 3366
rect 11545 3298 11685 3332
rect 11545 3264 11598 3298
rect 11632 3264 11685 3298
rect 11545 3230 11685 3264
rect 11545 3196 11598 3230
rect 11632 3196 11685 3230
rect 11545 3162 11685 3196
rect 11545 3128 11598 3162
rect 11632 3128 11685 3162
rect 11545 3058 11685 3128
rect 12537 4046 12677 4058
rect 12537 4012 12590 4046
rect 12624 4012 12677 4046
rect 12537 3978 12677 4012
rect 12537 3944 12590 3978
rect 12624 3944 12677 3978
rect 12537 3910 12677 3944
rect 12537 3876 12590 3910
rect 12624 3876 12677 3910
rect 12537 3842 12677 3876
rect 12537 3808 12590 3842
rect 12624 3808 12677 3842
rect 12537 3774 12677 3808
rect 12537 3740 12590 3774
rect 12624 3740 12677 3774
rect 12537 3706 12677 3740
rect 12537 3672 12590 3706
rect 12624 3672 12677 3706
rect 12537 3638 12677 3672
rect 12537 3604 12590 3638
rect 12624 3604 12677 3638
rect 12537 3570 12677 3604
rect 12537 3536 12590 3570
rect 12624 3536 12677 3570
rect 12537 3502 12677 3536
rect 12537 3468 12590 3502
rect 12624 3468 12677 3502
rect 12537 3434 12677 3468
rect 12537 3400 12590 3434
rect 12624 3400 12677 3434
rect 12537 3366 12677 3400
rect 12537 3332 12590 3366
rect 12624 3332 12677 3366
rect 12537 3298 12677 3332
rect 12537 3264 12590 3298
rect 12624 3264 12677 3298
rect 12537 3230 12677 3264
rect 12537 3196 12590 3230
rect 12624 3196 12677 3230
rect 12537 3162 12677 3196
rect 12537 3128 12590 3162
rect 12624 3128 12677 3162
rect 12537 3058 12677 3128
rect 13529 4046 13669 4058
rect 13529 4012 13582 4046
rect 13616 4012 13669 4046
rect 13529 3978 13669 4012
rect 13529 3944 13582 3978
rect 13616 3944 13669 3978
rect 13529 3910 13669 3944
rect 13529 3876 13582 3910
rect 13616 3876 13669 3910
rect 13529 3842 13669 3876
rect 13529 3808 13582 3842
rect 13616 3808 13669 3842
rect 13529 3774 13669 3808
rect 13529 3740 13582 3774
rect 13616 3740 13669 3774
rect 13529 3706 13669 3740
rect 13529 3672 13582 3706
rect 13616 3672 13669 3706
rect 13529 3638 13669 3672
rect 13529 3604 13582 3638
rect 13616 3604 13669 3638
rect 13529 3570 13669 3604
rect 13529 3536 13582 3570
rect 13616 3536 13669 3570
rect 13529 3502 13669 3536
rect 13529 3468 13582 3502
rect 13616 3468 13669 3502
rect 13529 3434 13669 3468
rect 13529 3400 13582 3434
rect 13616 3400 13669 3434
rect 13529 3366 13669 3400
rect 13529 3332 13582 3366
rect 13616 3332 13669 3366
rect 13529 3298 13669 3332
rect 13529 3264 13582 3298
rect 13616 3264 13669 3298
rect 13529 3230 13669 3264
rect 13529 3196 13582 3230
rect 13616 3196 13669 3230
rect 13529 3162 13669 3196
rect 13529 3128 13582 3162
rect 13616 3128 13669 3162
rect 13529 3058 13669 3128
rect 14435 4041 14667 4058
rect 14435 4034 14565 4041
rect 14435 4000 14454 4034
rect 14488 4007 14565 4034
rect 14599 4007 14633 4041
rect 14488 4000 14667 4007
rect 14435 3970 14667 4000
rect 14435 3966 14565 3970
rect 14435 3932 14454 3966
rect 14488 3936 14565 3966
rect 14599 3936 14633 3970
rect 14488 3932 14667 3936
rect 14435 3898 14667 3932
rect 14435 3864 14454 3898
rect 14488 3896 14667 3898
rect 14488 3864 14565 3896
rect 14435 3862 14565 3864
rect 14599 3862 14633 3896
rect 14435 3830 14667 3862
rect 14435 3796 14454 3830
rect 14488 3825 14667 3830
rect 14488 3796 14565 3825
rect 14435 3791 14565 3796
rect 14599 3791 14633 3825
rect 14435 3762 14667 3791
rect 14435 3728 14454 3762
rect 14488 3751 14667 3762
rect 14488 3728 14565 3751
rect 14435 3717 14565 3728
rect 14599 3717 14633 3751
rect 14435 3694 14667 3717
rect 14435 3660 14454 3694
rect 14488 3680 14667 3694
rect 14488 3660 14565 3680
rect 14435 3646 14565 3660
rect 14599 3646 14633 3680
rect 14435 3626 14667 3646
rect 14435 3592 14454 3626
rect 14488 3606 14667 3626
rect 14488 3592 14565 3606
rect 14435 3572 14565 3592
rect 14599 3572 14633 3606
rect 14435 3558 14667 3572
rect 14435 3524 14454 3558
rect 14488 3535 14667 3558
rect 14488 3524 14565 3535
rect 14435 3501 14565 3524
rect 14599 3501 14633 3535
rect 14435 3490 14667 3501
rect 14435 3456 14454 3490
rect 14488 3461 14667 3490
rect 14488 3456 14565 3461
rect 14435 3427 14565 3456
rect 14599 3427 14633 3461
rect 14435 3422 14667 3427
rect 14435 3388 14454 3422
rect 14488 3390 14667 3422
rect 14488 3388 14565 3390
rect 14435 3356 14565 3388
rect 14599 3356 14633 3390
rect 14435 3354 14667 3356
rect 14435 3320 14454 3354
rect 14488 3320 14667 3354
rect 14435 3316 14667 3320
rect 14435 3286 14565 3316
rect 14435 3252 14454 3286
rect 14488 3282 14565 3286
rect 14599 3282 14633 3316
rect 14488 3252 14667 3282
rect 14435 3245 14667 3252
rect 14435 3218 14565 3245
rect 14435 3184 14454 3218
rect 14488 3211 14565 3218
rect 14599 3211 14633 3245
rect 14488 3184 14667 3211
rect 14435 3151 14667 3184
rect 14435 3150 14565 3151
rect 14435 3116 14454 3150
rect 14488 3117 14565 3150
rect 14599 3117 14633 3151
rect 14488 3116 14667 3117
rect 14435 3066 14667 3116
rect 14435 3058 14565 3066
rect 657 3013 725 3058
rect 657 2457 725 2503
rect 1578 2935 1814 2969
rect 1578 2901 1645 2935
rect 1679 2901 1713 2935
rect 1747 2901 1814 2935
rect 1578 2855 1814 2901
rect 1578 2821 1645 2855
rect 1679 2821 1713 2855
rect 1747 2821 1814 2855
rect 1578 2775 1814 2821
rect 1578 2741 1645 2775
rect 1679 2741 1713 2775
rect 1747 2741 1814 2775
rect 1578 2695 1814 2741
rect 1578 2661 1645 2695
rect 1679 2661 1713 2695
rect 1747 2661 1814 2695
rect 1578 2614 1814 2661
rect 1578 2580 1645 2614
rect 1679 2580 1713 2614
rect 1747 2580 1814 2614
rect 1578 2546 1814 2580
rect 2570 2935 2806 2969
rect 2570 2901 2637 2935
rect 2671 2901 2705 2935
rect 2739 2901 2806 2935
rect 2570 2855 2806 2901
rect 2570 2821 2637 2855
rect 2671 2821 2705 2855
rect 2739 2821 2806 2855
rect 2570 2775 2806 2821
rect 2570 2741 2637 2775
rect 2671 2741 2705 2775
rect 2739 2741 2806 2775
rect 2570 2695 2806 2741
rect 2570 2661 2637 2695
rect 2671 2661 2705 2695
rect 2739 2661 2806 2695
rect 2570 2614 2806 2661
rect 2570 2580 2637 2614
rect 2671 2580 2705 2614
rect 2739 2580 2806 2614
rect 2570 2546 2806 2580
rect 3562 2935 3798 2969
rect 3562 2901 3629 2935
rect 3663 2901 3697 2935
rect 3731 2901 3798 2935
rect 3562 2855 3798 2901
rect 3562 2821 3629 2855
rect 3663 2821 3697 2855
rect 3731 2821 3798 2855
rect 3562 2775 3798 2821
rect 3562 2741 3629 2775
rect 3663 2741 3697 2775
rect 3731 2741 3798 2775
rect 3562 2695 3798 2741
rect 3562 2661 3629 2695
rect 3663 2661 3697 2695
rect 3731 2661 3798 2695
rect 3562 2614 3798 2661
rect 3562 2580 3629 2614
rect 3663 2580 3697 2614
rect 3731 2580 3798 2614
rect 3562 2546 3798 2580
rect 4554 2935 4790 2969
rect 4554 2901 4621 2935
rect 4655 2901 4689 2935
rect 4723 2901 4790 2935
rect 4554 2855 4790 2901
rect 4554 2821 4621 2855
rect 4655 2821 4689 2855
rect 4723 2821 4790 2855
rect 4554 2775 4790 2821
rect 4554 2741 4621 2775
rect 4655 2741 4689 2775
rect 4723 2741 4790 2775
rect 4554 2695 4790 2741
rect 4554 2661 4621 2695
rect 4655 2661 4689 2695
rect 4723 2661 4790 2695
rect 4554 2614 4790 2661
rect 4554 2580 4621 2614
rect 4655 2580 4689 2614
rect 4723 2580 4790 2614
rect 4554 2546 4790 2580
rect 5546 2935 5782 2969
rect 5546 2901 5613 2935
rect 5647 2901 5681 2935
rect 5715 2901 5782 2935
rect 5546 2855 5782 2901
rect 5546 2821 5613 2855
rect 5647 2821 5681 2855
rect 5715 2821 5782 2855
rect 5546 2775 5782 2821
rect 5546 2741 5613 2775
rect 5647 2741 5681 2775
rect 5715 2741 5782 2775
rect 5546 2695 5782 2741
rect 5546 2661 5613 2695
rect 5647 2661 5681 2695
rect 5715 2661 5782 2695
rect 5546 2614 5782 2661
rect 5546 2580 5613 2614
rect 5647 2580 5681 2614
rect 5715 2580 5782 2614
rect 5546 2546 5782 2580
rect 6538 2935 6774 2969
rect 6538 2901 6605 2935
rect 6639 2901 6673 2935
rect 6707 2901 6774 2935
rect 6538 2855 6774 2901
rect 6538 2821 6605 2855
rect 6639 2821 6673 2855
rect 6707 2821 6774 2855
rect 6538 2775 6774 2821
rect 6538 2741 6605 2775
rect 6639 2741 6673 2775
rect 6707 2741 6774 2775
rect 6538 2695 6774 2741
rect 6538 2661 6605 2695
rect 6639 2661 6673 2695
rect 6707 2661 6774 2695
rect 6538 2614 6774 2661
rect 6538 2580 6605 2614
rect 6639 2580 6673 2614
rect 6707 2580 6774 2614
rect 6538 2546 6774 2580
rect 7530 2935 7766 2969
rect 7530 2901 7597 2935
rect 7631 2901 7665 2935
rect 7699 2901 7766 2935
rect 7530 2855 7766 2901
rect 7530 2821 7597 2855
rect 7631 2821 7665 2855
rect 7699 2821 7766 2855
rect 7530 2775 7766 2821
rect 7530 2741 7597 2775
rect 7631 2741 7665 2775
rect 7699 2741 7766 2775
rect 7530 2695 7766 2741
rect 7530 2661 7597 2695
rect 7631 2661 7665 2695
rect 7699 2661 7766 2695
rect 7530 2614 7766 2661
rect 7530 2580 7597 2614
rect 7631 2580 7665 2614
rect 7699 2580 7766 2614
rect 7530 2546 7766 2580
rect 8522 2935 8758 2969
rect 8522 2901 8589 2935
rect 8623 2901 8657 2935
rect 8691 2901 8758 2935
rect 8522 2855 8758 2901
rect 8522 2821 8589 2855
rect 8623 2821 8657 2855
rect 8691 2821 8758 2855
rect 8522 2775 8758 2821
rect 8522 2741 8589 2775
rect 8623 2741 8657 2775
rect 8691 2741 8758 2775
rect 8522 2695 8758 2741
rect 8522 2661 8589 2695
rect 8623 2661 8657 2695
rect 8691 2661 8758 2695
rect 8522 2614 8758 2661
rect 8522 2580 8589 2614
rect 8623 2580 8657 2614
rect 8691 2580 8758 2614
rect 8522 2546 8758 2580
rect 9514 2935 9750 2969
rect 9514 2901 9581 2935
rect 9615 2901 9649 2935
rect 9683 2901 9750 2935
rect 9514 2855 9750 2901
rect 9514 2821 9581 2855
rect 9615 2821 9649 2855
rect 9683 2821 9750 2855
rect 9514 2775 9750 2821
rect 9514 2741 9581 2775
rect 9615 2741 9649 2775
rect 9683 2741 9750 2775
rect 9514 2695 9750 2741
rect 9514 2661 9581 2695
rect 9615 2661 9649 2695
rect 9683 2661 9750 2695
rect 9514 2614 9750 2661
rect 9514 2580 9581 2614
rect 9615 2580 9649 2614
rect 9683 2580 9750 2614
rect 9514 2546 9750 2580
rect 10506 2935 10742 2969
rect 10506 2901 10573 2935
rect 10607 2901 10641 2935
rect 10675 2901 10742 2935
rect 10506 2855 10742 2901
rect 10506 2821 10573 2855
rect 10607 2821 10641 2855
rect 10675 2821 10742 2855
rect 10506 2775 10742 2821
rect 10506 2741 10573 2775
rect 10607 2741 10641 2775
rect 10675 2741 10742 2775
rect 10506 2695 10742 2741
rect 10506 2661 10573 2695
rect 10607 2661 10641 2695
rect 10675 2661 10742 2695
rect 10506 2614 10742 2661
rect 10506 2580 10573 2614
rect 10607 2580 10641 2614
rect 10675 2580 10742 2614
rect 10506 2546 10742 2580
rect 11498 2935 11734 2969
rect 11498 2901 11565 2935
rect 11599 2901 11633 2935
rect 11667 2901 11734 2935
rect 11498 2855 11734 2901
rect 11498 2821 11565 2855
rect 11599 2821 11633 2855
rect 11667 2821 11734 2855
rect 11498 2775 11734 2821
rect 11498 2741 11565 2775
rect 11599 2741 11633 2775
rect 11667 2741 11734 2775
rect 11498 2695 11734 2741
rect 11498 2661 11565 2695
rect 11599 2661 11633 2695
rect 11667 2661 11734 2695
rect 11498 2614 11734 2661
rect 11498 2580 11565 2614
rect 11599 2580 11633 2614
rect 11667 2580 11734 2614
rect 11498 2546 11734 2580
rect 12490 2935 12726 2969
rect 12490 2901 12557 2935
rect 12591 2901 12625 2935
rect 12659 2901 12726 2935
rect 12490 2855 12726 2901
rect 12490 2821 12557 2855
rect 12591 2821 12625 2855
rect 12659 2821 12726 2855
rect 12490 2775 12726 2821
rect 12490 2741 12557 2775
rect 12591 2741 12625 2775
rect 12659 2741 12726 2775
rect 12490 2695 12726 2741
rect 12490 2661 12557 2695
rect 12591 2661 12625 2695
rect 12659 2661 12726 2695
rect 12490 2614 12726 2661
rect 12490 2580 12557 2614
rect 12591 2580 12625 2614
rect 12659 2580 12726 2614
rect 12490 2546 12726 2580
rect 13482 2935 13718 2969
rect 13482 2901 13549 2935
rect 13583 2901 13617 2935
rect 13651 2901 13718 2935
rect 13482 2855 13718 2901
rect 13482 2821 13549 2855
rect 13583 2821 13617 2855
rect 13651 2821 13718 2855
rect 13482 2775 13718 2821
rect 13482 2741 13549 2775
rect 13583 2741 13617 2775
rect 13651 2741 13718 2775
rect 13482 2695 13718 2741
rect 13482 2661 13549 2695
rect 13583 2661 13617 2695
rect 13651 2661 13718 2695
rect 13482 2614 13718 2661
rect 13482 2580 13549 2614
rect 13583 2580 13617 2614
rect 13651 2580 13718 2614
rect 13482 2546 13718 2580
rect 14497 3032 14565 3058
rect 14599 3032 14633 3066
rect 14497 2972 14667 3032
rect 14497 2485 14667 2530
rect 14497 2457 14565 2485
rect 657 2433 787 2457
rect 657 2399 734 2433
rect 768 2399 787 2433
rect 657 2367 787 2399
rect 555 2365 787 2367
rect 555 2331 734 2365
rect 768 2331 787 2365
rect 555 2327 787 2331
rect 589 2293 623 2327
rect 657 2297 787 2327
rect 657 2293 734 2297
rect 555 2263 734 2293
rect 768 2263 787 2297
rect 555 2250 787 2263
rect 589 2216 623 2250
rect 657 2229 787 2250
rect 657 2216 734 2229
rect 555 2195 734 2216
rect 768 2195 787 2229
rect 555 2161 787 2195
rect 555 2156 734 2161
rect 589 2122 623 2156
rect 657 2127 734 2156
rect 768 2127 787 2161
rect 657 2122 787 2127
rect 555 2093 787 2122
rect 555 2085 734 2093
rect 589 2051 623 2085
rect 657 2059 734 2085
rect 768 2059 787 2093
rect 657 2051 787 2059
rect 555 2025 787 2051
rect 555 2011 734 2025
rect 589 1977 623 2011
rect 657 1991 734 2011
rect 768 1991 787 2025
rect 657 1977 787 1991
rect 555 1957 787 1977
rect 555 1940 734 1957
rect 589 1906 623 1940
rect 657 1923 734 1940
rect 768 1923 787 1957
rect 657 1906 787 1923
rect 555 1889 787 1906
rect 555 1866 734 1889
rect 589 1832 623 1866
rect 657 1855 734 1866
rect 768 1855 787 1889
rect 657 1832 787 1855
rect 555 1821 787 1832
rect 555 1795 734 1821
rect 589 1761 623 1795
rect 657 1787 734 1795
rect 768 1787 787 1821
rect 657 1761 787 1787
rect 555 1753 787 1761
rect 555 1721 734 1753
rect 589 1687 623 1721
rect 657 1719 734 1721
rect 768 1719 787 1753
rect 657 1687 787 1719
rect 555 1685 787 1687
rect 555 1651 734 1685
rect 768 1651 787 1685
rect 555 1650 787 1651
rect 589 1616 623 1650
rect 657 1617 787 1650
rect 657 1616 734 1617
rect 555 1583 734 1616
rect 768 1583 787 1617
rect 555 1576 787 1583
rect 589 1542 623 1576
rect 657 1549 787 1576
rect 657 1542 734 1549
rect 555 1515 734 1542
rect 768 1515 787 1549
rect 555 1505 787 1515
rect 589 1471 623 1505
rect 657 1471 787 1505
rect 555 1457 787 1471
rect 1625 2445 1765 2457
rect 1625 2411 1678 2445
rect 1712 2411 1765 2445
rect 1625 2377 1765 2411
rect 1625 2343 1678 2377
rect 1712 2343 1765 2377
rect 1625 2309 1765 2343
rect 1625 2275 1678 2309
rect 1712 2275 1765 2309
rect 1625 2241 1765 2275
rect 1625 2207 1678 2241
rect 1712 2207 1765 2241
rect 1625 2173 1765 2207
rect 1625 2139 1678 2173
rect 1712 2139 1765 2173
rect 1625 2105 1765 2139
rect 1625 2071 1678 2105
rect 1712 2071 1765 2105
rect 1625 2037 1765 2071
rect 1625 2003 1678 2037
rect 1712 2003 1765 2037
rect 1625 1969 1765 2003
rect 1625 1935 1678 1969
rect 1712 1935 1765 1969
rect 1625 1901 1765 1935
rect 1625 1867 1678 1901
rect 1712 1867 1765 1901
rect 1625 1833 1765 1867
rect 1625 1799 1678 1833
rect 1712 1799 1765 1833
rect 1625 1765 1765 1799
rect 1625 1731 1678 1765
rect 1712 1731 1765 1765
rect 1625 1697 1765 1731
rect 1625 1663 1678 1697
rect 1712 1663 1765 1697
rect 1625 1629 1765 1663
rect 1625 1595 1678 1629
rect 1712 1595 1765 1629
rect 1625 1561 1765 1595
rect 1625 1527 1678 1561
rect 1712 1527 1765 1561
rect 1625 1457 1765 1527
rect 2617 2445 2757 2457
rect 2617 2411 2670 2445
rect 2704 2411 2757 2445
rect 2617 2377 2757 2411
rect 2617 2343 2670 2377
rect 2704 2343 2757 2377
rect 2617 2309 2757 2343
rect 2617 2275 2670 2309
rect 2704 2275 2757 2309
rect 2617 2241 2757 2275
rect 2617 2207 2670 2241
rect 2704 2207 2757 2241
rect 2617 2173 2757 2207
rect 2617 2139 2670 2173
rect 2704 2139 2757 2173
rect 2617 2105 2757 2139
rect 2617 2071 2670 2105
rect 2704 2071 2757 2105
rect 2617 2037 2757 2071
rect 2617 2003 2670 2037
rect 2704 2003 2757 2037
rect 2617 1969 2757 2003
rect 2617 1935 2670 1969
rect 2704 1935 2757 1969
rect 2617 1901 2757 1935
rect 2617 1867 2670 1901
rect 2704 1867 2757 1901
rect 2617 1833 2757 1867
rect 2617 1799 2670 1833
rect 2704 1799 2757 1833
rect 2617 1765 2757 1799
rect 2617 1731 2670 1765
rect 2704 1731 2757 1765
rect 2617 1697 2757 1731
rect 2617 1663 2670 1697
rect 2704 1663 2757 1697
rect 2617 1629 2757 1663
rect 2617 1595 2670 1629
rect 2704 1595 2757 1629
rect 2617 1561 2757 1595
rect 2617 1527 2670 1561
rect 2704 1527 2757 1561
rect 2617 1457 2757 1527
rect 3609 2445 3749 2457
rect 3609 2411 3662 2445
rect 3696 2411 3749 2445
rect 3609 2377 3749 2411
rect 3609 2343 3662 2377
rect 3696 2343 3749 2377
rect 3609 2309 3749 2343
rect 3609 2275 3662 2309
rect 3696 2275 3749 2309
rect 3609 2241 3749 2275
rect 3609 2207 3662 2241
rect 3696 2207 3749 2241
rect 3609 2173 3749 2207
rect 3609 2139 3662 2173
rect 3696 2139 3749 2173
rect 3609 2105 3749 2139
rect 3609 2071 3662 2105
rect 3696 2071 3749 2105
rect 3609 2037 3749 2071
rect 3609 2003 3662 2037
rect 3696 2003 3749 2037
rect 3609 1969 3749 2003
rect 3609 1935 3662 1969
rect 3696 1935 3749 1969
rect 3609 1901 3749 1935
rect 3609 1867 3662 1901
rect 3696 1867 3749 1901
rect 3609 1833 3749 1867
rect 3609 1799 3662 1833
rect 3696 1799 3749 1833
rect 3609 1765 3749 1799
rect 3609 1731 3662 1765
rect 3696 1731 3749 1765
rect 3609 1697 3749 1731
rect 3609 1663 3662 1697
rect 3696 1663 3749 1697
rect 3609 1629 3749 1663
rect 3609 1595 3662 1629
rect 3696 1595 3749 1629
rect 3609 1561 3749 1595
rect 3609 1527 3662 1561
rect 3696 1527 3749 1561
rect 3609 1457 3749 1527
rect 4601 2445 4741 2457
rect 4601 2411 4654 2445
rect 4688 2411 4741 2445
rect 4601 2377 4741 2411
rect 4601 2343 4654 2377
rect 4688 2343 4741 2377
rect 4601 2309 4741 2343
rect 4601 2275 4654 2309
rect 4688 2275 4741 2309
rect 4601 2241 4741 2275
rect 4601 2207 4654 2241
rect 4688 2207 4741 2241
rect 4601 2173 4741 2207
rect 4601 2139 4654 2173
rect 4688 2139 4741 2173
rect 4601 2105 4741 2139
rect 4601 2071 4654 2105
rect 4688 2071 4741 2105
rect 4601 2037 4741 2071
rect 4601 2003 4654 2037
rect 4688 2003 4741 2037
rect 4601 1969 4741 2003
rect 4601 1935 4654 1969
rect 4688 1935 4741 1969
rect 4601 1901 4741 1935
rect 4601 1867 4654 1901
rect 4688 1867 4741 1901
rect 4601 1833 4741 1867
rect 4601 1799 4654 1833
rect 4688 1799 4741 1833
rect 4601 1765 4741 1799
rect 4601 1731 4654 1765
rect 4688 1731 4741 1765
rect 4601 1697 4741 1731
rect 4601 1663 4654 1697
rect 4688 1663 4741 1697
rect 4601 1629 4741 1663
rect 4601 1595 4654 1629
rect 4688 1595 4741 1629
rect 4601 1561 4741 1595
rect 4601 1527 4654 1561
rect 4688 1527 4741 1561
rect 4601 1457 4741 1527
rect 5593 2445 5733 2457
rect 5593 2411 5646 2445
rect 5680 2411 5733 2445
rect 5593 2377 5733 2411
rect 5593 2343 5646 2377
rect 5680 2343 5733 2377
rect 5593 2309 5733 2343
rect 5593 2275 5646 2309
rect 5680 2275 5733 2309
rect 5593 2241 5733 2275
rect 5593 2207 5646 2241
rect 5680 2207 5733 2241
rect 5593 2173 5733 2207
rect 5593 2139 5646 2173
rect 5680 2139 5733 2173
rect 5593 2105 5733 2139
rect 5593 2071 5646 2105
rect 5680 2071 5733 2105
rect 5593 2037 5733 2071
rect 5593 2003 5646 2037
rect 5680 2003 5733 2037
rect 5593 1969 5733 2003
rect 5593 1935 5646 1969
rect 5680 1935 5733 1969
rect 5593 1901 5733 1935
rect 5593 1867 5646 1901
rect 5680 1867 5733 1901
rect 5593 1833 5733 1867
rect 5593 1799 5646 1833
rect 5680 1799 5733 1833
rect 5593 1765 5733 1799
rect 5593 1731 5646 1765
rect 5680 1731 5733 1765
rect 5593 1697 5733 1731
rect 5593 1663 5646 1697
rect 5680 1663 5733 1697
rect 5593 1629 5733 1663
rect 5593 1595 5646 1629
rect 5680 1595 5733 1629
rect 5593 1561 5733 1595
rect 5593 1527 5646 1561
rect 5680 1527 5733 1561
rect 5593 1457 5733 1527
rect 6585 2445 6725 2457
rect 6585 2411 6638 2445
rect 6672 2411 6725 2445
rect 6585 2377 6725 2411
rect 6585 2343 6638 2377
rect 6672 2343 6725 2377
rect 6585 2309 6725 2343
rect 6585 2275 6638 2309
rect 6672 2275 6725 2309
rect 6585 2241 6725 2275
rect 6585 2207 6638 2241
rect 6672 2207 6725 2241
rect 6585 2173 6725 2207
rect 6585 2139 6638 2173
rect 6672 2139 6725 2173
rect 6585 2105 6725 2139
rect 6585 2071 6638 2105
rect 6672 2071 6725 2105
rect 6585 2037 6725 2071
rect 6585 2003 6638 2037
rect 6672 2003 6725 2037
rect 6585 1969 6725 2003
rect 6585 1935 6638 1969
rect 6672 1935 6725 1969
rect 6585 1901 6725 1935
rect 6585 1867 6638 1901
rect 6672 1867 6725 1901
rect 6585 1833 6725 1867
rect 6585 1799 6638 1833
rect 6672 1799 6725 1833
rect 6585 1765 6725 1799
rect 6585 1731 6638 1765
rect 6672 1731 6725 1765
rect 6585 1697 6725 1731
rect 6585 1663 6638 1697
rect 6672 1663 6725 1697
rect 6585 1629 6725 1663
rect 6585 1595 6638 1629
rect 6672 1595 6725 1629
rect 6585 1561 6725 1595
rect 6585 1527 6638 1561
rect 6672 1527 6725 1561
rect 6585 1457 6725 1527
rect 7577 2445 7717 2457
rect 7577 2411 7630 2445
rect 7664 2411 7717 2445
rect 7577 2377 7717 2411
rect 7577 2343 7630 2377
rect 7664 2343 7717 2377
rect 7577 2309 7717 2343
rect 7577 2275 7630 2309
rect 7664 2275 7717 2309
rect 7577 2241 7717 2275
rect 7577 2207 7630 2241
rect 7664 2207 7717 2241
rect 7577 2173 7717 2207
rect 7577 2139 7630 2173
rect 7664 2139 7717 2173
rect 7577 2105 7717 2139
rect 7577 2071 7630 2105
rect 7664 2071 7717 2105
rect 7577 2037 7717 2071
rect 7577 2003 7630 2037
rect 7664 2003 7717 2037
rect 7577 1969 7717 2003
rect 7577 1935 7630 1969
rect 7664 1935 7717 1969
rect 7577 1901 7717 1935
rect 7577 1867 7630 1901
rect 7664 1867 7717 1901
rect 7577 1833 7717 1867
rect 7577 1799 7630 1833
rect 7664 1799 7717 1833
rect 7577 1765 7717 1799
rect 7577 1731 7630 1765
rect 7664 1731 7717 1765
rect 7577 1697 7717 1731
rect 7577 1663 7630 1697
rect 7664 1663 7717 1697
rect 7577 1629 7717 1663
rect 7577 1595 7630 1629
rect 7664 1595 7717 1629
rect 7577 1561 7717 1595
rect 7577 1527 7630 1561
rect 7664 1527 7717 1561
rect 7577 1457 7717 1527
rect 8569 2445 8709 2457
rect 8569 2411 8622 2445
rect 8656 2411 8709 2445
rect 8569 2377 8709 2411
rect 8569 2343 8622 2377
rect 8656 2343 8709 2377
rect 8569 2309 8709 2343
rect 8569 2275 8622 2309
rect 8656 2275 8709 2309
rect 8569 2241 8709 2275
rect 8569 2207 8622 2241
rect 8656 2207 8709 2241
rect 8569 2173 8709 2207
rect 8569 2139 8622 2173
rect 8656 2139 8709 2173
rect 8569 2105 8709 2139
rect 8569 2071 8622 2105
rect 8656 2071 8709 2105
rect 8569 2037 8709 2071
rect 8569 2003 8622 2037
rect 8656 2003 8709 2037
rect 8569 1969 8709 2003
rect 8569 1935 8622 1969
rect 8656 1935 8709 1969
rect 8569 1901 8709 1935
rect 8569 1867 8622 1901
rect 8656 1867 8709 1901
rect 8569 1833 8709 1867
rect 8569 1799 8622 1833
rect 8656 1799 8709 1833
rect 8569 1765 8709 1799
rect 8569 1731 8622 1765
rect 8656 1731 8709 1765
rect 8569 1697 8709 1731
rect 8569 1663 8622 1697
rect 8656 1663 8709 1697
rect 8569 1629 8709 1663
rect 8569 1595 8622 1629
rect 8656 1595 8709 1629
rect 8569 1561 8709 1595
rect 8569 1527 8622 1561
rect 8656 1527 8709 1561
rect 8569 1457 8709 1527
rect 9561 2445 9701 2457
rect 9561 2411 9614 2445
rect 9648 2411 9701 2445
rect 9561 2377 9701 2411
rect 9561 2343 9614 2377
rect 9648 2343 9701 2377
rect 9561 2309 9701 2343
rect 9561 2275 9614 2309
rect 9648 2275 9701 2309
rect 9561 2241 9701 2275
rect 9561 2207 9614 2241
rect 9648 2207 9701 2241
rect 9561 2173 9701 2207
rect 9561 2139 9614 2173
rect 9648 2139 9701 2173
rect 9561 2105 9701 2139
rect 9561 2071 9614 2105
rect 9648 2071 9701 2105
rect 9561 2037 9701 2071
rect 9561 2003 9614 2037
rect 9648 2003 9701 2037
rect 9561 1969 9701 2003
rect 9561 1935 9614 1969
rect 9648 1935 9701 1969
rect 9561 1901 9701 1935
rect 9561 1867 9614 1901
rect 9648 1867 9701 1901
rect 9561 1833 9701 1867
rect 9561 1799 9614 1833
rect 9648 1799 9701 1833
rect 9561 1765 9701 1799
rect 9561 1731 9614 1765
rect 9648 1731 9701 1765
rect 9561 1697 9701 1731
rect 9561 1663 9614 1697
rect 9648 1663 9701 1697
rect 9561 1629 9701 1663
rect 9561 1595 9614 1629
rect 9648 1595 9701 1629
rect 9561 1561 9701 1595
rect 9561 1527 9614 1561
rect 9648 1527 9701 1561
rect 9561 1457 9701 1527
rect 10553 2445 10693 2457
rect 10553 2411 10606 2445
rect 10640 2411 10693 2445
rect 10553 2377 10693 2411
rect 10553 2343 10606 2377
rect 10640 2343 10693 2377
rect 10553 2309 10693 2343
rect 10553 2275 10606 2309
rect 10640 2275 10693 2309
rect 10553 2241 10693 2275
rect 10553 2207 10606 2241
rect 10640 2207 10693 2241
rect 10553 2173 10693 2207
rect 10553 2139 10606 2173
rect 10640 2139 10693 2173
rect 10553 2105 10693 2139
rect 10553 2071 10606 2105
rect 10640 2071 10693 2105
rect 10553 2037 10693 2071
rect 10553 2003 10606 2037
rect 10640 2003 10693 2037
rect 10553 1969 10693 2003
rect 10553 1935 10606 1969
rect 10640 1935 10693 1969
rect 10553 1901 10693 1935
rect 10553 1867 10606 1901
rect 10640 1867 10693 1901
rect 10553 1833 10693 1867
rect 10553 1799 10606 1833
rect 10640 1799 10693 1833
rect 10553 1765 10693 1799
rect 10553 1731 10606 1765
rect 10640 1731 10693 1765
rect 10553 1697 10693 1731
rect 10553 1663 10606 1697
rect 10640 1663 10693 1697
rect 10553 1629 10693 1663
rect 10553 1595 10606 1629
rect 10640 1595 10693 1629
rect 10553 1561 10693 1595
rect 10553 1527 10606 1561
rect 10640 1527 10693 1561
rect 10553 1457 10693 1527
rect 11545 2445 11685 2457
rect 11545 2411 11598 2445
rect 11632 2411 11685 2445
rect 11545 2377 11685 2411
rect 11545 2343 11598 2377
rect 11632 2343 11685 2377
rect 11545 2309 11685 2343
rect 11545 2275 11598 2309
rect 11632 2275 11685 2309
rect 11545 2241 11685 2275
rect 11545 2207 11598 2241
rect 11632 2207 11685 2241
rect 11545 2173 11685 2207
rect 11545 2139 11598 2173
rect 11632 2139 11685 2173
rect 11545 2105 11685 2139
rect 11545 2071 11598 2105
rect 11632 2071 11685 2105
rect 11545 2037 11685 2071
rect 11545 2003 11598 2037
rect 11632 2003 11685 2037
rect 11545 1969 11685 2003
rect 11545 1935 11598 1969
rect 11632 1935 11685 1969
rect 11545 1901 11685 1935
rect 11545 1867 11598 1901
rect 11632 1867 11685 1901
rect 11545 1833 11685 1867
rect 11545 1799 11598 1833
rect 11632 1799 11685 1833
rect 11545 1765 11685 1799
rect 11545 1731 11598 1765
rect 11632 1731 11685 1765
rect 11545 1697 11685 1731
rect 11545 1663 11598 1697
rect 11632 1663 11685 1697
rect 11545 1629 11685 1663
rect 11545 1595 11598 1629
rect 11632 1595 11685 1629
rect 11545 1561 11685 1595
rect 11545 1527 11598 1561
rect 11632 1527 11685 1561
rect 11545 1457 11685 1527
rect 12537 2445 12677 2457
rect 12537 2411 12590 2445
rect 12624 2411 12677 2445
rect 12537 2377 12677 2411
rect 12537 2343 12590 2377
rect 12624 2343 12677 2377
rect 12537 2309 12677 2343
rect 12537 2275 12590 2309
rect 12624 2275 12677 2309
rect 12537 2241 12677 2275
rect 12537 2207 12590 2241
rect 12624 2207 12677 2241
rect 12537 2173 12677 2207
rect 12537 2139 12590 2173
rect 12624 2139 12677 2173
rect 12537 2105 12677 2139
rect 12537 2071 12590 2105
rect 12624 2071 12677 2105
rect 12537 2037 12677 2071
rect 12537 2003 12590 2037
rect 12624 2003 12677 2037
rect 12537 1969 12677 2003
rect 12537 1935 12590 1969
rect 12624 1935 12677 1969
rect 12537 1901 12677 1935
rect 12537 1867 12590 1901
rect 12624 1867 12677 1901
rect 12537 1833 12677 1867
rect 12537 1799 12590 1833
rect 12624 1799 12677 1833
rect 12537 1765 12677 1799
rect 12537 1731 12590 1765
rect 12624 1731 12677 1765
rect 12537 1697 12677 1731
rect 12537 1663 12590 1697
rect 12624 1663 12677 1697
rect 12537 1629 12677 1663
rect 12537 1595 12590 1629
rect 12624 1595 12677 1629
rect 12537 1561 12677 1595
rect 12537 1527 12590 1561
rect 12624 1527 12677 1561
rect 12537 1457 12677 1527
rect 13529 2445 13669 2457
rect 13529 2411 13582 2445
rect 13616 2411 13669 2445
rect 13529 2377 13669 2411
rect 13529 2343 13582 2377
rect 13616 2343 13669 2377
rect 13529 2309 13669 2343
rect 13529 2275 13582 2309
rect 13616 2275 13669 2309
rect 13529 2241 13669 2275
rect 13529 2207 13582 2241
rect 13616 2207 13669 2241
rect 13529 2173 13669 2207
rect 13529 2139 13582 2173
rect 13616 2139 13669 2173
rect 13529 2105 13669 2139
rect 13529 2071 13582 2105
rect 13616 2071 13669 2105
rect 13529 2037 13669 2071
rect 13529 2003 13582 2037
rect 13616 2003 13669 2037
rect 13529 1969 13669 2003
rect 13529 1935 13582 1969
rect 13616 1935 13669 1969
rect 13529 1901 13669 1935
rect 13529 1867 13582 1901
rect 13616 1867 13669 1901
rect 13529 1833 13669 1867
rect 13529 1799 13582 1833
rect 13616 1799 13669 1833
rect 13529 1765 13669 1799
rect 13529 1731 13582 1765
rect 13616 1731 13669 1765
rect 13529 1697 13669 1731
rect 13529 1663 13582 1697
rect 13616 1663 13669 1697
rect 13529 1629 13669 1663
rect 13529 1595 13582 1629
rect 13616 1595 13669 1629
rect 13529 1561 13669 1595
rect 13529 1527 13582 1561
rect 13616 1527 13669 1561
rect 13529 1457 13669 1527
rect 14435 2451 14565 2457
rect 14599 2451 14633 2485
rect 14435 2433 14667 2451
rect 14435 2399 14454 2433
rect 14488 2403 14667 2433
rect 14488 2399 14565 2403
rect 14435 2369 14565 2399
rect 14599 2369 14633 2403
rect 14435 2365 14667 2369
rect 14435 2331 14454 2365
rect 14488 2331 14667 2365
rect 14435 2327 14667 2331
rect 14435 2297 14565 2327
rect 14435 2263 14454 2297
rect 14488 2293 14565 2297
rect 14599 2293 14633 2327
rect 14488 2263 14667 2293
rect 14435 2250 14667 2263
rect 14435 2229 14565 2250
rect 14435 2195 14454 2229
rect 14488 2216 14565 2229
rect 14599 2216 14633 2250
rect 14488 2195 14667 2216
rect 14435 2161 14667 2195
rect 14435 2127 14454 2161
rect 14488 2156 14667 2161
rect 14488 2127 14565 2156
rect 14435 2122 14565 2127
rect 14599 2122 14633 2156
rect 14435 2093 14667 2122
rect 14435 2059 14454 2093
rect 14488 2085 14667 2093
rect 14488 2059 14565 2085
rect 14435 2051 14565 2059
rect 14599 2051 14633 2085
rect 14435 2025 14667 2051
rect 14435 1991 14454 2025
rect 14488 2011 14667 2025
rect 14488 1991 14565 2011
rect 14435 1977 14565 1991
rect 14599 1977 14633 2011
rect 14435 1957 14667 1977
rect 14435 1923 14454 1957
rect 14488 1940 14667 1957
rect 14488 1923 14565 1940
rect 14435 1906 14565 1923
rect 14599 1906 14633 1940
rect 14435 1889 14667 1906
rect 14435 1855 14454 1889
rect 14488 1866 14667 1889
rect 14488 1855 14565 1866
rect 14435 1832 14565 1855
rect 14599 1832 14633 1866
rect 14435 1821 14667 1832
rect 14435 1787 14454 1821
rect 14488 1795 14667 1821
rect 14488 1787 14565 1795
rect 14435 1761 14565 1787
rect 14599 1761 14633 1795
rect 14435 1753 14667 1761
rect 14435 1719 14454 1753
rect 14488 1721 14667 1753
rect 14488 1719 14565 1721
rect 14435 1687 14565 1719
rect 14599 1687 14633 1721
rect 14435 1685 14667 1687
rect 14435 1651 14454 1685
rect 14488 1651 14667 1685
rect 14435 1650 14667 1651
rect 14435 1617 14565 1650
rect 14435 1583 14454 1617
rect 14488 1616 14565 1617
rect 14599 1616 14633 1650
rect 14488 1583 14667 1616
rect 14435 1576 14667 1583
rect 14435 1549 14565 1576
rect 14435 1515 14454 1549
rect 14488 1542 14565 1549
rect 14599 1542 14633 1576
rect 14488 1515 14667 1542
rect 14435 1505 14667 1515
rect 14435 1471 14565 1505
rect 14599 1471 14633 1505
rect 14435 1457 14667 1471
rect 555 1375 725 1457
rect 589 1341 623 1375
rect 657 1341 691 1375
rect 555 1221 725 1341
rect 14497 1387 14667 1457
rect 14531 1353 14565 1387
rect 14599 1353 14633 1387
rect 14497 1319 14667 1353
rect 14497 1311 14633 1319
rect 14497 1308 14565 1311
rect 589 1187 623 1221
rect 657 1219 725 1221
rect 657 1187 691 1219
rect 555 1185 691 1187
rect 555 1150 725 1185
rect 555 1140 623 1150
rect 589 1116 623 1140
rect 657 1148 725 1150
rect 14531 1277 14565 1308
rect 14599 1285 14633 1311
rect 14599 1277 14667 1285
rect 14531 1274 14667 1277
rect 14497 1251 14667 1274
rect 14497 1234 14633 1251
rect 14497 1228 14565 1234
rect 14531 1200 14565 1228
rect 14599 1217 14633 1234
rect 14599 1200 14667 1217
rect 14531 1194 14667 1200
rect 14497 1183 14667 1194
rect 14497 1157 14633 1183
rect 14497 1148 14565 1157
rect 657 1116 691 1148
rect 589 1114 691 1116
rect 725 1114 760 1148
rect 794 1114 829 1148
rect 589 1106 829 1114
rect 555 1080 829 1106
rect 14531 1123 14565 1148
rect 14599 1149 14633 1157
rect 14599 1123 14667 1149
rect 14531 1115 14667 1123
rect 14531 1081 14633 1115
rect 14531 1080 14667 1081
rect 555 1046 623 1080
rect 657 1046 692 1080
rect 726 1046 761 1080
rect 14599 1046 14667 1080
rect 555 1012 761 1046
rect 14565 1012 14633 1046
rect 555 978 589 1012
rect 623 978 658 1012
rect 692 978 727 1012
rect 14565 978 14667 1012
<< mvnsubdiff >>
rect 232 5388 300 5422
rect 334 5388 369 5422
rect 403 5388 438 5422
rect 472 5388 507 5422
rect 541 5388 576 5422
rect 610 5388 645 5422
rect 679 5388 714 5422
rect 748 5388 783 5422
rect 817 5388 852 5422
rect 886 5388 921 5422
rect 955 5388 990 5422
rect 1024 5388 1059 5422
rect 1093 5388 1128 5422
rect 1162 5388 1197 5422
rect 1231 5388 1266 5422
rect 1300 5388 1335 5422
rect 1369 5388 1404 5422
rect 1438 5388 1473 5422
rect 1507 5388 1542 5422
rect 1576 5388 1611 5422
rect 1645 5388 1680 5422
rect 1714 5388 1749 5422
rect 1783 5388 1818 5422
rect 1852 5388 1887 5422
rect 1921 5388 1956 5422
rect 1990 5388 2025 5422
rect 2059 5388 2094 5422
rect 2128 5388 2163 5422
rect 2197 5388 2232 5422
rect 232 5354 2232 5388
rect 334 5320 369 5354
rect 403 5320 438 5354
rect 472 5320 507 5354
rect 541 5320 576 5354
rect 610 5320 645 5354
rect 679 5320 714 5354
rect 748 5320 783 5354
rect 817 5320 852 5354
rect 886 5320 921 5354
rect 955 5320 990 5354
rect 1024 5320 1059 5354
rect 1093 5320 1128 5354
rect 1162 5320 1197 5354
rect 1231 5320 1266 5354
rect 1300 5320 1335 5354
rect 1369 5320 1404 5354
rect 1438 5320 1473 5354
rect 1507 5320 1542 5354
rect 1576 5320 1611 5354
rect 1645 5320 1680 5354
rect 1714 5320 1749 5354
rect 1783 5320 1818 5354
rect 1852 5320 1887 5354
rect 1921 5320 1956 5354
rect 1990 5320 2025 5354
rect 2059 5320 2094 5354
rect 2128 5320 2163 5354
rect 2197 5320 2232 5354
rect 334 5286 2300 5320
rect 402 5252 437 5286
rect 471 5252 506 5286
rect 540 5252 575 5286
rect 609 5252 644 5286
rect 678 5252 713 5286
rect 747 5252 782 5286
rect 816 5252 851 5286
rect 885 5252 920 5286
rect 954 5252 989 5286
rect 1023 5252 1058 5286
rect 1092 5252 1127 5286
rect 1161 5252 1196 5286
rect 1230 5252 1265 5286
rect 1299 5252 1334 5286
rect 1368 5252 1403 5286
rect 1437 5252 1472 5286
rect 1506 5252 1541 5286
rect 1575 5252 1610 5286
rect 1644 5252 1679 5286
rect 1713 5252 1748 5286
rect 1782 5252 1817 5286
rect 1851 5252 1886 5286
rect 1920 5252 1955 5286
rect 1989 5252 2024 5286
rect 2058 5252 2093 5286
rect 2127 5252 2162 5286
rect 2196 5252 2231 5286
rect 2265 5252 2300 5286
rect 14914 5218 14990 5422
rect 334 729 402 764
rect 334 696 368 729
rect 232 695 368 696
rect 232 661 402 695
rect 266 627 300 661
rect 334 660 402 661
rect 14820 660 14990 696
rect 334 627 368 660
rect 232 592 368 627
rect 12982 626 13017 660
rect 13051 626 13086 660
rect 13120 626 13155 660
rect 13189 626 13224 660
rect 13258 626 13293 660
rect 13327 626 13362 660
rect 13396 626 13431 660
rect 13465 626 13500 660
rect 13534 626 13569 660
rect 13603 626 13638 660
rect 13672 626 13707 660
rect 13741 626 13776 660
rect 13810 626 13845 660
rect 13879 626 13914 660
rect 13948 626 13983 660
rect 14017 626 14052 660
rect 14086 626 14121 660
rect 14155 626 14190 660
rect 14224 626 14259 660
rect 14293 626 14328 660
rect 14362 626 14397 660
rect 14431 626 14466 660
rect 14500 626 14535 660
rect 14569 626 14604 660
rect 14638 626 14673 660
rect 14707 626 14742 660
rect 14776 626 14811 660
rect 14845 626 14880 660
rect 14914 626 14990 660
rect 12982 592 14990 626
rect 266 558 300 592
rect 232 490 300 558
rect 12982 558 13017 592
rect 13051 558 13086 592
rect 13120 558 13155 592
rect 13189 558 13224 592
rect 13258 558 13293 592
rect 13327 558 13362 592
rect 13396 558 13431 592
rect 13465 558 13500 592
rect 13534 558 13569 592
rect 13603 558 13638 592
rect 13672 558 13707 592
rect 13741 558 13776 592
rect 13810 558 13845 592
rect 13879 558 13914 592
rect 13948 558 13983 592
rect 14017 558 14052 592
rect 14086 558 14121 592
rect 14155 558 14190 592
rect 14224 558 14259 592
rect 14293 558 14328 592
rect 14362 558 14397 592
rect 14431 558 14466 592
rect 14500 558 14535 592
rect 14569 558 14604 592
rect 14638 558 14673 592
rect 14707 558 14742 592
rect 14776 558 14811 592
rect 14845 558 14880 592
rect 14914 579 14990 592
rect 14914 558 14948 579
rect 12982 524 14948 558
rect 12982 490 13017 524
rect 13051 490 13086 524
rect 13120 490 13155 524
rect 13189 490 13224 524
rect 13258 490 13293 524
rect 13327 490 13362 524
rect 13396 490 13431 524
rect 13465 490 13500 524
rect 13534 490 13569 524
rect 13603 490 13638 524
rect 13672 490 13707 524
rect 13741 490 13776 524
rect 13810 490 13845 524
rect 13879 490 13914 524
rect 13948 490 13983 524
rect 14017 490 14052 524
rect 14086 490 14121 524
rect 14155 490 14190 524
rect 14224 490 14259 524
rect 14293 490 14328 524
rect 14362 490 14397 524
rect 14431 490 14466 524
rect 14500 490 14535 524
rect 14569 490 14604 524
rect 14638 490 14673 524
rect 14707 490 14742 524
rect 14776 490 14811 524
rect 14845 490 14880 524
rect 14914 490 14948 524
<< mvpsubdiffcont >>
rect 657 4922 14495 4956
rect 14530 4922 14564 4956
rect 14599 4922 14633 4956
rect 555 4888 589 4922
rect 657 4888 14461 4922
rect 623 4854 14461 4888
rect 14496 4854 14530 4888
rect 14565 4854 14599 4888
rect 555 4816 589 4850
rect 623 4785 657 4819
rect 691 4786 14393 4854
rect 14428 4786 14462 4820
rect 14497 4786 14531 4820
rect 555 4744 589 4778
rect 623 4716 657 4750
rect 691 4717 725 4751
rect 555 4672 589 4706
rect 623 4647 657 4681
rect 691 4648 725 4682
rect 555 4600 589 4634
rect 555 4529 589 4563
rect 555 4458 589 4492
rect 555 4387 589 4421
rect 555 4316 589 4350
rect 555 4245 589 4279
rect 555 4174 589 4208
rect 555 4103 589 4137
rect 623 4103 725 4613
rect 14565 4784 14599 4818
rect 14633 4810 14667 4844
rect 14497 4716 14531 4750
rect 14565 4714 14599 4748
rect 14633 4737 14667 4771
rect 14497 4646 14531 4680
rect 14565 4644 14599 4678
rect 14633 4664 14667 4698
rect 14497 4576 14531 4610
rect 14565 4574 14599 4608
rect 14633 4591 14667 4625
rect 14497 4506 14531 4540
rect 14565 4504 14599 4538
rect 14633 4518 14667 4552
rect 14497 4436 14531 4470
rect 14565 4434 14599 4468
rect 14633 4445 14667 4479
rect 14497 4365 14531 4399
rect 14565 4364 14599 4398
rect 14633 4372 14667 4406
rect 14497 4294 14531 4328
rect 14565 4294 14599 4328
rect 14633 4299 14667 4333
rect 14497 4223 14531 4257
rect 14565 4223 14599 4257
rect 14633 4226 14667 4260
rect 14497 4152 14531 4186
rect 14565 4152 14599 4186
rect 14633 4152 14667 4186
rect 14565 4081 14599 4115
rect 14633 4081 14667 4115
rect 555 4007 589 4041
rect 623 4007 657 4041
rect 734 4000 768 4034
rect 555 3936 589 3970
rect 623 3936 657 3970
rect 734 3932 768 3966
rect 555 3862 589 3896
rect 623 3862 657 3896
rect 734 3864 768 3898
rect 555 3791 589 3825
rect 623 3791 657 3825
rect 734 3796 768 3830
rect 555 3717 589 3751
rect 623 3717 657 3751
rect 734 3728 768 3762
rect 555 3646 589 3680
rect 623 3646 657 3680
rect 734 3660 768 3694
rect 555 3572 589 3606
rect 623 3572 657 3606
rect 734 3592 768 3626
rect 555 3501 589 3535
rect 623 3501 657 3535
rect 734 3524 768 3558
rect 555 3427 589 3461
rect 623 3427 657 3461
rect 734 3456 768 3490
rect 555 3356 589 3390
rect 623 3356 657 3390
rect 734 3388 768 3422
rect 734 3320 768 3354
rect 555 3282 589 3316
rect 623 3282 657 3316
rect 734 3252 768 3286
rect 555 3211 589 3245
rect 623 3211 657 3245
rect 734 3184 768 3218
rect 555 3117 589 3151
rect 623 3117 657 3151
rect 734 3116 768 3150
rect 555 3013 657 3081
rect 1678 4012 1712 4046
rect 1678 3944 1712 3978
rect 1678 3876 1712 3910
rect 1678 3808 1712 3842
rect 1678 3740 1712 3774
rect 1678 3672 1712 3706
rect 1678 3604 1712 3638
rect 1678 3536 1712 3570
rect 1678 3468 1712 3502
rect 1678 3400 1712 3434
rect 1678 3332 1712 3366
rect 1678 3264 1712 3298
rect 1678 3196 1712 3230
rect 1678 3128 1712 3162
rect 2670 4012 2704 4046
rect 2670 3944 2704 3978
rect 2670 3876 2704 3910
rect 2670 3808 2704 3842
rect 2670 3740 2704 3774
rect 2670 3672 2704 3706
rect 2670 3604 2704 3638
rect 2670 3536 2704 3570
rect 2670 3468 2704 3502
rect 2670 3400 2704 3434
rect 2670 3332 2704 3366
rect 2670 3264 2704 3298
rect 2670 3196 2704 3230
rect 2670 3128 2704 3162
rect 3662 4012 3696 4046
rect 3662 3944 3696 3978
rect 3662 3876 3696 3910
rect 3662 3808 3696 3842
rect 3662 3740 3696 3774
rect 3662 3672 3696 3706
rect 3662 3604 3696 3638
rect 3662 3536 3696 3570
rect 3662 3468 3696 3502
rect 3662 3400 3696 3434
rect 3662 3332 3696 3366
rect 3662 3264 3696 3298
rect 3662 3196 3696 3230
rect 3662 3128 3696 3162
rect 4654 4012 4688 4046
rect 4654 3944 4688 3978
rect 4654 3876 4688 3910
rect 4654 3808 4688 3842
rect 4654 3740 4688 3774
rect 4654 3672 4688 3706
rect 4654 3604 4688 3638
rect 4654 3536 4688 3570
rect 4654 3468 4688 3502
rect 4654 3400 4688 3434
rect 4654 3332 4688 3366
rect 4654 3264 4688 3298
rect 4654 3196 4688 3230
rect 4654 3128 4688 3162
rect 5646 4012 5680 4046
rect 5646 3944 5680 3978
rect 5646 3876 5680 3910
rect 5646 3808 5680 3842
rect 5646 3740 5680 3774
rect 5646 3672 5680 3706
rect 5646 3604 5680 3638
rect 5646 3536 5680 3570
rect 5646 3468 5680 3502
rect 5646 3400 5680 3434
rect 5646 3332 5680 3366
rect 5646 3264 5680 3298
rect 5646 3196 5680 3230
rect 5646 3128 5680 3162
rect 6638 4012 6672 4046
rect 6638 3944 6672 3978
rect 6638 3876 6672 3910
rect 6638 3808 6672 3842
rect 6638 3740 6672 3774
rect 6638 3672 6672 3706
rect 6638 3604 6672 3638
rect 6638 3536 6672 3570
rect 6638 3468 6672 3502
rect 6638 3400 6672 3434
rect 6638 3332 6672 3366
rect 6638 3264 6672 3298
rect 6638 3196 6672 3230
rect 6638 3128 6672 3162
rect 7630 4012 7664 4046
rect 7630 3944 7664 3978
rect 7630 3876 7664 3910
rect 7630 3808 7664 3842
rect 7630 3740 7664 3774
rect 7630 3672 7664 3706
rect 7630 3604 7664 3638
rect 7630 3536 7664 3570
rect 7630 3468 7664 3502
rect 7630 3400 7664 3434
rect 7630 3332 7664 3366
rect 7630 3264 7664 3298
rect 7630 3196 7664 3230
rect 7630 3128 7664 3162
rect 8622 4012 8656 4046
rect 8622 3944 8656 3978
rect 8622 3876 8656 3910
rect 8622 3808 8656 3842
rect 8622 3740 8656 3774
rect 8622 3672 8656 3706
rect 8622 3604 8656 3638
rect 8622 3536 8656 3570
rect 8622 3468 8656 3502
rect 8622 3400 8656 3434
rect 8622 3332 8656 3366
rect 8622 3264 8656 3298
rect 8622 3196 8656 3230
rect 8622 3128 8656 3162
rect 9614 4012 9648 4046
rect 9614 3944 9648 3978
rect 9614 3876 9648 3910
rect 9614 3808 9648 3842
rect 9614 3740 9648 3774
rect 9614 3672 9648 3706
rect 9614 3604 9648 3638
rect 9614 3536 9648 3570
rect 9614 3468 9648 3502
rect 9614 3400 9648 3434
rect 9614 3332 9648 3366
rect 9614 3264 9648 3298
rect 9614 3196 9648 3230
rect 9614 3128 9648 3162
rect 10606 4012 10640 4046
rect 10606 3944 10640 3978
rect 10606 3876 10640 3910
rect 10606 3808 10640 3842
rect 10606 3740 10640 3774
rect 10606 3672 10640 3706
rect 10606 3604 10640 3638
rect 10606 3536 10640 3570
rect 10606 3468 10640 3502
rect 10606 3400 10640 3434
rect 10606 3332 10640 3366
rect 10606 3264 10640 3298
rect 10606 3196 10640 3230
rect 10606 3128 10640 3162
rect 11598 4012 11632 4046
rect 11598 3944 11632 3978
rect 11598 3876 11632 3910
rect 11598 3808 11632 3842
rect 11598 3740 11632 3774
rect 11598 3672 11632 3706
rect 11598 3604 11632 3638
rect 11598 3536 11632 3570
rect 11598 3468 11632 3502
rect 11598 3400 11632 3434
rect 11598 3332 11632 3366
rect 11598 3264 11632 3298
rect 11598 3196 11632 3230
rect 11598 3128 11632 3162
rect 12590 4012 12624 4046
rect 12590 3944 12624 3978
rect 12590 3876 12624 3910
rect 12590 3808 12624 3842
rect 12590 3740 12624 3774
rect 12590 3672 12624 3706
rect 12590 3604 12624 3638
rect 12590 3536 12624 3570
rect 12590 3468 12624 3502
rect 12590 3400 12624 3434
rect 12590 3332 12624 3366
rect 12590 3264 12624 3298
rect 12590 3196 12624 3230
rect 12590 3128 12624 3162
rect 13582 4012 13616 4046
rect 13582 3944 13616 3978
rect 13582 3876 13616 3910
rect 13582 3808 13616 3842
rect 13582 3740 13616 3774
rect 13582 3672 13616 3706
rect 13582 3604 13616 3638
rect 13582 3536 13616 3570
rect 13582 3468 13616 3502
rect 13582 3400 13616 3434
rect 13582 3332 13616 3366
rect 13582 3264 13616 3298
rect 13582 3196 13616 3230
rect 13582 3128 13616 3162
rect 14454 4000 14488 4034
rect 14565 4007 14599 4041
rect 14633 4007 14667 4041
rect 14454 3932 14488 3966
rect 14565 3936 14599 3970
rect 14633 3936 14667 3970
rect 14454 3864 14488 3898
rect 14565 3862 14599 3896
rect 14633 3862 14667 3896
rect 14454 3796 14488 3830
rect 14565 3791 14599 3825
rect 14633 3791 14667 3825
rect 14454 3728 14488 3762
rect 14565 3717 14599 3751
rect 14633 3717 14667 3751
rect 14454 3660 14488 3694
rect 14565 3646 14599 3680
rect 14633 3646 14667 3680
rect 14454 3592 14488 3626
rect 14565 3572 14599 3606
rect 14633 3572 14667 3606
rect 14454 3524 14488 3558
rect 14565 3501 14599 3535
rect 14633 3501 14667 3535
rect 14454 3456 14488 3490
rect 14565 3427 14599 3461
rect 14633 3427 14667 3461
rect 14454 3388 14488 3422
rect 14565 3356 14599 3390
rect 14633 3356 14667 3390
rect 14454 3320 14488 3354
rect 14454 3252 14488 3286
rect 14565 3282 14599 3316
rect 14633 3282 14667 3316
rect 14454 3184 14488 3218
rect 14565 3211 14599 3245
rect 14633 3211 14667 3245
rect 14454 3116 14488 3150
rect 14565 3117 14599 3151
rect 14633 3117 14667 3151
rect 555 2503 725 3013
rect 555 2367 657 2503
rect 1645 2901 1679 2935
rect 1713 2901 1747 2935
rect 1645 2821 1679 2855
rect 1713 2821 1747 2855
rect 1645 2741 1679 2775
rect 1713 2741 1747 2775
rect 1645 2661 1679 2695
rect 1713 2661 1747 2695
rect 1645 2580 1679 2614
rect 1713 2580 1747 2614
rect 2637 2901 2671 2935
rect 2705 2901 2739 2935
rect 2637 2821 2671 2855
rect 2705 2821 2739 2855
rect 2637 2741 2671 2775
rect 2705 2741 2739 2775
rect 2637 2661 2671 2695
rect 2705 2661 2739 2695
rect 2637 2580 2671 2614
rect 2705 2580 2739 2614
rect 3629 2901 3663 2935
rect 3697 2901 3731 2935
rect 3629 2821 3663 2855
rect 3697 2821 3731 2855
rect 3629 2741 3663 2775
rect 3697 2741 3731 2775
rect 3629 2661 3663 2695
rect 3697 2661 3731 2695
rect 3629 2580 3663 2614
rect 3697 2580 3731 2614
rect 4621 2901 4655 2935
rect 4689 2901 4723 2935
rect 4621 2821 4655 2855
rect 4689 2821 4723 2855
rect 4621 2741 4655 2775
rect 4689 2741 4723 2775
rect 4621 2661 4655 2695
rect 4689 2661 4723 2695
rect 4621 2580 4655 2614
rect 4689 2580 4723 2614
rect 5613 2901 5647 2935
rect 5681 2901 5715 2935
rect 5613 2821 5647 2855
rect 5681 2821 5715 2855
rect 5613 2741 5647 2775
rect 5681 2741 5715 2775
rect 5613 2661 5647 2695
rect 5681 2661 5715 2695
rect 5613 2580 5647 2614
rect 5681 2580 5715 2614
rect 6605 2901 6639 2935
rect 6673 2901 6707 2935
rect 6605 2821 6639 2855
rect 6673 2821 6707 2855
rect 6605 2741 6639 2775
rect 6673 2741 6707 2775
rect 6605 2661 6639 2695
rect 6673 2661 6707 2695
rect 6605 2580 6639 2614
rect 6673 2580 6707 2614
rect 7597 2901 7631 2935
rect 7665 2901 7699 2935
rect 7597 2821 7631 2855
rect 7665 2821 7699 2855
rect 7597 2741 7631 2775
rect 7665 2741 7699 2775
rect 7597 2661 7631 2695
rect 7665 2661 7699 2695
rect 7597 2580 7631 2614
rect 7665 2580 7699 2614
rect 8589 2901 8623 2935
rect 8657 2901 8691 2935
rect 8589 2821 8623 2855
rect 8657 2821 8691 2855
rect 8589 2741 8623 2775
rect 8657 2741 8691 2775
rect 8589 2661 8623 2695
rect 8657 2661 8691 2695
rect 8589 2580 8623 2614
rect 8657 2580 8691 2614
rect 9581 2901 9615 2935
rect 9649 2901 9683 2935
rect 9581 2821 9615 2855
rect 9649 2821 9683 2855
rect 9581 2741 9615 2775
rect 9649 2741 9683 2775
rect 9581 2661 9615 2695
rect 9649 2661 9683 2695
rect 9581 2580 9615 2614
rect 9649 2580 9683 2614
rect 10573 2901 10607 2935
rect 10641 2901 10675 2935
rect 10573 2821 10607 2855
rect 10641 2821 10675 2855
rect 10573 2741 10607 2775
rect 10641 2741 10675 2775
rect 10573 2661 10607 2695
rect 10641 2661 10675 2695
rect 10573 2580 10607 2614
rect 10641 2580 10675 2614
rect 11565 2901 11599 2935
rect 11633 2901 11667 2935
rect 11565 2821 11599 2855
rect 11633 2821 11667 2855
rect 11565 2741 11599 2775
rect 11633 2741 11667 2775
rect 11565 2661 11599 2695
rect 11633 2661 11667 2695
rect 11565 2580 11599 2614
rect 11633 2580 11667 2614
rect 12557 2901 12591 2935
rect 12625 2901 12659 2935
rect 12557 2821 12591 2855
rect 12625 2821 12659 2855
rect 12557 2741 12591 2775
rect 12625 2741 12659 2775
rect 12557 2661 12591 2695
rect 12625 2661 12659 2695
rect 12557 2580 12591 2614
rect 12625 2580 12659 2614
rect 13549 2901 13583 2935
rect 13617 2901 13651 2935
rect 13549 2821 13583 2855
rect 13617 2821 13651 2855
rect 13549 2741 13583 2775
rect 13617 2741 13651 2775
rect 13549 2661 13583 2695
rect 13617 2661 13651 2695
rect 13549 2580 13583 2614
rect 13617 2580 13651 2614
rect 14565 3032 14599 3066
rect 14633 3032 14667 3066
rect 14497 2530 14667 2972
rect 734 2399 768 2433
rect 734 2331 768 2365
rect 555 2293 589 2327
rect 623 2293 657 2327
rect 734 2263 768 2297
rect 555 2216 589 2250
rect 623 2216 657 2250
rect 734 2195 768 2229
rect 555 2122 589 2156
rect 623 2122 657 2156
rect 734 2127 768 2161
rect 555 2051 589 2085
rect 623 2051 657 2085
rect 734 2059 768 2093
rect 555 1977 589 2011
rect 623 1977 657 2011
rect 734 1991 768 2025
rect 555 1906 589 1940
rect 623 1906 657 1940
rect 734 1923 768 1957
rect 555 1832 589 1866
rect 623 1832 657 1866
rect 734 1855 768 1889
rect 555 1761 589 1795
rect 623 1761 657 1795
rect 734 1787 768 1821
rect 555 1687 589 1721
rect 623 1687 657 1721
rect 734 1719 768 1753
rect 734 1651 768 1685
rect 555 1616 589 1650
rect 623 1616 657 1650
rect 734 1583 768 1617
rect 555 1542 589 1576
rect 623 1542 657 1576
rect 734 1515 768 1549
rect 555 1471 589 1505
rect 623 1471 657 1505
rect 1678 2411 1712 2445
rect 1678 2343 1712 2377
rect 1678 2275 1712 2309
rect 1678 2207 1712 2241
rect 1678 2139 1712 2173
rect 1678 2071 1712 2105
rect 1678 2003 1712 2037
rect 1678 1935 1712 1969
rect 1678 1867 1712 1901
rect 1678 1799 1712 1833
rect 1678 1731 1712 1765
rect 1678 1663 1712 1697
rect 1678 1595 1712 1629
rect 1678 1527 1712 1561
rect 2670 2411 2704 2445
rect 2670 2343 2704 2377
rect 2670 2275 2704 2309
rect 2670 2207 2704 2241
rect 2670 2139 2704 2173
rect 2670 2071 2704 2105
rect 2670 2003 2704 2037
rect 2670 1935 2704 1969
rect 2670 1867 2704 1901
rect 2670 1799 2704 1833
rect 2670 1731 2704 1765
rect 2670 1663 2704 1697
rect 2670 1595 2704 1629
rect 2670 1527 2704 1561
rect 3662 2411 3696 2445
rect 3662 2343 3696 2377
rect 3662 2275 3696 2309
rect 3662 2207 3696 2241
rect 3662 2139 3696 2173
rect 3662 2071 3696 2105
rect 3662 2003 3696 2037
rect 3662 1935 3696 1969
rect 3662 1867 3696 1901
rect 3662 1799 3696 1833
rect 3662 1731 3696 1765
rect 3662 1663 3696 1697
rect 3662 1595 3696 1629
rect 3662 1527 3696 1561
rect 4654 2411 4688 2445
rect 4654 2343 4688 2377
rect 4654 2275 4688 2309
rect 4654 2207 4688 2241
rect 4654 2139 4688 2173
rect 4654 2071 4688 2105
rect 4654 2003 4688 2037
rect 4654 1935 4688 1969
rect 4654 1867 4688 1901
rect 4654 1799 4688 1833
rect 4654 1731 4688 1765
rect 4654 1663 4688 1697
rect 4654 1595 4688 1629
rect 4654 1527 4688 1561
rect 5646 2411 5680 2445
rect 5646 2343 5680 2377
rect 5646 2275 5680 2309
rect 5646 2207 5680 2241
rect 5646 2139 5680 2173
rect 5646 2071 5680 2105
rect 5646 2003 5680 2037
rect 5646 1935 5680 1969
rect 5646 1867 5680 1901
rect 5646 1799 5680 1833
rect 5646 1731 5680 1765
rect 5646 1663 5680 1697
rect 5646 1595 5680 1629
rect 5646 1527 5680 1561
rect 6638 2411 6672 2445
rect 6638 2343 6672 2377
rect 6638 2275 6672 2309
rect 6638 2207 6672 2241
rect 6638 2139 6672 2173
rect 6638 2071 6672 2105
rect 6638 2003 6672 2037
rect 6638 1935 6672 1969
rect 6638 1867 6672 1901
rect 6638 1799 6672 1833
rect 6638 1731 6672 1765
rect 6638 1663 6672 1697
rect 6638 1595 6672 1629
rect 6638 1527 6672 1561
rect 7630 2411 7664 2445
rect 7630 2343 7664 2377
rect 7630 2275 7664 2309
rect 7630 2207 7664 2241
rect 7630 2139 7664 2173
rect 7630 2071 7664 2105
rect 7630 2003 7664 2037
rect 7630 1935 7664 1969
rect 7630 1867 7664 1901
rect 7630 1799 7664 1833
rect 7630 1731 7664 1765
rect 7630 1663 7664 1697
rect 7630 1595 7664 1629
rect 7630 1527 7664 1561
rect 8622 2411 8656 2445
rect 8622 2343 8656 2377
rect 8622 2275 8656 2309
rect 8622 2207 8656 2241
rect 8622 2139 8656 2173
rect 8622 2071 8656 2105
rect 8622 2003 8656 2037
rect 8622 1935 8656 1969
rect 8622 1867 8656 1901
rect 8622 1799 8656 1833
rect 8622 1731 8656 1765
rect 8622 1663 8656 1697
rect 8622 1595 8656 1629
rect 8622 1527 8656 1561
rect 9614 2411 9648 2445
rect 9614 2343 9648 2377
rect 9614 2275 9648 2309
rect 9614 2207 9648 2241
rect 9614 2139 9648 2173
rect 9614 2071 9648 2105
rect 9614 2003 9648 2037
rect 9614 1935 9648 1969
rect 9614 1867 9648 1901
rect 9614 1799 9648 1833
rect 9614 1731 9648 1765
rect 9614 1663 9648 1697
rect 9614 1595 9648 1629
rect 9614 1527 9648 1561
rect 10606 2411 10640 2445
rect 10606 2343 10640 2377
rect 10606 2275 10640 2309
rect 10606 2207 10640 2241
rect 10606 2139 10640 2173
rect 10606 2071 10640 2105
rect 10606 2003 10640 2037
rect 10606 1935 10640 1969
rect 10606 1867 10640 1901
rect 10606 1799 10640 1833
rect 10606 1731 10640 1765
rect 10606 1663 10640 1697
rect 10606 1595 10640 1629
rect 10606 1527 10640 1561
rect 11598 2411 11632 2445
rect 11598 2343 11632 2377
rect 11598 2275 11632 2309
rect 11598 2207 11632 2241
rect 11598 2139 11632 2173
rect 11598 2071 11632 2105
rect 11598 2003 11632 2037
rect 11598 1935 11632 1969
rect 11598 1867 11632 1901
rect 11598 1799 11632 1833
rect 11598 1731 11632 1765
rect 11598 1663 11632 1697
rect 11598 1595 11632 1629
rect 11598 1527 11632 1561
rect 12590 2411 12624 2445
rect 12590 2343 12624 2377
rect 12590 2275 12624 2309
rect 12590 2207 12624 2241
rect 12590 2139 12624 2173
rect 12590 2071 12624 2105
rect 12590 2003 12624 2037
rect 12590 1935 12624 1969
rect 12590 1867 12624 1901
rect 12590 1799 12624 1833
rect 12590 1731 12624 1765
rect 12590 1663 12624 1697
rect 12590 1595 12624 1629
rect 12590 1527 12624 1561
rect 13582 2411 13616 2445
rect 13582 2343 13616 2377
rect 13582 2275 13616 2309
rect 13582 2207 13616 2241
rect 13582 2139 13616 2173
rect 13582 2071 13616 2105
rect 13582 2003 13616 2037
rect 13582 1935 13616 1969
rect 13582 1867 13616 1901
rect 13582 1799 13616 1833
rect 13582 1731 13616 1765
rect 13582 1663 13616 1697
rect 13582 1595 13616 1629
rect 13582 1527 13616 1561
rect 14565 2451 14599 2485
rect 14633 2451 14667 2485
rect 14454 2399 14488 2433
rect 14565 2369 14599 2403
rect 14633 2369 14667 2403
rect 14454 2331 14488 2365
rect 14454 2263 14488 2297
rect 14565 2293 14599 2327
rect 14633 2293 14667 2327
rect 14454 2195 14488 2229
rect 14565 2216 14599 2250
rect 14633 2216 14667 2250
rect 14454 2127 14488 2161
rect 14565 2122 14599 2156
rect 14633 2122 14667 2156
rect 14454 2059 14488 2093
rect 14565 2051 14599 2085
rect 14633 2051 14667 2085
rect 14454 1991 14488 2025
rect 14565 1977 14599 2011
rect 14633 1977 14667 2011
rect 14454 1923 14488 1957
rect 14565 1906 14599 1940
rect 14633 1906 14667 1940
rect 14454 1855 14488 1889
rect 14565 1832 14599 1866
rect 14633 1832 14667 1866
rect 14454 1787 14488 1821
rect 14565 1761 14599 1795
rect 14633 1761 14667 1795
rect 14454 1719 14488 1753
rect 14565 1687 14599 1721
rect 14633 1687 14667 1721
rect 14454 1651 14488 1685
rect 14454 1583 14488 1617
rect 14565 1616 14599 1650
rect 14633 1616 14667 1650
rect 14454 1515 14488 1549
rect 14565 1542 14599 1576
rect 14633 1542 14667 1576
rect 14565 1471 14599 1505
rect 14633 1471 14667 1505
rect 555 1341 589 1375
rect 623 1341 657 1375
rect 691 1341 725 1375
rect 14497 1353 14531 1387
rect 14565 1353 14599 1387
rect 14633 1353 14667 1387
rect 555 1187 589 1221
rect 623 1187 657 1221
rect 691 1185 725 1219
rect 555 1106 589 1140
rect 623 1116 657 1150
rect 14497 1274 14531 1308
rect 14565 1277 14599 1311
rect 14633 1285 14667 1319
rect 14497 1194 14531 1228
rect 14565 1200 14599 1234
rect 14633 1217 14667 1251
rect 691 1114 725 1148
rect 760 1114 794 1148
rect 829 1080 14531 1148
rect 14565 1123 14599 1157
rect 14633 1149 14667 1183
rect 14633 1081 14667 1115
rect 623 1046 657 1080
rect 692 1046 726 1080
rect 761 1046 14599 1080
rect 761 1012 14565 1046
rect 14633 1012 14667 1046
rect 589 978 623 1012
rect 658 978 692 1012
rect 727 978 14565 1012
<< mvnsubdiffcont >>
rect 300 5388 334 5422
rect 369 5388 403 5422
rect 438 5388 472 5422
rect 507 5388 541 5422
rect 576 5388 610 5422
rect 645 5388 679 5422
rect 714 5388 748 5422
rect 783 5388 817 5422
rect 852 5388 886 5422
rect 921 5388 955 5422
rect 990 5388 1024 5422
rect 1059 5388 1093 5422
rect 1128 5388 1162 5422
rect 1197 5388 1231 5422
rect 1266 5388 1300 5422
rect 1335 5388 1369 5422
rect 1404 5388 1438 5422
rect 1473 5388 1507 5422
rect 1542 5388 1576 5422
rect 1611 5388 1645 5422
rect 1680 5388 1714 5422
rect 1749 5388 1783 5422
rect 1818 5388 1852 5422
rect 1887 5388 1921 5422
rect 1956 5388 1990 5422
rect 2025 5388 2059 5422
rect 2094 5388 2128 5422
rect 2163 5388 2197 5422
rect 232 5286 334 5354
rect 369 5320 403 5354
rect 438 5320 472 5354
rect 507 5320 541 5354
rect 576 5320 610 5354
rect 645 5320 679 5354
rect 714 5320 748 5354
rect 783 5320 817 5354
rect 852 5320 886 5354
rect 921 5320 955 5354
rect 990 5320 1024 5354
rect 1059 5320 1093 5354
rect 1128 5320 1162 5354
rect 1197 5320 1231 5354
rect 1266 5320 1300 5354
rect 1335 5320 1369 5354
rect 1404 5320 1438 5354
rect 1473 5320 1507 5354
rect 1542 5320 1576 5354
rect 1611 5320 1645 5354
rect 1680 5320 1714 5354
rect 1749 5320 1783 5354
rect 1818 5320 1852 5354
rect 1887 5320 1921 5354
rect 1956 5320 1990 5354
rect 2025 5320 2059 5354
rect 2094 5320 2128 5354
rect 2163 5320 2197 5354
rect 2232 5320 14914 5422
rect 232 764 402 5286
rect 437 5252 471 5286
rect 506 5252 540 5286
rect 575 5252 609 5286
rect 644 5252 678 5286
rect 713 5252 747 5286
rect 782 5252 816 5286
rect 851 5252 885 5286
rect 920 5252 954 5286
rect 989 5252 1023 5286
rect 1058 5252 1092 5286
rect 1127 5252 1161 5286
rect 1196 5252 1230 5286
rect 1265 5252 1299 5286
rect 1334 5252 1368 5286
rect 1403 5252 1437 5286
rect 1472 5252 1506 5286
rect 1541 5252 1575 5286
rect 1610 5252 1644 5286
rect 1679 5252 1713 5286
rect 1748 5252 1782 5286
rect 1817 5252 1851 5286
rect 1886 5252 1920 5286
rect 1955 5252 1989 5286
rect 2024 5252 2058 5286
rect 2093 5252 2127 5286
rect 2162 5252 2196 5286
rect 2231 5252 2265 5286
rect 2300 5252 14914 5320
rect 14820 5218 14914 5252
rect 232 696 334 764
rect 368 695 402 729
rect 232 627 266 661
rect 300 627 334 661
rect 14820 696 14990 5218
rect 368 592 12982 660
rect 13017 626 13051 660
rect 13086 626 13120 660
rect 13155 626 13189 660
rect 13224 626 13258 660
rect 13293 626 13327 660
rect 13362 626 13396 660
rect 13431 626 13465 660
rect 13500 626 13534 660
rect 13569 626 13603 660
rect 13638 626 13672 660
rect 13707 626 13741 660
rect 13776 626 13810 660
rect 13845 626 13879 660
rect 13914 626 13948 660
rect 13983 626 14017 660
rect 14052 626 14086 660
rect 14121 626 14155 660
rect 14190 626 14224 660
rect 14259 626 14293 660
rect 14328 626 14362 660
rect 14397 626 14431 660
rect 14466 626 14500 660
rect 14535 626 14569 660
rect 14604 626 14638 660
rect 14673 626 14707 660
rect 14742 626 14776 660
rect 14811 626 14845 660
rect 14880 626 14914 660
rect 232 558 266 592
rect 300 490 12982 592
rect 13017 558 13051 592
rect 13086 558 13120 592
rect 13155 558 13189 592
rect 13224 558 13258 592
rect 13293 558 13327 592
rect 13362 558 13396 592
rect 13431 558 13465 592
rect 13500 558 13534 592
rect 13569 558 13603 592
rect 13638 558 13672 592
rect 13707 558 13741 592
rect 13776 558 13810 592
rect 13845 558 13879 592
rect 13914 558 13948 592
rect 13983 558 14017 592
rect 14052 558 14086 592
rect 14121 558 14155 592
rect 14190 558 14224 592
rect 14259 558 14293 592
rect 14328 558 14362 592
rect 14397 558 14431 592
rect 14466 558 14500 592
rect 14535 558 14569 592
rect 14604 558 14638 592
rect 14673 558 14707 592
rect 14742 558 14776 592
rect 14811 558 14845 592
rect 14880 558 14914 592
rect 13017 490 13051 524
rect 13086 490 13120 524
rect 13155 490 13189 524
rect 13224 490 13258 524
rect 13293 490 13327 524
rect 13362 490 13396 524
rect 13431 490 13465 524
rect 13500 490 13534 524
rect 13569 490 13603 524
rect 13638 490 13672 524
rect 13707 490 13741 524
rect 13776 490 13810 524
rect 13845 490 13879 524
rect 13914 490 13948 524
rect 13983 490 14017 524
rect 14052 490 14086 524
rect 14121 490 14155 524
rect 14190 490 14224 524
rect 14259 490 14293 524
rect 14328 490 14362 524
rect 14397 490 14431 524
rect 14466 490 14500 524
rect 14535 490 14569 524
rect 14604 490 14638 524
rect 14673 490 14707 524
rect 14742 490 14776 524
rect 14811 490 14845 524
rect 14880 490 14914 524
<< poly >>
rect 924 4214 1044 4230
rect 924 4180 967 4214
rect 1001 4180 1044 4214
rect 924 4140 1044 4180
rect 924 4106 967 4140
rect 1001 4106 1044 4140
rect 924 4058 1044 4106
rect 1354 4214 1474 4230
rect 1354 4180 1397 4214
rect 1431 4180 1474 4214
rect 1354 4140 1474 4180
rect 1354 4106 1397 4140
rect 1431 4106 1474 4140
rect 1354 4058 1474 4106
rect 1916 4214 2036 4230
rect 1916 4180 1959 4214
rect 1993 4180 2036 4214
rect 1916 4140 2036 4180
rect 1916 4106 1959 4140
rect 1993 4106 2036 4140
rect 1916 4058 2036 4106
rect 2346 4214 2466 4230
rect 2346 4180 2389 4214
rect 2423 4180 2466 4214
rect 2346 4140 2466 4180
rect 2346 4106 2389 4140
rect 2423 4106 2466 4140
rect 2346 4058 2466 4106
rect 2908 4214 3028 4230
rect 2908 4180 2951 4214
rect 2985 4180 3028 4214
rect 2908 4140 3028 4180
rect 2908 4106 2951 4140
rect 2985 4106 3028 4140
rect 2908 4058 3028 4106
rect 3338 4214 3458 4230
rect 3338 4180 3381 4214
rect 3415 4180 3458 4214
rect 3338 4140 3458 4180
rect 3338 4106 3381 4140
rect 3415 4106 3458 4140
rect 3338 4058 3458 4106
rect 3900 4214 4020 4230
rect 3900 4180 3943 4214
rect 3977 4180 4020 4214
rect 3900 4140 4020 4180
rect 3900 4106 3943 4140
rect 3977 4106 4020 4140
rect 3900 4058 4020 4106
rect 4330 4214 4450 4230
rect 4330 4180 4373 4214
rect 4407 4180 4450 4214
rect 4330 4140 4450 4180
rect 4330 4106 4373 4140
rect 4407 4106 4450 4140
rect 4330 4058 4450 4106
rect 4892 4214 5012 4230
rect 4892 4180 4935 4214
rect 4969 4180 5012 4214
rect 4892 4140 5012 4180
rect 4892 4106 4935 4140
rect 4969 4106 5012 4140
rect 4892 4058 5012 4106
rect 5322 4214 5442 4230
rect 5322 4180 5365 4214
rect 5399 4180 5442 4214
rect 5322 4140 5442 4180
rect 5322 4106 5365 4140
rect 5399 4106 5442 4140
rect 5322 4058 5442 4106
rect 5884 4214 6004 4230
rect 5884 4180 5927 4214
rect 5961 4180 6004 4214
rect 5884 4140 6004 4180
rect 5884 4106 5927 4140
rect 5961 4106 6004 4140
rect 5884 4058 6004 4106
rect 6314 4214 6434 4230
rect 6314 4180 6357 4214
rect 6391 4180 6434 4214
rect 6314 4140 6434 4180
rect 6314 4106 6357 4140
rect 6391 4106 6434 4140
rect 6314 4058 6434 4106
rect 6876 4214 6996 4230
rect 6876 4180 6919 4214
rect 6953 4180 6996 4214
rect 6876 4140 6996 4180
rect 6876 4106 6919 4140
rect 6953 4106 6996 4140
rect 6876 4058 6996 4106
rect 7306 4214 7426 4230
rect 7306 4180 7349 4214
rect 7383 4180 7426 4214
rect 7306 4140 7426 4180
rect 7306 4106 7349 4140
rect 7383 4106 7426 4140
rect 7306 4058 7426 4106
rect 7868 4214 7988 4230
rect 7868 4180 7911 4214
rect 7945 4180 7988 4214
rect 7868 4140 7988 4180
rect 7868 4106 7911 4140
rect 7945 4106 7988 4140
rect 7868 4058 7988 4106
rect 8298 4214 8418 4230
rect 8298 4180 8341 4214
rect 8375 4180 8418 4214
rect 8298 4140 8418 4180
rect 8298 4106 8341 4140
rect 8375 4106 8418 4140
rect 8298 4058 8418 4106
rect 8860 4214 8980 4230
rect 8860 4180 8903 4214
rect 8937 4180 8980 4214
rect 8860 4140 8980 4180
rect 8860 4106 8903 4140
rect 8937 4106 8980 4140
rect 8860 4058 8980 4106
rect 9290 4214 9410 4230
rect 9290 4180 9333 4214
rect 9367 4180 9410 4214
rect 9290 4140 9410 4180
rect 9290 4106 9333 4140
rect 9367 4106 9410 4140
rect 9290 4058 9410 4106
rect 9852 4214 9972 4230
rect 9852 4180 9895 4214
rect 9929 4180 9972 4214
rect 9852 4140 9972 4180
rect 9852 4106 9895 4140
rect 9929 4106 9972 4140
rect 9852 4058 9972 4106
rect 10282 4214 10402 4230
rect 10282 4180 10325 4214
rect 10359 4180 10402 4214
rect 10282 4140 10402 4180
rect 10282 4106 10325 4140
rect 10359 4106 10402 4140
rect 10282 4058 10402 4106
rect 10844 4214 10964 4230
rect 10844 4180 10887 4214
rect 10921 4180 10964 4214
rect 10844 4140 10964 4180
rect 10844 4106 10887 4140
rect 10921 4106 10964 4140
rect 10844 4058 10964 4106
rect 11274 4214 11394 4230
rect 11274 4180 11317 4214
rect 11351 4180 11394 4214
rect 11274 4140 11394 4180
rect 11274 4106 11317 4140
rect 11351 4106 11394 4140
rect 11274 4058 11394 4106
rect 11836 4214 11956 4230
rect 11836 4180 11879 4214
rect 11913 4180 11956 4214
rect 11836 4140 11956 4180
rect 11836 4106 11879 4140
rect 11913 4106 11956 4140
rect 11836 4058 11956 4106
rect 12266 4214 12386 4230
rect 12266 4180 12309 4214
rect 12343 4180 12386 4214
rect 12266 4140 12386 4180
rect 12266 4106 12309 4140
rect 12343 4106 12386 4140
rect 12266 4058 12386 4106
rect 12828 4214 12948 4230
rect 12828 4180 12871 4214
rect 12905 4180 12948 4214
rect 12828 4140 12948 4180
rect 12828 4106 12871 4140
rect 12905 4106 12948 4140
rect 12828 4058 12948 4106
rect 13258 4214 13378 4230
rect 13258 4180 13301 4214
rect 13335 4180 13378 4214
rect 13258 4140 13378 4180
rect 13258 4106 13301 4140
rect 13335 4106 13378 4140
rect 13258 4058 13378 4106
rect 13820 4214 13940 4230
rect 13820 4180 13863 4214
rect 13897 4180 13940 4214
rect 13820 4140 13940 4180
rect 13820 4106 13863 4140
rect 13897 4106 13940 4140
rect 13820 4058 13940 4106
rect 14178 4214 14298 4230
rect 14178 4180 14221 4214
rect 14255 4180 14298 4214
rect 14178 4140 14298 4180
rect 14178 4106 14221 4140
rect 14255 4106 14298 4140
rect 14178 4058 14298 4106
rect 924 3010 1044 3058
rect 924 2976 967 3010
rect 1001 2976 1044 3010
rect 924 2932 1044 2976
rect 924 2898 967 2932
rect 1001 2898 1044 2932
rect 924 2854 1044 2898
rect 924 2820 967 2854
rect 1001 2820 1044 2854
rect 924 2776 1044 2820
rect 924 2742 967 2776
rect 1001 2742 1044 2776
rect 924 2697 1044 2742
rect 924 2663 967 2697
rect 1001 2663 1044 2697
rect 924 2618 1044 2663
rect 924 2584 967 2618
rect 1001 2584 1044 2618
rect 924 2539 1044 2584
rect 924 2505 967 2539
rect 1001 2505 1044 2539
rect 924 2457 1044 2505
rect 1354 3010 1474 3058
rect 1354 2976 1397 3010
rect 1431 2976 1474 3010
rect 1354 2932 1474 2976
rect 1916 3010 2036 3058
rect 1916 2976 1959 3010
rect 1993 2976 2036 3010
rect 1354 2898 1397 2932
rect 1431 2898 1474 2932
rect 1354 2854 1474 2898
rect 1354 2820 1397 2854
rect 1431 2820 1474 2854
rect 1354 2776 1474 2820
rect 1354 2742 1397 2776
rect 1431 2742 1474 2776
rect 1354 2697 1474 2742
rect 1354 2663 1397 2697
rect 1431 2663 1474 2697
rect 1354 2618 1474 2663
rect 1354 2584 1397 2618
rect 1431 2584 1474 2618
rect 1354 2539 1474 2584
rect 1916 2932 2036 2976
rect 1916 2898 1959 2932
rect 1993 2898 2036 2932
rect 1916 2854 2036 2898
rect 1916 2820 1959 2854
rect 1993 2820 2036 2854
rect 1916 2776 2036 2820
rect 1916 2742 1959 2776
rect 1993 2742 2036 2776
rect 1916 2697 2036 2742
rect 1916 2663 1959 2697
rect 1993 2663 2036 2697
rect 1916 2618 2036 2663
rect 1916 2584 1959 2618
rect 1993 2584 2036 2618
rect 1354 2505 1397 2539
rect 1431 2505 1474 2539
rect 1354 2457 1474 2505
rect 1916 2539 2036 2584
rect 1916 2505 1959 2539
rect 1993 2505 2036 2539
rect 1916 2457 2036 2505
rect 2346 3010 2466 3058
rect 2346 2976 2389 3010
rect 2423 2976 2466 3010
rect 2346 2932 2466 2976
rect 2908 3010 3028 3058
rect 2908 2976 2951 3010
rect 2985 2976 3028 3010
rect 2346 2898 2389 2932
rect 2423 2898 2466 2932
rect 2346 2854 2466 2898
rect 2346 2820 2389 2854
rect 2423 2820 2466 2854
rect 2346 2776 2466 2820
rect 2346 2742 2389 2776
rect 2423 2742 2466 2776
rect 2346 2697 2466 2742
rect 2346 2663 2389 2697
rect 2423 2663 2466 2697
rect 2346 2618 2466 2663
rect 2346 2584 2389 2618
rect 2423 2584 2466 2618
rect 2346 2539 2466 2584
rect 2908 2932 3028 2976
rect 2908 2898 2951 2932
rect 2985 2898 3028 2932
rect 2908 2854 3028 2898
rect 2908 2820 2951 2854
rect 2985 2820 3028 2854
rect 2908 2776 3028 2820
rect 2908 2742 2951 2776
rect 2985 2742 3028 2776
rect 2908 2697 3028 2742
rect 2908 2663 2951 2697
rect 2985 2663 3028 2697
rect 2908 2618 3028 2663
rect 2908 2584 2951 2618
rect 2985 2584 3028 2618
rect 2346 2505 2389 2539
rect 2423 2505 2466 2539
rect 2346 2457 2466 2505
rect 2908 2539 3028 2584
rect 2908 2505 2951 2539
rect 2985 2505 3028 2539
rect 2908 2457 3028 2505
rect 3338 3010 3458 3058
rect 3338 2976 3381 3010
rect 3415 2976 3458 3010
rect 3338 2932 3458 2976
rect 3900 3010 4020 3058
rect 3900 2976 3943 3010
rect 3977 2976 4020 3010
rect 3338 2898 3381 2932
rect 3415 2898 3458 2932
rect 3338 2854 3458 2898
rect 3338 2820 3381 2854
rect 3415 2820 3458 2854
rect 3338 2776 3458 2820
rect 3338 2742 3381 2776
rect 3415 2742 3458 2776
rect 3338 2697 3458 2742
rect 3338 2663 3381 2697
rect 3415 2663 3458 2697
rect 3338 2618 3458 2663
rect 3338 2584 3381 2618
rect 3415 2584 3458 2618
rect 3338 2539 3458 2584
rect 3900 2932 4020 2976
rect 3900 2898 3943 2932
rect 3977 2898 4020 2932
rect 3900 2854 4020 2898
rect 3900 2820 3943 2854
rect 3977 2820 4020 2854
rect 3900 2776 4020 2820
rect 3900 2742 3943 2776
rect 3977 2742 4020 2776
rect 3900 2697 4020 2742
rect 3900 2663 3943 2697
rect 3977 2663 4020 2697
rect 3900 2618 4020 2663
rect 3900 2584 3943 2618
rect 3977 2584 4020 2618
rect 3338 2505 3381 2539
rect 3415 2505 3458 2539
rect 3338 2457 3458 2505
rect 3900 2539 4020 2584
rect 3900 2505 3943 2539
rect 3977 2505 4020 2539
rect 3900 2457 4020 2505
rect 4330 3010 4450 3058
rect 4330 2976 4373 3010
rect 4407 2976 4450 3010
rect 4330 2932 4450 2976
rect 4892 3010 5012 3058
rect 4892 2976 4935 3010
rect 4969 2976 5012 3010
rect 4330 2898 4373 2932
rect 4407 2898 4450 2932
rect 4330 2854 4450 2898
rect 4330 2820 4373 2854
rect 4407 2820 4450 2854
rect 4330 2776 4450 2820
rect 4330 2742 4373 2776
rect 4407 2742 4450 2776
rect 4330 2697 4450 2742
rect 4330 2663 4373 2697
rect 4407 2663 4450 2697
rect 4330 2618 4450 2663
rect 4330 2584 4373 2618
rect 4407 2584 4450 2618
rect 4330 2539 4450 2584
rect 4892 2932 5012 2976
rect 4892 2898 4935 2932
rect 4969 2898 5012 2932
rect 4892 2854 5012 2898
rect 4892 2820 4935 2854
rect 4969 2820 5012 2854
rect 4892 2776 5012 2820
rect 4892 2742 4935 2776
rect 4969 2742 5012 2776
rect 4892 2697 5012 2742
rect 4892 2663 4935 2697
rect 4969 2663 5012 2697
rect 4892 2618 5012 2663
rect 4892 2584 4935 2618
rect 4969 2584 5012 2618
rect 4330 2505 4373 2539
rect 4407 2505 4450 2539
rect 4330 2457 4450 2505
rect 4892 2539 5012 2584
rect 4892 2505 4935 2539
rect 4969 2505 5012 2539
rect 4892 2457 5012 2505
rect 5322 3010 5442 3058
rect 5322 2976 5365 3010
rect 5399 2976 5442 3010
rect 5322 2932 5442 2976
rect 5884 3010 6004 3058
rect 5884 2976 5927 3010
rect 5961 2976 6004 3010
rect 5322 2898 5365 2932
rect 5399 2898 5442 2932
rect 5322 2854 5442 2898
rect 5322 2820 5365 2854
rect 5399 2820 5442 2854
rect 5322 2776 5442 2820
rect 5322 2742 5365 2776
rect 5399 2742 5442 2776
rect 5322 2697 5442 2742
rect 5322 2663 5365 2697
rect 5399 2663 5442 2697
rect 5322 2618 5442 2663
rect 5322 2584 5365 2618
rect 5399 2584 5442 2618
rect 5322 2539 5442 2584
rect 5884 2932 6004 2976
rect 5884 2898 5927 2932
rect 5961 2898 6004 2932
rect 5884 2854 6004 2898
rect 5884 2820 5927 2854
rect 5961 2820 6004 2854
rect 5884 2776 6004 2820
rect 5884 2742 5927 2776
rect 5961 2742 6004 2776
rect 5884 2697 6004 2742
rect 5884 2663 5927 2697
rect 5961 2663 6004 2697
rect 5884 2618 6004 2663
rect 5884 2584 5927 2618
rect 5961 2584 6004 2618
rect 5322 2505 5365 2539
rect 5399 2505 5442 2539
rect 5322 2457 5442 2505
rect 5884 2539 6004 2584
rect 5884 2505 5927 2539
rect 5961 2505 6004 2539
rect 5884 2457 6004 2505
rect 6314 3010 6434 3058
rect 6314 2976 6357 3010
rect 6391 2976 6434 3010
rect 6314 2932 6434 2976
rect 6876 3010 6996 3058
rect 6876 2976 6919 3010
rect 6953 2976 6996 3010
rect 6314 2898 6357 2932
rect 6391 2898 6434 2932
rect 6314 2854 6434 2898
rect 6314 2820 6357 2854
rect 6391 2820 6434 2854
rect 6314 2776 6434 2820
rect 6314 2742 6357 2776
rect 6391 2742 6434 2776
rect 6314 2697 6434 2742
rect 6314 2663 6357 2697
rect 6391 2663 6434 2697
rect 6314 2618 6434 2663
rect 6314 2584 6357 2618
rect 6391 2584 6434 2618
rect 6314 2539 6434 2584
rect 6876 2932 6996 2976
rect 6876 2898 6919 2932
rect 6953 2898 6996 2932
rect 6876 2854 6996 2898
rect 6876 2820 6919 2854
rect 6953 2820 6996 2854
rect 6876 2776 6996 2820
rect 6876 2742 6919 2776
rect 6953 2742 6996 2776
rect 6876 2697 6996 2742
rect 6876 2663 6919 2697
rect 6953 2663 6996 2697
rect 6876 2618 6996 2663
rect 6876 2584 6919 2618
rect 6953 2584 6996 2618
rect 6314 2505 6357 2539
rect 6391 2505 6434 2539
rect 6314 2457 6434 2505
rect 6876 2539 6996 2584
rect 6876 2505 6919 2539
rect 6953 2505 6996 2539
rect 6876 2457 6996 2505
rect 7306 3010 7426 3058
rect 7306 2976 7349 3010
rect 7383 2976 7426 3010
rect 7306 2932 7426 2976
rect 7868 3010 7988 3058
rect 7868 2976 7911 3010
rect 7945 2976 7988 3010
rect 7306 2898 7349 2932
rect 7383 2898 7426 2932
rect 7306 2854 7426 2898
rect 7306 2820 7349 2854
rect 7383 2820 7426 2854
rect 7306 2776 7426 2820
rect 7306 2742 7349 2776
rect 7383 2742 7426 2776
rect 7306 2697 7426 2742
rect 7306 2663 7349 2697
rect 7383 2663 7426 2697
rect 7306 2618 7426 2663
rect 7306 2584 7349 2618
rect 7383 2584 7426 2618
rect 7306 2539 7426 2584
rect 7868 2932 7988 2976
rect 7868 2898 7911 2932
rect 7945 2898 7988 2932
rect 7868 2854 7988 2898
rect 7868 2820 7911 2854
rect 7945 2820 7988 2854
rect 7868 2776 7988 2820
rect 7868 2742 7911 2776
rect 7945 2742 7988 2776
rect 7868 2697 7988 2742
rect 7868 2663 7911 2697
rect 7945 2663 7988 2697
rect 7868 2618 7988 2663
rect 7868 2584 7911 2618
rect 7945 2584 7988 2618
rect 7306 2505 7349 2539
rect 7383 2505 7426 2539
rect 7306 2457 7426 2505
rect 7868 2539 7988 2584
rect 7868 2505 7911 2539
rect 7945 2505 7988 2539
rect 7868 2457 7988 2505
rect 8298 3010 8418 3058
rect 8298 2976 8341 3010
rect 8375 2976 8418 3010
rect 8298 2932 8418 2976
rect 8860 3010 8980 3058
rect 8860 2976 8903 3010
rect 8937 2976 8980 3010
rect 8298 2898 8341 2932
rect 8375 2898 8418 2932
rect 8298 2854 8418 2898
rect 8298 2820 8341 2854
rect 8375 2820 8418 2854
rect 8298 2776 8418 2820
rect 8298 2742 8341 2776
rect 8375 2742 8418 2776
rect 8298 2697 8418 2742
rect 8298 2663 8341 2697
rect 8375 2663 8418 2697
rect 8298 2618 8418 2663
rect 8298 2584 8341 2618
rect 8375 2584 8418 2618
rect 8298 2539 8418 2584
rect 8860 2932 8980 2976
rect 8860 2898 8903 2932
rect 8937 2898 8980 2932
rect 8860 2854 8980 2898
rect 8860 2820 8903 2854
rect 8937 2820 8980 2854
rect 8860 2776 8980 2820
rect 8860 2742 8903 2776
rect 8937 2742 8980 2776
rect 8860 2697 8980 2742
rect 8860 2663 8903 2697
rect 8937 2663 8980 2697
rect 8860 2618 8980 2663
rect 8860 2584 8903 2618
rect 8937 2584 8980 2618
rect 8298 2505 8341 2539
rect 8375 2505 8418 2539
rect 8298 2457 8418 2505
rect 8860 2539 8980 2584
rect 8860 2505 8903 2539
rect 8937 2505 8980 2539
rect 8860 2457 8980 2505
rect 9290 3010 9410 3058
rect 9290 2976 9333 3010
rect 9367 2976 9410 3010
rect 9290 2932 9410 2976
rect 9852 3010 9972 3058
rect 9852 2976 9895 3010
rect 9929 2976 9972 3010
rect 9290 2898 9333 2932
rect 9367 2898 9410 2932
rect 9290 2854 9410 2898
rect 9290 2820 9333 2854
rect 9367 2820 9410 2854
rect 9290 2776 9410 2820
rect 9290 2742 9333 2776
rect 9367 2742 9410 2776
rect 9290 2697 9410 2742
rect 9290 2663 9333 2697
rect 9367 2663 9410 2697
rect 9290 2618 9410 2663
rect 9290 2584 9333 2618
rect 9367 2584 9410 2618
rect 9290 2539 9410 2584
rect 9852 2932 9972 2976
rect 9852 2898 9895 2932
rect 9929 2898 9972 2932
rect 9852 2854 9972 2898
rect 9852 2820 9895 2854
rect 9929 2820 9972 2854
rect 9852 2776 9972 2820
rect 9852 2742 9895 2776
rect 9929 2742 9972 2776
rect 9852 2697 9972 2742
rect 9852 2663 9895 2697
rect 9929 2663 9972 2697
rect 9852 2618 9972 2663
rect 9852 2584 9895 2618
rect 9929 2584 9972 2618
rect 9290 2505 9333 2539
rect 9367 2505 9410 2539
rect 9290 2457 9410 2505
rect 9852 2539 9972 2584
rect 9852 2505 9895 2539
rect 9929 2505 9972 2539
rect 9852 2457 9972 2505
rect 10282 3010 10402 3058
rect 10282 2976 10325 3010
rect 10359 2976 10402 3010
rect 10282 2932 10402 2976
rect 10844 3010 10964 3058
rect 10844 2976 10887 3010
rect 10921 2976 10964 3010
rect 10282 2898 10325 2932
rect 10359 2898 10402 2932
rect 10282 2854 10402 2898
rect 10282 2820 10325 2854
rect 10359 2820 10402 2854
rect 10282 2776 10402 2820
rect 10282 2742 10325 2776
rect 10359 2742 10402 2776
rect 10282 2697 10402 2742
rect 10282 2663 10325 2697
rect 10359 2663 10402 2697
rect 10282 2618 10402 2663
rect 10282 2584 10325 2618
rect 10359 2584 10402 2618
rect 10282 2539 10402 2584
rect 10844 2932 10964 2976
rect 10844 2898 10887 2932
rect 10921 2898 10964 2932
rect 10844 2854 10964 2898
rect 10844 2820 10887 2854
rect 10921 2820 10964 2854
rect 10844 2776 10964 2820
rect 10844 2742 10887 2776
rect 10921 2742 10964 2776
rect 10844 2697 10964 2742
rect 10844 2663 10887 2697
rect 10921 2663 10964 2697
rect 10844 2618 10964 2663
rect 10844 2584 10887 2618
rect 10921 2584 10964 2618
rect 10282 2505 10325 2539
rect 10359 2505 10402 2539
rect 10282 2457 10402 2505
rect 10844 2539 10964 2584
rect 10844 2505 10887 2539
rect 10921 2505 10964 2539
rect 10844 2457 10964 2505
rect 11274 3010 11394 3058
rect 11274 2976 11317 3010
rect 11351 2976 11394 3010
rect 11274 2932 11394 2976
rect 11836 3010 11956 3058
rect 11836 2976 11879 3010
rect 11913 2976 11956 3010
rect 11274 2898 11317 2932
rect 11351 2898 11394 2932
rect 11274 2854 11394 2898
rect 11274 2820 11317 2854
rect 11351 2820 11394 2854
rect 11274 2776 11394 2820
rect 11274 2742 11317 2776
rect 11351 2742 11394 2776
rect 11274 2697 11394 2742
rect 11274 2663 11317 2697
rect 11351 2663 11394 2697
rect 11274 2618 11394 2663
rect 11274 2584 11317 2618
rect 11351 2584 11394 2618
rect 11274 2539 11394 2584
rect 11836 2932 11956 2976
rect 11836 2898 11879 2932
rect 11913 2898 11956 2932
rect 11836 2854 11956 2898
rect 11836 2820 11879 2854
rect 11913 2820 11956 2854
rect 11836 2776 11956 2820
rect 11836 2742 11879 2776
rect 11913 2742 11956 2776
rect 11836 2697 11956 2742
rect 11836 2663 11879 2697
rect 11913 2663 11956 2697
rect 11836 2618 11956 2663
rect 11836 2584 11879 2618
rect 11913 2584 11956 2618
rect 11274 2505 11317 2539
rect 11351 2505 11394 2539
rect 11274 2457 11394 2505
rect 11836 2539 11956 2584
rect 11836 2505 11879 2539
rect 11913 2505 11956 2539
rect 11836 2457 11956 2505
rect 12266 3010 12386 3058
rect 12266 2976 12309 3010
rect 12343 2976 12386 3010
rect 12266 2932 12386 2976
rect 12828 3010 12948 3058
rect 12828 2976 12871 3010
rect 12905 2976 12948 3010
rect 12266 2898 12309 2932
rect 12343 2898 12386 2932
rect 12266 2854 12386 2898
rect 12266 2820 12309 2854
rect 12343 2820 12386 2854
rect 12266 2776 12386 2820
rect 12266 2742 12309 2776
rect 12343 2742 12386 2776
rect 12266 2697 12386 2742
rect 12266 2663 12309 2697
rect 12343 2663 12386 2697
rect 12266 2618 12386 2663
rect 12266 2584 12309 2618
rect 12343 2584 12386 2618
rect 12266 2539 12386 2584
rect 12828 2932 12948 2976
rect 12828 2898 12871 2932
rect 12905 2898 12948 2932
rect 12828 2854 12948 2898
rect 12828 2820 12871 2854
rect 12905 2820 12948 2854
rect 12828 2776 12948 2820
rect 12828 2742 12871 2776
rect 12905 2742 12948 2776
rect 12828 2697 12948 2742
rect 12828 2663 12871 2697
rect 12905 2663 12948 2697
rect 12828 2618 12948 2663
rect 12828 2584 12871 2618
rect 12905 2584 12948 2618
rect 12266 2505 12309 2539
rect 12343 2505 12386 2539
rect 12266 2457 12386 2505
rect 12828 2539 12948 2584
rect 12828 2505 12871 2539
rect 12905 2505 12948 2539
rect 12828 2457 12948 2505
rect 13258 3010 13378 3058
rect 13258 2976 13301 3010
rect 13335 2976 13378 3010
rect 13258 2932 13378 2976
rect 13820 3010 13940 3058
rect 13820 2976 13863 3010
rect 13897 2976 13940 3010
rect 13258 2898 13301 2932
rect 13335 2898 13378 2932
rect 13258 2854 13378 2898
rect 13258 2820 13301 2854
rect 13335 2820 13378 2854
rect 13258 2776 13378 2820
rect 13258 2742 13301 2776
rect 13335 2742 13378 2776
rect 13258 2697 13378 2742
rect 13258 2663 13301 2697
rect 13335 2663 13378 2697
rect 13258 2618 13378 2663
rect 13258 2584 13301 2618
rect 13335 2584 13378 2618
rect 13258 2539 13378 2584
rect 13820 2932 13940 2976
rect 13820 2898 13863 2932
rect 13897 2898 13940 2932
rect 13820 2854 13940 2898
rect 13820 2820 13863 2854
rect 13897 2820 13940 2854
rect 13820 2776 13940 2820
rect 13820 2742 13863 2776
rect 13897 2742 13940 2776
rect 13820 2697 13940 2742
rect 13820 2663 13863 2697
rect 13897 2663 13940 2697
rect 13820 2618 13940 2663
rect 13820 2584 13863 2618
rect 13897 2584 13940 2618
rect 13258 2505 13301 2539
rect 13335 2505 13378 2539
rect 13258 2457 13378 2505
rect 13820 2539 13940 2584
rect 13820 2505 13863 2539
rect 13897 2505 13940 2539
rect 13820 2457 13940 2505
rect 14178 3010 14298 3058
rect 14178 2976 14221 3010
rect 14255 2976 14298 3010
rect 14178 2932 14298 2976
rect 14178 2898 14221 2932
rect 14255 2898 14298 2932
rect 14178 2854 14298 2898
rect 14178 2820 14221 2854
rect 14255 2820 14298 2854
rect 14178 2776 14298 2820
rect 14178 2742 14221 2776
rect 14255 2742 14298 2776
rect 14178 2697 14298 2742
rect 14178 2663 14221 2697
rect 14255 2663 14298 2697
rect 14178 2618 14298 2663
rect 14178 2584 14221 2618
rect 14255 2584 14298 2618
rect 14178 2539 14298 2584
rect 14178 2505 14221 2539
rect 14255 2505 14298 2539
rect 14178 2457 14298 2505
rect 924 1409 1044 1457
rect 924 1375 967 1409
rect 1001 1375 1044 1409
rect 924 1335 1044 1375
rect 924 1301 967 1335
rect 1001 1301 1044 1335
rect 924 1285 1044 1301
rect 1354 1409 1474 1457
rect 1354 1375 1397 1409
rect 1431 1375 1474 1409
rect 1354 1335 1474 1375
rect 1354 1301 1397 1335
rect 1431 1301 1474 1335
rect 1354 1285 1474 1301
rect 1916 1409 2036 1457
rect 1916 1375 1959 1409
rect 1993 1375 2036 1409
rect 1916 1335 2036 1375
rect 1916 1301 1959 1335
rect 1993 1301 2036 1335
rect 1916 1285 2036 1301
rect 2346 1409 2466 1457
rect 2346 1375 2389 1409
rect 2423 1375 2466 1409
rect 2346 1335 2466 1375
rect 2346 1301 2389 1335
rect 2423 1301 2466 1335
rect 2346 1285 2466 1301
rect 2908 1409 3028 1457
rect 2908 1375 2951 1409
rect 2985 1375 3028 1409
rect 2908 1335 3028 1375
rect 2908 1301 2951 1335
rect 2985 1301 3028 1335
rect 2908 1285 3028 1301
rect 3338 1409 3458 1457
rect 3338 1375 3381 1409
rect 3415 1375 3458 1409
rect 3338 1335 3458 1375
rect 3338 1301 3381 1335
rect 3415 1301 3458 1335
rect 3338 1285 3458 1301
rect 3900 1409 4020 1457
rect 3900 1375 3943 1409
rect 3977 1375 4020 1409
rect 3900 1335 4020 1375
rect 3900 1301 3943 1335
rect 3977 1301 4020 1335
rect 3900 1285 4020 1301
rect 4330 1409 4450 1457
rect 4330 1375 4373 1409
rect 4407 1375 4450 1409
rect 4330 1335 4450 1375
rect 4330 1301 4373 1335
rect 4407 1301 4450 1335
rect 4330 1285 4450 1301
rect 4892 1409 5012 1457
rect 4892 1375 4935 1409
rect 4969 1375 5012 1409
rect 4892 1335 5012 1375
rect 4892 1301 4935 1335
rect 4969 1301 5012 1335
rect 4892 1285 5012 1301
rect 5322 1409 5442 1457
rect 5322 1375 5365 1409
rect 5399 1375 5442 1409
rect 5322 1335 5442 1375
rect 5322 1301 5365 1335
rect 5399 1301 5442 1335
rect 5322 1285 5442 1301
rect 5884 1409 6004 1457
rect 5884 1375 5927 1409
rect 5961 1375 6004 1409
rect 5884 1335 6004 1375
rect 5884 1301 5927 1335
rect 5961 1301 6004 1335
rect 5884 1285 6004 1301
rect 6314 1409 6434 1457
rect 6314 1375 6357 1409
rect 6391 1375 6434 1409
rect 6314 1335 6434 1375
rect 6314 1301 6357 1335
rect 6391 1301 6434 1335
rect 6314 1285 6434 1301
rect 6876 1409 6996 1457
rect 6876 1375 6919 1409
rect 6953 1375 6996 1409
rect 6876 1335 6996 1375
rect 6876 1301 6919 1335
rect 6953 1301 6996 1335
rect 6876 1285 6996 1301
rect 7306 1409 7426 1457
rect 7306 1375 7349 1409
rect 7383 1375 7426 1409
rect 7306 1335 7426 1375
rect 7306 1301 7349 1335
rect 7383 1301 7426 1335
rect 7306 1285 7426 1301
rect 7868 1409 7988 1457
rect 7868 1375 7911 1409
rect 7945 1375 7988 1409
rect 7868 1335 7988 1375
rect 7868 1301 7911 1335
rect 7945 1301 7988 1335
rect 7868 1285 7988 1301
rect 8298 1409 8418 1457
rect 8298 1375 8341 1409
rect 8375 1375 8418 1409
rect 8298 1335 8418 1375
rect 8298 1301 8341 1335
rect 8375 1301 8418 1335
rect 8298 1285 8418 1301
rect 8860 1409 8980 1457
rect 8860 1375 8903 1409
rect 8937 1375 8980 1409
rect 8860 1335 8980 1375
rect 8860 1301 8903 1335
rect 8937 1301 8980 1335
rect 8860 1285 8980 1301
rect 9290 1409 9410 1457
rect 9290 1375 9333 1409
rect 9367 1375 9410 1409
rect 9290 1335 9410 1375
rect 9290 1301 9333 1335
rect 9367 1301 9410 1335
rect 9290 1285 9410 1301
rect 9852 1409 9972 1457
rect 9852 1375 9895 1409
rect 9929 1375 9972 1409
rect 9852 1335 9972 1375
rect 9852 1301 9895 1335
rect 9929 1301 9972 1335
rect 9852 1285 9972 1301
rect 10282 1409 10402 1457
rect 10282 1375 10325 1409
rect 10359 1375 10402 1409
rect 10282 1335 10402 1375
rect 10282 1301 10325 1335
rect 10359 1301 10402 1335
rect 10282 1285 10402 1301
rect 10844 1409 10964 1457
rect 10844 1375 10887 1409
rect 10921 1375 10964 1409
rect 10844 1335 10964 1375
rect 10844 1301 10887 1335
rect 10921 1301 10964 1335
rect 10844 1285 10964 1301
rect 11274 1409 11394 1457
rect 11274 1375 11317 1409
rect 11351 1375 11394 1409
rect 11274 1335 11394 1375
rect 11274 1301 11317 1335
rect 11351 1301 11394 1335
rect 11274 1285 11394 1301
rect 11836 1409 11956 1457
rect 11836 1375 11879 1409
rect 11913 1375 11956 1409
rect 11836 1335 11956 1375
rect 11836 1301 11879 1335
rect 11913 1301 11956 1335
rect 11836 1285 11956 1301
rect 12266 1409 12386 1457
rect 12266 1375 12309 1409
rect 12343 1375 12386 1409
rect 12266 1335 12386 1375
rect 12266 1301 12309 1335
rect 12343 1301 12386 1335
rect 12266 1285 12386 1301
rect 12828 1409 12948 1457
rect 12828 1375 12871 1409
rect 12905 1375 12948 1409
rect 12828 1335 12948 1375
rect 12828 1301 12871 1335
rect 12905 1301 12948 1335
rect 12828 1285 12948 1301
rect 13258 1409 13378 1457
rect 13258 1375 13301 1409
rect 13335 1375 13378 1409
rect 13258 1335 13378 1375
rect 13258 1301 13301 1335
rect 13335 1301 13378 1335
rect 13258 1285 13378 1301
rect 13820 1409 13940 1457
rect 13820 1375 13863 1409
rect 13897 1375 13940 1409
rect 13820 1335 13940 1375
rect 13820 1301 13863 1335
rect 13897 1301 13940 1335
rect 13820 1285 13940 1301
rect 14178 1409 14298 1457
rect 14178 1375 14221 1409
rect 14255 1375 14298 1409
rect 14178 1335 14298 1375
rect 14178 1301 14221 1335
rect 14255 1301 14298 1335
rect 14178 1285 14298 1301
<< polycont >>
rect 967 4180 1001 4214
rect 967 4106 1001 4140
rect 1397 4180 1431 4214
rect 1397 4106 1431 4140
rect 1959 4180 1993 4214
rect 1959 4106 1993 4140
rect 2389 4180 2423 4214
rect 2389 4106 2423 4140
rect 2951 4180 2985 4214
rect 2951 4106 2985 4140
rect 3381 4180 3415 4214
rect 3381 4106 3415 4140
rect 3943 4180 3977 4214
rect 3943 4106 3977 4140
rect 4373 4180 4407 4214
rect 4373 4106 4407 4140
rect 4935 4180 4969 4214
rect 4935 4106 4969 4140
rect 5365 4180 5399 4214
rect 5365 4106 5399 4140
rect 5927 4180 5961 4214
rect 5927 4106 5961 4140
rect 6357 4180 6391 4214
rect 6357 4106 6391 4140
rect 6919 4180 6953 4214
rect 6919 4106 6953 4140
rect 7349 4180 7383 4214
rect 7349 4106 7383 4140
rect 7911 4180 7945 4214
rect 7911 4106 7945 4140
rect 8341 4180 8375 4214
rect 8341 4106 8375 4140
rect 8903 4180 8937 4214
rect 8903 4106 8937 4140
rect 9333 4180 9367 4214
rect 9333 4106 9367 4140
rect 9895 4180 9929 4214
rect 9895 4106 9929 4140
rect 10325 4180 10359 4214
rect 10325 4106 10359 4140
rect 10887 4180 10921 4214
rect 10887 4106 10921 4140
rect 11317 4180 11351 4214
rect 11317 4106 11351 4140
rect 11879 4180 11913 4214
rect 11879 4106 11913 4140
rect 12309 4180 12343 4214
rect 12309 4106 12343 4140
rect 12871 4180 12905 4214
rect 12871 4106 12905 4140
rect 13301 4180 13335 4214
rect 13301 4106 13335 4140
rect 13863 4180 13897 4214
rect 13863 4106 13897 4140
rect 14221 4180 14255 4214
rect 14221 4106 14255 4140
rect 967 2976 1001 3010
rect 967 2898 1001 2932
rect 967 2820 1001 2854
rect 967 2742 1001 2776
rect 967 2663 1001 2697
rect 967 2584 1001 2618
rect 967 2505 1001 2539
rect 1397 2976 1431 3010
rect 1959 2976 1993 3010
rect 1397 2898 1431 2932
rect 1397 2820 1431 2854
rect 1397 2742 1431 2776
rect 1397 2663 1431 2697
rect 1397 2584 1431 2618
rect 1959 2898 1993 2932
rect 1959 2820 1993 2854
rect 1959 2742 1993 2776
rect 1959 2663 1993 2697
rect 1959 2584 1993 2618
rect 1397 2505 1431 2539
rect 1959 2505 1993 2539
rect 2389 2976 2423 3010
rect 2951 2976 2985 3010
rect 2389 2898 2423 2932
rect 2389 2820 2423 2854
rect 2389 2742 2423 2776
rect 2389 2663 2423 2697
rect 2389 2584 2423 2618
rect 2951 2898 2985 2932
rect 2951 2820 2985 2854
rect 2951 2742 2985 2776
rect 2951 2663 2985 2697
rect 2951 2584 2985 2618
rect 2389 2505 2423 2539
rect 2951 2505 2985 2539
rect 3381 2976 3415 3010
rect 3943 2976 3977 3010
rect 3381 2898 3415 2932
rect 3381 2820 3415 2854
rect 3381 2742 3415 2776
rect 3381 2663 3415 2697
rect 3381 2584 3415 2618
rect 3943 2898 3977 2932
rect 3943 2820 3977 2854
rect 3943 2742 3977 2776
rect 3943 2663 3977 2697
rect 3943 2584 3977 2618
rect 3381 2505 3415 2539
rect 3943 2505 3977 2539
rect 4373 2976 4407 3010
rect 4935 2976 4969 3010
rect 4373 2898 4407 2932
rect 4373 2820 4407 2854
rect 4373 2742 4407 2776
rect 4373 2663 4407 2697
rect 4373 2584 4407 2618
rect 4935 2898 4969 2932
rect 4935 2820 4969 2854
rect 4935 2742 4969 2776
rect 4935 2663 4969 2697
rect 4935 2584 4969 2618
rect 4373 2505 4407 2539
rect 4935 2505 4969 2539
rect 5365 2976 5399 3010
rect 5927 2976 5961 3010
rect 5365 2898 5399 2932
rect 5365 2820 5399 2854
rect 5365 2742 5399 2776
rect 5365 2663 5399 2697
rect 5365 2584 5399 2618
rect 5927 2898 5961 2932
rect 5927 2820 5961 2854
rect 5927 2742 5961 2776
rect 5927 2663 5961 2697
rect 5927 2584 5961 2618
rect 5365 2505 5399 2539
rect 5927 2505 5961 2539
rect 6357 2976 6391 3010
rect 6919 2976 6953 3010
rect 6357 2898 6391 2932
rect 6357 2820 6391 2854
rect 6357 2742 6391 2776
rect 6357 2663 6391 2697
rect 6357 2584 6391 2618
rect 6919 2898 6953 2932
rect 6919 2820 6953 2854
rect 6919 2742 6953 2776
rect 6919 2663 6953 2697
rect 6919 2584 6953 2618
rect 6357 2505 6391 2539
rect 6919 2505 6953 2539
rect 7349 2976 7383 3010
rect 7911 2976 7945 3010
rect 7349 2898 7383 2932
rect 7349 2820 7383 2854
rect 7349 2742 7383 2776
rect 7349 2663 7383 2697
rect 7349 2584 7383 2618
rect 7911 2898 7945 2932
rect 7911 2820 7945 2854
rect 7911 2742 7945 2776
rect 7911 2663 7945 2697
rect 7911 2584 7945 2618
rect 7349 2505 7383 2539
rect 7911 2505 7945 2539
rect 8341 2976 8375 3010
rect 8903 2976 8937 3010
rect 8341 2898 8375 2932
rect 8341 2820 8375 2854
rect 8341 2742 8375 2776
rect 8341 2663 8375 2697
rect 8341 2584 8375 2618
rect 8903 2898 8937 2932
rect 8903 2820 8937 2854
rect 8903 2742 8937 2776
rect 8903 2663 8937 2697
rect 8903 2584 8937 2618
rect 8341 2505 8375 2539
rect 8903 2505 8937 2539
rect 9333 2976 9367 3010
rect 9895 2976 9929 3010
rect 9333 2898 9367 2932
rect 9333 2820 9367 2854
rect 9333 2742 9367 2776
rect 9333 2663 9367 2697
rect 9333 2584 9367 2618
rect 9895 2898 9929 2932
rect 9895 2820 9929 2854
rect 9895 2742 9929 2776
rect 9895 2663 9929 2697
rect 9895 2584 9929 2618
rect 9333 2505 9367 2539
rect 9895 2505 9929 2539
rect 10325 2976 10359 3010
rect 10887 2976 10921 3010
rect 10325 2898 10359 2932
rect 10325 2820 10359 2854
rect 10325 2742 10359 2776
rect 10325 2663 10359 2697
rect 10325 2584 10359 2618
rect 10887 2898 10921 2932
rect 10887 2820 10921 2854
rect 10887 2742 10921 2776
rect 10887 2663 10921 2697
rect 10887 2584 10921 2618
rect 10325 2505 10359 2539
rect 10887 2505 10921 2539
rect 11317 2976 11351 3010
rect 11879 2976 11913 3010
rect 11317 2898 11351 2932
rect 11317 2820 11351 2854
rect 11317 2742 11351 2776
rect 11317 2663 11351 2697
rect 11317 2584 11351 2618
rect 11879 2898 11913 2932
rect 11879 2820 11913 2854
rect 11879 2742 11913 2776
rect 11879 2663 11913 2697
rect 11879 2584 11913 2618
rect 11317 2505 11351 2539
rect 11879 2505 11913 2539
rect 12309 2976 12343 3010
rect 12871 2976 12905 3010
rect 12309 2898 12343 2932
rect 12309 2820 12343 2854
rect 12309 2742 12343 2776
rect 12309 2663 12343 2697
rect 12309 2584 12343 2618
rect 12871 2898 12905 2932
rect 12871 2820 12905 2854
rect 12871 2742 12905 2776
rect 12871 2663 12905 2697
rect 12871 2584 12905 2618
rect 12309 2505 12343 2539
rect 12871 2505 12905 2539
rect 13301 2976 13335 3010
rect 13863 2976 13897 3010
rect 13301 2898 13335 2932
rect 13301 2820 13335 2854
rect 13301 2742 13335 2776
rect 13301 2663 13335 2697
rect 13301 2584 13335 2618
rect 13863 2898 13897 2932
rect 13863 2820 13897 2854
rect 13863 2742 13897 2776
rect 13863 2663 13897 2697
rect 13863 2584 13897 2618
rect 13301 2505 13335 2539
rect 13863 2505 13897 2539
rect 14221 2976 14255 3010
rect 14221 2898 14255 2932
rect 14221 2820 14255 2854
rect 14221 2742 14255 2776
rect 14221 2663 14255 2697
rect 14221 2584 14255 2618
rect 14221 2505 14255 2539
rect 967 1375 1001 1409
rect 967 1301 1001 1335
rect 1397 1375 1431 1409
rect 1397 1301 1431 1335
rect 1959 1375 1993 1409
rect 1959 1301 1993 1335
rect 2389 1375 2423 1409
rect 2389 1301 2423 1335
rect 2951 1375 2985 1409
rect 2951 1301 2985 1335
rect 3381 1375 3415 1409
rect 3381 1301 3415 1335
rect 3943 1375 3977 1409
rect 3943 1301 3977 1335
rect 4373 1375 4407 1409
rect 4373 1301 4407 1335
rect 4935 1375 4969 1409
rect 4935 1301 4969 1335
rect 5365 1375 5399 1409
rect 5365 1301 5399 1335
rect 5927 1375 5961 1409
rect 5927 1301 5961 1335
rect 6357 1375 6391 1409
rect 6357 1301 6391 1335
rect 6919 1375 6953 1409
rect 6919 1301 6953 1335
rect 7349 1375 7383 1409
rect 7349 1301 7383 1335
rect 7911 1375 7945 1409
rect 7911 1301 7945 1335
rect 8341 1375 8375 1409
rect 8341 1301 8375 1335
rect 8903 1375 8937 1409
rect 8903 1301 8937 1335
rect 9333 1375 9367 1409
rect 9333 1301 9367 1335
rect 9895 1375 9929 1409
rect 9895 1301 9929 1335
rect 10325 1375 10359 1409
rect 10325 1301 10359 1335
rect 10887 1375 10921 1409
rect 10887 1301 10921 1335
rect 11317 1375 11351 1409
rect 11317 1301 11351 1335
rect 11879 1375 11913 1409
rect 11879 1301 11913 1335
rect 12309 1375 12343 1409
rect 12309 1301 12343 1335
rect 12871 1375 12905 1409
rect 12871 1301 12905 1335
rect 13301 1375 13335 1409
rect 13301 1301 13335 1335
rect 13863 1375 13897 1409
rect 13863 1301 13897 1335
rect 14221 1375 14255 1409
rect 14221 1301 14255 1335
<< locali >>
rect 233 5425 305 5459
rect 339 5425 377 5459
rect 411 5425 449 5459
rect 483 5425 521 5459
rect 555 5425 593 5459
rect 627 5425 665 5459
rect 699 5425 737 5459
rect 771 5425 809 5459
rect 843 5425 881 5459
rect 915 5425 953 5459
rect 987 5425 1025 5459
rect 1059 5425 1097 5459
rect 1131 5425 1169 5459
rect 1203 5425 1241 5459
rect 1275 5425 1313 5459
rect 1347 5425 1385 5459
rect 1419 5425 1457 5459
rect 1491 5425 1529 5459
rect 1563 5425 1601 5459
rect 1635 5425 1673 5459
rect 1707 5425 1745 5459
rect 1779 5425 1817 5459
rect 1851 5425 1889 5459
rect 1923 5425 1961 5459
rect 1995 5425 2033 5459
rect 2067 5425 2105 5459
rect 2139 5425 2177 5459
rect 2211 5425 2249 5459
rect 2283 5425 2321 5459
rect 2355 5425 2393 5459
rect 2427 5425 2465 5459
rect 2499 5425 2537 5459
rect 2571 5425 2609 5459
rect 2643 5425 2681 5459
rect 2715 5425 2753 5459
rect 2787 5425 2825 5459
rect 2859 5425 2897 5459
rect 2931 5425 2969 5459
rect 3003 5425 3041 5459
rect 3075 5425 3113 5459
rect 3147 5425 3185 5459
rect 3219 5425 3257 5459
rect 3291 5425 3329 5459
rect 3363 5425 3401 5459
rect 3435 5425 3473 5459
rect 3507 5425 3545 5459
rect 3579 5425 3617 5459
rect 3651 5425 3689 5459
rect 3723 5425 3761 5459
rect 3795 5425 3833 5459
rect 3867 5425 3905 5459
rect 3939 5425 3977 5459
rect 4011 5425 4049 5459
rect 4083 5425 4121 5459
rect 4155 5425 4193 5459
rect 4227 5425 4265 5459
rect 4299 5425 4337 5459
rect 4371 5425 4409 5459
rect 4443 5425 4481 5459
rect 4515 5425 4553 5459
rect 4587 5425 4625 5459
rect 4659 5425 4697 5459
rect 4731 5425 4769 5459
rect 4803 5425 4841 5459
rect 4875 5425 4913 5459
rect 4947 5425 4985 5459
rect 5019 5425 5057 5459
rect 5091 5425 5129 5459
rect 5163 5425 5201 5459
rect 5235 5425 5273 5459
rect 5307 5425 5345 5459
rect 5379 5425 5417 5459
rect 5451 5425 5489 5459
rect 5523 5425 5561 5459
rect 5595 5425 5633 5459
rect 5667 5425 5705 5459
rect 5739 5425 5777 5459
rect 5811 5425 5849 5459
rect 5883 5425 5921 5459
rect 5955 5425 5993 5459
rect 6027 5425 6065 5459
rect 6099 5425 6137 5459
rect 6171 5425 6209 5459
rect 6243 5425 6281 5459
rect 6315 5425 6353 5459
rect 6387 5425 6425 5459
rect 6459 5425 6497 5459
rect 6531 5425 6569 5459
rect 6603 5425 6641 5459
rect 6675 5425 6713 5459
rect 6747 5425 6785 5459
rect 6819 5425 6857 5459
rect 6891 5425 6929 5459
rect 6963 5425 7001 5459
rect 7035 5425 7073 5459
rect 7107 5425 7145 5459
rect 7179 5425 7217 5459
rect 7251 5425 7289 5459
rect 7323 5425 7361 5459
rect 7395 5425 7433 5459
rect 7467 5425 7505 5459
rect 7539 5425 7577 5459
rect 7611 5425 7649 5459
rect 7683 5425 7721 5459
rect 7755 5425 7793 5459
rect 7827 5425 7865 5459
rect 7899 5425 7937 5459
rect 7971 5425 8009 5459
rect 8043 5425 8081 5459
rect 8115 5425 8153 5459
rect 8187 5425 8225 5459
rect 8259 5425 8297 5459
rect 8331 5425 8369 5459
rect 8403 5425 8441 5459
rect 8475 5425 8513 5459
rect 8547 5425 8585 5459
rect 8619 5425 8657 5459
rect 8691 5425 8729 5459
rect 8763 5425 8801 5459
rect 8835 5425 8873 5459
rect 8907 5425 8945 5459
rect 8979 5425 9017 5459
rect 9051 5425 9089 5459
rect 9123 5425 9161 5459
rect 9195 5425 9233 5459
rect 9267 5425 9305 5459
rect 9339 5425 9377 5459
rect 9411 5425 9449 5459
rect 9483 5425 9521 5459
rect 9555 5425 9593 5459
rect 9627 5425 9665 5459
rect 9699 5425 9737 5459
rect 9771 5425 9809 5459
rect 9843 5425 9881 5459
rect 9915 5425 9953 5459
rect 9987 5425 10025 5459
rect 10059 5425 10097 5459
rect 10131 5425 10169 5459
rect 10203 5425 10241 5459
rect 10275 5425 10313 5459
rect 10347 5425 10385 5459
rect 10419 5425 10457 5459
rect 10491 5425 10529 5459
rect 10563 5425 10601 5459
rect 10635 5425 10673 5459
rect 10707 5425 10745 5459
rect 10779 5425 10817 5459
rect 10851 5425 10889 5459
rect 10923 5425 10961 5459
rect 10995 5425 11033 5459
rect 11067 5425 11105 5459
rect 11139 5425 11177 5459
rect 11211 5425 11249 5459
rect 11283 5425 11321 5459
rect 11355 5425 11393 5459
rect 11427 5425 11466 5459
rect 11500 5425 11539 5459
rect 11573 5425 11612 5459
rect 11646 5425 11685 5459
rect 11719 5425 11758 5459
rect 11792 5425 11831 5459
rect 11865 5425 11904 5459
rect 11938 5425 11977 5459
rect 12011 5425 12050 5459
rect 12084 5425 12123 5459
rect 12157 5425 12196 5459
rect 12230 5425 12269 5459
rect 12303 5425 12342 5459
rect 12376 5425 12415 5459
rect 12449 5425 12488 5459
rect 12522 5425 12561 5459
rect 12595 5425 12634 5459
rect 12668 5425 12707 5459
rect 12741 5425 12780 5459
rect 12814 5425 12853 5459
rect 12887 5425 12926 5459
rect 12960 5425 12999 5459
rect 13033 5425 13072 5459
rect 13106 5425 13145 5459
rect 13179 5425 13218 5459
rect 13252 5425 13291 5459
rect 13325 5425 13364 5459
rect 13398 5425 13437 5459
rect 13471 5425 13510 5459
rect 13544 5425 13583 5459
rect 13617 5425 13656 5459
rect 13690 5425 13729 5459
rect 13763 5425 13802 5459
rect 13836 5425 13875 5459
rect 13909 5425 13948 5459
rect 13982 5425 14021 5459
rect 14055 5425 14094 5459
rect 14128 5425 14167 5459
rect 14201 5425 14240 5459
rect 14274 5425 14313 5459
rect 14347 5425 14386 5459
rect 14420 5425 14459 5459
rect 14493 5425 14532 5459
rect 14566 5425 14605 5459
rect 14639 5425 14678 5459
rect 14712 5425 14751 5459
rect 14785 5425 14824 5459
rect 14858 5425 14897 5459
rect 14931 5425 15003 5459
rect 233 5422 15003 5425
rect 232 5388 300 5422
rect 334 5388 369 5422
rect 403 5388 438 5422
rect 472 5388 507 5422
rect 541 5388 576 5422
rect 610 5388 645 5422
rect 679 5388 714 5422
rect 748 5388 783 5422
rect 817 5388 852 5422
rect 886 5388 921 5422
rect 955 5388 990 5422
rect 1024 5388 1059 5422
rect 1093 5388 1128 5422
rect 1162 5388 1197 5422
rect 1231 5388 1266 5422
rect 1300 5388 1335 5422
rect 1369 5388 1404 5422
rect 1438 5388 1473 5422
rect 1507 5388 1542 5422
rect 1576 5388 1611 5422
rect 1645 5388 1680 5422
rect 1714 5388 1749 5422
rect 1783 5388 1818 5422
rect 1852 5388 1887 5422
rect 1921 5388 1956 5422
rect 1990 5388 2025 5422
rect 2059 5388 2094 5422
rect 2128 5388 2163 5422
rect 2197 5388 2232 5422
rect 232 5387 2232 5388
rect 232 5354 233 5387
rect 267 5354 2232 5387
rect 334 5289 369 5354
rect 403 5320 438 5354
rect 472 5323 507 5354
rect 541 5323 576 5354
rect 610 5323 645 5354
rect 679 5323 714 5354
rect 748 5323 783 5354
rect 817 5323 852 5354
rect 886 5323 921 5354
rect 955 5323 990 5354
rect 1024 5323 1059 5354
rect 1093 5323 1128 5354
rect 1162 5323 1197 5354
rect 475 5320 507 5323
rect 547 5320 576 5323
rect 619 5320 645 5323
rect 691 5320 714 5323
rect 763 5320 783 5323
rect 835 5320 852 5323
rect 907 5320 921 5323
rect 979 5320 990 5323
rect 1051 5320 1059 5323
rect 1123 5320 1128 5323
rect 1195 5320 1197 5323
rect 1231 5323 1266 5354
rect 1300 5323 1335 5354
rect 1369 5323 1404 5354
rect 1438 5323 1473 5354
rect 1507 5323 1542 5354
rect 1576 5323 1611 5354
rect 1645 5323 1680 5354
rect 1714 5323 1749 5354
rect 1783 5323 1818 5354
rect 1852 5323 1887 5354
rect 1921 5323 1956 5354
rect 1231 5320 1233 5323
rect 1300 5320 1305 5323
rect 1369 5320 1377 5323
rect 1438 5320 1449 5323
rect 1507 5320 1521 5323
rect 1576 5320 1593 5323
rect 1645 5320 1665 5323
rect 1714 5320 1737 5323
rect 1783 5320 1809 5323
rect 1852 5320 1881 5323
rect 1921 5320 1953 5323
rect 1990 5320 2025 5354
rect 2059 5320 2094 5354
rect 2128 5323 2163 5354
rect 2197 5323 2232 5354
rect 14914 5387 15003 5422
rect 14914 5353 14969 5387
rect 2131 5320 2163 5323
rect 2203 5320 2232 5323
rect 403 5289 441 5320
rect 475 5289 513 5320
rect 547 5289 585 5320
rect 619 5289 657 5320
rect 691 5289 729 5320
rect 763 5289 801 5320
rect 835 5289 873 5320
rect 907 5289 945 5320
rect 979 5289 1017 5320
rect 1051 5289 1089 5320
rect 1123 5289 1161 5320
rect 1195 5289 1233 5320
rect 1267 5289 1305 5320
rect 1339 5289 1377 5320
rect 1411 5289 1449 5320
rect 1483 5289 1521 5320
rect 1555 5289 1593 5320
rect 1627 5289 1665 5320
rect 1699 5289 1737 5320
rect 1771 5289 1809 5320
rect 1843 5289 1881 5320
rect 1915 5289 1953 5320
rect 1987 5289 2025 5320
rect 2059 5289 2097 5320
rect 2131 5289 2169 5320
rect 2203 5289 2241 5320
rect 2275 5289 2300 5320
rect 14914 5315 15003 5353
rect 334 5286 2300 5289
rect 402 5252 437 5286
rect 471 5252 506 5286
rect 540 5252 575 5286
rect 609 5252 644 5286
rect 678 5252 713 5286
rect 747 5252 782 5286
rect 816 5252 851 5286
rect 885 5252 920 5286
rect 954 5252 989 5286
rect 1023 5252 1058 5286
rect 1092 5252 1127 5286
rect 1161 5252 1196 5286
rect 1230 5252 1265 5286
rect 1299 5252 1334 5286
rect 1368 5252 1403 5286
rect 1437 5252 1472 5286
rect 1506 5252 1541 5286
rect 1575 5252 1610 5286
rect 1644 5252 1679 5286
rect 1713 5252 1748 5286
rect 1782 5252 1817 5286
rect 1851 5252 1886 5286
rect 1920 5252 1955 5286
rect 1989 5252 2024 5286
rect 2058 5252 2093 5286
rect 2127 5252 2162 5286
rect 2196 5252 2231 5286
rect 2265 5252 2300 5286
rect 14914 5281 14969 5315
rect 402 5250 403 5252
rect 402 5177 403 5216
rect 402 5104 403 5143
rect 402 5031 403 5070
rect 402 4958 403 4997
rect 14914 5243 15003 5281
rect 14914 5218 14969 5243
rect 14990 5171 15003 5209
rect 14990 5099 15003 5137
rect 14990 5027 15003 5065
rect 402 4885 403 4924
rect 402 4812 403 4851
rect 402 4739 403 4778
rect 402 4666 403 4705
rect 402 4593 403 4632
rect 402 4520 403 4559
rect 402 4447 403 4486
rect 402 4374 403 4413
rect 402 4301 403 4340
rect 402 4228 403 4267
rect 402 4155 403 4194
rect 402 4082 403 4121
rect 402 4009 403 4048
rect 402 3936 403 3975
rect 402 3863 403 3902
rect 402 3790 403 3829
rect 402 3717 403 3756
rect 402 3644 403 3683
rect 402 3571 403 3610
rect 402 3498 403 3537
rect 402 3425 403 3464
rect 402 3352 403 3391
rect 402 3279 403 3318
rect 402 3206 403 3245
rect 402 3133 403 3172
rect 402 3060 403 3099
rect 402 2987 403 3026
rect 402 2914 403 2953
rect 402 2841 403 2880
rect 402 2768 403 2807
rect 402 2695 403 2734
rect 402 2622 403 2661
rect 402 2549 403 2588
rect 402 2476 403 2515
rect 402 2403 403 2442
rect 402 2330 403 2369
rect 402 2257 403 2296
rect 402 2184 403 2223
rect 402 2111 403 2150
rect 402 2038 403 2077
rect 402 1965 403 2004
rect 402 1892 403 1931
rect 402 1819 403 1858
rect 402 1746 403 1785
rect 402 1673 403 1712
rect 402 1600 403 1639
rect 402 1527 403 1566
rect 402 1454 403 1493
rect 402 1381 403 1420
rect 402 1308 403 1347
rect 402 1235 403 1274
rect 402 1162 403 1201
rect 402 1089 403 1128
rect 402 1016 403 1055
rect 402 944 403 982
rect 555 4922 657 4956
rect 589 4888 657 4922
rect 555 4854 623 4888
rect 555 4850 691 4854
rect 589 4819 691 4850
rect 589 4816 623 4819
rect 555 4785 623 4816
rect 657 4786 691 4819
rect 14495 4922 14530 4956
rect 14564 4922 14599 4956
rect 14633 4922 14667 4956
rect 14461 4888 14667 4922
rect 14461 4854 14496 4888
rect 14530 4854 14565 4888
rect 14599 4854 14667 4888
rect 14393 4852 14667 4854
rect 14393 4818 14402 4852
rect 14436 4844 14667 4852
rect 14436 4820 14633 4844
rect 14393 4786 14428 4818
rect 14462 4786 14497 4820
rect 14531 4818 14633 4820
rect 14531 4786 14565 4818
rect 657 4785 822 4786
rect 555 4778 822 4785
rect 589 4774 822 4778
rect 589 4751 733 4774
rect 589 4750 691 4751
rect 589 4744 623 4750
rect 555 4710 587 4744
rect 621 4716 623 4744
rect 657 4744 691 4750
rect 657 4716 659 4744
rect 725 4740 733 4751
rect 767 4740 822 4774
rect 725 4717 822 4740
rect 621 4710 659 4716
rect 693 4710 822 4717
rect 555 4706 822 4710
rect 589 4701 822 4706
rect 589 4682 733 4701
rect 589 4681 691 4682
rect 589 4672 623 4681
rect 555 4670 623 4672
rect 555 4636 587 4670
rect 621 4647 623 4670
rect 657 4670 691 4681
rect 657 4647 659 4670
rect 725 4667 733 4682
rect 767 4667 822 4701
rect 725 4648 822 4667
rect 621 4636 659 4647
rect 693 4636 822 4648
rect 555 4634 822 4636
rect 589 4628 822 4634
rect 589 4613 733 4628
rect 589 4600 623 4613
rect 555 4596 623 4600
rect 555 4563 587 4596
rect 621 4562 623 4596
rect 725 4594 733 4613
rect 767 4594 822 4628
rect 589 4529 623 4562
rect 555 4522 623 4529
rect 725 4555 822 4594
rect 555 4492 587 4522
rect 621 4488 623 4522
rect 725 4521 733 4555
rect 767 4521 822 4555
rect 589 4458 623 4488
rect 555 4449 623 4458
rect 725 4482 822 4521
rect 14400 4784 14565 4786
rect 14599 4810 14633 4818
rect 14599 4784 14667 4810
rect 14400 4774 14667 4784
rect 14400 4740 14431 4774
rect 14465 4771 14667 4774
rect 14465 4750 14633 4771
rect 14465 4740 14497 4750
rect 14531 4748 14633 4750
rect 14531 4743 14565 4748
rect 14599 4743 14633 4748
rect 14400 4716 14497 4740
rect 14400 4709 14510 4716
rect 14544 4714 14565 4743
rect 14616 4737 14633 4743
rect 14544 4709 14582 4714
rect 14616 4709 14667 4737
rect 14400 4701 14667 4709
rect 14400 4667 14431 4701
rect 14465 4698 14667 4701
rect 14465 4680 14633 4698
rect 14465 4667 14497 4680
rect 14531 4678 14633 4680
rect 14531 4670 14565 4678
rect 14599 4670 14633 4678
rect 14400 4646 14497 4667
rect 14400 4636 14510 4646
rect 14544 4644 14565 4670
rect 14616 4664 14633 4670
rect 14544 4636 14582 4644
rect 14616 4636 14667 4664
rect 14400 4628 14667 4636
rect 14400 4594 14431 4628
rect 14465 4625 14667 4628
rect 14465 4610 14633 4625
rect 14465 4594 14497 4610
rect 14531 4608 14633 4610
rect 14531 4597 14565 4608
rect 14599 4597 14633 4608
rect 14400 4576 14497 4594
rect 14400 4563 14510 4576
rect 14544 4574 14565 4597
rect 14616 4591 14633 4597
rect 14544 4563 14582 4574
rect 14616 4563 14667 4591
rect 14400 4555 14667 4563
rect 14400 4521 14431 4555
rect 14465 4552 14667 4555
rect 14465 4540 14633 4552
rect 14465 4521 14497 4540
rect 14531 4538 14633 4540
rect 14531 4524 14565 4538
rect 14599 4524 14633 4538
rect 14400 4506 14497 4521
rect 555 4421 587 4449
rect 621 4415 623 4449
rect 725 4448 733 4482
rect 767 4448 822 4482
rect 589 4387 623 4415
rect 555 4376 623 4387
rect 725 4409 822 4448
rect 555 4350 587 4376
rect 621 4342 623 4376
rect 725 4375 733 4409
rect 767 4375 822 4409
rect 589 4316 623 4342
rect 555 4303 623 4316
rect 725 4336 822 4375
rect 555 4279 587 4303
rect 621 4269 623 4303
rect 725 4302 733 4336
rect 767 4302 822 4336
rect 589 4245 623 4269
rect 555 4230 623 4245
rect 725 4263 822 4302
rect 555 4208 587 4230
rect 621 4196 623 4230
rect 725 4229 733 4263
rect 767 4229 822 4263
rect 589 4174 623 4196
rect 555 4157 623 4174
rect 725 4190 822 4229
rect 555 4137 587 4157
rect 621 4123 623 4157
rect 725 4156 733 4190
rect 767 4156 822 4190
rect 589 4103 623 4123
rect 725 4117 822 4156
rect 725 4103 733 4117
rect 555 4084 733 4103
rect 555 4050 587 4084
rect 621 4050 659 4084
rect 693 4083 733 4084
rect 767 4083 822 4117
rect 693 4062 822 4083
rect 924 4388 931 4494
rect 1037 4388 1044 4494
rect 924 4214 1044 4388
rect 924 4180 967 4214
rect 1001 4180 1044 4214
rect 924 4140 1044 4180
rect 924 4106 967 4140
rect 1001 4106 1044 4140
rect 693 4050 836 4062
rect 555 4046 836 4050
rect 555 4044 802 4046
rect 555 4041 733 4044
rect 589 4011 623 4041
rect 621 4007 623 4011
rect 657 4011 733 4041
rect 767 4034 802 4044
rect 657 4007 659 4011
rect 555 3977 587 4007
rect 621 3977 659 4007
rect 693 4010 733 4011
rect 768 4012 802 4034
rect 693 4000 734 4010
rect 768 4000 836 4012
rect 693 3978 836 4000
rect 693 3977 802 3978
rect 555 3971 802 3977
rect 555 3970 733 3971
rect 589 3938 623 3970
rect 621 3936 623 3938
rect 657 3938 733 3970
rect 767 3966 802 3971
rect 657 3936 659 3938
rect 555 3904 587 3936
rect 621 3904 659 3936
rect 693 3937 733 3938
rect 768 3944 802 3966
rect 693 3932 734 3937
rect 768 3932 836 3944
rect 693 3910 836 3932
rect 693 3904 802 3910
rect 555 3898 802 3904
rect 555 3896 733 3898
rect 589 3865 623 3896
rect 621 3862 623 3865
rect 657 3865 733 3896
rect 657 3862 659 3865
rect 555 3831 587 3862
rect 621 3831 659 3862
rect 693 3864 733 3865
rect 768 3876 802 3898
rect 768 3864 836 3876
rect 693 3842 836 3864
rect 693 3831 802 3842
rect 555 3830 802 3831
rect 555 3825 734 3830
rect 589 3792 623 3825
rect 621 3791 623 3792
rect 657 3792 733 3825
rect 768 3808 802 3830
rect 768 3796 836 3808
rect 657 3791 659 3792
rect 555 3758 587 3791
rect 621 3758 659 3791
rect 693 3791 733 3792
rect 767 3791 836 3796
rect 693 3774 836 3791
rect 693 3762 802 3774
rect 693 3758 734 3762
rect 555 3752 734 3758
rect 555 3751 733 3752
rect 589 3719 623 3751
rect 621 3717 623 3719
rect 657 3719 733 3751
rect 768 3740 802 3762
rect 768 3728 836 3740
rect 657 3717 659 3719
rect 555 3685 587 3717
rect 621 3685 659 3717
rect 693 3718 733 3719
rect 767 3718 836 3728
rect 693 3706 836 3718
rect 693 3694 802 3706
rect 693 3685 734 3694
rect 555 3680 734 3685
rect 589 3646 623 3680
rect 657 3679 734 3680
rect 657 3646 733 3679
rect 768 3672 802 3694
rect 768 3660 836 3672
rect 555 3612 587 3646
rect 621 3612 659 3646
rect 693 3645 733 3646
rect 767 3645 836 3660
rect 693 3638 836 3645
rect 693 3626 802 3638
rect 693 3612 734 3626
rect 555 3606 734 3612
rect 589 3573 623 3606
rect 621 3572 623 3573
rect 657 3573 733 3606
rect 768 3604 802 3626
rect 768 3592 836 3604
rect 657 3572 659 3573
rect 555 3539 587 3572
rect 621 3539 659 3572
rect 693 3572 733 3573
rect 767 3572 836 3592
rect 693 3570 836 3572
rect 693 3558 802 3570
rect 693 3539 734 3558
rect 555 3535 734 3539
rect 589 3501 623 3535
rect 657 3533 734 3535
rect 768 3536 802 3558
rect 657 3501 733 3533
rect 768 3524 836 3536
rect 555 3500 733 3501
rect 555 3466 587 3500
rect 621 3466 659 3500
rect 693 3499 733 3500
rect 767 3502 836 3524
rect 767 3499 802 3502
rect 693 3490 802 3499
rect 693 3466 734 3490
rect 555 3461 734 3466
rect 589 3427 623 3461
rect 657 3460 734 3461
rect 768 3468 802 3490
rect 657 3427 733 3460
rect 768 3456 836 3468
rect 555 3393 587 3427
rect 621 3393 659 3427
rect 693 3426 733 3427
rect 767 3434 836 3456
rect 767 3426 802 3434
rect 693 3422 802 3426
rect 693 3393 734 3422
rect 555 3390 734 3393
rect 589 3356 623 3390
rect 657 3388 734 3390
rect 768 3400 802 3422
rect 768 3388 836 3400
rect 657 3387 836 3388
rect 657 3356 733 3387
rect 555 3354 733 3356
rect 767 3366 836 3387
rect 767 3354 802 3366
rect 555 3320 587 3354
rect 621 3320 659 3354
rect 693 3353 733 3354
rect 693 3320 734 3353
rect 768 3332 802 3354
rect 768 3320 836 3332
rect 555 3316 836 3320
rect 589 3282 623 3316
rect 657 3314 836 3316
rect 657 3282 733 3314
rect 767 3298 836 3314
rect 767 3286 802 3298
rect 555 3281 733 3282
rect 555 3247 587 3281
rect 621 3247 659 3281
rect 693 3280 733 3281
rect 693 3252 734 3280
rect 768 3264 802 3286
rect 768 3252 836 3264
rect 693 3247 836 3252
rect 555 3245 836 3247
rect 589 3211 623 3245
rect 657 3241 836 3245
rect 657 3211 733 3241
rect 767 3230 836 3241
rect 767 3218 802 3230
rect 555 3208 733 3211
rect 555 3174 587 3208
rect 621 3174 659 3208
rect 693 3207 733 3208
rect 693 3184 734 3207
rect 768 3196 802 3218
rect 768 3184 836 3196
rect 693 3174 836 3184
rect 555 3168 836 3174
rect 555 3151 733 3168
rect 589 3135 623 3151
rect 621 3117 623 3135
rect 657 3135 733 3151
rect 767 3162 836 3168
rect 767 3150 802 3162
rect 657 3117 659 3135
rect 555 3101 587 3117
rect 621 3101 659 3117
rect 693 3134 733 3135
rect 693 3116 734 3134
rect 768 3128 802 3150
rect 768 3116 836 3128
rect 693 3101 836 3116
rect 555 3100 836 3101
rect 555 3095 822 3100
rect 555 3081 733 3095
rect 657 3062 733 3081
rect 657 3028 659 3062
rect 693 3061 733 3062
rect 767 3061 822 3095
rect 693 3028 822 3061
rect 657 3022 822 3028
rect 657 3013 733 3022
rect 725 2988 733 3013
rect 767 2988 822 3022
rect 725 2949 822 2988
rect 725 2915 733 2949
rect 767 2915 822 2949
rect 725 2876 822 2915
rect 725 2842 733 2876
rect 767 2842 822 2876
rect 725 2803 822 2842
rect 725 2769 733 2803
rect 767 2769 822 2803
rect 725 2730 822 2769
rect 725 2696 733 2730
rect 767 2696 822 2730
rect 725 2657 822 2696
rect 725 2623 733 2657
rect 767 2623 822 2657
rect 725 2584 822 2623
rect 725 2550 733 2584
rect 767 2550 822 2584
rect 725 2511 822 2550
rect 725 2503 733 2511
rect 657 2478 733 2503
rect 657 2444 659 2478
rect 693 2477 733 2478
rect 767 2477 822 2511
rect 693 2461 822 2477
rect 924 3010 1044 4106
rect 1354 4388 1361 4494
rect 1467 4388 1474 4494
rect 1354 4214 1474 4388
rect 1354 4180 1397 4214
rect 1431 4180 1474 4214
rect 1354 4140 1474 4180
rect 1354 4106 1397 4140
rect 1431 4106 1474 4140
rect 924 2976 967 3010
rect 1001 2976 1044 3010
rect 924 2932 1044 2976
rect 924 2898 967 2932
rect 1001 2898 1044 2932
rect 924 2854 1044 2898
rect 924 2820 967 2854
rect 1001 2820 1044 2854
rect 924 2776 1044 2820
rect 924 2742 967 2776
rect 1001 2742 1044 2776
rect 924 2697 1044 2742
rect 924 2663 967 2697
rect 1001 2663 1044 2697
rect 924 2618 1044 2663
rect 924 2584 967 2618
rect 1001 2584 1044 2618
rect 924 2539 1044 2584
rect 924 2505 967 2539
rect 1001 2505 1044 2539
rect 693 2445 836 2461
rect 693 2444 802 2445
rect 657 2438 802 2444
rect 657 2405 733 2438
rect 767 2433 802 2438
rect 657 2371 659 2405
rect 693 2404 733 2405
rect 768 2411 802 2433
rect 693 2399 734 2404
rect 768 2399 836 2411
rect 693 2377 836 2399
rect 693 2371 802 2377
rect 657 2367 802 2371
rect 555 2365 802 2367
rect 555 2332 733 2365
rect 555 2327 587 2332
rect 621 2327 659 2332
rect 621 2298 623 2327
rect 589 2293 623 2298
rect 657 2298 659 2327
rect 693 2331 733 2332
rect 768 2343 802 2365
rect 768 2331 836 2343
rect 693 2309 836 2331
rect 693 2298 802 2309
rect 657 2297 802 2298
rect 657 2293 734 2297
rect 555 2292 734 2293
rect 555 2259 733 2292
rect 768 2275 802 2297
rect 768 2263 836 2275
rect 555 2250 587 2259
rect 621 2250 659 2259
rect 621 2225 623 2250
rect 589 2216 623 2225
rect 657 2225 659 2250
rect 693 2258 733 2259
rect 767 2258 836 2263
rect 693 2241 836 2258
rect 693 2229 802 2241
rect 693 2225 734 2229
rect 657 2219 734 2225
rect 657 2216 733 2219
rect 555 2186 733 2216
rect 768 2207 802 2229
rect 768 2195 836 2207
rect 555 2156 587 2186
rect 621 2156 659 2186
rect 621 2152 623 2156
rect 589 2122 623 2152
rect 657 2152 659 2156
rect 693 2185 733 2186
rect 767 2185 836 2195
rect 693 2173 836 2185
rect 693 2161 802 2173
rect 693 2152 734 2161
rect 657 2146 734 2152
rect 657 2122 733 2146
rect 768 2139 802 2161
rect 768 2127 836 2139
rect 555 2113 733 2122
rect 555 2085 587 2113
rect 621 2085 659 2113
rect 621 2079 623 2085
rect 589 2051 623 2079
rect 657 2079 659 2085
rect 693 2112 733 2113
rect 767 2112 836 2127
rect 693 2105 836 2112
rect 693 2093 802 2105
rect 693 2079 734 2093
rect 657 2073 734 2079
rect 657 2051 733 2073
rect 768 2071 802 2093
rect 768 2059 836 2071
rect 555 2040 733 2051
rect 555 2011 587 2040
rect 621 2011 659 2040
rect 621 2006 623 2011
rect 589 1977 623 2006
rect 657 2006 659 2011
rect 693 2039 733 2040
rect 767 2039 836 2059
rect 693 2037 836 2039
rect 693 2025 802 2037
rect 693 2006 734 2025
rect 657 2000 734 2006
rect 768 2003 802 2025
rect 657 1977 733 2000
rect 768 1991 836 2003
rect 555 1967 733 1977
rect 555 1940 587 1967
rect 621 1940 659 1967
rect 621 1933 623 1940
rect 589 1906 623 1933
rect 657 1933 659 1940
rect 693 1966 733 1967
rect 767 1969 836 1991
rect 767 1966 802 1969
rect 693 1957 802 1966
rect 693 1933 734 1957
rect 657 1927 734 1933
rect 768 1935 802 1957
rect 657 1906 733 1927
rect 768 1923 836 1935
rect 555 1894 733 1906
rect 555 1866 587 1894
rect 621 1866 659 1894
rect 621 1860 623 1866
rect 589 1832 623 1860
rect 657 1860 659 1866
rect 693 1893 733 1894
rect 767 1901 836 1923
rect 767 1893 802 1901
rect 693 1889 802 1893
rect 693 1860 734 1889
rect 657 1855 734 1860
rect 768 1867 802 1889
rect 768 1855 836 1867
rect 657 1854 836 1855
rect 657 1832 733 1854
rect 555 1821 733 1832
rect 767 1833 836 1854
rect 767 1821 802 1833
rect 555 1795 587 1821
rect 621 1795 659 1821
rect 621 1787 623 1795
rect 589 1761 623 1787
rect 657 1787 659 1795
rect 693 1820 733 1821
rect 693 1787 734 1820
rect 768 1799 802 1821
rect 768 1787 836 1799
rect 657 1781 836 1787
rect 657 1761 733 1781
rect 555 1748 733 1761
rect 767 1765 836 1781
rect 767 1753 802 1765
rect 555 1721 587 1748
rect 621 1721 659 1748
rect 621 1714 623 1721
rect 589 1687 623 1714
rect 657 1714 659 1721
rect 693 1747 733 1748
rect 693 1719 734 1747
rect 768 1731 802 1753
rect 768 1719 836 1731
rect 693 1714 836 1719
rect 657 1708 836 1714
rect 657 1687 733 1708
rect 555 1675 733 1687
rect 767 1697 836 1708
rect 767 1685 802 1697
rect 555 1650 587 1675
rect 621 1650 659 1675
rect 621 1641 623 1650
rect 589 1616 623 1641
rect 657 1641 659 1650
rect 693 1674 733 1675
rect 693 1651 734 1674
rect 768 1663 802 1685
rect 768 1651 836 1663
rect 693 1641 836 1651
rect 657 1635 836 1641
rect 657 1616 733 1635
rect 767 1629 836 1635
rect 767 1617 802 1629
rect 555 1602 733 1616
rect 555 1576 587 1602
rect 621 1576 659 1602
rect 621 1568 623 1576
rect 589 1542 623 1568
rect 657 1568 659 1576
rect 693 1601 733 1602
rect 693 1583 734 1601
rect 768 1595 802 1617
rect 768 1583 836 1595
rect 693 1568 836 1583
rect 657 1562 836 1568
rect 657 1542 733 1562
rect 767 1561 836 1562
rect 767 1549 802 1561
rect 555 1529 733 1542
rect 555 1505 587 1529
rect 621 1505 659 1529
rect 621 1495 623 1505
rect 589 1471 623 1495
rect 657 1495 659 1505
rect 693 1528 733 1529
rect 693 1515 734 1528
rect 768 1527 802 1549
rect 768 1515 836 1527
rect 693 1499 836 1515
rect 693 1495 822 1499
rect 657 1489 822 1495
rect 657 1471 733 1489
rect 555 1455 733 1471
rect 767 1455 822 1489
rect 555 1419 822 1455
rect 555 1385 587 1419
rect 621 1385 659 1419
rect 693 1416 822 1419
rect 693 1385 733 1416
rect 555 1382 733 1385
rect 767 1382 822 1416
rect 555 1375 822 1382
rect 589 1341 623 1375
rect 657 1341 691 1375
rect 725 1342 822 1375
rect 725 1341 733 1342
rect 555 1330 733 1341
rect 555 1296 587 1330
rect 621 1296 659 1330
rect 693 1308 733 1330
rect 767 1308 822 1342
rect 693 1296 822 1308
rect 555 1268 822 1296
rect 924 1409 1044 2505
rect 1109 4028 1110 4062
rect 1144 4046 1182 4062
rect 1144 4028 1146 4046
rect 1109 4012 1146 4028
rect 1180 4028 1182 4046
rect 1216 4046 1254 4062
rect 1216 4028 1218 4046
rect 1180 4012 1218 4028
rect 1252 4028 1254 4046
rect 1288 4028 1289 4062
rect 1252 4012 1289 4028
rect 1109 3988 1289 4012
rect 1109 3954 1110 3988
rect 1144 3978 1182 3988
rect 1144 3954 1146 3978
rect 1109 3944 1146 3954
rect 1180 3954 1182 3978
rect 1216 3978 1254 3988
rect 1216 3954 1218 3978
rect 1180 3944 1218 3954
rect 1252 3954 1254 3978
rect 1288 3954 1289 3988
rect 1252 3944 1289 3954
rect 1109 3914 1289 3944
rect 1109 3880 1110 3914
rect 1144 3910 1182 3914
rect 1144 3880 1146 3910
rect 1109 3876 1146 3880
rect 1180 3880 1182 3910
rect 1216 3910 1254 3914
rect 1216 3880 1218 3910
rect 1180 3876 1218 3880
rect 1252 3880 1254 3910
rect 1288 3880 1289 3914
rect 1252 3876 1289 3880
rect 1109 3842 1289 3876
rect 1109 3840 1146 3842
rect 1109 3806 1110 3840
rect 1144 3808 1146 3840
rect 1180 3840 1218 3842
rect 1180 3808 1182 3840
rect 1144 3806 1182 3808
rect 1216 3808 1218 3840
rect 1252 3840 1289 3842
rect 1252 3808 1254 3840
rect 1216 3806 1254 3808
rect 1288 3806 1289 3840
rect 1109 3774 1289 3806
rect 1109 3766 1146 3774
rect 1109 3732 1110 3766
rect 1144 3740 1146 3766
rect 1180 3766 1218 3774
rect 1180 3740 1182 3766
rect 1144 3732 1182 3740
rect 1216 3740 1218 3766
rect 1252 3766 1289 3774
rect 1252 3740 1254 3766
rect 1216 3732 1254 3740
rect 1288 3732 1289 3766
rect 1109 3706 1289 3732
rect 1109 3692 1146 3706
rect 1109 3658 1110 3692
rect 1144 3672 1146 3692
rect 1180 3692 1218 3706
rect 1180 3672 1182 3692
rect 1144 3658 1182 3672
rect 1216 3672 1218 3692
rect 1252 3692 1289 3706
rect 1252 3672 1254 3692
rect 1216 3658 1254 3672
rect 1288 3658 1289 3692
rect 1109 3638 1289 3658
rect 1109 3618 1146 3638
rect 1109 3584 1110 3618
rect 1144 3604 1146 3618
rect 1180 3618 1218 3638
rect 1180 3604 1182 3618
rect 1144 3584 1182 3604
rect 1216 3604 1218 3618
rect 1252 3618 1289 3638
rect 1252 3604 1254 3618
rect 1216 3584 1254 3604
rect 1288 3584 1289 3618
rect 1109 3570 1289 3584
rect 1109 3544 1146 3570
rect 1109 3510 1110 3544
rect 1144 3536 1146 3544
rect 1180 3544 1218 3570
rect 1180 3536 1182 3544
rect 1144 3510 1182 3536
rect 1216 3536 1218 3544
rect 1252 3544 1289 3570
rect 1252 3536 1254 3544
rect 1216 3510 1254 3536
rect 1288 3510 1289 3544
rect 1109 3502 1289 3510
rect 1109 3470 1146 3502
rect 1109 3436 1110 3470
rect 1144 3468 1146 3470
rect 1180 3470 1218 3502
rect 1180 3468 1182 3470
rect 1144 3436 1182 3468
rect 1216 3468 1218 3470
rect 1252 3470 1289 3502
rect 1252 3468 1254 3470
rect 1216 3436 1254 3468
rect 1288 3436 1289 3470
rect 1109 3434 1289 3436
rect 1109 3400 1146 3434
rect 1180 3400 1218 3434
rect 1252 3400 1289 3434
rect 1109 3396 1289 3400
rect 1109 3362 1110 3396
rect 1144 3366 1182 3396
rect 1144 3362 1146 3366
rect 1109 3332 1146 3362
rect 1180 3362 1182 3366
rect 1216 3366 1254 3396
rect 1216 3362 1218 3366
rect 1180 3332 1218 3362
rect 1252 3362 1254 3366
rect 1288 3362 1289 3396
rect 1252 3332 1289 3362
rect 1109 3322 1289 3332
rect 1109 3288 1110 3322
rect 1144 3298 1182 3322
rect 1144 3288 1146 3298
rect 1109 3264 1146 3288
rect 1180 3288 1182 3298
rect 1216 3298 1254 3322
rect 1216 3288 1218 3298
rect 1180 3264 1218 3288
rect 1252 3288 1254 3298
rect 1288 3288 1289 3322
rect 1252 3264 1289 3288
rect 1109 3248 1289 3264
rect 1109 3214 1110 3248
rect 1144 3230 1182 3248
rect 1144 3214 1146 3230
rect 1109 3196 1146 3214
rect 1180 3214 1182 3230
rect 1216 3230 1254 3248
rect 1216 3214 1218 3230
rect 1180 3196 1218 3214
rect 1252 3214 1254 3230
rect 1288 3214 1289 3248
rect 1252 3196 1289 3214
rect 1109 3174 1289 3196
rect 1109 3140 1110 3174
rect 1144 3162 1182 3174
rect 1144 3140 1146 3162
rect 1109 3128 1146 3140
rect 1180 3140 1182 3162
rect 1216 3162 1254 3174
rect 1216 3140 1218 3162
rect 1180 3128 1218 3140
rect 1252 3140 1254 3162
rect 1288 3140 1289 3174
rect 1252 3128 1289 3140
rect 1109 3100 1289 3128
rect 1109 3066 1110 3100
rect 1144 3066 1182 3100
rect 1216 3066 1254 3100
rect 1288 3066 1289 3100
rect 1109 3026 1289 3066
rect 1109 2992 1110 3026
rect 1144 2992 1182 3026
rect 1216 2992 1254 3026
rect 1288 2992 1289 3026
rect 1109 2952 1289 2992
rect 1109 2918 1110 2952
rect 1144 2918 1182 2952
rect 1216 2918 1254 2952
rect 1288 2918 1289 2952
rect 1109 2878 1289 2918
rect 1109 2844 1110 2878
rect 1144 2844 1182 2878
rect 1216 2844 1254 2878
rect 1288 2844 1289 2878
rect 1109 2804 1289 2844
rect 1109 2770 1110 2804
rect 1144 2770 1182 2804
rect 1216 2770 1254 2804
rect 1288 2770 1289 2804
rect 1109 2730 1289 2770
rect 1109 2696 1110 2730
rect 1144 2696 1182 2730
rect 1216 2696 1254 2730
rect 1288 2696 1289 2730
rect 1109 2656 1289 2696
rect 1109 2622 1110 2656
rect 1144 2622 1182 2656
rect 1216 2622 1254 2656
rect 1288 2622 1289 2656
rect 1109 2582 1289 2622
rect 1109 2548 1110 2582
rect 1144 2548 1182 2582
rect 1216 2548 1254 2582
rect 1288 2548 1289 2582
rect 1109 2508 1289 2548
rect 1109 2474 1110 2508
rect 1144 2474 1182 2508
rect 1216 2474 1254 2508
rect 1288 2474 1289 2508
rect 1109 2445 1289 2474
rect 1109 2434 1146 2445
rect 1109 2400 1110 2434
rect 1144 2411 1146 2434
rect 1180 2434 1218 2445
rect 1180 2411 1182 2434
rect 1144 2400 1182 2411
rect 1216 2411 1218 2434
rect 1252 2434 1289 2445
rect 1252 2411 1254 2434
rect 1216 2400 1254 2411
rect 1288 2400 1289 2434
rect 1109 2377 1289 2400
rect 1109 2360 1146 2377
rect 1109 2326 1110 2360
rect 1144 2343 1146 2360
rect 1180 2360 1218 2377
rect 1180 2343 1182 2360
rect 1144 2326 1182 2343
rect 1216 2343 1218 2360
rect 1252 2360 1289 2377
rect 1252 2343 1254 2360
rect 1216 2326 1254 2343
rect 1288 2326 1289 2360
rect 1109 2309 1289 2326
rect 1109 2286 1146 2309
rect 1109 2252 1110 2286
rect 1144 2275 1146 2286
rect 1180 2286 1218 2309
rect 1180 2275 1182 2286
rect 1144 2252 1182 2275
rect 1216 2275 1218 2286
rect 1252 2286 1289 2309
rect 1252 2275 1254 2286
rect 1216 2252 1254 2275
rect 1288 2252 1289 2286
rect 1109 2241 1289 2252
rect 1109 2212 1146 2241
rect 1109 2178 1110 2212
rect 1144 2207 1146 2212
rect 1180 2212 1218 2241
rect 1180 2207 1182 2212
rect 1144 2178 1182 2207
rect 1216 2207 1218 2212
rect 1252 2212 1289 2241
rect 1252 2207 1254 2212
rect 1216 2178 1254 2207
rect 1288 2178 1289 2212
rect 1109 2173 1289 2178
rect 1109 2139 1146 2173
rect 1180 2139 1218 2173
rect 1252 2139 1289 2173
rect 1109 2138 1289 2139
rect 1109 2104 1110 2138
rect 1144 2105 1182 2138
rect 1144 2104 1146 2105
rect 1109 2071 1146 2104
rect 1180 2104 1182 2105
rect 1216 2105 1254 2138
rect 1216 2104 1218 2105
rect 1180 2071 1218 2104
rect 1252 2104 1254 2105
rect 1288 2104 1289 2138
rect 1252 2071 1289 2104
rect 1109 2064 1289 2071
rect 1109 2030 1110 2064
rect 1144 2037 1182 2064
rect 1144 2030 1146 2037
rect 1109 2003 1146 2030
rect 1180 2030 1182 2037
rect 1216 2037 1254 2064
rect 1216 2030 1218 2037
rect 1180 2003 1218 2030
rect 1252 2030 1254 2037
rect 1288 2030 1289 2064
rect 1252 2003 1289 2030
rect 1109 1990 1289 2003
rect 1109 1956 1110 1990
rect 1144 1969 1182 1990
rect 1144 1956 1146 1969
rect 1109 1935 1146 1956
rect 1180 1956 1182 1969
rect 1216 1969 1254 1990
rect 1216 1956 1218 1969
rect 1180 1935 1218 1956
rect 1252 1956 1254 1969
rect 1288 1956 1289 1990
rect 1252 1935 1289 1956
rect 1109 1916 1289 1935
rect 1109 1882 1110 1916
rect 1144 1901 1182 1916
rect 1144 1882 1146 1901
rect 1109 1867 1146 1882
rect 1180 1882 1182 1901
rect 1216 1901 1254 1916
rect 1216 1882 1218 1901
rect 1180 1867 1218 1882
rect 1252 1882 1254 1901
rect 1288 1882 1289 1916
rect 1252 1867 1289 1882
rect 1109 1842 1289 1867
rect 1109 1808 1110 1842
rect 1144 1833 1182 1842
rect 1144 1808 1146 1833
rect 1109 1799 1146 1808
rect 1180 1808 1182 1833
rect 1216 1833 1254 1842
rect 1216 1808 1218 1833
rect 1180 1799 1218 1808
rect 1252 1808 1254 1833
rect 1288 1808 1289 1842
rect 1252 1799 1289 1808
rect 1109 1768 1289 1799
rect 1109 1734 1110 1768
rect 1144 1765 1182 1768
rect 1144 1734 1146 1765
rect 1109 1731 1146 1734
rect 1180 1734 1182 1765
rect 1216 1765 1254 1768
rect 1216 1734 1218 1765
rect 1180 1731 1218 1734
rect 1252 1734 1254 1765
rect 1288 1734 1289 1768
rect 1252 1731 1289 1734
rect 1109 1697 1289 1731
rect 1109 1694 1146 1697
rect 1109 1660 1110 1694
rect 1144 1663 1146 1694
rect 1180 1694 1218 1697
rect 1180 1663 1182 1694
rect 1144 1660 1182 1663
rect 1216 1663 1218 1694
rect 1252 1694 1289 1697
rect 1252 1663 1254 1694
rect 1216 1660 1254 1663
rect 1288 1660 1289 1694
rect 1109 1629 1289 1660
rect 1109 1620 1146 1629
rect 1109 1586 1110 1620
rect 1144 1595 1146 1620
rect 1180 1620 1218 1629
rect 1180 1595 1182 1620
rect 1144 1586 1182 1595
rect 1216 1595 1218 1620
rect 1252 1620 1289 1629
rect 1252 1595 1254 1620
rect 1216 1586 1254 1595
rect 1288 1586 1289 1620
rect 1109 1561 1289 1586
rect 1109 1545 1146 1561
rect 1109 1511 1110 1545
rect 1144 1527 1146 1545
rect 1180 1545 1218 1561
rect 1180 1527 1182 1545
rect 1144 1511 1182 1527
rect 1216 1527 1218 1545
rect 1252 1545 1289 1561
rect 1252 1527 1254 1545
rect 1216 1511 1254 1527
rect 1288 1511 1289 1545
rect 1354 3010 1474 4106
rect 1916 4388 1923 4494
rect 2029 4388 2036 4494
rect 1916 4214 2036 4388
rect 1916 4180 1959 4214
rect 1993 4180 2036 4214
rect 1916 4140 2036 4180
rect 1916 4106 1959 4140
rect 1993 4106 2036 4140
rect 1354 2976 1397 3010
rect 1431 2976 1474 3010
rect 1354 2932 1474 2976
rect 1354 2898 1397 2932
rect 1431 2898 1474 2932
rect 1354 2854 1474 2898
rect 1354 2820 1397 2854
rect 1431 2820 1474 2854
rect 1354 2776 1474 2820
rect 1354 2742 1397 2776
rect 1431 2742 1474 2776
rect 1354 2697 1474 2742
rect 1354 2663 1397 2697
rect 1431 2663 1474 2697
rect 1354 2618 1474 2663
rect 1354 2584 1397 2618
rect 1431 2584 1474 2618
rect 1354 2539 1474 2584
rect 1354 2505 1397 2539
rect 1431 2505 1474 2539
rect 1146 1491 1252 1511
rect 924 1375 967 1409
rect 1001 1375 1044 1409
rect 924 1335 1044 1375
rect 924 1301 967 1335
rect 1001 1301 1044 1335
rect 924 1285 1044 1301
rect 1354 1409 1474 2505
rect 1576 4050 1678 4062
rect 1712 4050 1814 4062
rect 1576 4046 1606 4050
rect 1784 4046 1814 4050
rect 1576 3978 1606 4012
rect 1784 3978 1814 4012
rect 1576 3910 1606 3944
rect 1784 3910 1814 3944
rect 1576 3842 1606 3876
rect 1784 3842 1814 3876
rect 1576 3774 1606 3808
rect 1784 3774 1814 3808
rect 1576 3706 1606 3740
rect 1784 3706 1814 3740
rect 1576 3638 1606 3672
rect 1784 3638 1814 3672
rect 1576 3570 1606 3604
rect 1784 3570 1814 3604
rect 1576 3502 1606 3536
rect 1784 3502 1814 3536
rect 1576 3434 1606 3468
rect 1784 3434 1814 3468
rect 1576 3366 1606 3400
rect 1784 3366 1814 3400
rect 1576 3298 1606 3332
rect 1784 3298 1814 3332
rect 1576 3230 1606 3264
rect 1784 3230 1814 3264
rect 1576 3162 1606 3196
rect 1784 3162 1814 3196
rect 1576 3080 1606 3128
rect 1640 3080 1750 3092
rect 1784 3080 1814 3128
rect 1576 3040 1814 3080
rect 1576 2574 1606 3040
rect 1784 2574 1814 3040
rect 1576 2535 1814 2574
rect 1576 2501 1606 2535
rect 1640 2501 1678 2535
rect 1712 2501 1750 2535
rect 1784 2501 1814 2535
rect 1576 2461 1814 2501
rect 1576 2449 1678 2461
rect 1712 2449 1814 2461
rect 1576 2445 1606 2449
rect 1784 2445 1814 2449
rect 1576 2377 1606 2411
rect 1784 2377 1814 2411
rect 1576 2309 1606 2343
rect 1784 2309 1814 2343
rect 1576 2241 1606 2275
rect 1784 2241 1814 2275
rect 1576 2173 1606 2207
rect 1784 2173 1814 2207
rect 1576 2105 1606 2139
rect 1784 2105 1814 2139
rect 1576 2037 1606 2071
rect 1784 2037 1814 2071
rect 1576 1969 1606 2003
rect 1784 1969 1814 2003
rect 1576 1901 1606 1935
rect 1784 1901 1814 1935
rect 1576 1833 1606 1867
rect 1784 1833 1814 1867
rect 1576 1765 1606 1799
rect 1784 1765 1814 1799
rect 1576 1697 1606 1731
rect 1784 1697 1814 1731
rect 1576 1629 1606 1663
rect 1784 1629 1814 1663
rect 1576 1561 1606 1595
rect 1784 1561 1814 1595
rect 1576 1479 1606 1527
rect 1640 1479 1750 1491
rect 1784 1479 1814 1527
rect 1576 1464 1814 1479
rect 1916 3010 2036 4106
rect 2346 4388 2353 4494
rect 2459 4388 2466 4494
rect 2346 4214 2466 4388
rect 2346 4180 2389 4214
rect 2423 4180 2466 4214
rect 2346 4140 2466 4180
rect 2346 4106 2389 4140
rect 2423 4106 2466 4140
rect 1916 2976 1959 3010
rect 1993 2976 2036 3010
rect 1916 2932 2036 2976
rect 1916 2898 1959 2932
rect 1993 2898 2036 2932
rect 1916 2854 2036 2898
rect 1916 2820 1959 2854
rect 1993 2820 2036 2854
rect 1916 2776 2036 2820
rect 1916 2742 1959 2776
rect 1993 2742 2036 2776
rect 1916 2697 2036 2742
rect 1916 2663 1959 2697
rect 1993 2663 2036 2697
rect 1916 2618 2036 2663
rect 1916 2584 1959 2618
rect 1993 2584 2036 2618
rect 1916 2539 2036 2584
rect 1916 2505 1959 2539
rect 1993 2505 2036 2539
rect 1354 1375 1397 1409
rect 1431 1375 1474 1409
rect 1354 1335 1474 1375
rect 1354 1301 1397 1335
rect 1431 1301 1474 1335
rect 1354 1285 1474 1301
rect 1916 1409 2036 2505
rect 2101 4028 2102 4062
rect 2136 4046 2174 4062
rect 2136 4028 2138 4046
rect 2101 4012 2138 4028
rect 2172 4028 2174 4046
rect 2208 4046 2246 4062
rect 2208 4028 2210 4046
rect 2172 4012 2210 4028
rect 2244 4028 2246 4046
rect 2280 4028 2281 4062
rect 2244 4012 2281 4028
rect 2101 3988 2281 4012
rect 2101 3954 2102 3988
rect 2136 3978 2174 3988
rect 2136 3954 2138 3978
rect 2101 3944 2138 3954
rect 2172 3954 2174 3978
rect 2208 3978 2246 3988
rect 2208 3954 2210 3978
rect 2172 3944 2210 3954
rect 2244 3954 2246 3978
rect 2280 3954 2281 3988
rect 2244 3944 2281 3954
rect 2101 3914 2281 3944
rect 2101 3880 2102 3914
rect 2136 3910 2174 3914
rect 2136 3880 2138 3910
rect 2101 3876 2138 3880
rect 2172 3880 2174 3910
rect 2208 3910 2246 3914
rect 2208 3880 2210 3910
rect 2172 3876 2210 3880
rect 2244 3880 2246 3910
rect 2280 3880 2281 3914
rect 2244 3876 2281 3880
rect 2101 3842 2281 3876
rect 2101 3840 2138 3842
rect 2101 3806 2102 3840
rect 2136 3808 2138 3840
rect 2172 3840 2210 3842
rect 2172 3808 2174 3840
rect 2136 3806 2174 3808
rect 2208 3808 2210 3840
rect 2244 3840 2281 3842
rect 2244 3808 2246 3840
rect 2208 3806 2246 3808
rect 2280 3806 2281 3840
rect 2101 3774 2281 3806
rect 2101 3766 2138 3774
rect 2101 3732 2102 3766
rect 2136 3740 2138 3766
rect 2172 3766 2210 3774
rect 2172 3740 2174 3766
rect 2136 3732 2174 3740
rect 2208 3740 2210 3766
rect 2244 3766 2281 3774
rect 2244 3740 2246 3766
rect 2208 3732 2246 3740
rect 2280 3732 2281 3766
rect 2101 3706 2281 3732
rect 2101 3692 2138 3706
rect 2101 3658 2102 3692
rect 2136 3672 2138 3692
rect 2172 3692 2210 3706
rect 2172 3672 2174 3692
rect 2136 3658 2174 3672
rect 2208 3672 2210 3692
rect 2244 3692 2281 3706
rect 2244 3672 2246 3692
rect 2208 3658 2246 3672
rect 2280 3658 2281 3692
rect 2101 3638 2281 3658
rect 2101 3618 2138 3638
rect 2101 3584 2102 3618
rect 2136 3604 2138 3618
rect 2172 3618 2210 3638
rect 2172 3604 2174 3618
rect 2136 3584 2174 3604
rect 2208 3604 2210 3618
rect 2244 3618 2281 3638
rect 2244 3604 2246 3618
rect 2208 3584 2246 3604
rect 2280 3584 2281 3618
rect 2101 3570 2281 3584
rect 2101 3544 2138 3570
rect 2101 3510 2102 3544
rect 2136 3536 2138 3544
rect 2172 3544 2210 3570
rect 2172 3536 2174 3544
rect 2136 3510 2174 3536
rect 2208 3536 2210 3544
rect 2244 3544 2281 3570
rect 2244 3536 2246 3544
rect 2208 3510 2246 3536
rect 2280 3510 2281 3544
rect 2101 3502 2281 3510
rect 2101 3470 2138 3502
rect 2101 3436 2102 3470
rect 2136 3468 2138 3470
rect 2172 3470 2210 3502
rect 2172 3468 2174 3470
rect 2136 3436 2174 3468
rect 2208 3468 2210 3470
rect 2244 3470 2281 3502
rect 2244 3468 2246 3470
rect 2208 3436 2246 3468
rect 2280 3436 2281 3470
rect 2101 3434 2281 3436
rect 2101 3400 2138 3434
rect 2172 3400 2210 3434
rect 2244 3400 2281 3434
rect 2101 3396 2281 3400
rect 2101 3362 2102 3396
rect 2136 3366 2174 3396
rect 2136 3362 2138 3366
rect 2101 3332 2138 3362
rect 2172 3362 2174 3366
rect 2208 3366 2246 3396
rect 2208 3362 2210 3366
rect 2172 3332 2210 3362
rect 2244 3362 2246 3366
rect 2280 3362 2281 3396
rect 2244 3332 2281 3362
rect 2101 3322 2281 3332
rect 2101 3288 2102 3322
rect 2136 3298 2174 3322
rect 2136 3288 2138 3298
rect 2101 3264 2138 3288
rect 2172 3288 2174 3298
rect 2208 3298 2246 3322
rect 2208 3288 2210 3298
rect 2172 3264 2210 3288
rect 2244 3288 2246 3298
rect 2280 3288 2281 3322
rect 2244 3264 2281 3288
rect 2101 3248 2281 3264
rect 2101 3214 2102 3248
rect 2136 3230 2174 3248
rect 2136 3214 2138 3230
rect 2101 3196 2138 3214
rect 2172 3214 2174 3230
rect 2208 3230 2246 3248
rect 2208 3214 2210 3230
rect 2172 3196 2210 3214
rect 2244 3214 2246 3230
rect 2280 3214 2281 3248
rect 2244 3196 2281 3214
rect 2101 3174 2281 3196
rect 2101 3140 2102 3174
rect 2136 3162 2174 3174
rect 2136 3140 2138 3162
rect 2101 3128 2138 3140
rect 2172 3140 2174 3162
rect 2208 3162 2246 3174
rect 2208 3140 2210 3162
rect 2172 3128 2210 3140
rect 2244 3140 2246 3162
rect 2280 3140 2281 3174
rect 2244 3128 2281 3140
rect 2101 3100 2281 3128
rect 2101 3066 2102 3100
rect 2136 3066 2174 3100
rect 2208 3066 2246 3100
rect 2280 3066 2281 3100
rect 2101 3026 2281 3066
rect 2101 2992 2102 3026
rect 2136 2992 2174 3026
rect 2208 2992 2246 3026
rect 2280 2992 2281 3026
rect 2101 2952 2281 2992
rect 2101 2918 2102 2952
rect 2136 2918 2174 2952
rect 2208 2918 2246 2952
rect 2280 2918 2281 2952
rect 2101 2878 2281 2918
rect 2101 2844 2102 2878
rect 2136 2844 2174 2878
rect 2208 2844 2246 2878
rect 2280 2844 2281 2878
rect 2101 2804 2281 2844
rect 2101 2770 2102 2804
rect 2136 2770 2174 2804
rect 2208 2770 2246 2804
rect 2280 2770 2281 2804
rect 2101 2730 2281 2770
rect 2101 2696 2102 2730
rect 2136 2696 2174 2730
rect 2208 2696 2246 2730
rect 2280 2696 2281 2730
rect 2101 2656 2281 2696
rect 2101 2622 2102 2656
rect 2136 2622 2174 2656
rect 2208 2622 2246 2656
rect 2280 2622 2281 2656
rect 2101 2582 2281 2622
rect 2101 2548 2102 2582
rect 2136 2548 2174 2582
rect 2208 2548 2246 2582
rect 2280 2548 2281 2582
rect 2101 2508 2281 2548
rect 2101 2474 2102 2508
rect 2136 2474 2174 2508
rect 2208 2474 2246 2508
rect 2280 2474 2281 2508
rect 2101 2445 2281 2474
rect 2101 2434 2138 2445
rect 2101 2400 2102 2434
rect 2136 2411 2138 2434
rect 2172 2434 2210 2445
rect 2172 2411 2174 2434
rect 2136 2400 2174 2411
rect 2208 2411 2210 2434
rect 2244 2434 2281 2445
rect 2244 2411 2246 2434
rect 2208 2400 2246 2411
rect 2280 2400 2281 2434
rect 2101 2377 2281 2400
rect 2101 2360 2138 2377
rect 2101 2326 2102 2360
rect 2136 2343 2138 2360
rect 2172 2360 2210 2377
rect 2172 2343 2174 2360
rect 2136 2326 2174 2343
rect 2208 2343 2210 2360
rect 2244 2360 2281 2377
rect 2244 2343 2246 2360
rect 2208 2326 2246 2343
rect 2280 2326 2281 2360
rect 2101 2309 2281 2326
rect 2101 2286 2138 2309
rect 2101 2252 2102 2286
rect 2136 2275 2138 2286
rect 2172 2286 2210 2309
rect 2172 2275 2174 2286
rect 2136 2252 2174 2275
rect 2208 2275 2210 2286
rect 2244 2286 2281 2309
rect 2244 2275 2246 2286
rect 2208 2252 2246 2275
rect 2280 2252 2281 2286
rect 2101 2241 2281 2252
rect 2101 2212 2138 2241
rect 2101 2178 2102 2212
rect 2136 2207 2138 2212
rect 2172 2212 2210 2241
rect 2172 2207 2174 2212
rect 2136 2178 2174 2207
rect 2208 2207 2210 2212
rect 2244 2212 2281 2241
rect 2244 2207 2246 2212
rect 2208 2178 2246 2207
rect 2280 2178 2281 2212
rect 2101 2173 2281 2178
rect 2101 2139 2138 2173
rect 2172 2139 2210 2173
rect 2244 2139 2281 2173
rect 2101 2138 2281 2139
rect 2101 2104 2102 2138
rect 2136 2105 2174 2138
rect 2136 2104 2138 2105
rect 2101 2071 2138 2104
rect 2172 2104 2174 2105
rect 2208 2105 2246 2138
rect 2208 2104 2210 2105
rect 2172 2071 2210 2104
rect 2244 2104 2246 2105
rect 2280 2104 2281 2138
rect 2244 2071 2281 2104
rect 2101 2064 2281 2071
rect 2101 2030 2102 2064
rect 2136 2037 2174 2064
rect 2136 2030 2138 2037
rect 2101 2003 2138 2030
rect 2172 2030 2174 2037
rect 2208 2037 2246 2064
rect 2208 2030 2210 2037
rect 2172 2003 2210 2030
rect 2244 2030 2246 2037
rect 2280 2030 2281 2064
rect 2244 2003 2281 2030
rect 2101 1990 2281 2003
rect 2101 1956 2102 1990
rect 2136 1969 2174 1990
rect 2136 1956 2138 1969
rect 2101 1935 2138 1956
rect 2172 1956 2174 1969
rect 2208 1969 2246 1990
rect 2208 1956 2210 1969
rect 2172 1935 2210 1956
rect 2244 1956 2246 1969
rect 2280 1956 2281 1990
rect 2244 1935 2281 1956
rect 2101 1916 2281 1935
rect 2101 1882 2102 1916
rect 2136 1901 2174 1916
rect 2136 1882 2138 1901
rect 2101 1867 2138 1882
rect 2172 1882 2174 1901
rect 2208 1901 2246 1916
rect 2208 1882 2210 1901
rect 2172 1867 2210 1882
rect 2244 1882 2246 1901
rect 2280 1882 2281 1916
rect 2244 1867 2281 1882
rect 2101 1842 2281 1867
rect 2101 1808 2102 1842
rect 2136 1833 2174 1842
rect 2136 1808 2138 1833
rect 2101 1799 2138 1808
rect 2172 1808 2174 1833
rect 2208 1833 2246 1842
rect 2208 1808 2210 1833
rect 2172 1799 2210 1808
rect 2244 1808 2246 1833
rect 2280 1808 2281 1842
rect 2244 1799 2281 1808
rect 2101 1768 2281 1799
rect 2101 1734 2102 1768
rect 2136 1765 2174 1768
rect 2136 1734 2138 1765
rect 2101 1731 2138 1734
rect 2172 1734 2174 1765
rect 2208 1765 2246 1768
rect 2208 1734 2210 1765
rect 2172 1731 2210 1734
rect 2244 1734 2246 1765
rect 2280 1734 2281 1768
rect 2244 1731 2281 1734
rect 2101 1697 2281 1731
rect 2101 1694 2138 1697
rect 2101 1660 2102 1694
rect 2136 1663 2138 1694
rect 2172 1694 2210 1697
rect 2172 1663 2174 1694
rect 2136 1660 2174 1663
rect 2208 1663 2210 1694
rect 2244 1694 2281 1697
rect 2244 1663 2246 1694
rect 2208 1660 2246 1663
rect 2280 1660 2281 1694
rect 2101 1629 2281 1660
rect 2101 1620 2138 1629
rect 2101 1586 2102 1620
rect 2136 1595 2138 1620
rect 2172 1620 2210 1629
rect 2172 1595 2174 1620
rect 2136 1586 2174 1595
rect 2208 1595 2210 1620
rect 2244 1620 2281 1629
rect 2244 1595 2246 1620
rect 2208 1586 2246 1595
rect 2280 1586 2281 1620
rect 2101 1561 2281 1586
rect 2101 1545 2138 1561
rect 2101 1511 2102 1545
rect 2136 1527 2138 1545
rect 2172 1545 2210 1561
rect 2172 1527 2174 1545
rect 2136 1511 2174 1527
rect 2208 1527 2210 1545
rect 2244 1545 2281 1561
rect 2244 1527 2246 1545
rect 2208 1511 2246 1527
rect 2280 1511 2281 1545
rect 2346 3010 2466 4106
rect 2908 4388 2915 4494
rect 3021 4388 3028 4494
rect 2908 4214 3028 4388
rect 2908 4180 2951 4214
rect 2985 4180 3028 4214
rect 2908 4140 3028 4180
rect 2908 4106 2951 4140
rect 2985 4106 3028 4140
rect 2346 2976 2389 3010
rect 2423 2976 2466 3010
rect 2346 2932 2466 2976
rect 2346 2898 2389 2932
rect 2423 2898 2466 2932
rect 2346 2854 2466 2898
rect 2346 2820 2389 2854
rect 2423 2820 2466 2854
rect 2346 2776 2466 2820
rect 2346 2742 2389 2776
rect 2423 2742 2466 2776
rect 2346 2697 2466 2742
rect 2346 2663 2389 2697
rect 2423 2663 2466 2697
rect 2346 2618 2466 2663
rect 2346 2584 2389 2618
rect 2423 2584 2466 2618
rect 2346 2539 2466 2584
rect 2346 2505 2389 2539
rect 2423 2505 2466 2539
rect 2138 1491 2244 1511
rect 1916 1375 1959 1409
rect 1993 1375 2036 1409
rect 1916 1335 2036 1375
rect 1916 1301 1959 1335
rect 1993 1301 2036 1335
rect 1916 1285 2036 1301
rect 2346 1409 2466 2505
rect 2568 4050 2670 4062
rect 2704 4050 2806 4062
rect 2568 4046 2598 4050
rect 2776 4046 2806 4050
rect 2568 3978 2598 4012
rect 2776 3978 2806 4012
rect 2568 3910 2598 3944
rect 2776 3910 2806 3944
rect 2568 3842 2598 3876
rect 2776 3842 2806 3876
rect 2568 3774 2598 3808
rect 2776 3774 2806 3808
rect 2568 3706 2598 3740
rect 2776 3706 2806 3740
rect 2568 3638 2598 3672
rect 2776 3638 2806 3672
rect 2568 3570 2598 3604
rect 2776 3570 2806 3604
rect 2568 3502 2598 3536
rect 2776 3502 2806 3536
rect 2568 3434 2598 3468
rect 2776 3434 2806 3468
rect 2568 3366 2598 3400
rect 2776 3366 2806 3400
rect 2568 3298 2598 3332
rect 2776 3298 2806 3332
rect 2568 3230 2598 3264
rect 2776 3230 2806 3264
rect 2568 3162 2598 3196
rect 2776 3162 2806 3196
rect 2568 3080 2598 3128
rect 2632 3080 2742 3092
rect 2776 3080 2806 3128
rect 2568 3040 2806 3080
rect 2568 2574 2598 3040
rect 2776 2574 2806 3040
rect 2568 2535 2806 2574
rect 2568 2501 2598 2535
rect 2632 2501 2670 2535
rect 2704 2501 2742 2535
rect 2776 2501 2806 2535
rect 2568 2461 2806 2501
rect 2568 2449 2670 2461
rect 2704 2449 2806 2461
rect 2568 2445 2598 2449
rect 2776 2445 2806 2449
rect 2568 2377 2598 2411
rect 2776 2377 2806 2411
rect 2568 2309 2598 2343
rect 2776 2309 2806 2343
rect 2568 2241 2598 2275
rect 2776 2241 2806 2275
rect 2568 2173 2598 2207
rect 2776 2173 2806 2207
rect 2568 2105 2598 2139
rect 2776 2105 2806 2139
rect 2568 2037 2598 2071
rect 2776 2037 2806 2071
rect 2568 1969 2598 2003
rect 2776 1969 2806 2003
rect 2568 1901 2598 1935
rect 2776 1901 2806 1935
rect 2568 1833 2598 1867
rect 2776 1833 2806 1867
rect 2568 1765 2598 1799
rect 2776 1765 2806 1799
rect 2568 1697 2598 1731
rect 2776 1697 2806 1731
rect 2568 1629 2598 1663
rect 2776 1629 2806 1663
rect 2568 1561 2598 1595
rect 2776 1561 2806 1595
rect 2568 1479 2598 1527
rect 2632 1479 2742 1491
rect 2776 1479 2806 1527
rect 2568 1464 2806 1479
rect 2908 3010 3028 4106
rect 3338 4388 3345 4494
rect 3451 4388 3458 4494
rect 3338 4214 3458 4388
rect 3338 4180 3381 4214
rect 3415 4180 3458 4214
rect 3338 4140 3458 4180
rect 3338 4106 3381 4140
rect 3415 4106 3458 4140
rect 2908 2976 2951 3010
rect 2985 2976 3028 3010
rect 2908 2932 3028 2976
rect 2908 2898 2951 2932
rect 2985 2898 3028 2932
rect 2908 2854 3028 2898
rect 2908 2820 2951 2854
rect 2985 2820 3028 2854
rect 2908 2776 3028 2820
rect 2908 2742 2951 2776
rect 2985 2742 3028 2776
rect 2908 2697 3028 2742
rect 2908 2663 2951 2697
rect 2985 2663 3028 2697
rect 2908 2618 3028 2663
rect 2908 2584 2951 2618
rect 2985 2584 3028 2618
rect 2908 2539 3028 2584
rect 2908 2505 2951 2539
rect 2985 2505 3028 2539
rect 2346 1375 2389 1409
rect 2423 1375 2466 1409
rect 2346 1335 2466 1375
rect 2346 1301 2389 1335
rect 2423 1301 2466 1335
rect 2346 1285 2466 1301
rect 2908 1409 3028 2505
rect 3093 4028 3094 4062
rect 3128 4046 3166 4062
rect 3128 4028 3130 4046
rect 3093 4012 3130 4028
rect 3164 4028 3166 4046
rect 3200 4046 3238 4062
rect 3200 4028 3202 4046
rect 3164 4012 3202 4028
rect 3236 4028 3238 4046
rect 3272 4028 3273 4062
rect 3236 4012 3273 4028
rect 3093 3988 3273 4012
rect 3093 3954 3094 3988
rect 3128 3978 3166 3988
rect 3128 3954 3130 3978
rect 3093 3944 3130 3954
rect 3164 3954 3166 3978
rect 3200 3978 3238 3988
rect 3200 3954 3202 3978
rect 3164 3944 3202 3954
rect 3236 3954 3238 3978
rect 3272 3954 3273 3988
rect 3236 3944 3273 3954
rect 3093 3914 3273 3944
rect 3093 3880 3094 3914
rect 3128 3910 3166 3914
rect 3128 3880 3130 3910
rect 3093 3876 3130 3880
rect 3164 3880 3166 3910
rect 3200 3910 3238 3914
rect 3200 3880 3202 3910
rect 3164 3876 3202 3880
rect 3236 3880 3238 3910
rect 3272 3880 3273 3914
rect 3236 3876 3273 3880
rect 3093 3842 3273 3876
rect 3093 3840 3130 3842
rect 3093 3806 3094 3840
rect 3128 3808 3130 3840
rect 3164 3840 3202 3842
rect 3164 3808 3166 3840
rect 3128 3806 3166 3808
rect 3200 3808 3202 3840
rect 3236 3840 3273 3842
rect 3236 3808 3238 3840
rect 3200 3806 3238 3808
rect 3272 3806 3273 3840
rect 3093 3774 3273 3806
rect 3093 3766 3130 3774
rect 3093 3732 3094 3766
rect 3128 3740 3130 3766
rect 3164 3766 3202 3774
rect 3164 3740 3166 3766
rect 3128 3732 3166 3740
rect 3200 3740 3202 3766
rect 3236 3766 3273 3774
rect 3236 3740 3238 3766
rect 3200 3732 3238 3740
rect 3272 3732 3273 3766
rect 3093 3706 3273 3732
rect 3093 3692 3130 3706
rect 3093 3658 3094 3692
rect 3128 3672 3130 3692
rect 3164 3692 3202 3706
rect 3164 3672 3166 3692
rect 3128 3658 3166 3672
rect 3200 3672 3202 3692
rect 3236 3692 3273 3706
rect 3236 3672 3238 3692
rect 3200 3658 3238 3672
rect 3272 3658 3273 3692
rect 3093 3638 3273 3658
rect 3093 3618 3130 3638
rect 3093 3584 3094 3618
rect 3128 3604 3130 3618
rect 3164 3618 3202 3638
rect 3164 3604 3166 3618
rect 3128 3584 3166 3604
rect 3200 3604 3202 3618
rect 3236 3618 3273 3638
rect 3236 3604 3238 3618
rect 3200 3584 3238 3604
rect 3272 3584 3273 3618
rect 3093 3570 3273 3584
rect 3093 3544 3130 3570
rect 3093 3510 3094 3544
rect 3128 3536 3130 3544
rect 3164 3544 3202 3570
rect 3164 3536 3166 3544
rect 3128 3510 3166 3536
rect 3200 3536 3202 3544
rect 3236 3544 3273 3570
rect 3236 3536 3238 3544
rect 3200 3510 3238 3536
rect 3272 3510 3273 3544
rect 3093 3502 3273 3510
rect 3093 3470 3130 3502
rect 3093 3436 3094 3470
rect 3128 3468 3130 3470
rect 3164 3470 3202 3502
rect 3164 3468 3166 3470
rect 3128 3436 3166 3468
rect 3200 3468 3202 3470
rect 3236 3470 3273 3502
rect 3236 3468 3238 3470
rect 3200 3436 3238 3468
rect 3272 3436 3273 3470
rect 3093 3434 3273 3436
rect 3093 3400 3130 3434
rect 3164 3400 3202 3434
rect 3236 3400 3273 3434
rect 3093 3396 3273 3400
rect 3093 3362 3094 3396
rect 3128 3366 3166 3396
rect 3128 3362 3130 3366
rect 3093 3332 3130 3362
rect 3164 3362 3166 3366
rect 3200 3366 3238 3396
rect 3200 3362 3202 3366
rect 3164 3332 3202 3362
rect 3236 3362 3238 3366
rect 3272 3362 3273 3396
rect 3236 3332 3273 3362
rect 3093 3322 3273 3332
rect 3093 3288 3094 3322
rect 3128 3298 3166 3322
rect 3128 3288 3130 3298
rect 3093 3264 3130 3288
rect 3164 3288 3166 3298
rect 3200 3298 3238 3322
rect 3200 3288 3202 3298
rect 3164 3264 3202 3288
rect 3236 3288 3238 3298
rect 3272 3288 3273 3322
rect 3236 3264 3273 3288
rect 3093 3248 3273 3264
rect 3093 3214 3094 3248
rect 3128 3230 3166 3248
rect 3128 3214 3130 3230
rect 3093 3196 3130 3214
rect 3164 3214 3166 3230
rect 3200 3230 3238 3248
rect 3200 3214 3202 3230
rect 3164 3196 3202 3214
rect 3236 3214 3238 3230
rect 3272 3214 3273 3248
rect 3236 3196 3273 3214
rect 3093 3174 3273 3196
rect 3093 3140 3094 3174
rect 3128 3162 3166 3174
rect 3128 3140 3130 3162
rect 3093 3128 3130 3140
rect 3164 3140 3166 3162
rect 3200 3162 3238 3174
rect 3200 3140 3202 3162
rect 3164 3128 3202 3140
rect 3236 3140 3238 3162
rect 3272 3140 3273 3174
rect 3236 3128 3273 3140
rect 3093 3100 3273 3128
rect 3093 3066 3094 3100
rect 3128 3066 3166 3100
rect 3200 3066 3238 3100
rect 3272 3066 3273 3100
rect 3093 3026 3273 3066
rect 3093 2992 3094 3026
rect 3128 2992 3166 3026
rect 3200 2992 3238 3026
rect 3272 2992 3273 3026
rect 3093 2952 3273 2992
rect 3093 2918 3094 2952
rect 3128 2918 3166 2952
rect 3200 2918 3238 2952
rect 3272 2918 3273 2952
rect 3093 2878 3273 2918
rect 3093 2844 3094 2878
rect 3128 2844 3166 2878
rect 3200 2844 3238 2878
rect 3272 2844 3273 2878
rect 3093 2804 3273 2844
rect 3093 2770 3094 2804
rect 3128 2770 3166 2804
rect 3200 2770 3238 2804
rect 3272 2770 3273 2804
rect 3093 2730 3273 2770
rect 3093 2696 3094 2730
rect 3128 2696 3166 2730
rect 3200 2696 3238 2730
rect 3272 2696 3273 2730
rect 3093 2656 3273 2696
rect 3093 2622 3094 2656
rect 3128 2622 3166 2656
rect 3200 2622 3238 2656
rect 3272 2622 3273 2656
rect 3093 2582 3273 2622
rect 3093 2548 3094 2582
rect 3128 2548 3166 2582
rect 3200 2548 3238 2582
rect 3272 2548 3273 2582
rect 3093 2508 3273 2548
rect 3093 2474 3094 2508
rect 3128 2474 3166 2508
rect 3200 2474 3238 2508
rect 3272 2474 3273 2508
rect 3093 2445 3273 2474
rect 3093 2434 3130 2445
rect 3093 2400 3094 2434
rect 3128 2411 3130 2434
rect 3164 2434 3202 2445
rect 3164 2411 3166 2434
rect 3128 2400 3166 2411
rect 3200 2411 3202 2434
rect 3236 2434 3273 2445
rect 3236 2411 3238 2434
rect 3200 2400 3238 2411
rect 3272 2400 3273 2434
rect 3093 2377 3273 2400
rect 3093 2360 3130 2377
rect 3093 2326 3094 2360
rect 3128 2343 3130 2360
rect 3164 2360 3202 2377
rect 3164 2343 3166 2360
rect 3128 2326 3166 2343
rect 3200 2343 3202 2360
rect 3236 2360 3273 2377
rect 3236 2343 3238 2360
rect 3200 2326 3238 2343
rect 3272 2326 3273 2360
rect 3093 2309 3273 2326
rect 3093 2286 3130 2309
rect 3093 2252 3094 2286
rect 3128 2275 3130 2286
rect 3164 2286 3202 2309
rect 3164 2275 3166 2286
rect 3128 2252 3166 2275
rect 3200 2275 3202 2286
rect 3236 2286 3273 2309
rect 3236 2275 3238 2286
rect 3200 2252 3238 2275
rect 3272 2252 3273 2286
rect 3093 2241 3273 2252
rect 3093 2212 3130 2241
rect 3093 2178 3094 2212
rect 3128 2207 3130 2212
rect 3164 2212 3202 2241
rect 3164 2207 3166 2212
rect 3128 2178 3166 2207
rect 3200 2207 3202 2212
rect 3236 2212 3273 2241
rect 3236 2207 3238 2212
rect 3200 2178 3238 2207
rect 3272 2178 3273 2212
rect 3093 2173 3273 2178
rect 3093 2139 3130 2173
rect 3164 2139 3202 2173
rect 3236 2139 3273 2173
rect 3093 2138 3273 2139
rect 3093 2104 3094 2138
rect 3128 2105 3166 2138
rect 3128 2104 3130 2105
rect 3093 2071 3130 2104
rect 3164 2104 3166 2105
rect 3200 2105 3238 2138
rect 3200 2104 3202 2105
rect 3164 2071 3202 2104
rect 3236 2104 3238 2105
rect 3272 2104 3273 2138
rect 3236 2071 3273 2104
rect 3093 2064 3273 2071
rect 3093 2030 3094 2064
rect 3128 2037 3166 2064
rect 3128 2030 3130 2037
rect 3093 2003 3130 2030
rect 3164 2030 3166 2037
rect 3200 2037 3238 2064
rect 3200 2030 3202 2037
rect 3164 2003 3202 2030
rect 3236 2030 3238 2037
rect 3272 2030 3273 2064
rect 3236 2003 3273 2030
rect 3093 1990 3273 2003
rect 3093 1956 3094 1990
rect 3128 1969 3166 1990
rect 3128 1956 3130 1969
rect 3093 1935 3130 1956
rect 3164 1956 3166 1969
rect 3200 1969 3238 1990
rect 3200 1956 3202 1969
rect 3164 1935 3202 1956
rect 3236 1956 3238 1969
rect 3272 1956 3273 1990
rect 3236 1935 3273 1956
rect 3093 1916 3273 1935
rect 3093 1882 3094 1916
rect 3128 1901 3166 1916
rect 3128 1882 3130 1901
rect 3093 1867 3130 1882
rect 3164 1882 3166 1901
rect 3200 1901 3238 1916
rect 3200 1882 3202 1901
rect 3164 1867 3202 1882
rect 3236 1882 3238 1901
rect 3272 1882 3273 1916
rect 3236 1867 3273 1882
rect 3093 1842 3273 1867
rect 3093 1808 3094 1842
rect 3128 1833 3166 1842
rect 3128 1808 3130 1833
rect 3093 1799 3130 1808
rect 3164 1808 3166 1833
rect 3200 1833 3238 1842
rect 3200 1808 3202 1833
rect 3164 1799 3202 1808
rect 3236 1808 3238 1833
rect 3272 1808 3273 1842
rect 3236 1799 3273 1808
rect 3093 1768 3273 1799
rect 3093 1734 3094 1768
rect 3128 1765 3166 1768
rect 3128 1734 3130 1765
rect 3093 1731 3130 1734
rect 3164 1734 3166 1765
rect 3200 1765 3238 1768
rect 3200 1734 3202 1765
rect 3164 1731 3202 1734
rect 3236 1734 3238 1765
rect 3272 1734 3273 1768
rect 3236 1731 3273 1734
rect 3093 1697 3273 1731
rect 3093 1694 3130 1697
rect 3093 1660 3094 1694
rect 3128 1663 3130 1694
rect 3164 1694 3202 1697
rect 3164 1663 3166 1694
rect 3128 1660 3166 1663
rect 3200 1663 3202 1694
rect 3236 1694 3273 1697
rect 3236 1663 3238 1694
rect 3200 1660 3238 1663
rect 3272 1660 3273 1694
rect 3093 1629 3273 1660
rect 3093 1620 3130 1629
rect 3093 1586 3094 1620
rect 3128 1595 3130 1620
rect 3164 1620 3202 1629
rect 3164 1595 3166 1620
rect 3128 1586 3166 1595
rect 3200 1595 3202 1620
rect 3236 1620 3273 1629
rect 3236 1595 3238 1620
rect 3200 1586 3238 1595
rect 3272 1586 3273 1620
rect 3093 1561 3273 1586
rect 3093 1545 3130 1561
rect 3093 1511 3094 1545
rect 3128 1527 3130 1545
rect 3164 1545 3202 1561
rect 3164 1527 3166 1545
rect 3128 1511 3166 1527
rect 3200 1527 3202 1545
rect 3236 1545 3273 1561
rect 3236 1527 3238 1545
rect 3200 1511 3238 1527
rect 3272 1511 3273 1545
rect 3338 3010 3458 4106
rect 3900 4388 3907 4494
rect 4013 4388 4020 4494
rect 3900 4214 4020 4388
rect 3900 4180 3943 4214
rect 3977 4180 4020 4214
rect 3900 4140 4020 4180
rect 3900 4106 3943 4140
rect 3977 4106 4020 4140
rect 3338 2976 3381 3010
rect 3415 2976 3458 3010
rect 3338 2932 3458 2976
rect 3338 2898 3381 2932
rect 3415 2898 3458 2932
rect 3338 2854 3458 2898
rect 3338 2820 3381 2854
rect 3415 2820 3458 2854
rect 3338 2776 3458 2820
rect 3338 2742 3381 2776
rect 3415 2742 3458 2776
rect 3338 2697 3458 2742
rect 3338 2663 3381 2697
rect 3415 2663 3458 2697
rect 3338 2618 3458 2663
rect 3338 2584 3381 2618
rect 3415 2584 3458 2618
rect 3338 2539 3458 2584
rect 3338 2505 3381 2539
rect 3415 2505 3458 2539
rect 3130 1491 3236 1511
rect 2908 1375 2951 1409
rect 2985 1375 3028 1409
rect 2908 1335 3028 1375
rect 2908 1301 2951 1335
rect 2985 1301 3028 1335
rect 2908 1285 3028 1301
rect 3338 1409 3458 2505
rect 3560 4050 3662 4062
rect 3696 4050 3798 4062
rect 3560 4046 3590 4050
rect 3768 4046 3798 4050
rect 3560 3978 3590 4012
rect 3768 3978 3798 4012
rect 3560 3910 3590 3944
rect 3768 3910 3798 3944
rect 3560 3842 3590 3876
rect 3768 3842 3798 3876
rect 3560 3774 3590 3808
rect 3768 3774 3798 3808
rect 3560 3706 3590 3740
rect 3768 3706 3798 3740
rect 3560 3638 3590 3672
rect 3768 3638 3798 3672
rect 3560 3570 3590 3604
rect 3768 3570 3798 3604
rect 3560 3502 3590 3536
rect 3768 3502 3798 3536
rect 3560 3434 3590 3468
rect 3768 3434 3798 3468
rect 3560 3366 3590 3400
rect 3768 3366 3798 3400
rect 3560 3298 3590 3332
rect 3768 3298 3798 3332
rect 3560 3230 3590 3264
rect 3768 3230 3798 3264
rect 3560 3162 3590 3196
rect 3768 3162 3798 3196
rect 3560 3080 3590 3128
rect 3624 3080 3734 3092
rect 3768 3080 3798 3128
rect 3560 3040 3798 3080
rect 3560 2574 3590 3040
rect 3768 2574 3798 3040
rect 3560 2535 3798 2574
rect 3560 2501 3590 2535
rect 3624 2501 3662 2535
rect 3696 2501 3734 2535
rect 3768 2501 3798 2535
rect 3560 2461 3798 2501
rect 3560 2449 3662 2461
rect 3696 2449 3798 2461
rect 3560 2445 3590 2449
rect 3768 2445 3798 2449
rect 3560 2377 3590 2411
rect 3768 2377 3798 2411
rect 3560 2309 3590 2343
rect 3768 2309 3798 2343
rect 3560 2241 3590 2275
rect 3768 2241 3798 2275
rect 3560 2173 3590 2207
rect 3768 2173 3798 2207
rect 3560 2105 3590 2139
rect 3768 2105 3798 2139
rect 3560 2037 3590 2071
rect 3768 2037 3798 2071
rect 3560 1969 3590 2003
rect 3768 1969 3798 2003
rect 3560 1901 3590 1935
rect 3768 1901 3798 1935
rect 3560 1833 3590 1867
rect 3768 1833 3798 1867
rect 3560 1765 3590 1799
rect 3768 1765 3798 1799
rect 3560 1697 3590 1731
rect 3768 1697 3798 1731
rect 3560 1629 3590 1663
rect 3768 1629 3798 1663
rect 3560 1561 3590 1595
rect 3768 1561 3798 1595
rect 3560 1479 3590 1527
rect 3624 1479 3734 1491
rect 3768 1479 3798 1527
rect 3560 1464 3798 1479
rect 3900 3010 4020 4106
rect 4330 4388 4337 4494
rect 4443 4388 4450 4494
rect 4330 4214 4450 4388
rect 4330 4180 4373 4214
rect 4407 4180 4450 4214
rect 4330 4140 4450 4180
rect 4330 4106 4373 4140
rect 4407 4106 4450 4140
rect 3900 2976 3943 3010
rect 3977 2976 4020 3010
rect 3900 2932 4020 2976
rect 3900 2898 3943 2932
rect 3977 2898 4020 2932
rect 3900 2854 4020 2898
rect 3900 2820 3943 2854
rect 3977 2820 4020 2854
rect 3900 2776 4020 2820
rect 3900 2742 3943 2776
rect 3977 2742 4020 2776
rect 3900 2697 4020 2742
rect 3900 2663 3943 2697
rect 3977 2663 4020 2697
rect 3900 2618 4020 2663
rect 3900 2584 3943 2618
rect 3977 2584 4020 2618
rect 3900 2539 4020 2584
rect 3900 2505 3943 2539
rect 3977 2505 4020 2539
rect 3338 1375 3381 1409
rect 3415 1375 3458 1409
rect 3338 1335 3458 1375
rect 3338 1301 3381 1335
rect 3415 1301 3458 1335
rect 3338 1285 3458 1301
rect 3900 1409 4020 2505
rect 4085 4028 4086 4062
rect 4120 4046 4158 4062
rect 4120 4028 4122 4046
rect 4085 4012 4122 4028
rect 4156 4028 4158 4046
rect 4192 4046 4230 4062
rect 4192 4028 4194 4046
rect 4156 4012 4194 4028
rect 4228 4028 4230 4046
rect 4264 4028 4265 4062
rect 4228 4012 4265 4028
rect 4085 3988 4265 4012
rect 4085 3954 4086 3988
rect 4120 3978 4158 3988
rect 4120 3954 4122 3978
rect 4085 3944 4122 3954
rect 4156 3954 4158 3978
rect 4192 3978 4230 3988
rect 4192 3954 4194 3978
rect 4156 3944 4194 3954
rect 4228 3954 4230 3978
rect 4264 3954 4265 3988
rect 4228 3944 4265 3954
rect 4085 3914 4265 3944
rect 4085 3880 4086 3914
rect 4120 3910 4158 3914
rect 4120 3880 4122 3910
rect 4085 3876 4122 3880
rect 4156 3880 4158 3910
rect 4192 3910 4230 3914
rect 4192 3880 4194 3910
rect 4156 3876 4194 3880
rect 4228 3880 4230 3910
rect 4264 3880 4265 3914
rect 4228 3876 4265 3880
rect 4085 3842 4265 3876
rect 4085 3840 4122 3842
rect 4085 3806 4086 3840
rect 4120 3808 4122 3840
rect 4156 3840 4194 3842
rect 4156 3808 4158 3840
rect 4120 3806 4158 3808
rect 4192 3808 4194 3840
rect 4228 3840 4265 3842
rect 4228 3808 4230 3840
rect 4192 3806 4230 3808
rect 4264 3806 4265 3840
rect 4085 3774 4265 3806
rect 4085 3766 4122 3774
rect 4085 3732 4086 3766
rect 4120 3740 4122 3766
rect 4156 3766 4194 3774
rect 4156 3740 4158 3766
rect 4120 3732 4158 3740
rect 4192 3740 4194 3766
rect 4228 3766 4265 3774
rect 4228 3740 4230 3766
rect 4192 3732 4230 3740
rect 4264 3732 4265 3766
rect 4085 3706 4265 3732
rect 4085 3692 4122 3706
rect 4085 3658 4086 3692
rect 4120 3672 4122 3692
rect 4156 3692 4194 3706
rect 4156 3672 4158 3692
rect 4120 3658 4158 3672
rect 4192 3672 4194 3692
rect 4228 3692 4265 3706
rect 4228 3672 4230 3692
rect 4192 3658 4230 3672
rect 4264 3658 4265 3692
rect 4085 3638 4265 3658
rect 4085 3618 4122 3638
rect 4085 3584 4086 3618
rect 4120 3604 4122 3618
rect 4156 3618 4194 3638
rect 4156 3604 4158 3618
rect 4120 3584 4158 3604
rect 4192 3604 4194 3618
rect 4228 3618 4265 3638
rect 4228 3604 4230 3618
rect 4192 3584 4230 3604
rect 4264 3584 4265 3618
rect 4085 3570 4265 3584
rect 4085 3544 4122 3570
rect 4085 3510 4086 3544
rect 4120 3536 4122 3544
rect 4156 3544 4194 3570
rect 4156 3536 4158 3544
rect 4120 3510 4158 3536
rect 4192 3536 4194 3544
rect 4228 3544 4265 3570
rect 4228 3536 4230 3544
rect 4192 3510 4230 3536
rect 4264 3510 4265 3544
rect 4085 3502 4265 3510
rect 4085 3470 4122 3502
rect 4085 3436 4086 3470
rect 4120 3468 4122 3470
rect 4156 3470 4194 3502
rect 4156 3468 4158 3470
rect 4120 3436 4158 3468
rect 4192 3468 4194 3470
rect 4228 3470 4265 3502
rect 4228 3468 4230 3470
rect 4192 3436 4230 3468
rect 4264 3436 4265 3470
rect 4085 3434 4265 3436
rect 4085 3400 4122 3434
rect 4156 3400 4194 3434
rect 4228 3400 4265 3434
rect 4085 3396 4265 3400
rect 4085 3362 4086 3396
rect 4120 3366 4158 3396
rect 4120 3362 4122 3366
rect 4085 3332 4122 3362
rect 4156 3362 4158 3366
rect 4192 3366 4230 3396
rect 4192 3362 4194 3366
rect 4156 3332 4194 3362
rect 4228 3362 4230 3366
rect 4264 3362 4265 3396
rect 4228 3332 4265 3362
rect 4085 3322 4265 3332
rect 4085 3288 4086 3322
rect 4120 3298 4158 3322
rect 4120 3288 4122 3298
rect 4085 3264 4122 3288
rect 4156 3288 4158 3298
rect 4192 3298 4230 3322
rect 4192 3288 4194 3298
rect 4156 3264 4194 3288
rect 4228 3288 4230 3298
rect 4264 3288 4265 3322
rect 4228 3264 4265 3288
rect 4085 3248 4265 3264
rect 4085 3214 4086 3248
rect 4120 3230 4158 3248
rect 4120 3214 4122 3230
rect 4085 3196 4122 3214
rect 4156 3214 4158 3230
rect 4192 3230 4230 3248
rect 4192 3214 4194 3230
rect 4156 3196 4194 3214
rect 4228 3214 4230 3230
rect 4264 3214 4265 3248
rect 4228 3196 4265 3214
rect 4085 3174 4265 3196
rect 4085 3140 4086 3174
rect 4120 3162 4158 3174
rect 4120 3140 4122 3162
rect 4085 3128 4122 3140
rect 4156 3140 4158 3162
rect 4192 3162 4230 3174
rect 4192 3140 4194 3162
rect 4156 3128 4194 3140
rect 4228 3140 4230 3162
rect 4264 3140 4265 3174
rect 4228 3128 4265 3140
rect 4085 3100 4265 3128
rect 4085 3066 4086 3100
rect 4120 3066 4158 3100
rect 4192 3066 4230 3100
rect 4264 3066 4265 3100
rect 4085 3026 4265 3066
rect 4085 2992 4086 3026
rect 4120 2992 4158 3026
rect 4192 2992 4230 3026
rect 4264 2992 4265 3026
rect 4085 2952 4265 2992
rect 4085 2918 4086 2952
rect 4120 2918 4158 2952
rect 4192 2918 4230 2952
rect 4264 2918 4265 2952
rect 4085 2878 4265 2918
rect 4085 2844 4086 2878
rect 4120 2844 4158 2878
rect 4192 2844 4230 2878
rect 4264 2844 4265 2878
rect 4085 2804 4265 2844
rect 4085 2770 4086 2804
rect 4120 2770 4158 2804
rect 4192 2770 4230 2804
rect 4264 2770 4265 2804
rect 4085 2730 4265 2770
rect 4085 2696 4086 2730
rect 4120 2696 4158 2730
rect 4192 2696 4230 2730
rect 4264 2696 4265 2730
rect 4085 2656 4265 2696
rect 4085 2622 4086 2656
rect 4120 2622 4158 2656
rect 4192 2622 4230 2656
rect 4264 2622 4265 2656
rect 4085 2582 4265 2622
rect 4085 2548 4086 2582
rect 4120 2548 4158 2582
rect 4192 2548 4230 2582
rect 4264 2548 4265 2582
rect 4085 2508 4265 2548
rect 4085 2474 4086 2508
rect 4120 2474 4158 2508
rect 4192 2474 4230 2508
rect 4264 2474 4265 2508
rect 4085 2445 4265 2474
rect 4085 2434 4122 2445
rect 4085 2400 4086 2434
rect 4120 2411 4122 2434
rect 4156 2434 4194 2445
rect 4156 2411 4158 2434
rect 4120 2400 4158 2411
rect 4192 2411 4194 2434
rect 4228 2434 4265 2445
rect 4228 2411 4230 2434
rect 4192 2400 4230 2411
rect 4264 2400 4265 2434
rect 4085 2377 4265 2400
rect 4085 2360 4122 2377
rect 4085 2326 4086 2360
rect 4120 2343 4122 2360
rect 4156 2360 4194 2377
rect 4156 2343 4158 2360
rect 4120 2326 4158 2343
rect 4192 2343 4194 2360
rect 4228 2360 4265 2377
rect 4228 2343 4230 2360
rect 4192 2326 4230 2343
rect 4264 2326 4265 2360
rect 4085 2309 4265 2326
rect 4085 2286 4122 2309
rect 4085 2252 4086 2286
rect 4120 2275 4122 2286
rect 4156 2286 4194 2309
rect 4156 2275 4158 2286
rect 4120 2252 4158 2275
rect 4192 2275 4194 2286
rect 4228 2286 4265 2309
rect 4228 2275 4230 2286
rect 4192 2252 4230 2275
rect 4264 2252 4265 2286
rect 4085 2241 4265 2252
rect 4085 2212 4122 2241
rect 4085 2178 4086 2212
rect 4120 2207 4122 2212
rect 4156 2212 4194 2241
rect 4156 2207 4158 2212
rect 4120 2178 4158 2207
rect 4192 2207 4194 2212
rect 4228 2212 4265 2241
rect 4228 2207 4230 2212
rect 4192 2178 4230 2207
rect 4264 2178 4265 2212
rect 4085 2173 4265 2178
rect 4085 2139 4122 2173
rect 4156 2139 4194 2173
rect 4228 2139 4265 2173
rect 4085 2138 4265 2139
rect 4085 2104 4086 2138
rect 4120 2105 4158 2138
rect 4120 2104 4122 2105
rect 4085 2071 4122 2104
rect 4156 2104 4158 2105
rect 4192 2105 4230 2138
rect 4192 2104 4194 2105
rect 4156 2071 4194 2104
rect 4228 2104 4230 2105
rect 4264 2104 4265 2138
rect 4228 2071 4265 2104
rect 4085 2064 4265 2071
rect 4085 2030 4086 2064
rect 4120 2037 4158 2064
rect 4120 2030 4122 2037
rect 4085 2003 4122 2030
rect 4156 2030 4158 2037
rect 4192 2037 4230 2064
rect 4192 2030 4194 2037
rect 4156 2003 4194 2030
rect 4228 2030 4230 2037
rect 4264 2030 4265 2064
rect 4228 2003 4265 2030
rect 4085 1990 4265 2003
rect 4085 1956 4086 1990
rect 4120 1969 4158 1990
rect 4120 1956 4122 1969
rect 4085 1935 4122 1956
rect 4156 1956 4158 1969
rect 4192 1969 4230 1990
rect 4192 1956 4194 1969
rect 4156 1935 4194 1956
rect 4228 1956 4230 1969
rect 4264 1956 4265 1990
rect 4228 1935 4265 1956
rect 4085 1916 4265 1935
rect 4085 1882 4086 1916
rect 4120 1901 4158 1916
rect 4120 1882 4122 1901
rect 4085 1867 4122 1882
rect 4156 1882 4158 1901
rect 4192 1901 4230 1916
rect 4192 1882 4194 1901
rect 4156 1867 4194 1882
rect 4228 1882 4230 1901
rect 4264 1882 4265 1916
rect 4228 1867 4265 1882
rect 4085 1842 4265 1867
rect 4085 1808 4086 1842
rect 4120 1833 4158 1842
rect 4120 1808 4122 1833
rect 4085 1799 4122 1808
rect 4156 1808 4158 1833
rect 4192 1833 4230 1842
rect 4192 1808 4194 1833
rect 4156 1799 4194 1808
rect 4228 1808 4230 1833
rect 4264 1808 4265 1842
rect 4228 1799 4265 1808
rect 4085 1768 4265 1799
rect 4085 1734 4086 1768
rect 4120 1765 4158 1768
rect 4120 1734 4122 1765
rect 4085 1731 4122 1734
rect 4156 1734 4158 1765
rect 4192 1765 4230 1768
rect 4192 1734 4194 1765
rect 4156 1731 4194 1734
rect 4228 1734 4230 1765
rect 4264 1734 4265 1768
rect 4228 1731 4265 1734
rect 4085 1697 4265 1731
rect 4085 1694 4122 1697
rect 4085 1660 4086 1694
rect 4120 1663 4122 1694
rect 4156 1694 4194 1697
rect 4156 1663 4158 1694
rect 4120 1660 4158 1663
rect 4192 1663 4194 1694
rect 4228 1694 4265 1697
rect 4228 1663 4230 1694
rect 4192 1660 4230 1663
rect 4264 1660 4265 1694
rect 4085 1629 4265 1660
rect 4085 1620 4122 1629
rect 4085 1586 4086 1620
rect 4120 1595 4122 1620
rect 4156 1620 4194 1629
rect 4156 1595 4158 1620
rect 4120 1586 4158 1595
rect 4192 1595 4194 1620
rect 4228 1620 4265 1629
rect 4228 1595 4230 1620
rect 4192 1586 4230 1595
rect 4264 1586 4265 1620
rect 4085 1561 4265 1586
rect 4085 1545 4122 1561
rect 4085 1511 4086 1545
rect 4120 1527 4122 1545
rect 4156 1545 4194 1561
rect 4156 1527 4158 1545
rect 4120 1511 4158 1527
rect 4192 1527 4194 1545
rect 4228 1545 4265 1561
rect 4228 1527 4230 1545
rect 4192 1511 4230 1527
rect 4264 1511 4265 1545
rect 4330 3010 4450 4106
rect 4892 4388 4899 4494
rect 5005 4388 5012 4494
rect 4892 4214 5012 4388
rect 4892 4180 4935 4214
rect 4969 4180 5012 4214
rect 4892 4140 5012 4180
rect 4892 4106 4935 4140
rect 4969 4106 5012 4140
rect 4330 2976 4373 3010
rect 4407 2976 4450 3010
rect 4330 2932 4450 2976
rect 4330 2898 4373 2932
rect 4407 2898 4450 2932
rect 4330 2854 4450 2898
rect 4330 2820 4373 2854
rect 4407 2820 4450 2854
rect 4330 2776 4450 2820
rect 4330 2742 4373 2776
rect 4407 2742 4450 2776
rect 4330 2697 4450 2742
rect 4330 2663 4373 2697
rect 4407 2663 4450 2697
rect 4330 2618 4450 2663
rect 4330 2584 4373 2618
rect 4407 2584 4450 2618
rect 4330 2539 4450 2584
rect 4330 2505 4373 2539
rect 4407 2505 4450 2539
rect 4122 1491 4228 1511
rect 3900 1375 3943 1409
rect 3977 1375 4020 1409
rect 3900 1335 4020 1375
rect 3900 1301 3943 1335
rect 3977 1301 4020 1335
rect 3900 1285 4020 1301
rect 4330 1409 4450 2505
rect 4552 4050 4654 4062
rect 4688 4050 4790 4062
rect 4552 4046 4582 4050
rect 4760 4046 4790 4050
rect 4552 3978 4582 4012
rect 4760 3978 4790 4012
rect 4552 3910 4582 3944
rect 4760 3910 4790 3944
rect 4552 3842 4582 3876
rect 4760 3842 4790 3876
rect 4552 3774 4582 3808
rect 4760 3774 4790 3808
rect 4552 3706 4582 3740
rect 4760 3706 4790 3740
rect 4552 3638 4582 3672
rect 4760 3638 4790 3672
rect 4552 3570 4582 3604
rect 4760 3570 4790 3604
rect 4552 3502 4582 3536
rect 4760 3502 4790 3536
rect 4552 3434 4582 3468
rect 4760 3434 4790 3468
rect 4552 3366 4582 3400
rect 4760 3366 4790 3400
rect 4552 3298 4582 3332
rect 4760 3298 4790 3332
rect 4552 3230 4582 3264
rect 4760 3230 4790 3264
rect 4552 3162 4582 3196
rect 4760 3162 4790 3196
rect 4552 3080 4582 3128
rect 4616 3080 4726 3092
rect 4760 3080 4790 3128
rect 4552 3040 4790 3080
rect 4552 2574 4582 3040
rect 4760 2574 4790 3040
rect 4552 2535 4790 2574
rect 4552 2501 4582 2535
rect 4616 2501 4654 2535
rect 4688 2501 4726 2535
rect 4760 2501 4790 2535
rect 4552 2461 4790 2501
rect 4552 2449 4654 2461
rect 4688 2449 4790 2461
rect 4552 2445 4582 2449
rect 4760 2445 4790 2449
rect 4552 2377 4582 2411
rect 4760 2377 4790 2411
rect 4552 2309 4582 2343
rect 4760 2309 4790 2343
rect 4552 2241 4582 2275
rect 4760 2241 4790 2275
rect 4552 2173 4582 2207
rect 4760 2173 4790 2207
rect 4552 2105 4582 2139
rect 4760 2105 4790 2139
rect 4552 2037 4582 2071
rect 4760 2037 4790 2071
rect 4552 1969 4582 2003
rect 4760 1969 4790 2003
rect 4552 1901 4582 1935
rect 4760 1901 4790 1935
rect 4552 1833 4582 1867
rect 4760 1833 4790 1867
rect 4552 1765 4582 1799
rect 4760 1765 4790 1799
rect 4552 1697 4582 1731
rect 4760 1697 4790 1731
rect 4552 1629 4582 1663
rect 4760 1629 4790 1663
rect 4552 1561 4582 1595
rect 4760 1561 4790 1595
rect 4552 1479 4582 1527
rect 4616 1479 4726 1491
rect 4760 1479 4790 1527
rect 4552 1464 4790 1479
rect 4892 3010 5012 4106
rect 5322 4388 5329 4494
rect 5435 4388 5442 4494
rect 5322 4214 5442 4388
rect 5322 4180 5365 4214
rect 5399 4180 5442 4214
rect 5322 4140 5442 4180
rect 5322 4106 5365 4140
rect 5399 4106 5442 4140
rect 4892 2976 4935 3010
rect 4969 2976 5012 3010
rect 4892 2932 5012 2976
rect 4892 2898 4935 2932
rect 4969 2898 5012 2932
rect 4892 2854 5012 2898
rect 4892 2820 4935 2854
rect 4969 2820 5012 2854
rect 4892 2776 5012 2820
rect 4892 2742 4935 2776
rect 4969 2742 5012 2776
rect 4892 2697 5012 2742
rect 4892 2663 4935 2697
rect 4969 2663 5012 2697
rect 4892 2618 5012 2663
rect 4892 2584 4935 2618
rect 4969 2584 5012 2618
rect 4892 2539 5012 2584
rect 4892 2505 4935 2539
rect 4969 2505 5012 2539
rect 4330 1375 4373 1409
rect 4407 1375 4450 1409
rect 4330 1335 4450 1375
rect 4330 1301 4373 1335
rect 4407 1301 4450 1335
rect 4330 1285 4450 1301
rect 4892 1409 5012 2505
rect 5077 4028 5078 4062
rect 5112 4046 5150 4062
rect 5112 4028 5114 4046
rect 5077 4012 5114 4028
rect 5148 4028 5150 4046
rect 5184 4046 5222 4062
rect 5184 4028 5186 4046
rect 5148 4012 5186 4028
rect 5220 4028 5222 4046
rect 5256 4028 5257 4062
rect 5220 4012 5257 4028
rect 5077 3988 5257 4012
rect 5077 3954 5078 3988
rect 5112 3978 5150 3988
rect 5112 3954 5114 3978
rect 5077 3944 5114 3954
rect 5148 3954 5150 3978
rect 5184 3978 5222 3988
rect 5184 3954 5186 3978
rect 5148 3944 5186 3954
rect 5220 3954 5222 3978
rect 5256 3954 5257 3988
rect 5220 3944 5257 3954
rect 5077 3914 5257 3944
rect 5077 3880 5078 3914
rect 5112 3910 5150 3914
rect 5112 3880 5114 3910
rect 5077 3876 5114 3880
rect 5148 3880 5150 3910
rect 5184 3910 5222 3914
rect 5184 3880 5186 3910
rect 5148 3876 5186 3880
rect 5220 3880 5222 3910
rect 5256 3880 5257 3914
rect 5220 3876 5257 3880
rect 5077 3842 5257 3876
rect 5077 3840 5114 3842
rect 5077 3806 5078 3840
rect 5112 3808 5114 3840
rect 5148 3840 5186 3842
rect 5148 3808 5150 3840
rect 5112 3806 5150 3808
rect 5184 3808 5186 3840
rect 5220 3840 5257 3842
rect 5220 3808 5222 3840
rect 5184 3806 5222 3808
rect 5256 3806 5257 3840
rect 5077 3774 5257 3806
rect 5077 3766 5114 3774
rect 5077 3732 5078 3766
rect 5112 3740 5114 3766
rect 5148 3766 5186 3774
rect 5148 3740 5150 3766
rect 5112 3732 5150 3740
rect 5184 3740 5186 3766
rect 5220 3766 5257 3774
rect 5220 3740 5222 3766
rect 5184 3732 5222 3740
rect 5256 3732 5257 3766
rect 5077 3706 5257 3732
rect 5077 3692 5114 3706
rect 5077 3658 5078 3692
rect 5112 3672 5114 3692
rect 5148 3692 5186 3706
rect 5148 3672 5150 3692
rect 5112 3658 5150 3672
rect 5184 3672 5186 3692
rect 5220 3692 5257 3706
rect 5220 3672 5222 3692
rect 5184 3658 5222 3672
rect 5256 3658 5257 3692
rect 5077 3638 5257 3658
rect 5077 3618 5114 3638
rect 5077 3584 5078 3618
rect 5112 3604 5114 3618
rect 5148 3618 5186 3638
rect 5148 3604 5150 3618
rect 5112 3584 5150 3604
rect 5184 3604 5186 3618
rect 5220 3618 5257 3638
rect 5220 3604 5222 3618
rect 5184 3584 5222 3604
rect 5256 3584 5257 3618
rect 5077 3570 5257 3584
rect 5077 3544 5114 3570
rect 5077 3510 5078 3544
rect 5112 3536 5114 3544
rect 5148 3544 5186 3570
rect 5148 3536 5150 3544
rect 5112 3510 5150 3536
rect 5184 3536 5186 3544
rect 5220 3544 5257 3570
rect 5220 3536 5222 3544
rect 5184 3510 5222 3536
rect 5256 3510 5257 3544
rect 5077 3502 5257 3510
rect 5077 3470 5114 3502
rect 5077 3436 5078 3470
rect 5112 3468 5114 3470
rect 5148 3470 5186 3502
rect 5148 3468 5150 3470
rect 5112 3436 5150 3468
rect 5184 3468 5186 3470
rect 5220 3470 5257 3502
rect 5220 3468 5222 3470
rect 5184 3436 5222 3468
rect 5256 3436 5257 3470
rect 5077 3434 5257 3436
rect 5077 3400 5114 3434
rect 5148 3400 5186 3434
rect 5220 3400 5257 3434
rect 5077 3396 5257 3400
rect 5077 3362 5078 3396
rect 5112 3366 5150 3396
rect 5112 3362 5114 3366
rect 5077 3332 5114 3362
rect 5148 3362 5150 3366
rect 5184 3366 5222 3396
rect 5184 3362 5186 3366
rect 5148 3332 5186 3362
rect 5220 3362 5222 3366
rect 5256 3362 5257 3396
rect 5220 3332 5257 3362
rect 5077 3322 5257 3332
rect 5077 3288 5078 3322
rect 5112 3298 5150 3322
rect 5112 3288 5114 3298
rect 5077 3264 5114 3288
rect 5148 3288 5150 3298
rect 5184 3298 5222 3322
rect 5184 3288 5186 3298
rect 5148 3264 5186 3288
rect 5220 3288 5222 3298
rect 5256 3288 5257 3322
rect 5220 3264 5257 3288
rect 5077 3248 5257 3264
rect 5077 3214 5078 3248
rect 5112 3230 5150 3248
rect 5112 3214 5114 3230
rect 5077 3196 5114 3214
rect 5148 3214 5150 3230
rect 5184 3230 5222 3248
rect 5184 3214 5186 3230
rect 5148 3196 5186 3214
rect 5220 3214 5222 3230
rect 5256 3214 5257 3248
rect 5220 3196 5257 3214
rect 5077 3174 5257 3196
rect 5077 3140 5078 3174
rect 5112 3162 5150 3174
rect 5112 3140 5114 3162
rect 5077 3128 5114 3140
rect 5148 3140 5150 3162
rect 5184 3162 5222 3174
rect 5184 3140 5186 3162
rect 5148 3128 5186 3140
rect 5220 3140 5222 3162
rect 5256 3140 5257 3174
rect 5220 3128 5257 3140
rect 5077 3100 5257 3128
rect 5077 3066 5078 3100
rect 5112 3066 5150 3100
rect 5184 3066 5222 3100
rect 5256 3066 5257 3100
rect 5077 3026 5257 3066
rect 5077 2992 5078 3026
rect 5112 2992 5150 3026
rect 5184 2992 5222 3026
rect 5256 2992 5257 3026
rect 5077 2952 5257 2992
rect 5077 2918 5078 2952
rect 5112 2918 5150 2952
rect 5184 2918 5222 2952
rect 5256 2918 5257 2952
rect 5077 2878 5257 2918
rect 5077 2844 5078 2878
rect 5112 2844 5150 2878
rect 5184 2844 5222 2878
rect 5256 2844 5257 2878
rect 5077 2804 5257 2844
rect 5077 2770 5078 2804
rect 5112 2770 5150 2804
rect 5184 2770 5222 2804
rect 5256 2770 5257 2804
rect 5077 2730 5257 2770
rect 5077 2696 5078 2730
rect 5112 2696 5150 2730
rect 5184 2696 5222 2730
rect 5256 2696 5257 2730
rect 5077 2656 5257 2696
rect 5077 2622 5078 2656
rect 5112 2622 5150 2656
rect 5184 2622 5222 2656
rect 5256 2622 5257 2656
rect 5077 2582 5257 2622
rect 5077 2548 5078 2582
rect 5112 2548 5150 2582
rect 5184 2548 5222 2582
rect 5256 2548 5257 2582
rect 5077 2508 5257 2548
rect 5077 2474 5078 2508
rect 5112 2474 5150 2508
rect 5184 2474 5222 2508
rect 5256 2474 5257 2508
rect 5077 2445 5257 2474
rect 5077 2434 5114 2445
rect 5077 2400 5078 2434
rect 5112 2411 5114 2434
rect 5148 2434 5186 2445
rect 5148 2411 5150 2434
rect 5112 2400 5150 2411
rect 5184 2411 5186 2434
rect 5220 2434 5257 2445
rect 5220 2411 5222 2434
rect 5184 2400 5222 2411
rect 5256 2400 5257 2434
rect 5077 2377 5257 2400
rect 5077 2360 5114 2377
rect 5077 2326 5078 2360
rect 5112 2343 5114 2360
rect 5148 2360 5186 2377
rect 5148 2343 5150 2360
rect 5112 2326 5150 2343
rect 5184 2343 5186 2360
rect 5220 2360 5257 2377
rect 5220 2343 5222 2360
rect 5184 2326 5222 2343
rect 5256 2326 5257 2360
rect 5077 2309 5257 2326
rect 5077 2286 5114 2309
rect 5077 2252 5078 2286
rect 5112 2275 5114 2286
rect 5148 2286 5186 2309
rect 5148 2275 5150 2286
rect 5112 2252 5150 2275
rect 5184 2275 5186 2286
rect 5220 2286 5257 2309
rect 5220 2275 5222 2286
rect 5184 2252 5222 2275
rect 5256 2252 5257 2286
rect 5077 2241 5257 2252
rect 5077 2212 5114 2241
rect 5077 2178 5078 2212
rect 5112 2207 5114 2212
rect 5148 2212 5186 2241
rect 5148 2207 5150 2212
rect 5112 2178 5150 2207
rect 5184 2207 5186 2212
rect 5220 2212 5257 2241
rect 5220 2207 5222 2212
rect 5184 2178 5222 2207
rect 5256 2178 5257 2212
rect 5077 2173 5257 2178
rect 5077 2139 5114 2173
rect 5148 2139 5186 2173
rect 5220 2139 5257 2173
rect 5077 2138 5257 2139
rect 5077 2104 5078 2138
rect 5112 2105 5150 2138
rect 5112 2104 5114 2105
rect 5077 2071 5114 2104
rect 5148 2104 5150 2105
rect 5184 2105 5222 2138
rect 5184 2104 5186 2105
rect 5148 2071 5186 2104
rect 5220 2104 5222 2105
rect 5256 2104 5257 2138
rect 5220 2071 5257 2104
rect 5077 2064 5257 2071
rect 5077 2030 5078 2064
rect 5112 2037 5150 2064
rect 5112 2030 5114 2037
rect 5077 2003 5114 2030
rect 5148 2030 5150 2037
rect 5184 2037 5222 2064
rect 5184 2030 5186 2037
rect 5148 2003 5186 2030
rect 5220 2030 5222 2037
rect 5256 2030 5257 2064
rect 5220 2003 5257 2030
rect 5077 1990 5257 2003
rect 5077 1956 5078 1990
rect 5112 1969 5150 1990
rect 5112 1956 5114 1969
rect 5077 1935 5114 1956
rect 5148 1956 5150 1969
rect 5184 1969 5222 1990
rect 5184 1956 5186 1969
rect 5148 1935 5186 1956
rect 5220 1956 5222 1969
rect 5256 1956 5257 1990
rect 5220 1935 5257 1956
rect 5077 1916 5257 1935
rect 5077 1882 5078 1916
rect 5112 1901 5150 1916
rect 5112 1882 5114 1901
rect 5077 1867 5114 1882
rect 5148 1882 5150 1901
rect 5184 1901 5222 1916
rect 5184 1882 5186 1901
rect 5148 1867 5186 1882
rect 5220 1882 5222 1901
rect 5256 1882 5257 1916
rect 5220 1867 5257 1882
rect 5077 1842 5257 1867
rect 5077 1808 5078 1842
rect 5112 1833 5150 1842
rect 5112 1808 5114 1833
rect 5077 1799 5114 1808
rect 5148 1808 5150 1833
rect 5184 1833 5222 1842
rect 5184 1808 5186 1833
rect 5148 1799 5186 1808
rect 5220 1808 5222 1833
rect 5256 1808 5257 1842
rect 5220 1799 5257 1808
rect 5077 1768 5257 1799
rect 5077 1734 5078 1768
rect 5112 1765 5150 1768
rect 5112 1734 5114 1765
rect 5077 1731 5114 1734
rect 5148 1734 5150 1765
rect 5184 1765 5222 1768
rect 5184 1734 5186 1765
rect 5148 1731 5186 1734
rect 5220 1734 5222 1765
rect 5256 1734 5257 1768
rect 5220 1731 5257 1734
rect 5077 1697 5257 1731
rect 5077 1694 5114 1697
rect 5077 1660 5078 1694
rect 5112 1663 5114 1694
rect 5148 1694 5186 1697
rect 5148 1663 5150 1694
rect 5112 1660 5150 1663
rect 5184 1663 5186 1694
rect 5220 1694 5257 1697
rect 5220 1663 5222 1694
rect 5184 1660 5222 1663
rect 5256 1660 5257 1694
rect 5077 1629 5257 1660
rect 5077 1620 5114 1629
rect 5077 1586 5078 1620
rect 5112 1595 5114 1620
rect 5148 1620 5186 1629
rect 5148 1595 5150 1620
rect 5112 1586 5150 1595
rect 5184 1595 5186 1620
rect 5220 1620 5257 1629
rect 5220 1595 5222 1620
rect 5184 1586 5222 1595
rect 5256 1586 5257 1620
rect 5077 1561 5257 1586
rect 5077 1545 5114 1561
rect 5077 1511 5078 1545
rect 5112 1527 5114 1545
rect 5148 1545 5186 1561
rect 5148 1527 5150 1545
rect 5112 1511 5150 1527
rect 5184 1527 5186 1545
rect 5220 1545 5257 1561
rect 5220 1527 5222 1545
rect 5184 1511 5222 1527
rect 5256 1511 5257 1545
rect 5322 3010 5442 4106
rect 5884 4388 5891 4494
rect 5997 4388 6004 4494
rect 5884 4214 6004 4388
rect 5884 4180 5927 4214
rect 5961 4180 6004 4214
rect 5884 4140 6004 4180
rect 5884 4106 5927 4140
rect 5961 4106 6004 4140
rect 5322 2976 5365 3010
rect 5399 2976 5442 3010
rect 5322 2932 5442 2976
rect 5322 2898 5365 2932
rect 5399 2898 5442 2932
rect 5322 2854 5442 2898
rect 5322 2820 5365 2854
rect 5399 2820 5442 2854
rect 5322 2776 5442 2820
rect 5322 2742 5365 2776
rect 5399 2742 5442 2776
rect 5322 2697 5442 2742
rect 5322 2663 5365 2697
rect 5399 2663 5442 2697
rect 5322 2618 5442 2663
rect 5322 2584 5365 2618
rect 5399 2584 5442 2618
rect 5322 2539 5442 2584
rect 5322 2505 5365 2539
rect 5399 2505 5442 2539
rect 5114 1491 5220 1511
rect 4892 1375 4935 1409
rect 4969 1375 5012 1409
rect 4892 1335 5012 1375
rect 4892 1301 4935 1335
rect 4969 1301 5012 1335
rect 4892 1285 5012 1301
rect 5322 1409 5442 2505
rect 5544 4050 5646 4062
rect 5680 4050 5782 4062
rect 5544 4046 5574 4050
rect 5752 4046 5782 4050
rect 5544 3978 5574 4012
rect 5752 3978 5782 4012
rect 5544 3910 5574 3944
rect 5752 3910 5782 3944
rect 5544 3842 5574 3876
rect 5752 3842 5782 3876
rect 5544 3774 5574 3808
rect 5752 3774 5782 3808
rect 5544 3706 5574 3740
rect 5752 3706 5782 3740
rect 5544 3638 5574 3672
rect 5752 3638 5782 3672
rect 5544 3570 5574 3604
rect 5752 3570 5782 3604
rect 5544 3502 5574 3536
rect 5752 3502 5782 3536
rect 5544 3434 5574 3468
rect 5752 3434 5782 3468
rect 5544 3366 5574 3400
rect 5752 3366 5782 3400
rect 5544 3298 5574 3332
rect 5752 3298 5782 3332
rect 5544 3230 5574 3264
rect 5752 3230 5782 3264
rect 5544 3162 5574 3196
rect 5752 3162 5782 3196
rect 5544 3080 5574 3128
rect 5608 3080 5718 3092
rect 5752 3080 5782 3128
rect 5544 3040 5782 3080
rect 5544 2574 5574 3040
rect 5752 2574 5782 3040
rect 5544 2535 5782 2574
rect 5544 2501 5574 2535
rect 5608 2501 5646 2535
rect 5680 2501 5718 2535
rect 5752 2501 5782 2535
rect 5544 2461 5782 2501
rect 5544 2449 5646 2461
rect 5680 2449 5782 2461
rect 5544 2445 5574 2449
rect 5752 2445 5782 2449
rect 5544 2377 5574 2411
rect 5752 2377 5782 2411
rect 5544 2309 5574 2343
rect 5752 2309 5782 2343
rect 5544 2241 5574 2275
rect 5752 2241 5782 2275
rect 5544 2173 5574 2207
rect 5752 2173 5782 2207
rect 5544 2105 5574 2139
rect 5752 2105 5782 2139
rect 5544 2037 5574 2071
rect 5752 2037 5782 2071
rect 5544 1969 5574 2003
rect 5752 1969 5782 2003
rect 5544 1901 5574 1935
rect 5752 1901 5782 1935
rect 5544 1833 5574 1867
rect 5752 1833 5782 1867
rect 5544 1765 5574 1799
rect 5752 1765 5782 1799
rect 5544 1697 5574 1731
rect 5752 1697 5782 1731
rect 5544 1629 5574 1663
rect 5752 1629 5782 1663
rect 5544 1561 5574 1595
rect 5752 1561 5782 1595
rect 5544 1479 5574 1527
rect 5608 1479 5718 1491
rect 5752 1479 5782 1527
rect 5544 1464 5782 1479
rect 5884 3010 6004 4106
rect 6314 4388 6321 4494
rect 6427 4388 6434 4494
rect 6974 4388 6996 4494
rect 6314 4214 6434 4388
rect 6314 4180 6357 4214
rect 6391 4180 6434 4214
rect 6314 4140 6434 4180
rect 6314 4106 6357 4140
rect 6391 4106 6434 4140
rect 5884 2976 5927 3010
rect 5961 2976 6004 3010
rect 5884 2932 6004 2976
rect 5884 2898 5927 2932
rect 5961 2898 6004 2932
rect 5884 2854 6004 2898
rect 5884 2820 5927 2854
rect 5961 2820 6004 2854
rect 5884 2776 6004 2820
rect 5884 2742 5927 2776
rect 5961 2742 6004 2776
rect 5884 2697 6004 2742
rect 5884 2663 5927 2697
rect 5961 2663 6004 2697
rect 5884 2618 6004 2663
rect 5884 2584 5927 2618
rect 5961 2584 6004 2618
rect 5884 2539 6004 2584
rect 5884 2505 5927 2539
rect 5961 2505 6004 2539
rect 5322 1375 5365 1409
rect 5399 1375 5442 1409
rect 5322 1335 5442 1375
rect 5322 1301 5365 1335
rect 5399 1301 5442 1335
rect 5322 1285 5442 1301
rect 5884 1409 6004 2505
rect 6069 4028 6070 4062
rect 6104 4046 6142 4062
rect 6104 4028 6106 4046
rect 6069 4012 6106 4028
rect 6140 4028 6142 4046
rect 6176 4046 6214 4062
rect 6176 4028 6178 4046
rect 6140 4012 6178 4028
rect 6212 4028 6214 4046
rect 6248 4028 6249 4062
rect 6212 4012 6249 4028
rect 6069 3988 6249 4012
rect 6069 3954 6070 3988
rect 6104 3978 6142 3988
rect 6104 3954 6106 3978
rect 6069 3944 6106 3954
rect 6140 3954 6142 3978
rect 6176 3978 6214 3988
rect 6176 3954 6178 3978
rect 6140 3944 6178 3954
rect 6212 3954 6214 3978
rect 6248 3954 6249 3988
rect 6212 3944 6249 3954
rect 6069 3914 6249 3944
rect 6069 3880 6070 3914
rect 6104 3910 6142 3914
rect 6104 3880 6106 3910
rect 6069 3876 6106 3880
rect 6140 3880 6142 3910
rect 6176 3910 6214 3914
rect 6176 3880 6178 3910
rect 6140 3876 6178 3880
rect 6212 3880 6214 3910
rect 6248 3880 6249 3914
rect 6212 3876 6249 3880
rect 6069 3842 6249 3876
rect 6069 3840 6106 3842
rect 6069 3806 6070 3840
rect 6104 3808 6106 3840
rect 6140 3840 6178 3842
rect 6140 3808 6142 3840
rect 6104 3806 6142 3808
rect 6176 3808 6178 3840
rect 6212 3840 6249 3842
rect 6212 3808 6214 3840
rect 6176 3806 6214 3808
rect 6248 3806 6249 3840
rect 6069 3774 6249 3806
rect 6069 3766 6106 3774
rect 6069 3732 6070 3766
rect 6104 3740 6106 3766
rect 6140 3766 6178 3774
rect 6140 3740 6142 3766
rect 6104 3732 6142 3740
rect 6176 3740 6178 3766
rect 6212 3766 6249 3774
rect 6212 3740 6214 3766
rect 6176 3732 6214 3740
rect 6248 3732 6249 3766
rect 6069 3706 6249 3732
rect 6069 3692 6106 3706
rect 6069 3658 6070 3692
rect 6104 3672 6106 3692
rect 6140 3692 6178 3706
rect 6140 3672 6142 3692
rect 6104 3658 6142 3672
rect 6176 3672 6178 3692
rect 6212 3692 6249 3706
rect 6212 3672 6214 3692
rect 6176 3658 6214 3672
rect 6248 3658 6249 3692
rect 6069 3638 6249 3658
rect 6069 3618 6106 3638
rect 6069 3584 6070 3618
rect 6104 3604 6106 3618
rect 6140 3618 6178 3638
rect 6140 3604 6142 3618
rect 6104 3584 6142 3604
rect 6176 3604 6178 3618
rect 6212 3618 6249 3638
rect 6212 3604 6214 3618
rect 6176 3584 6214 3604
rect 6248 3584 6249 3618
rect 6069 3570 6249 3584
rect 6069 3544 6106 3570
rect 6069 3510 6070 3544
rect 6104 3536 6106 3544
rect 6140 3544 6178 3570
rect 6140 3536 6142 3544
rect 6104 3510 6142 3536
rect 6176 3536 6178 3544
rect 6212 3544 6249 3570
rect 6212 3536 6214 3544
rect 6176 3510 6214 3536
rect 6248 3510 6249 3544
rect 6069 3502 6249 3510
rect 6069 3470 6106 3502
rect 6069 3436 6070 3470
rect 6104 3468 6106 3470
rect 6140 3470 6178 3502
rect 6140 3468 6142 3470
rect 6104 3436 6142 3468
rect 6176 3468 6178 3470
rect 6212 3470 6249 3502
rect 6212 3468 6214 3470
rect 6176 3436 6214 3468
rect 6248 3436 6249 3470
rect 6069 3434 6249 3436
rect 6069 3400 6106 3434
rect 6140 3400 6178 3434
rect 6212 3400 6249 3434
rect 6069 3396 6249 3400
rect 6069 3362 6070 3396
rect 6104 3366 6142 3396
rect 6104 3362 6106 3366
rect 6069 3332 6106 3362
rect 6140 3362 6142 3366
rect 6176 3366 6214 3396
rect 6176 3362 6178 3366
rect 6140 3332 6178 3362
rect 6212 3362 6214 3366
rect 6248 3362 6249 3396
rect 6212 3332 6249 3362
rect 6069 3322 6249 3332
rect 6069 3288 6070 3322
rect 6104 3298 6142 3322
rect 6104 3288 6106 3298
rect 6069 3264 6106 3288
rect 6140 3288 6142 3298
rect 6176 3298 6214 3322
rect 6176 3288 6178 3298
rect 6140 3264 6178 3288
rect 6212 3288 6214 3298
rect 6248 3288 6249 3322
rect 6212 3264 6249 3288
rect 6069 3248 6249 3264
rect 6069 3214 6070 3248
rect 6104 3230 6142 3248
rect 6104 3214 6106 3230
rect 6069 3196 6106 3214
rect 6140 3214 6142 3230
rect 6176 3230 6214 3248
rect 6176 3214 6178 3230
rect 6140 3196 6178 3214
rect 6212 3214 6214 3230
rect 6248 3214 6249 3248
rect 6212 3196 6249 3214
rect 6069 3174 6249 3196
rect 6069 3140 6070 3174
rect 6104 3162 6142 3174
rect 6104 3140 6106 3162
rect 6069 3128 6106 3140
rect 6140 3140 6142 3162
rect 6176 3162 6214 3174
rect 6176 3140 6178 3162
rect 6140 3128 6178 3140
rect 6212 3140 6214 3162
rect 6248 3140 6249 3174
rect 6212 3128 6249 3140
rect 6069 3100 6249 3128
rect 6069 3066 6070 3100
rect 6104 3066 6142 3100
rect 6176 3066 6214 3100
rect 6248 3066 6249 3100
rect 6069 3026 6249 3066
rect 6069 2992 6070 3026
rect 6104 2992 6142 3026
rect 6176 2992 6214 3026
rect 6248 2992 6249 3026
rect 6069 2952 6249 2992
rect 6069 2918 6070 2952
rect 6104 2918 6142 2952
rect 6176 2918 6214 2952
rect 6248 2918 6249 2952
rect 6069 2878 6249 2918
rect 6069 2844 6070 2878
rect 6104 2844 6142 2878
rect 6176 2844 6214 2878
rect 6248 2844 6249 2878
rect 6069 2804 6249 2844
rect 6069 2770 6070 2804
rect 6104 2770 6142 2804
rect 6176 2770 6214 2804
rect 6248 2770 6249 2804
rect 6069 2730 6249 2770
rect 6069 2696 6070 2730
rect 6104 2696 6142 2730
rect 6176 2696 6214 2730
rect 6248 2696 6249 2730
rect 6069 2656 6249 2696
rect 6069 2622 6070 2656
rect 6104 2622 6142 2656
rect 6176 2622 6214 2656
rect 6248 2622 6249 2656
rect 6069 2582 6249 2622
rect 6069 2548 6070 2582
rect 6104 2548 6142 2582
rect 6176 2548 6214 2582
rect 6248 2548 6249 2582
rect 6069 2508 6249 2548
rect 6069 2474 6070 2508
rect 6104 2474 6142 2508
rect 6176 2474 6214 2508
rect 6248 2474 6249 2508
rect 6069 2445 6249 2474
rect 6069 2434 6106 2445
rect 6069 2400 6070 2434
rect 6104 2411 6106 2434
rect 6140 2434 6178 2445
rect 6140 2411 6142 2434
rect 6104 2400 6142 2411
rect 6176 2411 6178 2434
rect 6212 2434 6249 2445
rect 6212 2411 6214 2434
rect 6176 2400 6214 2411
rect 6248 2400 6249 2434
rect 6069 2377 6249 2400
rect 6069 2360 6106 2377
rect 6069 2326 6070 2360
rect 6104 2343 6106 2360
rect 6140 2360 6178 2377
rect 6140 2343 6142 2360
rect 6104 2326 6142 2343
rect 6176 2343 6178 2360
rect 6212 2360 6249 2377
rect 6212 2343 6214 2360
rect 6176 2326 6214 2343
rect 6248 2326 6249 2360
rect 6069 2309 6249 2326
rect 6069 2286 6106 2309
rect 6069 2252 6070 2286
rect 6104 2275 6106 2286
rect 6140 2286 6178 2309
rect 6140 2275 6142 2286
rect 6104 2252 6142 2275
rect 6176 2275 6178 2286
rect 6212 2286 6249 2309
rect 6212 2275 6214 2286
rect 6176 2252 6214 2275
rect 6248 2252 6249 2286
rect 6069 2241 6249 2252
rect 6069 2212 6106 2241
rect 6069 2178 6070 2212
rect 6104 2207 6106 2212
rect 6140 2212 6178 2241
rect 6140 2207 6142 2212
rect 6104 2178 6142 2207
rect 6176 2207 6178 2212
rect 6212 2212 6249 2241
rect 6212 2207 6214 2212
rect 6176 2178 6214 2207
rect 6248 2178 6249 2212
rect 6069 2173 6249 2178
rect 6069 2139 6106 2173
rect 6140 2139 6178 2173
rect 6212 2139 6249 2173
rect 6069 2138 6249 2139
rect 6069 2104 6070 2138
rect 6104 2105 6142 2138
rect 6104 2104 6106 2105
rect 6069 2071 6106 2104
rect 6140 2104 6142 2105
rect 6176 2105 6214 2138
rect 6176 2104 6178 2105
rect 6140 2071 6178 2104
rect 6212 2104 6214 2105
rect 6248 2104 6249 2138
rect 6212 2071 6249 2104
rect 6069 2064 6249 2071
rect 6069 2030 6070 2064
rect 6104 2037 6142 2064
rect 6104 2030 6106 2037
rect 6069 2003 6106 2030
rect 6140 2030 6142 2037
rect 6176 2037 6214 2064
rect 6176 2030 6178 2037
rect 6140 2003 6178 2030
rect 6212 2030 6214 2037
rect 6248 2030 6249 2064
rect 6212 2003 6249 2030
rect 6069 1990 6249 2003
rect 6069 1956 6070 1990
rect 6104 1969 6142 1990
rect 6104 1956 6106 1969
rect 6069 1935 6106 1956
rect 6140 1956 6142 1969
rect 6176 1969 6214 1990
rect 6176 1956 6178 1969
rect 6140 1935 6178 1956
rect 6212 1956 6214 1969
rect 6248 1956 6249 1990
rect 6212 1935 6249 1956
rect 6069 1916 6249 1935
rect 6069 1882 6070 1916
rect 6104 1901 6142 1916
rect 6104 1882 6106 1901
rect 6069 1867 6106 1882
rect 6140 1882 6142 1901
rect 6176 1901 6214 1916
rect 6176 1882 6178 1901
rect 6140 1867 6178 1882
rect 6212 1882 6214 1901
rect 6248 1882 6249 1916
rect 6212 1867 6249 1882
rect 6069 1842 6249 1867
rect 6069 1808 6070 1842
rect 6104 1833 6142 1842
rect 6104 1808 6106 1833
rect 6069 1799 6106 1808
rect 6140 1808 6142 1833
rect 6176 1833 6214 1842
rect 6176 1808 6178 1833
rect 6140 1799 6178 1808
rect 6212 1808 6214 1833
rect 6248 1808 6249 1842
rect 6212 1799 6249 1808
rect 6069 1768 6249 1799
rect 6069 1734 6070 1768
rect 6104 1765 6142 1768
rect 6104 1734 6106 1765
rect 6069 1731 6106 1734
rect 6140 1734 6142 1765
rect 6176 1765 6214 1768
rect 6176 1734 6178 1765
rect 6140 1731 6178 1734
rect 6212 1734 6214 1765
rect 6248 1734 6249 1768
rect 6212 1731 6249 1734
rect 6069 1697 6249 1731
rect 6069 1694 6106 1697
rect 6069 1660 6070 1694
rect 6104 1663 6106 1694
rect 6140 1694 6178 1697
rect 6140 1663 6142 1694
rect 6104 1660 6142 1663
rect 6176 1663 6178 1694
rect 6212 1694 6249 1697
rect 6212 1663 6214 1694
rect 6176 1660 6214 1663
rect 6248 1660 6249 1694
rect 6069 1629 6249 1660
rect 6069 1620 6106 1629
rect 6069 1586 6070 1620
rect 6104 1595 6106 1620
rect 6140 1620 6178 1629
rect 6140 1595 6142 1620
rect 6104 1586 6142 1595
rect 6176 1595 6178 1620
rect 6212 1620 6249 1629
rect 6212 1595 6214 1620
rect 6176 1586 6214 1595
rect 6248 1586 6249 1620
rect 6069 1561 6249 1586
rect 6069 1545 6106 1561
rect 6069 1511 6070 1545
rect 6104 1527 6106 1545
rect 6140 1545 6178 1561
rect 6140 1527 6142 1545
rect 6104 1511 6142 1527
rect 6176 1527 6178 1545
rect 6212 1545 6249 1561
rect 6212 1527 6214 1545
rect 6176 1511 6214 1527
rect 6248 1511 6249 1545
rect 6314 3010 6434 4106
rect 6876 4214 6996 4388
rect 6876 4180 6919 4214
rect 6953 4180 6996 4214
rect 6876 4140 6996 4180
rect 6876 4106 6919 4140
rect 6953 4106 6996 4140
rect 6314 2976 6357 3010
rect 6391 2976 6434 3010
rect 6314 2932 6434 2976
rect 6314 2898 6357 2932
rect 6391 2898 6434 2932
rect 6314 2854 6434 2898
rect 6314 2820 6357 2854
rect 6391 2820 6434 2854
rect 6314 2776 6434 2820
rect 6314 2742 6357 2776
rect 6391 2742 6434 2776
rect 6314 2697 6434 2742
rect 6314 2663 6357 2697
rect 6391 2663 6434 2697
rect 6314 2618 6434 2663
rect 6314 2584 6357 2618
rect 6391 2584 6434 2618
rect 6314 2539 6434 2584
rect 6314 2505 6357 2539
rect 6391 2505 6434 2539
rect 6106 1491 6212 1511
rect 5884 1375 5927 1409
rect 5961 1375 6004 1409
rect 5884 1335 6004 1375
rect 5884 1301 5927 1335
rect 5961 1301 6004 1335
rect 5884 1285 6004 1301
rect 6314 1409 6434 2505
rect 6536 4050 6638 4062
rect 6672 4050 6774 4062
rect 6536 4046 6566 4050
rect 6744 4046 6774 4050
rect 6536 3978 6566 4012
rect 6744 3978 6774 4012
rect 6536 3910 6566 3944
rect 6744 3910 6774 3944
rect 6536 3842 6566 3876
rect 6744 3842 6774 3876
rect 6536 3774 6566 3808
rect 6744 3774 6774 3808
rect 6536 3706 6566 3740
rect 6744 3706 6774 3740
rect 6536 3638 6566 3672
rect 6744 3638 6774 3672
rect 6536 3570 6566 3604
rect 6744 3570 6774 3604
rect 6536 3502 6566 3536
rect 6744 3502 6774 3536
rect 6536 3434 6566 3468
rect 6744 3434 6774 3468
rect 6536 3366 6566 3400
rect 6744 3366 6774 3400
rect 6536 3298 6566 3332
rect 6744 3298 6774 3332
rect 6536 3230 6566 3264
rect 6744 3230 6774 3264
rect 6536 3162 6566 3196
rect 6744 3162 6774 3196
rect 6536 3080 6566 3128
rect 6600 3080 6710 3092
rect 6744 3080 6774 3128
rect 6536 3040 6774 3080
rect 6536 2574 6566 3040
rect 6744 2574 6774 3040
rect 6536 2535 6774 2574
rect 6536 2501 6566 2535
rect 6600 2501 6638 2535
rect 6672 2501 6710 2535
rect 6744 2501 6774 2535
rect 6536 2461 6774 2501
rect 6536 2449 6638 2461
rect 6672 2449 6774 2461
rect 6536 2445 6566 2449
rect 6744 2445 6774 2449
rect 6536 2377 6566 2411
rect 6744 2377 6774 2411
rect 6536 2309 6566 2343
rect 6744 2309 6774 2343
rect 6536 2241 6566 2275
rect 6744 2241 6774 2275
rect 6536 2173 6566 2207
rect 6744 2173 6774 2207
rect 6536 2105 6566 2139
rect 6744 2105 6774 2139
rect 6536 2037 6566 2071
rect 6744 2037 6774 2071
rect 6536 1969 6566 2003
rect 6744 1969 6774 2003
rect 6536 1901 6566 1935
rect 6744 1901 6774 1935
rect 6536 1833 6566 1867
rect 6744 1833 6774 1867
rect 6536 1765 6566 1799
rect 6744 1765 6774 1799
rect 6536 1697 6566 1731
rect 6744 1697 6774 1731
rect 6536 1629 6566 1663
rect 6744 1629 6774 1663
rect 6536 1561 6566 1595
rect 6744 1561 6774 1595
rect 6536 1479 6566 1527
rect 6600 1479 6710 1491
rect 6744 1479 6774 1527
rect 6536 1464 6774 1479
rect 6876 3010 6996 4106
rect 7306 4388 7313 4494
rect 7419 4388 7426 4494
rect 7306 4214 7426 4388
rect 7306 4180 7349 4214
rect 7383 4180 7426 4214
rect 7306 4140 7426 4180
rect 7306 4106 7349 4140
rect 7383 4106 7426 4140
rect 6876 2976 6919 3010
rect 6953 2976 6996 3010
rect 6876 2932 6996 2976
rect 6876 2898 6919 2932
rect 6953 2898 6996 2932
rect 6876 2854 6996 2898
rect 6876 2820 6919 2854
rect 6953 2820 6996 2854
rect 6876 2776 6996 2820
rect 6876 2742 6919 2776
rect 6953 2742 6996 2776
rect 6876 2697 6996 2742
rect 6876 2663 6919 2697
rect 6953 2663 6996 2697
rect 6876 2618 6996 2663
rect 6876 2584 6919 2618
rect 6953 2584 6996 2618
rect 6876 2539 6996 2584
rect 6876 2505 6919 2539
rect 6953 2505 6996 2539
rect 6314 1375 6357 1409
rect 6391 1375 6434 1409
rect 6314 1335 6434 1375
rect 6314 1301 6357 1335
rect 6391 1301 6434 1335
rect 6314 1285 6434 1301
rect 6876 1409 6996 2505
rect 7061 4028 7062 4062
rect 7096 4046 7134 4062
rect 7096 4028 7098 4046
rect 7061 4012 7098 4028
rect 7132 4028 7134 4046
rect 7168 4046 7206 4062
rect 7168 4028 7170 4046
rect 7132 4012 7170 4028
rect 7204 4028 7206 4046
rect 7240 4028 7241 4062
rect 7204 4012 7241 4028
rect 7061 3988 7241 4012
rect 7061 3954 7062 3988
rect 7096 3978 7134 3988
rect 7096 3954 7098 3978
rect 7061 3944 7098 3954
rect 7132 3954 7134 3978
rect 7168 3978 7206 3988
rect 7168 3954 7170 3978
rect 7132 3944 7170 3954
rect 7204 3954 7206 3978
rect 7240 3954 7241 3988
rect 7204 3944 7241 3954
rect 7061 3914 7241 3944
rect 7061 3880 7062 3914
rect 7096 3910 7134 3914
rect 7096 3880 7098 3910
rect 7061 3876 7098 3880
rect 7132 3880 7134 3910
rect 7168 3910 7206 3914
rect 7168 3880 7170 3910
rect 7132 3876 7170 3880
rect 7204 3880 7206 3910
rect 7240 3880 7241 3914
rect 7204 3876 7241 3880
rect 7061 3842 7241 3876
rect 7061 3840 7098 3842
rect 7061 3806 7062 3840
rect 7096 3808 7098 3840
rect 7132 3840 7170 3842
rect 7132 3808 7134 3840
rect 7096 3806 7134 3808
rect 7168 3808 7170 3840
rect 7204 3840 7241 3842
rect 7204 3808 7206 3840
rect 7168 3806 7206 3808
rect 7240 3806 7241 3840
rect 7061 3774 7241 3806
rect 7061 3766 7098 3774
rect 7061 3732 7062 3766
rect 7096 3740 7098 3766
rect 7132 3766 7170 3774
rect 7132 3740 7134 3766
rect 7096 3732 7134 3740
rect 7168 3740 7170 3766
rect 7204 3766 7241 3774
rect 7204 3740 7206 3766
rect 7168 3732 7206 3740
rect 7240 3732 7241 3766
rect 7061 3706 7241 3732
rect 7061 3692 7098 3706
rect 7061 3658 7062 3692
rect 7096 3672 7098 3692
rect 7132 3692 7170 3706
rect 7132 3672 7134 3692
rect 7096 3658 7134 3672
rect 7168 3672 7170 3692
rect 7204 3692 7241 3706
rect 7204 3672 7206 3692
rect 7168 3658 7206 3672
rect 7240 3658 7241 3692
rect 7061 3638 7241 3658
rect 7061 3618 7098 3638
rect 7061 3584 7062 3618
rect 7096 3604 7098 3618
rect 7132 3618 7170 3638
rect 7132 3604 7134 3618
rect 7096 3584 7134 3604
rect 7168 3604 7170 3618
rect 7204 3618 7241 3638
rect 7204 3604 7206 3618
rect 7168 3584 7206 3604
rect 7240 3584 7241 3618
rect 7061 3570 7241 3584
rect 7061 3544 7098 3570
rect 7061 3510 7062 3544
rect 7096 3536 7098 3544
rect 7132 3544 7170 3570
rect 7132 3536 7134 3544
rect 7096 3510 7134 3536
rect 7168 3536 7170 3544
rect 7204 3544 7241 3570
rect 7204 3536 7206 3544
rect 7168 3510 7206 3536
rect 7240 3510 7241 3544
rect 7061 3502 7241 3510
rect 7061 3470 7098 3502
rect 7061 3436 7062 3470
rect 7096 3468 7098 3470
rect 7132 3470 7170 3502
rect 7132 3468 7134 3470
rect 7096 3436 7134 3468
rect 7168 3468 7170 3470
rect 7204 3470 7241 3502
rect 7204 3468 7206 3470
rect 7168 3436 7206 3468
rect 7240 3436 7241 3470
rect 7061 3434 7241 3436
rect 7061 3400 7098 3434
rect 7132 3400 7170 3434
rect 7204 3400 7241 3434
rect 7061 3396 7241 3400
rect 7061 3362 7062 3396
rect 7096 3366 7134 3396
rect 7096 3362 7098 3366
rect 7061 3332 7098 3362
rect 7132 3362 7134 3366
rect 7168 3366 7206 3396
rect 7168 3362 7170 3366
rect 7132 3332 7170 3362
rect 7204 3362 7206 3366
rect 7240 3362 7241 3396
rect 7204 3332 7241 3362
rect 7061 3322 7241 3332
rect 7061 3288 7062 3322
rect 7096 3298 7134 3322
rect 7096 3288 7098 3298
rect 7061 3264 7098 3288
rect 7132 3288 7134 3298
rect 7168 3298 7206 3322
rect 7168 3288 7170 3298
rect 7132 3264 7170 3288
rect 7204 3288 7206 3298
rect 7240 3288 7241 3322
rect 7204 3264 7241 3288
rect 7061 3248 7241 3264
rect 7061 3214 7062 3248
rect 7096 3230 7134 3248
rect 7096 3214 7098 3230
rect 7061 3196 7098 3214
rect 7132 3214 7134 3230
rect 7168 3230 7206 3248
rect 7168 3214 7170 3230
rect 7132 3196 7170 3214
rect 7204 3214 7206 3230
rect 7240 3214 7241 3248
rect 7204 3196 7241 3214
rect 7061 3174 7241 3196
rect 7061 3140 7062 3174
rect 7096 3162 7134 3174
rect 7096 3140 7098 3162
rect 7061 3128 7098 3140
rect 7132 3140 7134 3162
rect 7168 3162 7206 3174
rect 7168 3140 7170 3162
rect 7132 3128 7170 3140
rect 7204 3140 7206 3162
rect 7240 3140 7241 3174
rect 7204 3128 7241 3140
rect 7061 3100 7241 3128
rect 7061 3066 7062 3100
rect 7096 3066 7134 3100
rect 7168 3066 7206 3100
rect 7240 3066 7241 3100
rect 7061 3026 7241 3066
rect 7061 2992 7062 3026
rect 7096 2992 7134 3026
rect 7168 2992 7206 3026
rect 7240 2992 7241 3026
rect 7061 2952 7241 2992
rect 7061 2918 7062 2952
rect 7096 2918 7134 2952
rect 7168 2918 7206 2952
rect 7240 2918 7241 2952
rect 7061 2878 7241 2918
rect 7061 2844 7062 2878
rect 7096 2844 7134 2878
rect 7168 2844 7206 2878
rect 7240 2844 7241 2878
rect 7061 2804 7241 2844
rect 7061 2770 7062 2804
rect 7096 2770 7134 2804
rect 7168 2770 7206 2804
rect 7240 2770 7241 2804
rect 7061 2730 7241 2770
rect 7061 2696 7062 2730
rect 7096 2696 7134 2730
rect 7168 2696 7206 2730
rect 7240 2696 7241 2730
rect 7061 2656 7241 2696
rect 7061 2622 7062 2656
rect 7096 2622 7134 2656
rect 7168 2622 7206 2656
rect 7240 2622 7241 2656
rect 7061 2582 7241 2622
rect 7061 2548 7062 2582
rect 7096 2548 7134 2582
rect 7168 2548 7206 2582
rect 7240 2548 7241 2582
rect 7061 2508 7241 2548
rect 7061 2474 7062 2508
rect 7096 2474 7134 2508
rect 7168 2474 7206 2508
rect 7240 2474 7241 2508
rect 7061 2445 7241 2474
rect 7061 2434 7098 2445
rect 7061 2400 7062 2434
rect 7096 2411 7098 2434
rect 7132 2434 7170 2445
rect 7132 2411 7134 2434
rect 7096 2400 7134 2411
rect 7168 2411 7170 2434
rect 7204 2434 7241 2445
rect 7204 2411 7206 2434
rect 7168 2400 7206 2411
rect 7240 2400 7241 2434
rect 7061 2377 7241 2400
rect 7061 2360 7098 2377
rect 7061 2326 7062 2360
rect 7096 2343 7098 2360
rect 7132 2360 7170 2377
rect 7132 2343 7134 2360
rect 7096 2326 7134 2343
rect 7168 2343 7170 2360
rect 7204 2360 7241 2377
rect 7204 2343 7206 2360
rect 7168 2326 7206 2343
rect 7240 2326 7241 2360
rect 7061 2309 7241 2326
rect 7061 2286 7098 2309
rect 7061 2252 7062 2286
rect 7096 2275 7098 2286
rect 7132 2286 7170 2309
rect 7132 2275 7134 2286
rect 7096 2252 7134 2275
rect 7168 2275 7170 2286
rect 7204 2286 7241 2309
rect 7204 2275 7206 2286
rect 7168 2252 7206 2275
rect 7240 2252 7241 2286
rect 7061 2241 7241 2252
rect 7061 2212 7098 2241
rect 7061 2178 7062 2212
rect 7096 2207 7098 2212
rect 7132 2212 7170 2241
rect 7132 2207 7134 2212
rect 7096 2178 7134 2207
rect 7168 2207 7170 2212
rect 7204 2212 7241 2241
rect 7204 2207 7206 2212
rect 7168 2178 7206 2207
rect 7240 2178 7241 2212
rect 7061 2173 7241 2178
rect 7061 2139 7098 2173
rect 7132 2139 7170 2173
rect 7204 2139 7241 2173
rect 7061 2138 7241 2139
rect 7061 2104 7062 2138
rect 7096 2105 7134 2138
rect 7096 2104 7098 2105
rect 7061 2071 7098 2104
rect 7132 2104 7134 2105
rect 7168 2105 7206 2138
rect 7168 2104 7170 2105
rect 7132 2071 7170 2104
rect 7204 2104 7206 2105
rect 7240 2104 7241 2138
rect 7204 2071 7241 2104
rect 7061 2064 7241 2071
rect 7061 2030 7062 2064
rect 7096 2037 7134 2064
rect 7096 2030 7098 2037
rect 7061 2003 7098 2030
rect 7132 2030 7134 2037
rect 7168 2037 7206 2064
rect 7168 2030 7170 2037
rect 7132 2003 7170 2030
rect 7204 2030 7206 2037
rect 7240 2030 7241 2064
rect 7204 2003 7241 2030
rect 7061 1990 7241 2003
rect 7061 1956 7062 1990
rect 7096 1969 7134 1990
rect 7096 1956 7098 1969
rect 7061 1935 7098 1956
rect 7132 1956 7134 1969
rect 7168 1969 7206 1990
rect 7168 1956 7170 1969
rect 7132 1935 7170 1956
rect 7204 1956 7206 1969
rect 7240 1956 7241 1990
rect 7204 1935 7241 1956
rect 7061 1916 7241 1935
rect 7061 1882 7062 1916
rect 7096 1901 7134 1916
rect 7096 1882 7098 1901
rect 7061 1867 7098 1882
rect 7132 1882 7134 1901
rect 7168 1901 7206 1916
rect 7168 1882 7170 1901
rect 7132 1867 7170 1882
rect 7204 1882 7206 1901
rect 7240 1882 7241 1916
rect 7204 1867 7241 1882
rect 7061 1842 7241 1867
rect 7061 1808 7062 1842
rect 7096 1833 7134 1842
rect 7096 1808 7098 1833
rect 7061 1799 7098 1808
rect 7132 1808 7134 1833
rect 7168 1833 7206 1842
rect 7168 1808 7170 1833
rect 7132 1799 7170 1808
rect 7204 1808 7206 1833
rect 7240 1808 7241 1842
rect 7204 1799 7241 1808
rect 7061 1768 7241 1799
rect 7061 1734 7062 1768
rect 7096 1765 7134 1768
rect 7096 1734 7098 1765
rect 7061 1731 7098 1734
rect 7132 1734 7134 1765
rect 7168 1765 7206 1768
rect 7168 1734 7170 1765
rect 7132 1731 7170 1734
rect 7204 1734 7206 1765
rect 7240 1734 7241 1768
rect 7204 1731 7241 1734
rect 7061 1697 7241 1731
rect 7061 1694 7098 1697
rect 7061 1660 7062 1694
rect 7096 1663 7098 1694
rect 7132 1694 7170 1697
rect 7132 1663 7134 1694
rect 7096 1660 7134 1663
rect 7168 1663 7170 1694
rect 7204 1694 7241 1697
rect 7204 1663 7206 1694
rect 7168 1660 7206 1663
rect 7240 1660 7241 1694
rect 7061 1629 7241 1660
rect 7061 1620 7098 1629
rect 7061 1586 7062 1620
rect 7096 1595 7098 1620
rect 7132 1620 7170 1629
rect 7132 1595 7134 1620
rect 7096 1586 7134 1595
rect 7168 1595 7170 1620
rect 7204 1620 7241 1629
rect 7204 1595 7206 1620
rect 7168 1586 7206 1595
rect 7240 1586 7241 1620
rect 7061 1561 7241 1586
rect 7061 1545 7098 1561
rect 7061 1511 7062 1545
rect 7096 1527 7098 1545
rect 7132 1545 7170 1561
rect 7132 1527 7134 1545
rect 7096 1511 7134 1527
rect 7168 1527 7170 1545
rect 7204 1545 7241 1561
rect 7204 1527 7206 1545
rect 7168 1511 7206 1527
rect 7240 1511 7241 1545
rect 7306 3010 7426 4106
rect 7868 4388 7875 4494
rect 7981 4388 7988 4494
rect 7868 4214 7988 4388
rect 7868 4180 7911 4214
rect 7945 4180 7988 4214
rect 7868 4140 7988 4180
rect 7868 4106 7911 4140
rect 7945 4106 7988 4140
rect 7306 2976 7349 3010
rect 7383 2976 7426 3010
rect 7306 2932 7426 2976
rect 7306 2898 7349 2932
rect 7383 2898 7426 2932
rect 7306 2854 7426 2898
rect 7306 2820 7349 2854
rect 7383 2820 7426 2854
rect 7306 2776 7426 2820
rect 7306 2742 7349 2776
rect 7383 2742 7426 2776
rect 7306 2697 7426 2742
rect 7306 2663 7349 2697
rect 7383 2663 7426 2697
rect 7306 2618 7426 2663
rect 7306 2584 7349 2618
rect 7383 2584 7426 2618
rect 7306 2539 7426 2584
rect 7306 2505 7349 2539
rect 7383 2505 7426 2539
rect 7098 1491 7204 1511
rect 6876 1375 6919 1409
rect 6953 1375 6996 1409
rect 6876 1335 6996 1375
rect 6876 1301 6919 1335
rect 6953 1301 6996 1335
rect 6876 1285 6996 1301
rect 7306 1409 7426 2505
rect 7528 4050 7630 4062
rect 7664 4050 7766 4062
rect 7528 4046 7558 4050
rect 7736 4046 7766 4050
rect 7528 3978 7558 4012
rect 7736 3978 7766 4012
rect 7528 3910 7558 3944
rect 7736 3910 7766 3944
rect 7528 3842 7558 3876
rect 7736 3842 7766 3876
rect 7528 3774 7558 3808
rect 7736 3774 7766 3808
rect 7528 3706 7558 3740
rect 7736 3706 7766 3740
rect 7528 3638 7558 3672
rect 7736 3638 7766 3672
rect 7528 3570 7558 3604
rect 7736 3570 7766 3604
rect 7528 3502 7558 3536
rect 7736 3502 7766 3536
rect 7528 3434 7558 3468
rect 7736 3434 7766 3468
rect 7528 3366 7558 3400
rect 7736 3366 7766 3400
rect 7528 3298 7558 3332
rect 7736 3298 7766 3332
rect 7528 3230 7558 3264
rect 7736 3230 7766 3264
rect 7528 3162 7558 3196
rect 7736 3162 7766 3196
rect 7528 3080 7558 3128
rect 7592 3080 7702 3092
rect 7736 3080 7766 3128
rect 7528 3040 7766 3080
rect 7528 2574 7558 3040
rect 7736 2574 7766 3040
rect 7528 2535 7766 2574
rect 7528 2501 7558 2535
rect 7592 2501 7630 2535
rect 7664 2501 7702 2535
rect 7736 2501 7766 2535
rect 7528 2461 7766 2501
rect 7528 2449 7630 2461
rect 7664 2449 7766 2461
rect 7528 2445 7558 2449
rect 7736 2445 7766 2449
rect 7528 2377 7558 2411
rect 7736 2377 7766 2411
rect 7528 2309 7558 2343
rect 7736 2309 7766 2343
rect 7528 2241 7558 2275
rect 7736 2241 7766 2275
rect 7528 2173 7558 2207
rect 7736 2173 7766 2207
rect 7528 2105 7558 2139
rect 7736 2105 7766 2139
rect 7528 2037 7558 2071
rect 7736 2037 7766 2071
rect 7528 1969 7558 2003
rect 7736 1969 7766 2003
rect 7528 1901 7558 1935
rect 7736 1901 7766 1935
rect 7528 1833 7558 1867
rect 7736 1833 7766 1867
rect 7528 1765 7558 1799
rect 7736 1765 7766 1799
rect 7528 1697 7558 1731
rect 7736 1697 7766 1731
rect 7528 1629 7558 1663
rect 7736 1629 7766 1663
rect 7528 1561 7558 1595
rect 7736 1561 7766 1595
rect 7528 1479 7558 1527
rect 7592 1479 7702 1491
rect 7736 1479 7766 1527
rect 7528 1464 7766 1479
rect 7868 3010 7988 4106
rect 8298 4388 8305 4494
rect 8411 4388 8418 4494
rect 8298 4214 8418 4388
rect 8298 4180 8341 4214
rect 8375 4180 8418 4214
rect 8298 4140 8418 4180
rect 8298 4106 8341 4140
rect 8375 4106 8418 4140
rect 7868 2976 7911 3010
rect 7945 2976 7988 3010
rect 7868 2932 7988 2976
rect 7868 2898 7911 2932
rect 7945 2898 7988 2932
rect 7868 2854 7988 2898
rect 7868 2820 7911 2854
rect 7945 2820 7988 2854
rect 7868 2776 7988 2820
rect 7868 2742 7911 2776
rect 7945 2742 7988 2776
rect 7868 2697 7988 2742
rect 7868 2663 7911 2697
rect 7945 2663 7988 2697
rect 7868 2618 7988 2663
rect 7868 2584 7911 2618
rect 7945 2584 7988 2618
rect 7868 2539 7988 2584
rect 7868 2505 7911 2539
rect 7945 2505 7988 2539
rect 7306 1375 7349 1409
rect 7383 1375 7426 1409
rect 7306 1335 7426 1375
rect 7306 1301 7349 1335
rect 7383 1301 7426 1335
rect 7306 1285 7426 1301
rect 7868 1409 7988 2505
rect 8053 4028 8054 4062
rect 8088 4046 8126 4062
rect 8088 4028 8090 4046
rect 8053 4012 8090 4028
rect 8124 4028 8126 4046
rect 8160 4046 8198 4062
rect 8160 4028 8162 4046
rect 8124 4012 8162 4028
rect 8196 4028 8198 4046
rect 8232 4028 8233 4062
rect 8196 4012 8233 4028
rect 8053 3988 8233 4012
rect 8053 3954 8054 3988
rect 8088 3978 8126 3988
rect 8088 3954 8090 3978
rect 8053 3944 8090 3954
rect 8124 3954 8126 3978
rect 8160 3978 8198 3988
rect 8160 3954 8162 3978
rect 8124 3944 8162 3954
rect 8196 3954 8198 3978
rect 8232 3954 8233 3988
rect 8196 3944 8233 3954
rect 8053 3914 8233 3944
rect 8053 3880 8054 3914
rect 8088 3910 8126 3914
rect 8088 3880 8090 3910
rect 8053 3876 8090 3880
rect 8124 3880 8126 3910
rect 8160 3910 8198 3914
rect 8160 3880 8162 3910
rect 8124 3876 8162 3880
rect 8196 3880 8198 3910
rect 8232 3880 8233 3914
rect 8196 3876 8233 3880
rect 8053 3842 8233 3876
rect 8053 3840 8090 3842
rect 8053 3806 8054 3840
rect 8088 3808 8090 3840
rect 8124 3840 8162 3842
rect 8124 3808 8126 3840
rect 8088 3806 8126 3808
rect 8160 3808 8162 3840
rect 8196 3840 8233 3842
rect 8196 3808 8198 3840
rect 8160 3806 8198 3808
rect 8232 3806 8233 3840
rect 8053 3774 8233 3806
rect 8053 3766 8090 3774
rect 8053 3732 8054 3766
rect 8088 3740 8090 3766
rect 8124 3766 8162 3774
rect 8124 3740 8126 3766
rect 8088 3732 8126 3740
rect 8160 3740 8162 3766
rect 8196 3766 8233 3774
rect 8196 3740 8198 3766
rect 8160 3732 8198 3740
rect 8232 3732 8233 3766
rect 8053 3706 8233 3732
rect 8053 3692 8090 3706
rect 8053 3658 8054 3692
rect 8088 3672 8090 3692
rect 8124 3692 8162 3706
rect 8124 3672 8126 3692
rect 8088 3658 8126 3672
rect 8160 3672 8162 3692
rect 8196 3692 8233 3706
rect 8196 3672 8198 3692
rect 8160 3658 8198 3672
rect 8232 3658 8233 3692
rect 8053 3638 8233 3658
rect 8053 3618 8090 3638
rect 8053 3584 8054 3618
rect 8088 3604 8090 3618
rect 8124 3618 8162 3638
rect 8124 3604 8126 3618
rect 8088 3584 8126 3604
rect 8160 3604 8162 3618
rect 8196 3618 8233 3638
rect 8196 3604 8198 3618
rect 8160 3584 8198 3604
rect 8232 3584 8233 3618
rect 8053 3570 8233 3584
rect 8053 3544 8090 3570
rect 8053 3510 8054 3544
rect 8088 3536 8090 3544
rect 8124 3544 8162 3570
rect 8124 3536 8126 3544
rect 8088 3510 8126 3536
rect 8160 3536 8162 3544
rect 8196 3544 8233 3570
rect 8196 3536 8198 3544
rect 8160 3510 8198 3536
rect 8232 3510 8233 3544
rect 8053 3502 8233 3510
rect 8053 3470 8090 3502
rect 8053 3436 8054 3470
rect 8088 3468 8090 3470
rect 8124 3470 8162 3502
rect 8124 3468 8126 3470
rect 8088 3436 8126 3468
rect 8160 3468 8162 3470
rect 8196 3470 8233 3502
rect 8196 3468 8198 3470
rect 8160 3436 8198 3468
rect 8232 3436 8233 3470
rect 8053 3434 8233 3436
rect 8053 3400 8090 3434
rect 8124 3400 8162 3434
rect 8196 3400 8233 3434
rect 8053 3396 8233 3400
rect 8053 3362 8054 3396
rect 8088 3366 8126 3396
rect 8088 3362 8090 3366
rect 8053 3332 8090 3362
rect 8124 3362 8126 3366
rect 8160 3366 8198 3396
rect 8160 3362 8162 3366
rect 8124 3332 8162 3362
rect 8196 3362 8198 3366
rect 8232 3362 8233 3396
rect 8196 3332 8233 3362
rect 8053 3322 8233 3332
rect 8053 3288 8054 3322
rect 8088 3298 8126 3322
rect 8088 3288 8090 3298
rect 8053 3264 8090 3288
rect 8124 3288 8126 3298
rect 8160 3298 8198 3322
rect 8160 3288 8162 3298
rect 8124 3264 8162 3288
rect 8196 3288 8198 3298
rect 8232 3288 8233 3322
rect 8196 3264 8233 3288
rect 8053 3248 8233 3264
rect 8053 3214 8054 3248
rect 8088 3230 8126 3248
rect 8088 3214 8090 3230
rect 8053 3196 8090 3214
rect 8124 3214 8126 3230
rect 8160 3230 8198 3248
rect 8160 3214 8162 3230
rect 8124 3196 8162 3214
rect 8196 3214 8198 3230
rect 8232 3214 8233 3248
rect 8196 3196 8233 3214
rect 8053 3174 8233 3196
rect 8053 3140 8054 3174
rect 8088 3162 8126 3174
rect 8088 3140 8090 3162
rect 8053 3128 8090 3140
rect 8124 3140 8126 3162
rect 8160 3162 8198 3174
rect 8160 3140 8162 3162
rect 8124 3128 8162 3140
rect 8196 3140 8198 3162
rect 8232 3140 8233 3174
rect 8196 3128 8233 3140
rect 8053 3100 8233 3128
rect 8053 3066 8054 3100
rect 8088 3066 8126 3100
rect 8160 3066 8198 3100
rect 8232 3066 8233 3100
rect 8053 3026 8233 3066
rect 8053 2992 8054 3026
rect 8088 2992 8126 3026
rect 8160 2992 8198 3026
rect 8232 2992 8233 3026
rect 8053 2952 8233 2992
rect 8053 2918 8054 2952
rect 8088 2918 8126 2952
rect 8160 2918 8198 2952
rect 8232 2918 8233 2952
rect 8053 2878 8233 2918
rect 8053 2844 8054 2878
rect 8088 2844 8126 2878
rect 8160 2844 8198 2878
rect 8232 2844 8233 2878
rect 8053 2804 8233 2844
rect 8053 2770 8054 2804
rect 8088 2770 8126 2804
rect 8160 2770 8198 2804
rect 8232 2770 8233 2804
rect 8053 2730 8233 2770
rect 8053 2696 8054 2730
rect 8088 2696 8126 2730
rect 8160 2696 8198 2730
rect 8232 2696 8233 2730
rect 8053 2656 8233 2696
rect 8053 2622 8054 2656
rect 8088 2622 8126 2656
rect 8160 2622 8198 2656
rect 8232 2622 8233 2656
rect 8053 2582 8233 2622
rect 8053 2548 8054 2582
rect 8088 2548 8126 2582
rect 8160 2548 8198 2582
rect 8232 2548 8233 2582
rect 8053 2508 8233 2548
rect 8053 2474 8054 2508
rect 8088 2474 8126 2508
rect 8160 2474 8198 2508
rect 8232 2474 8233 2508
rect 8053 2445 8233 2474
rect 8053 2434 8090 2445
rect 8053 2400 8054 2434
rect 8088 2411 8090 2434
rect 8124 2434 8162 2445
rect 8124 2411 8126 2434
rect 8088 2400 8126 2411
rect 8160 2411 8162 2434
rect 8196 2434 8233 2445
rect 8196 2411 8198 2434
rect 8160 2400 8198 2411
rect 8232 2400 8233 2434
rect 8053 2377 8233 2400
rect 8053 2360 8090 2377
rect 8053 2326 8054 2360
rect 8088 2343 8090 2360
rect 8124 2360 8162 2377
rect 8124 2343 8126 2360
rect 8088 2326 8126 2343
rect 8160 2343 8162 2360
rect 8196 2360 8233 2377
rect 8196 2343 8198 2360
rect 8160 2326 8198 2343
rect 8232 2326 8233 2360
rect 8053 2309 8233 2326
rect 8053 2286 8090 2309
rect 8053 2252 8054 2286
rect 8088 2275 8090 2286
rect 8124 2286 8162 2309
rect 8124 2275 8126 2286
rect 8088 2252 8126 2275
rect 8160 2275 8162 2286
rect 8196 2286 8233 2309
rect 8196 2275 8198 2286
rect 8160 2252 8198 2275
rect 8232 2252 8233 2286
rect 8053 2241 8233 2252
rect 8053 2212 8090 2241
rect 8053 2178 8054 2212
rect 8088 2207 8090 2212
rect 8124 2212 8162 2241
rect 8124 2207 8126 2212
rect 8088 2178 8126 2207
rect 8160 2207 8162 2212
rect 8196 2212 8233 2241
rect 8196 2207 8198 2212
rect 8160 2178 8198 2207
rect 8232 2178 8233 2212
rect 8053 2173 8233 2178
rect 8053 2139 8090 2173
rect 8124 2139 8162 2173
rect 8196 2139 8233 2173
rect 8053 2138 8233 2139
rect 8053 2104 8054 2138
rect 8088 2105 8126 2138
rect 8088 2104 8090 2105
rect 8053 2071 8090 2104
rect 8124 2104 8126 2105
rect 8160 2105 8198 2138
rect 8160 2104 8162 2105
rect 8124 2071 8162 2104
rect 8196 2104 8198 2105
rect 8232 2104 8233 2138
rect 8196 2071 8233 2104
rect 8053 2064 8233 2071
rect 8053 2030 8054 2064
rect 8088 2037 8126 2064
rect 8088 2030 8090 2037
rect 8053 2003 8090 2030
rect 8124 2030 8126 2037
rect 8160 2037 8198 2064
rect 8160 2030 8162 2037
rect 8124 2003 8162 2030
rect 8196 2030 8198 2037
rect 8232 2030 8233 2064
rect 8196 2003 8233 2030
rect 8053 1990 8233 2003
rect 8053 1956 8054 1990
rect 8088 1969 8126 1990
rect 8088 1956 8090 1969
rect 8053 1935 8090 1956
rect 8124 1956 8126 1969
rect 8160 1969 8198 1990
rect 8160 1956 8162 1969
rect 8124 1935 8162 1956
rect 8196 1956 8198 1969
rect 8232 1956 8233 1990
rect 8196 1935 8233 1956
rect 8053 1916 8233 1935
rect 8053 1882 8054 1916
rect 8088 1901 8126 1916
rect 8088 1882 8090 1901
rect 8053 1867 8090 1882
rect 8124 1882 8126 1901
rect 8160 1901 8198 1916
rect 8160 1882 8162 1901
rect 8124 1867 8162 1882
rect 8196 1882 8198 1901
rect 8232 1882 8233 1916
rect 8196 1867 8233 1882
rect 8053 1842 8233 1867
rect 8053 1808 8054 1842
rect 8088 1833 8126 1842
rect 8088 1808 8090 1833
rect 8053 1799 8090 1808
rect 8124 1808 8126 1833
rect 8160 1833 8198 1842
rect 8160 1808 8162 1833
rect 8124 1799 8162 1808
rect 8196 1808 8198 1833
rect 8232 1808 8233 1842
rect 8196 1799 8233 1808
rect 8053 1768 8233 1799
rect 8053 1734 8054 1768
rect 8088 1765 8126 1768
rect 8088 1734 8090 1765
rect 8053 1731 8090 1734
rect 8124 1734 8126 1765
rect 8160 1765 8198 1768
rect 8160 1734 8162 1765
rect 8124 1731 8162 1734
rect 8196 1734 8198 1765
rect 8232 1734 8233 1768
rect 8196 1731 8233 1734
rect 8053 1697 8233 1731
rect 8053 1694 8090 1697
rect 8053 1660 8054 1694
rect 8088 1663 8090 1694
rect 8124 1694 8162 1697
rect 8124 1663 8126 1694
rect 8088 1660 8126 1663
rect 8160 1663 8162 1694
rect 8196 1694 8233 1697
rect 8196 1663 8198 1694
rect 8160 1660 8198 1663
rect 8232 1660 8233 1694
rect 8053 1629 8233 1660
rect 8053 1620 8090 1629
rect 8053 1586 8054 1620
rect 8088 1595 8090 1620
rect 8124 1620 8162 1629
rect 8124 1595 8126 1620
rect 8088 1586 8126 1595
rect 8160 1595 8162 1620
rect 8196 1620 8233 1629
rect 8196 1595 8198 1620
rect 8160 1586 8198 1595
rect 8232 1586 8233 1620
rect 8053 1561 8233 1586
rect 8053 1545 8090 1561
rect 8053 1511 8054 1545
rect 8088 1527 8090 1545
rect 8124 1545 8162 1561
rect 8124 1527 8126 1545
rect 8088 1511 8126 1527
rect 8160 1527 8162 1545
rect 8196 1545 8233 1561
rect 8196 1527 8198 1545
rect 8160 1511 8198 1527
rect 8232 1511 8233 1545
rect 8298 3010 8418 4106
rect 8860 4388 8867 4494
rect 8973 4388 8980 4494
rect 8860 4214 8980 4388
rect 8860 4180 8903 4214
rect 8937 4180 8980 4214
rect 8860 4140 8980 4180
rect 8860 4106 8903 4140
rect 8937 4106 8980 4140
rect 8298 2976 8341 3010
rect 8375 2976 8418 3010
rect 8298 2932 8418 2976
rect 8298 2898 8341 2932
rect 8375 2898 8418 2932
rect 8298 2854 8418 2898
rect 8298 2820 8341 2854
rect 8375 2820 8418 2854
rect 8298 2776 8418 2820
rect 8298 2742 8341 2776
rect 8375 2742 8418 2776
rect 8298 2697 8418 2742
rect 8298 2663 8341 2697
rect 8375 2663 8418 2697
rect 8298 2618 8418 2663
rect 8298 2584 8341 2618
rect 8375 2584 8418 2618
rect 8298 2539 8418 2584
rect 8298 2505 8341 2539
rect 8375 2505 8418 2539
rect 8090 1491 8196 1511
rect 7868 1375 7911 1409
rect 7945 1375 7988 1409
rect 7868 1335 7988 1375
rect 7868 1301 7911 1335
rect 7945 1301 7988 1335
rect 7868 1285 7988 1301
rect 8298 1409 8418 2505
rect 8520 4050 8622 4062
rect 8656 4050 8758 4062
rect 8520 4046 8550 4050
rect 8728 4046 8758 4050
rect 8520 3978 8550 4012
rect 8728 3978 8758 4012
rect 8520 3910 8550 3944
rect 8728 3910 8758 3944
rect 8520 3842 8550 3876
rect 8728 3842 8758 3876
rect 8520 3774 8550 3808
rect 8728 3774 8758 3808
rect 8520 3706 8550 3740
rect 8728 3706 8758 3740
rect 8520 3638 8550 3672
rect 8728 3638 8758 3672
rect 8520 3570 8550 3604
rect 8728 3570 8758 3604
rect 8520 3502 8550 3536
rect 8728 3502 8758 3536
rect 8520 3434 8550 3468
rect 8728 3434 8758 3468
rect 8520 3366 8550 3400
rect 8728 3366 8758 3400
rect 8520 3298 8550 3332
rect 8728 3298 8758 3332
rect 8520 3230 8550 3264
rect 8728 3230 8758 3264
rect 8520 3162 8550 3196
rect 8728 3162 8758 3196
rect 8520 3080 8550 3128
rect 8584 3080 8694 3092
rect 8728 3080 8758 3128
rect 8520 3040 8758 3080
rect 8520 2574 8550 3040
rect 8728 2574 8758 3040
rect 8520 2535 8758 2574
rect 8520 2501 8550 2535
rect 8584 2501 8622 2535
rect 8656 2501 8694 2535
rect 8728 2501 8758 2535
rect 8520 2461 8758 2501
rect 8520 2449 8622 2461
rect 8656 2449 8758 2461
rect 8520 2445 8550 2449
rect 8728 2445 8758 2449
rect 8520 2377 8550 2411
rect 8728 2377 8758 2411
rect 8520 2309 8550 2343
rect 8728 2309 8758 2343
rect 8520 2241 8550 2275
rect 8728 2241 8758 2275
rect 8520 2173 8550 2207
rect 8728 2173 8758 2207
rect 8520 2105 8550 2139
rect 8728 2105 8758 2139
rect 8520 2037 8550 2071
rect 8728 2037 8758 2071
rect 8520 1969 8550 2003
rect 8728 1969 8758 2003
rect 8520 1901 8550 1935
rect 8728 1901 8758 1935
rect 8520 1833 8550 1867
rect 8728 1833 8758 1867
rect 8520 1765 8550 1799
rect 8728 1765 8758 1799
rect 8520 1697 8550 1731
rect 8728 1697 8758 1731
rect 8520 1629 8550 1663
rect 8728 1629 8758 1663
rect 8520 1561 8550 1595
rect 8728 1561 8758 1595
rect 8520 1479 8550 1527
rect 8584 1479 8694 1491
rect 8728 1479 8758 1527
rect 8520 1464 8758 1479
rect 8860 3010 8980 4106
rect 9290 4388 9297 4494
rect 9403 4388 9410 4494
rect 9290 4214 9410 4388
rect 9290 4180 9333 4214
rect 9367 4180 9410 4214
rect 9290 4140 9410 4180
rect 9290 4106 9333 4140
rect 9367 4106 9410 4140
rect 8860 2976 8903 3010
rect 8937 2976 8980 3010
rect 8860 2932 8980 2976
rect 8860 2898 8903 2932
rect 8937 2898 8980 2932
rect 8860 2854 8980 2898
rect 8860 2820 8903 2854
rect 8937 2820 8980 2854
rect 8860 2776 8980 2820
rect 8860 2742 8903 2776
rect 8937 2742 8980 2776
rect 8860 2697 8980 2742
rect 8860 2663 8903 2697
rect 8937 2663 8980 2697
rect 8860 2618 8980 2663
rect 8860 2584 8903 2618
rect 8937 2584 8980 2618
rect 8860 2539 8980 2584
rect 8860 2505 8903 2539
rect 8937 2505 8980 2539
rect 8298 1375 8341 1409
rect 8375 1375 8418 1409
rect 8298 1335 8418 1375
rect 8298 1301 8341 1335
rect 8375 1301 8418 1335
rect 8298 1285 8418 1301
rect 8860 1409 8980 2505
rect 9045 4028 9046 4062
rect 9080 4046 9118 4062
rect 9080 4028 9082 4046
rect 9045 4012 9082 4028
rect 9116 4028 9118 4046
rect 9152 4046 9190 4062
rect 9152 4028 9154 4046
rect 9116 4012 9154 4028
rect 9188 4028 9190 4046
rect 9224 4028 9225 4062
rect 9188 4012 9225 4028
rect 9045 3988 9225 4012
rect 9045 3954 9046 3988
rect 9080 3978 9118 3988
rect 9080 3954 9082 3978
rect 9045 3944 9082 3954
rect 9116 3954 9118 3978
rect 9152 3978 9190 3988
rect 9152 3954 9154 3978
rect 9116 3944 9154 3954
rect 9188 3954 9190 3978
rect 9224 3954 9225 3988
rect 9188 3944 9225 3954
rect 9045 3914 9225 3944
rect 9045 3880 9046 3914
rect 9080 3910 9118 3914
rect 9080 3880 9082 3910
rect 9045 3876 9082 3880
rect 9116 3880 9118 3910
rect 9152 3910 9190 3914
rect 9152 3880 9154 3910
rect 9116 3876 9154 3880
rect 9188 3880 9190 3910
rect 9224 3880 9225 3914
rect 9188 3876 9225 3880
rect 9045 3842 9225 3876
rect 9045 3840 9082 3842
rect 9045 3806 9046 3840
rect 9080 3808 9082 3840
rect 9116 3840 9154 3842
rect 9116 3808 9118 3840
rect 9080 3806 9118 3808
rect 9152 3808 9154 3840
rect 9188 3840 9225 3842
rect 9188 3808 9190 3840
rect 9152 3806 9190 3808
rect 9224 3806 9225 3840
rect 9045 3774 9225 3806
rect 9045 3766 9082 3774
rect 9045 3732 9046 3766
rect 9080 3740 9082 3766
rect 9116 3766 9154 3774
rect 9116 3740 9118 3766
rect 9080 3732 9118 3740
rect 9152 3740 9154 3766
rect 9188 3766 9225 3774
rect 9188 3740 9190 3766
rect 9152 3732 9190 3740
rect 9224 3732 9225 3766
rect 9045 3706 9225 3732
rect 9045 3692 9082 3706
rect 9045 3658 9046 3692
rect 9080 3672 9082 3692
rect 9116 3692 9154 3706
rect 9116 3672 9118 3692
rect 9080 3658 9118 3672
rect 9152 3672 9154 3692
rect 9188 3692 9225 3706
rect 9188 3672 9190 3692
rect 9152 3658 9190 3672
rect 9224 3658 9225 3692
rect 9045 3638 9225 3658
rect 9045 3618 9082 3638
rect 9045 3584 9046 3618
rect 9080 3604 9082 3618
rect 9116 3618 9154 3638
rect 9116 3604 9118 3618
rect 9080 3584 9118 3604
rect 9152 3604 9154 3618
rect 9188 3618 9225 3638
rect 9188 3604 9190 3618
rect 9152 3584 9190 3604
rect 9224 3584 9225 3618
rect 9045 3570 9225 3584
rect 9045 3544 9082 3570
rect 9045 3510 9046 3544
rect 9080 3536 9082 3544
rect 9116 3544 9154 3570
rect 9116 3536 9118 3544
rect 9080 3510 9118 3536
rect 9152 3536 9154 3544
rect 9188 3544 9225 3570
rect 9188 3536 9190 3544
rect 9152 3510 9190 3536
rect 9224 3510 9225 3544
rect 9045 3502 9225 3510
rect 9045 3470 9082 3502
rect 9045 3436 9046 3470
rect 9080 3468 9082 3470
rect 9116 3470 9154 3502
rect 9116 3468 9118 3470
rect 9080 3436 9118 3468
rect 9152 3468 9154 3470
rect 9188 3470 9225 3502
rect 9188 3468 9190 3470
rect 9152 3436 9190 3468
rect 9224 3436 9225 3470
rect 9045 3434 9225 3436
rect 9045 3400 9082 3434
rect 9116 3400 9154 3434
rect 9188 3400 9225 3434
rect 9045 3396 9225 3400
rect 9045 3362 9046 3396
rect 9080 3366 9118 3396
rect 9080 3362 9082 3366
rect 9045 3332 9082 3362
rect 9116 3362 9118 3366
rect 9152 3366 9190 3396
rect 9152 3362 9154 3366
rect 9116 3332 9154 3362
rect 9188 3362 9190 3366
rect 9224 3362 9225 3396
rect 9188 3332 9225 3362
rect 9045 3322 9225 3332
rect 9045 3288 9046 3322
rect 9080 3298 9118 3322
rect 9080 3288 9082 3298
rect 9045 3264 9082 3288
rect 9116 3288 9118 3298
rect 9152 3298 9190 3322
rect 9152 3288 9154 3298
rect 9116 3264 9154 3288
rect 9188 3288 9190 3298
rect 9224 3288 9225 3322
rect 9188 3264 9225 3288
rect 9045 3248 9225 3264
rect 9045 3214 9046 3248
rect 9080 3230 9118 3248
rect 9080 3214 9082 3230
rect 9045 3196 9082 3214
rect 9116 3214 9118 3230
rect 9152 3230 9190 3248
rect 9152 3214 9154 3230
rect 9116 3196 9154 3214
rect 9188 3214 9190 3230
rect 9224 3214 9225 3248
rect 9188 3196 9225 3214
rect 9045 3174 9225 3196
rect 9045 3140 9046 3174
rect 9080 3162 9118 3174
rect 9080 3140 9082 3162
rect 9045 3128 9082 3140
rect 9116 3140 9118 3162
rect 9152 3162 9190 3174
rect 9152 3140 9154 3162
rect 9116 3128 9154 3140
rect 9188 3140 9190 3162
rect 9224 3140 9225 3174
rect 9188 3128 9225 3140
rect 9045 3100 9225 3128
rect 9045 3066 9046 3100
rect 9080 3066 9118 3100
rect 9152 3066 9190 3100
rect 9224 3066 9225 3100
rect 9045 3026 9225 3066
rect 9045 2992 9046 3026
rect 9080 2992 9118 3026
rect 9152 2992 9190 3026
rect 9224 2992 9225 3026
rect 9045 2952 9225 2992
rect 9045 2918 9046 2952
rect 9080 2918 9118 2952
rect 9152 2918 9190 2952
rect 9224 2918 9225 2952
rect 9045 2878 9225 2918
rect 9045 2844 9046 2878
rect 9080 2844 9118 2878
rect 9152 2844 9190 2878
rect 9224 2844 9225 2878
rect 9045 2804 9225 2844
rect 9045 2770 9046 2804
rect 9080 2770 9118 2804
rect 9152 2770 9190 2804
rect 9224 2770 9225 2804
rect 9045 2730 9225 2770
rect 9045 2696 9046 2730
rect 9080 2696 9118 2730
rect 9152 2696 9190 2730
rect 9224 2696 9225 2730
rect 9045 2656 9225 2696
rect 9045 2622 9046 2656
rect 9080 2622 9118 2656
rect 9152 2622 9190 2656
rect 9224 2622 9225 2656
rect 9045 2582 9225 2622
rect 9045 2548 9046 2582
rect 9080 2548 9118 2582
rect 9152 2548 9190 2582
rect 9224 2548 9225 2582
rect 9045 2508 9225 2548
rect 9045 2474 9046 2508
rect 9080 2474 9118 2508
rect 9152 2474 9190 2508
rect 9224 2474 9225 2508
rect 9045 2445 9225 2474
rect 9045 2434 9082 2445
rect 9045 2400 9046 2434
rect 9080 2411 9082 2434
rect 9116 2434 9154 2445
rect 9116 2411 9118 2434
rect 9080 2400 9118 2411
rect 9152 2411 9154 2434
rect 9188 2434 9225 2445
rect 9188 2411 9190 2434
rect 9152 2400 9190 2411
rect 9224 2400 9225 2434
rect 9045 2377 9225 2400
rect 9045 2360 9082 2377
rect 9045 2326 9046 2360
rect 9080 2343 9082 2360
rect 9116 2360 9154 2377
rect 9116 2343 9118 2360
rect 9080 2326 9118 2343
rect 9152 2343 9154 2360
rect 9188 2360 9225 2377
rect 9188 2343 9190 2360
rect 9152 2326 9190 2343
rect 9224 2326 9225 2360
rect 9045 2309 9225 2326
rect 9045 2286 9082 2309
rect 9045 2252 9046 2286
rect 9080 2275 9082 2286
rect 9116 2286 9154 2309
rect 9116 2275 9118 2286
rect 9080 2252 9118 2275
rect 9152 2275 9154 2286
rect 9188 2286 9225 2309
rect 9188 2275 9190 2286
rect 9152 2252 9190 2275
rect 9224 2252 9225 2286
rect 9045 2241 9225 2252
rect 9045 2212 9082 2241
rect 9045 2178 9046 2212
rect 9080 2207 9082 2212
rect 9116 2212 9154 2241
rect 9116 2207 9118 2212
rect 9080 2178 9118 2207
rect 9152 2207 9154 2212
rect 9188 2212 9225 2241
rect 9188 2207 9190 2212
rect 9152 2178 9190 2207
rect 9224 2178 9225 2212
rect 9045 2173 9225 2178
rect 9045 2139 9082 2173
rect 9116 2139 9154 2173
rect 9188 2139 9225 2173
rect 9045 2138 9225 2139
rect 9045 2104 9046 2138
rect 9080 2105 9118 2138
rect 9080 2104 9082 2105
rect 9045 2071 9082 2104
rect 9116 2104 9118 2105
rect 9152 2105 9190 2138
rect 9152 2104 9154 2105
rect 9116 2071 9154 2104
rect 9188 2104 9190 2105
rect 9224 2104 9225 2138
rect 9188 2071 9225 2104
rect 9045 2064 9225 2071
rect 9045 2030 9046 2064
rect 9080 2037 9118 2064
rect 9080 2030 9082 2037
rect 9045 2003 9082 2030
rect 9116 2030 9118 2037
rect 9152 2037 9190 2064
rect 9152 2030 9154 2037
rect 9116 2003 9154 2030
rect 9188 2030 9190 2037
rect 9224 2030 9225 2064
rect 9188 2003 9225 2030
rect 9045 1990 9225 2003
rect 9045 1956 9046 1990
rect 9080 1969 9118 1990
rect 9080 1956 9082 1969
rect 9045 1935 9082 1956
rect 9116 1956 9118 1969
rect 9152 1969 9190 1990
rect 9152 1956 9154 1969
rect 9116 1935 9154 1956
rect 9188 1956 9190 1969
rect 9224 1956 9225 1990
rect 9188 1935 9225 1956
rect 9045 1916 9225 1935
rect 9045 1882 9046 1916
rect 9080 1901 9118 1916
rect 9080 1882 9082 1901
rect 9045 1867 9082 1882
rect 9116 1882 9118 1901
rect 9152 1901 9190 1916
rect 9152 1882 9154 1901
rect 9116 1867 9154 1882
rect 9188 1882 9190 1901
rect 9224 1882 9225 1916
rect 9188 1867 9225 1882
rect 9045 1842 9225 1867
rect 9045 1808 9046 1842
rect 9080 1833 9118 1842
rect 9080 1808 9082 1833
rect 9045 1799 9082 1808
rect 9116 1808 9118 1833
rect 9152 1833 9190 1842
rect 9152 1808 9154 1833
rect 9116 1799 9154 1808
rect 9188 1808 9190 1833
rect 9224 1808 9225 1842
rect 9188 1799 9225 1808
rect 9045 1768 9225 1799
rect 9045 1734 9046 1768
rect 9080 1765 9118 1768
rect 9080 1734 9082 1765
rect 9045 1731 9082 1734
rect 9116 1734 9118 1765
rect 9152 1765 9190 1768
rect 9152 1734 9154 1765
rect 9116 1731 9154 1734
rect 9188 1734 9190 1765
rect 9224 1734 9225 1768
rect 9188 1731 9225 1734
rect 9045 1697 9225 1731
rect 9045 1694 9082 1697
rect 9045 1660 9046 1694
rect 9080 1663 9082 1694
rect 9116 1694 9154 1697
rect 9116 1663 9118 1694
rect 9080 1660 9118 1663
rect 9152 1663 9154 1694
rect 9188 1694 9225 1697
rect 9188 1663 9190 1694
rect 9152 1660 9190 1663
rect 9224 1660 9225 1694
rect 9045 1629 9225 1660
rect 9045 1620 9082 1629
rect 9045 1586 9046 1620
rect 9080 1595 9082 1620
rect 9116 1620 9154 1629
rect 9116 1595 9118 1620
rect 9080 1586 9118 1595
rect 9152 1595 9154 1620
rect 9188 1620 9225 1629
rect 9188 1595 9190 1620
rect 9152 1586 9190 1595
rect 9224 1586 9225 1620
rect 9045 1561 9225 1586
rect 9045 1545 9082 1561
rect 9045 1511 9046 1545
rect 9080 1527 9082 1545
rect 9116 1545 9154 1561
rect 9116 1527 9118 1545
rect 9080 1511 9118 1527
rect 9152 1527 9154 1545
rect 9188 1545 9225 1561
rect 9188 1527 9190 1545
rect 9152 1511 9190 1527
rect 9224 1511 9225 1545
rect 9290 3010 9410 4106
rect 9852 4388 9859 4494
rect 9965 4388 9972 4494
rect 9852 4214 9972 4388
rect 9852 4180 9895 4214
rect 9929 4180 9972 4214
rect 9852 4140 9972 4180
rect 9852 4106 9895 4140
rect 9929 4106 9972 4140
rect 9290 2976 9333 3010
rect 9367 2976 9410 3010
rect 9290 2932 9410 2976
rect 9290 2898 9333 2932
rect 9367 2898 9410 2932
rect 9290 2854 9410 2898
rect 9290 2820 9333 2854
rect 9367 2820 9410 2854
rect 9290 2776 9410 2820
rect 9290 2742 9333 2776
rect 9367 2742 9410 2776
rect 9290 2697 9410 2742
rect 9290 2663 9333 2697
rect 9367 2663 9410 2697
rect 9290 2618 9410 2663
rect 9290 2584 9333 2618
rect 9367 2584 9410 2618
rect 9290 2539 9410 2584
rect 9290 2505 9333 2539
rect 9367 2505 9410 2539
rect 9082 1491 9188 1511
rect 8860 1375 8903 1409
rect 8937 1375 8980 1409
rect 8860 1335 8980 1375
rect 8860 1301 8903 1335
rect 8937 1301 8980 1335
rect 8860 1285 8980 1301
rect 9290 1409 9410 2505
rect 9512 4050 9614 4062
rect 9648 4050 9750 4062
rect 9512 4046 9542 4050
rect 9720 4046 9750 4050
rect 9512 3978 9542 4012
rect 9720 3978 9750 4012
rect 9512 3910 9542 3944
rect 9720 3910 9750 3944
rect 9512 3842 9542 3876
rect 9720 3842 9750 3876
rect 9512 3774 9542 3808
rect 9720 3774 9750 3808
rect 9512 3706 9542 3740
rect 9720 3706 9750 3740
rect 9512 3638 9542 3672
rect 9720 3638 9750 3672
rect 9512 3570 9542 3604
rect 9720 3570 9750 3604
rect 9512 3502 9542 3536
rect 9720 3502 9750 3536
rect 9512 3434 9542 3468
rect 9720 3434 9750 3468
rect 9512 3366 9542 3400
rect 9720 3366 9750 3400
rect 9512 3298 9542 3332
rect 9720 3298 9750 3332
rect 9512 3230 9542 3264
rect 9720 3230 9750 3264
rect 9512 3162 9542 3196
rect 9720 3162 9750 3196
rect 9512 3080 9542 3128
rect 9576 3080 9686 3092
rect 9720 3080 9750 3128
rect 9512 3040 9750 3080
rect 9512 2574 9542 3040
rect 9720 2574 9750 3040
rect 9512 2535 9750 2574
rect 9512 2501 9542 2535
rect 9576 2501 9614 2535
rect 9648 2501 9686 2535
rect 9720 2501 9750 2535
rect 9512 2461 9750 2501
rect 9512 2449 9614 2461
rect 9648 2449 9750 2461
rect 9512 2445 9542 2449
rect 9720 2445 9750 2449
rect 9512 2377 9542 2411
rect 9720 2377 9750 2411
rect 9512 2309 9542 2343
rect 9720 2309 9750 2343
rect 9512 2241 9542 2275
rect 9720 2241 9750 2275
rect 9512 2173 9542 2207
rect 9720 2173 9750 2207
rect 9512 2105 9542 2139
rect 9720 2105 9750 2139
rect 9512 2037 9542 2071
rect 9720 2037 9750 2071
rect 9512 1969 9542 2003
rect 9720 1969 9750 2003
rect 9512 1901 9542 1935
rect 9720 1901 9750 1935
rect 9512 1833 9542 1867
rect 9720 1833 9750 1867
rect 9512 1765 9542 1799
rect 9720 1765 9750 1799
rect 9512 1697 9542 1731
rect 9720 1697 9750 1731
rect 9512 1629 9542 1663
rect 9720 1629 9750 1663
rect 9512 1561 9542 1595
rect 9720 1561 9750 1595
rect 9512 1479 9542 1527
rect 9576 1479 9686 1491
rect 9720 1479 9750 1527
rect 9512 1464 9750 1479
rect 9852 3010 9972 4106
rect 10282 4388 10289 4494
rect 10395 4388 10402 4494
rect 10282 4214 10402 4388
rect 10282 4180 10325 4214
rect 10359 4180 10402 4214
rect 10282 4140 10402 4180
rect 10282 4106 10325 4140
rect 10359 4106 10402 4140
rect 9852 2976 9895 3010
rect 9929 2976 9972 3010
rect 9852 2932 9972 2976
rect 9852 2898 9895 2932
rect 9929 2898 9972 2932
rect 9852 2854 9972 2898
rect 9852 2820 9895 2854
rect 9929 2820 9972 2854
rect 9852 2776 9972 2820
rect 9852 2742 9895 2776
rect 9929 2742 9972 2776
rect 9852 2697 9972 2742
rect 9852 2663 9895 2697
rect 9929 2663 9972 2697
rect 9852 2618 9972 2663
rect 9852 2584 9895 2618
rect 9929 2584 9972 2618
rect 9852 2539 9972 2584
rect 9852 2505 9895 2539
rect 9929 2505 9972 2539
rect 9290 1375 9333 1409
rect 9367 1375 9410 1409
rect 9290 1335 9410 1375
rect 9290 1301 9333 1335
rect 9367 1301 9410 1335
rect 9290 1285 9410 1301
rect 9852 1409 9972 2505
rect 10037 4028 10038 4062
rect 10072 4046 10110 4062
rect 10072 4028 10074 4046
rect 10037 4012 10074 4028
rect 10108 4028 10110 4046
rect 10144 4046 10182 4062
rect 10144 4028 10146 4046
rect 10108 4012 10146 4028
rect 10180 4028 10182 4046
rect 10216 4028 10217 4062
rect 10180 4012 10217 4028
rect 10037 3988 10217 4012
rect 10037 3954 10038 3988
rect 10072 3978 10110 3988
rect 10072 3954 10074 3978
rect 10037 3944 10074 3954
rect 10108 3954 10110 3978
rect 10144 3978 10182 3988
rect 10144 3954 10146 3978
rect 10108 3944 10146 3954
rect 10180 3954 10182 3978
rect 10216 3954 10217 3988
rect 10180 3944 10217 3954
rect 10037 3914 10217 3944
rect 10037 3880 10038 3914
rect 10072 3910 10110 3914
rect 10072 3880 10074 3910
rect 10037 3876 10074 3880
rect 10108 3880 10110 3910
rect 10144 3910 10182 3914
rect 10144 3880 10146 3910
rect 10108 3876 10146 3880
rect 10180 3880 10182 3910
rect 10216 3880 10217 3914
rect 10180 3876 10217 3880
rect 10037 3842 10217 3876
rect 10037 3840 10074 3842
rect 10037 3806 10038 3840
rect 10072 3808 10074 3840
rect 10108 3840 10146 3842
rect 10108 3808 10110 3840
rect 10072 3806 10110 3808
rect 10144 3808 10146 3840
rect 10180 3840 10217 3842
rect 10180 3808 10182 3840
rect 10144 3806 10182 3808
rect 10216 3806 10217 3840
rect 10037 3774 10217 3806
rect 10037 3766 10074 3774
rect 10037 3732 10038 3766
rect 10072 3740 10074 3766
rect 10108 3766 10146 3774
rect 10108 3740 10110 3766
rect 10072 3732 10110 3740
rect 10144 3740 10146 3766
rect 10180 3766 10217 3774
rect 10180 3740 10182 3766
rect 10144 3732 10182 3740
rect 10216 3732 10217 3766
rect 10037 3706 10217 3732
rect 10037 3692 10074 3706
rect 10037 3658 10038 3692
rect 10072 3672 10074 3692
rect 10108 3692 10146 3706
rect 10108 3672 10110 3692
rect 10072 3658 10110 3672
rect 10144 3672 10146 3692
rect 10180 3692 10217 3706
rect 10180 3672 10182 3692
rect 10144 3658 10182 3672
rect 10216 3658 10217 3692
rect 10037 3638 10217 3658
rect 10037 3618 10074 3638
rect 10037 3584 10038 3618
rect 10072 3604 10074 3618
rect 10108 3618 10146 3638
rect 10108 3604 10110 3618
rect 10072 3584 10110 3604
rect 10144 3604 10146 3618
rect 10180 3618 10217 3638
rect 10180 3604 10182 3618
rect 10144 3584 10182 3604
rect 10216 3584 10217 3618
rect 10037 3570 10217 3584
rect 10037 3544 10074 3570
rect 10037 3510 10038 3544
rect 10072 3536 10074 3544
rect 10108 3544 10146 3570
rect 10108 3536 10110 3544
rect 10072 3510 10110 3536
rect 10144 3536 10146 3544
rect 10180 3544 10217 3570
rect 10180 3536 10182 3544
rect 10144 3510 10182 3536
rect 10216 3510 10217 3544
rect 10037 3502 10217 3510
rect 10037 3470 10074 3502
rect 10037 3436 10038 3470
rect 10072 3468 10074 3470
rect 10108 3470 10146 3502
rect 10108 3468 10110 3470
rect 10072 3436 10110 3468
rect 10144 3468 10146 3470
rect 10180 3470 10217 3502
rect 10180 3468 10182 3470
rect 10144 3436 10182 3468
rect 10216 3436 10217 3470
rect 10037 3434 10217 3436
rect 10037 3400 10074 3434
rect 10108 3400 10146 3434
rect 10180 3400 10217 3434
rect 10037 3396 10217 3400
rect 10037 3362 10038 3396
rect 10072 3366 10110 3396
rect 10072 3362 10074 3366
rect 10037 3332 10074 3362
rect 10108 3362 10110 3366
rect 10144 3366 10182 3396
rect 10144 3362 10146 3366
rect 10108 3332 10146 3362
rect 10180 3362 10182 3366
rect 10216 3362 10217 3396
rect 10180 3332 10217 3362
rect 10037 3322 10217 3332
rect 10037 3288 10038 3322
rect 10072 3298 10110 3322
rect 10072 3288 10074 3298
rect 10037 3264 10074 3288
rect 10108 3288 10110 3298
rect 10144 3298 10182 3322
rect 10144 3288 10146 3298
rect 10108 3264 10146 3288
rect 10180 3288 10182 3298
rect 10216 3288 10217 3322
rect 10180 3264 10217 3288
rect 10037 3248 10217 3264
rect 10037 3214 10038 3248
rect 10072 3230 10110 3248
rect 10072 3214 10074 3230
rect 10037 3196 10074 3214
rect 10108 3214 10110 3230
rect 10144 3230 10182 3248
rect 10144 3214 10146 3230
rect 10108 3196 10146 3214
rect 10180 3214 10182 3230
rect 10216 3214 10217 3248
rect 10180 3196 10217 3214
rect 10037 3174 10217 3196
rect 10037 3140 10038 3174
rect 10072 3162 10110 3174
rect 10072 3140 10074 3162
rect 10037 3128 10074 3140
rect 10108 3140 10110 3162
rect 10144 3162 10182 3174
rect 10144 3140 10146 3162
rect 10108 3128 10146 3140
rect 10180 3140 10182 3162
rect 10216 3140 10217 3174
rect 10180 3128 10217 3140
rect 10037 3100 10217 3128
rect 10037 3066 10038 3100
rect 10072 3066 10110 3100
rect 10144 3066 10182 3100
rect 10216 3066 10217 3100
rect 10037 3026 10217 3066
rect 10037 2992 10038 3026
rect 10072 2992 10110 3026
rect 10144 2992 10182 3026
rect 10216 2992 10217 3026
rect 10037 2952 10217 2992
rect 10037 2918 10038 2952
rect 10072 2918 10110 2952
rect 10144 2918 10182 2952
rect 10216 2918 10217 2952
rect 10037 2878 10217 2918
rect 10037 2844 10038 2878
rect 10072 2844 10110 2878
rect 10144 2844 10182 2878
rect 10216 2844 10217 2878
rect 10037 2804 10217 2844
rect 10037 2770 10038 2804
rect 10072 2770 10110 2804
rect 10144 2770 10182 2804
rect 10216 2770 10217 2804
rect 10037 2730 10217 2770
rect 10037 2696 10038 2730
rect 10072 2696 10110 2730
rect 10144 2696 10182 2730
rect 10216 2696 10217 2730
rect 10037 2656 10217 2696
rect 10037 2622 10038 2656
rect 10072 2622 10110 2656
rect 10144 2622 10182 2656
rect 10216 2622 10217 2656
rect 10037 2582 10217 2622
rect 10037 2548 10038 2582
rect 10072 2548 10110 2582
rect 10144 2548 10182 2582
rect 10216 2548 10217 2582
rect 10037 2508 10217 2548
rect 10037 2474 10038 2508
rect 10072 2474 10110 2508
rect 10144 2474 10182 2508
rect 10216 2474 10217 2508
rect 10037 2445 10217 2474
rect 10037 2434 10074 2445
rect 10037 2400 10038 2434
rect 10072 2411 10074 2434
rect 10108 2434 10146 2445
rect 10108 2411 10110 2434
rect 10072 2400 10110 2411
rect 10144 2411 10146 2434
rect 10180 2434 10217 2445
rect 10180 2411 10182 2434
rect 10144 2400 10182 2411
rect 10216 2400 10217 2434
rect 10037 2377 10217 2400
rect 10037 2360 10074 2377
rect 10037 2326 10038 2360
rect 10072 2343 10074 2360
rect 10108 2360 10146 2377
rect 10108 2343 10110 2360
rect 10072 2326 10110 2343
rect 10144 2343 10146 2360
rect 10180 2360 10217 2377
rect 10180 2343 10182 2360
rect 10144 2326 10182 2343
rect 10216 2326 10217 2360
rect 10037 2309 10217 2326
rect 10037 2286 10074 2309
rect 10037 2252 10038 2286
rect 10072 2275 10074 2286
rect 10108 2286 10146 2309
rect 10108 2275 10110 2286
rect 10072 2252 10110 2275
rect 10144 2275 10146 2286
rect 10180 2286 10217 2309
rect 10180 2275 10182 2286
rect 10144 2252 10182 2275
rect 10216 2252 10217 2286
rect 10037 2241 10217 2252
rect 10037 2212 10074 2241
rect 10037 2178 10038 2212
rect 10072 2207 10074 2212
rect 10108 2212 10146 2241
rect 10108 2207 10110 2212
rect 10072 2178 10110 2207
rect 10144 2207 10146 2212
rect 10180 2212 10217 2241
rect 10180 2207 10182 2212
rect 10144 2178 10182 2207
rect 10216 2178 10217 2212
rect 10037 2173 10217 2178
rect 10037 2139 10074 2173
rect 10108 2139 10146 2173
rect 10180 2139 10217 2173
rect 10037 2138 10217 2139
rect 10037 2104 10038 2138
rect 10072 2105 10110 2138
rect 10072 2104 10074 2105
rect 10037 2071 10074 2104
rect 10108 2104 10110 2105
rect 10144 2105 10182 2138
rect 10144 2104 10146 2105
rect 10108 2071 10146 2104
rect 10180 2104 10182 2105
rect 10216 2104 10217 2138
rect 10180 2071 10217 2104
rect 10037 2064 10217 2071
rect 10037 2030 10038 2064
rect 10072 2037 10110 2064
rect 10072 2030 10074 2037
rect 10037 2003 10074 2030
rect 10108 2030 10110 2037
rect 10144 2037 10182 2064
rect 10144 2030 10146 2037
rect 10108 2003 10146 2030
rect 10180 2030 10182 2037
rect 10216 2030 10217 2064
rect 10180 2003 10217 2030
rect 10037 1990 10217 2003
rect 10037 1956 10038 1990
rect 10072 1969 10110 1990
rect 10072 1956 10074 1969
rect 10037 1935 10074 1956
rect 10108 1956 10110 1969
rect 10144 1969 10182 1990
rect 10144 1956 10146 1969
rect 10108 1935 10146 1956
rect 10180 1956 10182 1969
rect 10216 1956 10217 1990
rect 10180 1935 10217 1956
rect 10037 1916 10217 1935
rect 10037 1882 10038 1916
rect 10072 1901 10110 1916
rect 10072 1882 10074 1901
rect 10037 1867 10074 1882
rect 10108 1882 10110 1901
rect 10144 1901 10182 1916
rect 10144 1882 10146 1901
rect 10108 1867 10146 1882
rect 10180 1882 10182 1901
rect 10216 1882 10217 1916
rect 10180 1867 10217 1882
rect 10037 1842 10217 1867
rect 10037 1808 10038 1842
rect 10072 1833 10110 1842
rect 10072 1808 10074 1833
rect 10037 1799 10074 1808
rect 10108 1808 10110 1833
rect 10144 1833 10182 1842
rect 10144 1808 10146 1833
rect 10108 1799 10146 1808
rect 10180 1808 10182 1833
rect 10216 1808 10217 1842
rect 10180 1799 10217 1808
rect 10037 1768 10217 1799
rect 10037 1734 10038 1768
rect 10072 1765 10110 1768
rect 10072 1734 10074 1765
rect 10037 1731 10074 1734
rect 10108 1734 10110 1765
rect 10144 1765 10182 1768
rect 10144 1734 10146 1765
rect 10108 1731 10146 1734
rect 10180 1734 10182 1765
rect 10216 1734 10217 1768
rect 10180 1731 10217 1734
rect 10037 1697 10217 1731
rect 10037 1694 10074 1697
rect 10037 1660 10038 1694
rect 10072 1663 10074 1694
rect 10108 1694 10146 1697
rect 10108 1663 10110 1694
rect 10072 1660 10110 1663
rect 10144 1663 10146 1694
rect 10180 1694 10217 1697
rect 10180 1663 10182 1694
rect 10144 1660 10182 1663
rect 10216 1660 10217 1694
rect 10037 1629 10217 1660
rect 10037 1620 10074 1629
rect 10037 1586 10038 1620
rect 10072 1595 10074 1620
rect 10108 1620 10146 1629
rect 10108 1595 10110 1620
rect 10072 1586 10110 1595
rect 10144 1595 10146 1620
rect 10180 1620 10217 1629
rect 10180 1595 10182 1620
rect 10144 1586 10182 1595
rect 10216 1586 10217 1620
rect 10037 1561 10217 1586
rect 10037 1545 10074 1561
rect 10037 1511 10038 1545
rect 10072 1527 10074 1545
rect 10108 1545 10146 1561
rect 10108 1527 10110 1545
rect 10072 1511 10110 1527
rect 10144 1527 10146 1545
rect 10180 1545 10217 1561
rect 10180 1527 10182 1545
rect 10144 1511 10182 1527
rect 10216 1511 10217 1545
rect 10282 3010 10402 4106
rect 10844 4388 10851 4494
rect 10957 4388 10964 4494
rect 10844 4214 10964 4388
rect 10844 4180 10887 4214
rect 10921 4180 10964 4214
rect 10844 4140 10964 4180
rect 10844 4106 10887 4140
rect 10921 4106 10964 4140
rect 10282 2976 10325 3010
rect 10359 2976 10402 3010
rect 10282 2932 10402 2976
rect 10282 2898 10325 2932
rect 10359 2898 10402 2932
rect 10282 2854 10402 2898
rect 10282 2820 10325 2854
rect 10359 2820 10402 2854
rect 10282 2776 10402 2820
rect 10282 2742 10325 2776
rect 10359 2742 10402 2776
rect 10282 2697 10402 2742
rect 10282 2663 10325 2697
rect 10359 2663 10402 2697
rect 10282 2618 10402 2663
rect 10282 2584 10325 2618
rect 10359 2584 10402 2618
rect 10282 2539 10402 2584
rect 10282 2505 10325 2539
rect 10359 2505 10402 2539
rect 10074 1491 10180 1511
rect 9852 1375 9895 1409
rect 9929 1375 9972 1409
rect 9852 1335 9972 1375
rect 9852 1301 9895 1335
rect 9929 1301 9972 1335
rect 9852 1285 9972 1301
rect 10282 1409 10402 2505
rect 10504 4050 10606 4062
rect 10640 4050 10742 4062
rect 10504 4046 10534 4050
rect 10712 4046 10742 4050
rect 10504 3978 10534 4012
rect 10712 3978 10742 4012
rect 10504 3910 10534 3944
rect 10712 3910 10742 3944
rect 10504 3842 10534 3876
rect 10712 3842 10742 3876
rect 10504 3774 10534 3808
rect 10712 3774 10742 3808
rect 10504 3706 10534 3740
rect 10712 3706 10742 3740
rect 10504 3638 10534 3672
rect 10712 3638 10742 3672
rect 10504 3570 10534 3604
rect 10712 3570 10742 3604
rect 10504 3502 10534 3536
rect 10712 3502 10742 3536
rect 10504 3434 10534 3468
rect 10712 3434 10742 3468
rect 10504 3366 10534 3400
rect 10712 3366 10742 3400
rect 10504 3298 10534 3332
rect 10712 3298 10742 3332
rect 10504 3230 10534 3264
rect 10712 3230 10742 3264
rect 10504 3162 10534 3196
rect 10712 3162 10742 3196
rect 10504 3080 10534 3128
rect 10568 3080 10678 3092
rect 10712 3080 10742 3128
rect 10504 3037 10742 3080
rect 10504 3003 10534 3037
rect 10568 3003 10606 3037
rect 10640 3003 10678 3037
rect 10712 3003 10742 3037
rect 10504 2954 10742 3003
rect 10504 2920 10534 2954
rect 10568 2935 10606 2954
rect 10640 2935 10678 2954
rect 10568 2920 10573 2935
rect 10640 2920 10641 2935
rect 10504 2901 10573 2920
rect 10607 2901 10641 2920
rect 10675 2920 10678 2935
rect 10712 2920 10742 2954
rect 10675 2901 10742 2920
rect 10504 2871 10742 2901
rect 10504 2837 10534 2871
rect 10568 2855 10606 2871
rect 10640 2855 10678 2871
rect 10568 2837 10573 2855
rect 10640 2837 10641 2855
rect 10504 2821 10573 2837
rect 10607 2821 10641 2837
rect 10675 2837 10678 2855
rect 10712 2837 10742 2871
rect 10675 2821 10742 2837
rect 10504 2787 10742 2821
rect 10504 2753 10534 2787
rect 10568 2775 10606 2787
rect 10640 2775 10678 2787
rect 10568 2753 10573 2775
rect 10640 2753 10641 2775
rect 10504 2741 10573 2753
rect 10607 2741 10641 2753
rect 10675 2753 10678 2775
rect 10712 2753 10742 2787
rect 10675 2741 10742 2753
rect 10504 2703 10742 2741
rect 10504 2669 10534 2703
rect 10568 2695 10606 2703
rect 10640 2695 10678 2703
rect 10568 2669 10573 2695
rect 10640 2669 10641 2695
rect 10504 2661 10573 2669
rect 10607 2661 10641 2669
rect 10675 2669 10678 2695
rect 10712 2669 10742 2703
rect 10675 2661 10742 2669
rect 10504 2619 10742 2661
rect 10504 2585 10534 2619
rect 10568 2614 10606 2619
rect 10640 2614 10678 2619
rect 10568 2585 10573 2614
rect 10640 2585 10641 2614
rect 10504 2580 10573 2585
rect 10607 2580 10641 2585
rect 10675 2585 10678 2614
rect 10712 2585 10742 2619
rect 10675 2580 10742 2585
rect 10504 2535 10742 2580
rect 10504 2501 10534 2535
rect 10568 2501 10606 2535
rect 10640 2501 10678 2535
rect 10712 2501 10742 2535
rect 10504 2461 10742 2501
rect 10504 2449 10606 2461
rect 10640 2449 10742 2461
rect 10504 2445 10534 2449
rect 10712 2445 10742 2449
rect 10504 2377 10534 2411
rect 10712 2377 10742 2411
rect 10504 2309 10534 2343
rect 10712 2309 10742 2343
rect 10504 2241 10534 2275
rect 10712 2241 10742 2275
rect 10504 2173 10534 2207
rect 10712 2173 10742 2207
rect 10504 2105 10534 2139
rect 10712 2105 10742 2139
rect 10504 2037 10534 2071
rect 10712 2037 10742 2071
rect 10504 1969 10534 2003
rect 10712 1969 10742 2003
rect 10504 1901 10534 1935
rect 10712 1901 10742 1935
rect 10504 1833 10534 1867
rect 10712 1833 10742 1867
rect 10504 1765 10534 1799
rect 10712 1765 10742 1799
rect 10504 1697 10534 1731
rect 10712 1697 10742 1731
rect 10504 1629 10534 1663
rect 10712 1629 10742 1663
rect 10504 1561 10534 1595
rect 10712 1561 10742 1595
rect 10504 1479 10534 1527
rect 10568 1479 10678 1491
rect 10712 1479 10742 1527
rect 10504 1464 10742 1479
rect 10844 3010 10964 4106
rect 11274 4388 11281 4494
rect 11387 4388 11394 4494
rect 11274 4214 11394 4388
rect 11274 4180 11317 4214
rect 11351 4180 11394 4214
rect 11274 4140 11394 4180
rect 11274 4106 11317 4140
rect 11351 4106 11394 4140
rect 10844 2976 10887 3010
rect 10921 2976 10964 3010
rect 10844 2932 10964 2976
rect 10844 2898 10887 2932
rect 10921 2898 10964 2932
rect 10844 2854 10964 2898
rect 10844 2820 10887 2854
rect 10921 2820 10964 2854
rect 10844 2776 10964 2820
rect 10844 2742 10887 2776
rect 10921 2742 10964 2776
rect 10844 2697 10964 2742
rect 10844 2663 10887 2697
rect 10921 2663 10964 2697
rect 10844 2618 10964 2663
rect 10844 2584 10887 2618
rect 10921 2584 10964 2618
rect 10844 2539 10964 2584
rect 10844 2505 10887 2539
rect 10921 2505 10964 2539
rect 10282 1375 10325 1409
rect 10359 1375 10402 1409
rect 10282 1335 10402 1375
rect 10282 1301 10325 1335
rect 10359 1301 10402 1335
rect 10282 1285 10402 1301
rect 10844 1409 10964 2505
rect 11029 4028 11030 4062
rect 11064 4046 11102 4062
rect 11064 4028 11066 4046
rect 11029 4012 11066 4028
rect 11100 4028 11102 4046
rect 11136 4046 11174 4062
rect 11136 4028 11138 4046
rect 11100 4012 11138 4028
rect 11172 4028 11174 4046
rect 11208 4028 11209 4062
rect 11172 4012 11209 4028
rect 11029 3988 11209 4012
rect 11029 3954 11030 3988
rect 11064 3978 11102 3988
rect 11064 3954 11066 3978
rect 11029 3944 11066 3954
rect 11100 3954 11102 3978
rect 11136 3978 11174 3988
rect 11136 3954 11138 3978
rect 11100 3944 11138 3954
rect 11172 3954 11174 3978
rect 11208 3954 11209 3988
rect 11172 3944 11209 3954
rect 11029 3914 11209 3944
rect 11029 3880 11030 3914
rect 11064 3910 11102 3914
rect 11064 3880 11066 3910
rect 11029 3876 11066 3880
rect 11100 3880 11102 3910
rect 11136 3910 11174 3914
rect 11136 3880 11138 3910
rect 11100 3876 11138 3880
rect 11172 3880 11174 3910
rect 11208 3880 11209 3914
rect 11172 3876 11209 3880
rect 11029 3842 11209 3876
rect 11029 3840 11066 3842
rect 11029 3806 11030 3840
rect 11064 3808 11066 3840
rect 11100 3840 11138 3842
rect 11100 3808 11102 3840
rect 11064 3806 11102 3808
rect 11136 3808 11138 3840
rect 11172 3840 11209 3842
rect 11172 3808 11174 3840
rect 11136 3806 11174 3808
rect 11208 3806 11209 3840
rect 11029 3774 11209 3806
rect 11029 3766 11066 3774
rect 11029 3732 11030 3766
rect 11064 3740 11066 3766
rect 11100 3766 11138 3774
rect 11100 3740 11102 3766
rect 11064 3732 11102 3740
rect 11136 3740 11138 3766
rect 11172 3766 11209 3774
rect 11172 3740 11174 3766
rect 11136 3732 11174 3740
rect 11208 3732 11209 3766
rect 11029 3706 11209 3732
rect 11029 3692 11066 3706
rect 11029 3658 11030 3692
rect 11064 3672 11066 3692
rect 11100 3692 11138 3706
rect 11100 3672 11102 3692
rect 11064 3658 11102 3672
rect 11136 3672 11138 3692
rect 11172 3692 11209 3706
rect 11172 3672 11174 3692
rect 11136 3658 11174 3672
rect 11208 3658 11209 3692
rect 11029 3638 11209 3658
rect 11029 3618 11066 3638
rect 11029 3584 11030 3618
rect 11064 3604 11066 3618
rect 11100 3618 11138 3638
rect 11100 3604 11102 3618
rect 11064 3584 11102 3604
rect 11136 3604 11138 3618
rect 11172 3618 11209 3638
rect 11172 3604 11174 3618
rect 11136 3584 11174 3604
rect 11208 3584 11209 3618
rect 11029 3570 11209 3584
rect 11029 3544 11066 3570
rect 11029 3510 11030 3544
rect 11064 3536 11066 3544
rect 11100 3544 11138 3570
rect 11100 3536 11102 3544
rect 11064 3510 11102 3536
rect 11136 3536 11138 3544
rect 11172 3544 11209 3570
rect 11172 3536 11174 3544
rect 11136 3510 11174 3536
rect 11208 3510 11209 3544
rect 11029 3502 11209 3510
rect 11029 3470 11066 3502
rect 11029 3436 11030 3470
rect 11064 3468 11066 3470
rect 11100 3470 11138 3502
rect 11100 3468 11102 3470
rect 11064 3436 11102 3468
rect 11136 3468 11138 3470
rect 11172 3470 11209 3502
rect 11172 3468 11174 3470
rect 11136 3436 11174 3468
rect 11208 3436 11209 3470
rect 11029 3434 11209 3436
rect 11029 3400 11066 3434
rect 11100 3400 11138 3434
rect 11172 3400 11209 3434
rect 11029 3396 11209 3400
rect 11029 3362 11030 3396
rect 11064 3366 11102 3396
rect 11064 3362 11066 3366
rect 11029 3332 11066 3362
rect 11100 3362 11102 3366
rect 11136 3366 11174 3396
rect 11136 3362 11138 3366
rect 11100 3332 11138 3362
rect 11172 3362 11174 3366
rect 11208 3362 11209 3396
rect 11172 3332 11209 3362
rect 11029 3322 11209 3332
rect 11029 3288 11030 3322
rect 11064 3298 11102 3322
rect 11064 3288 11066 3298
rect 11029 3264 11066 3288
rect 11100 3288 11102 3298
rect 11136 3298 11174 3322
rect 11136 3288 11138 3298
rect 11100 3264 11138 3288
rect 11172 3288 11174 3298
rect 11208 3288 11209 3322
rect 11172 3264 11209 3288
rect 11029 3248 11209 3264
rect 11029 3214 11030 3248
rect 11064 3230 11102 3248
rect 11064 3214 11066 3230
rect 11029 3196 11066 3214
rect 11100 3214 11102 3230
rect 11136 3230 11174 3248
rect 11136 3214 11138 3230
rect 11100 3196 11138 3214
rect 11172 3214 11174 3230
rect 11208 3214 11209 3248
rect 11172 3196 11209 3214
rect 11029 3174 11209 3196
rect 11029 3140 11030 3174
rect 11064 3162 11102 3174
rect 11064 3140 11066 3162
rect 11029 3128 11066 3140
rect 11100 3140 11102 3162
rect 11136 3162 11174 3174
rect 11136 3140 11138 3162
rect 11100 3128 11138 3140
rect 11172 3140 11174 3162
rect 11208 3140 11209 3174
rect 11172 3128 11209 3140
rect 11029 3100 11209 3128
rect 11029 3066 11030 3100
rect 11064 3066 11102 3100
rect 11136 3066 11174 3100
rect 11208 3066 11209 3100
rect 11029 3026 11209 3066
rect 11029 2992 11030 3026
rect 11064 2992 11102 3026
rect 11136 2992 11174 3026
rect 11208 2992 11209 3026
rect 11029 2952 11209 2992
rect 11029 2918 11030 2952
rect 11064 2918 11102 2952
rect 11136 2918 11174 2952
rect 11208 2918 11209 2952
rect 11029 2878 11209 2918
rect 11029 2844 11030 2878
rect 11064 2844 11102 2878
rect 11136 2844 11174 2878
rect 11208 2844 11209 2878
rect 11029 2804 11209 2844
rect 11029 2770 11030 2804
rect 11064 2770 11102 2804
rect 11136 2770 11174 2804
rect 11208 2770 11209 2804
rect 11029 2730 11209 2770
rect 11029 2696 11030 2730
rect 11064 2696 11102 2730
rect 11136 2696 11174 2730
rect 11208 2696 11209 2730
rect 11029 2656 11209 2696
rect 11029 2622 11030 2656
rect 11064 2622 11102 2656
rect 11136 2622 11174 2656
rect 11208 2622 11209 2656
rect 11029 2582 11209 2622
rect 11029 2548 11030 2582
rect 11064 2548 11102 2582
rect 11136 2548 11174 2582
rect 11208 2548 11209 2582
rect 11029 2508 11209 2548
rect 11029 2474 11030 2508
rect 11064 2474 11102 2508
rect 11136 2474 11174 2508
rect 11208 2474 11209 2508
rect 11029 2445 11209 2474
rect 11029 2434 11066 2445
rect 11029 2400 11030 2434
rect 11064 2411 11066 2434
rect 11100 2434 11138 2445
rect 11100 2411 11102 2434
rect 11064 2400 11102 2411
rect 11136 2411 11138 2434
rect 11172 2434 11209 2445
rect 11172 2411 11174 2434
rect 11136 2400 11174 2411
rect 11208 2400 11209 2434
rect 11029 2377 11209 2400
rect 11029 2360 11066 2377
rect 11029 2326 11030 2360
rect 11064 2343 11066 2360
rect 11100 2360 11138 2377
rect 11100 2343 11102 2360
rect 11064 2326 11102 2343
rect 11136 2343 11138 2360
rect 11172 2360 11209 2377
rect 11172 2343 11174 2360
rect 11136 2326 11174 2343
rect 11208 2326 11209 2360
rect 11029 2309 11209 2326
rect 11029 2286 11066 2309
rect 11029 2252 11030 2286
rect 11064 2275 11066 2286
rect 11100 2286 11138 2309
rect 11100 2275 11102 2286
rect 11064 2252 11102 2275
rect 11136 2275 11138 2286
rect 11172 2286 11209 2309
rect 11172 2275 11174 2286
rect 11136 2252 11174 2275
rect 11208 2252 11209 2286
rect 11029 2241 11209 2252
rect 11029 2212 11066 2241
rect 11029 2178 11030 2212
rect 11064 2207 11066 2212
rect 11100 2212 11138 2241
rect 11100 2207 11102 2212
rect 11064 2178 11102 2207
rect 11136 2207 11138 2212
rect 11172 2212 11209 2241
rect 11172 2207 11174 2212
rect 11136 2178 11174 2207
rect 11208 2178 11209 2212
rect 11029 2173 11209 2178
rect 11029 2139 11066 2173
rect 11100 2139 11138 2173
rect 11172 2139 11209 2173
rect 11029 2138 11209 2139
rect 11029 2104 11030 2138
rect 11064 2105 11102 2138
rect 11064 2104 11066 2105
rect 11029 2071 11066 2104
rect 11100 2104 11102 2105
rect 11136 2105 11174 2138
rect 11136 2104 11138 2105
rect 11100 2071 11138 2104
rect 11172 2104 11174 2105
rect 11208 2104 11209 2138
rect 11172 2071 11209 2104
rect 11029 2064 11209 2071
rect 11029 2030 11030 2064
rect 11064 2037 11102 2064
rect 11064 2030 11066 2037
rect 11029 2003 11066 2030
rect 11100 2030 11102 2037
rect 11136 2037 11174 2064
rect 11136 2030 11138 2037
rect 11100 2003 11138 2030
rect 11172 2030 11174 2037
rect 11208 2030 11209 2064
rect 11172 2003 11209 2030
rect 11029 1990 11209 2003
rect 11029 1956 11030 1990
rect 11064 1969 11102 1990
rect 11064 1956 11066 1969
rect 11029 1935 11066 1956
rect 11100 1956 11102 1969
rect 11136 1969 11174 1990
rect 11136 1956 11138 1969
rect 11100 1935 11138 1956
rect 11172 1956 11174 1969
rect 11208 1956 11209 1990
rect 11172 1935 11209 1956
rect 11029 1916 11209 1935
rect 11029 1882 11030 1916
rect 11064 1901 11102 1916
rect 11064 1882 11066 1901
rect 11029 1867 11066 1882
rect 11100 1882 11102 1901
rect 11136 1901 11174 1916
rect 11136 1882 11138 1901
rect 11100 1867 11138 1882
rect 11172 1882 11174 1901
rect 11208 1882 11209 1916
rect 11172 1867 11209 1882
rect 11029 1842 11209 1867
rect 11029 1808 11030 1842
rect 11064 1833 11102 1842
rect 11064 1808 11066 1833
rect 11029 1799 11066 1808
rect 11100 1808 11102 1833
rect 11136 1833 11174 1842
rect 11136 1808 11138 1833
rect 11100 1799 11138 1808
rect 11172 1808 11174 1833
rect 11208 1808 11209 1842
rect 11172 1799 11209 1808
rect 11029 1768 11209 1799
rect 11029 1734 11030 1768
rect 11064 1765 11102 1768
rect 11064 1734 11066 1765
rect 11029 1731 11066 1734
rect 11100 1734 11102 1765
rect 11136 1765 11174 1768
rect 11136 1734 11138 1765
rect 11100 1731 11138 1734
rect 11172 1734 11174 1765
rect 11208 1734 11209 1768
rect 11172 1731 11209 1734
rect 11029 1697 11209 1731
rect 11029 1694 11066 1697
rect 11029 1660 11030 1694
rect 11064 1663 11066 1694
rect 11100 1694 11138 1697
rect 11100 1663 11102 1694
rect 11064 1660 11102 1663
rect 11136 1663 11138 1694
rect 11172 1694 11209 1697
rect 11172 1663 11174 1694
rect 11136 1660 11174 1663
rect 11208 1660 11209 1694
rect 11029 1629 11209 1660
rect 11029 1620 11066 1629
rect 11029 1586 11030 1620
rect 11064 1595 11066 1620
rect 11100 1620 11138 1629
rect 11100 1595 11102 1620
rect 11064 1586 11102 1595
rect 11136 1595 11138 1620
rect 11172 1620 11209 1629
rect 11172 1595 11174 1620
rect 11136 1586 11174 1595
rect 11208 1586 11209 1620
rect 11029 1561 11209 1586
rect 11029 1545 11066 1561
rect 11029 1511 11030 1545
rect 11064 1527 11066 1545
rect 11100 1545 11138 1561
rect 11100 1527 11102 1545
rect 11064 1511 11102 1527
rect 11136 1527 11138 1545
rect 11172 1545 11209 1561
rect 11172 1527 11174 1545
rect 11136 1511 11174 1527
rect 11208 1511 11209 1545
rect 11274 3010 11394 4106
rect 11836 4388 11843 4494
rect 11949 4388 11956 4494
rect 11836 4214 11956 4388
rect 11836 4180 11879 4214
rect 11913 4180 11956 4214
rect 11836 4140 11956 4180
rect 11836 4106 11879 4140
rect 11913 4106 11956 4140
rect 11274 2976 11317 3010
rect 11351 2976 11394 3010
rect 11274 2932 11394 2976
rect 11274 2898 11317 2932
rect 11351 2898 11394 2932
rect 11274 2854 11394 2898
rect 11274 2820 11317 2854
rect 11351 2820 11394 2854
rect 11274 2776 11394 2820
rect 11274 2742 11317 2776
rect 11351 2742 11394 2776
rect 11274 2697 11394 2742
rect 11274 2663 11317 2697
rect 11351 2663 11394 2697
rect 11274 2618 11394 2663
rect 11274 2584 11317 2618
rect 11351 2584 11394 2618
rect 11274 2539 11394 2584
rect 11274 2505 11317 2539
rect 11351 2505 11394 2539
rect 11066 1491 11172 1511
rect 10844 1375 10887 1409
rect 10921 1375 10964 1409
rect 10844 1335 10964 1375
rect 10844 1301 10887 1335
rect 10921 1301 10964 1335
rect 10844 1285 10964 1301
rect 11274 1409 11394 2505
rect 11496 4050 11598 4062
rect 11632 4050 11734 4062
rect 11496 4046 11526 4050
rect 11704 4046 11734 4050
rect 11496 3978 11526 4012
rect 11704 3978 11734 4012
rect 11496 3910 11526 3944
rect 11704 3910 11734 3944
rect 11496 3842 11526 3876
rect 11704 3842 11734 3876
rect 11496 3774 11526 3808
rect 11704 3774 11734 3808
rect 11496 3706 11526 3740
rect 11704 3706 11734 3740
rect 11496 3638 11526 3672
rect 11704 3638 11734 3672
rect 11496 3570 11526 3604
rect 11704 3570 11734 3604
rect 11496 3502 11526 3536
rect 11704 3502 11734 3536
rect 11496 3434 11526 3468
rect 11704 3434 11734 3468
rect 11496 3366 11526 3400
rect 11704 3366 11734 3400
rect 11496 3298 11526 3332
rect 11704 3298 11734 3332
rect 11496 3230 11526 3264
rect 11704 3230 11734 3264
rect 11496 3162 11526 3196
rect 11704 3162 11734 3196
rect 11496 3080 11526 3128
rect 11560 3080 11670 3092
rect 11704 3080 11734 3128
rect 11496 3037 11734 3080
rect 11496 3003 11526 3037
rect 11560 3003 11598 3037
rect 11632 3003 11670 3037
rect 11704 3003 11734 3037
rect 11496 2954 11734 3003
rect 11496 2920 11526 2954
rect 11560 2935 11598 2954
rect 11632 2935 11670 2954
rect 11560 2920 11565 2935
rect 11632 2920 11633 2935
rect 11496 2901 11565 2920
rect 11599 2901 11633 2920
rect 11667 2920 11670 2935
rect 11704 2920 11734 2954
rect 11667 2901 11734 2920
rect 11496 2871 11734 2901
rect 11496 2837 11526 2871
rect 11560 2855 11598 2871
rect 11632 2855 11670 2871
rect 11560 2837 11565 2855
rect 11632 2837 11633 2855
rect 11496 2821 11565 2837
rect 11599 2821 11633 2837
rect 11667 2837 11670 2855
rect 11704 2837 11734 2871
rect 11667 2821 11734 2837
rect 11496 2787 11734 2821
rect 11496 2753 11526 2787
rect 11560 2775 11598 2787
rect 11632 2775 11670 2787
rect 11560 2753 11565 2775
rect 11632 2753 11633 2775
rect 11496 2741 11565 2753
rect 11599 2741 11633 2753
rect 11667 2753 11670 2775
rect 11704 2753 11734 2787
rect 11667 2741 11734 2753
rect 11496 2703 11734 2741
rect 11496 2669 11526 2703
rect 11560 2695 11598 2703
rect 11632 2695 11670 2703
rect 11560 2669 11565 2695
rect 11632 2669 11633 2695
rect 11496 2661 11565 2669
rect 11599 2661 11633 2669
rect 11667 2669 11670 2695
rect 11704 2669 11734 2703
rect 11667 2661 11734 2669
rect 11496 2619 11734 2661
rect 11496 2585 11526 2619
rect 11560 2614 11598 2619
rect 11632 2614 11670 2619
rect 11560 2585 11565 2614
rect 11632 2585 11633 2614
rect 11496 2580 11565 2585
rect 11599 2580 11633 2585
rect 11667 2585 11670 2614
rect 11704 2585 11734 2619
rect 11667 2580 11734 2585
rect 11496 2535 11734 2580
rect 11496 2501 11526 2535
rect 11560 2501 11598 2535
rect 11632 2501 11670 2535
rect 11704 2501 11734 2535
rect 11496 2461 11734 2501
rect 11496 2449 11598 2461
rect 11632 2449 11734 2461
rect 11496 2445 11526 2449
rect 11704 2445 11734 2449
rect 11496 2377 11526 2411
rect 11704 2377 11734 2411
rect 11496 2309 11526 2343
rect 11704 2309 11734 2343
rect 11496 2241 11526 2275
rect 11704 2241 11734 2275
rect 11496 2173 11526 2207
rect 11704 2173 11734 2207
rect 11496 2105 11526 2139
rect 11704 2105 11734 2139
rect 11496 2037 11526 2071
rect 11704 2037 11734 2071
rect 11496 1969 11526 2003
rect 11704 1969 11734 2003
rect 11496 1901 11526 1935
rect 11704 1901 11734 1935
rect 11496 1833 11526 1867
rect 11704 1833 11734 1867
rect 11496 1765 11526 1799
rect 11704 1765 11734 1799
rect 11496 1697 11526 1731
rect 11704 1697 11734 1731
rect 11496 1629 11526 1663
rect 11704 1629 11734 1663
rect 11496 1561 11526 1595
rect 11704 1561 11734 1595
rect 11496 1479 11526 1527
rect 11560 1479 11670 1491
rect 11704 1479 11734 1527
rect 11496 1464 11734 1479
rect 11836 3010 11956 4106
rect 12266 4388 12273 4494
rect 12379 4388 12386 4494
rect 12266 4214 12386 4388
rect 12266 4180 12309 4214
rect 12343 4180 12386 4214
rect 12266 4140 12386 4180
rect 12266 4106 12309 4140
rect 12343 4106 12386 4140
rect 11836 2976 11879 3010
rect 11913 2976 11956 3010
rect 11836 2932 11956 2976
rect 11836 2898 11879 2932
rect 11913 2898 11956 2932
rect 11836 2854 11956 2898
rect 11836 2820 11879 2854
rect 11913 2820 11956 2854
rect 11836 2776 11956 2820
rect 11836 2742 11879 2776
rect 11913 2742 11956 2776
rect 11836 2697 11956 2742
rect 11836 2663 11879 2697
rect 11913 2663 11956 2697
rect 11836 2618 11956 2663
rect 11836 2584 11879 2618
rect 11913 2584 11956 2618
rect 11836 2539 11956 2584
rect 11836 2505 11879 2539
rect 11913 2505 11956 2539
rect 11274 1375 11317 1409
rect 11351 1375 11394 1409
rect 11274 1335 11394 1375
rect 11274 1301 11317 1335
rect 11351 1301 11394 1335
rect 11274 1285 11394 1301
rect 11836 1409 11956 2505
rect 12021 4028 12022 4062
rect 12056 4046 12094 4062
rect 12056 4028 12058 4046
rect 12021 4012 12058 4028
rect 12092 4028 12094 4046
rect 12128 4046 12166 4062
rect 12128 4028 12130 4046
rect 12092 4012 12130 4028
rect 12164 4028 12166 4046
rect 12200 4028 12201 4062
rect 12164 4012 12201 4028
rect 12021 3988 12201 4012
rect 12021 3954 12022 3988
rect 12056 3978 12094 3988
rect 12056 3954 12058 3978
rect 12021 3944 12058 3954
rect 12092 3954 12094 3978
rect 12128 3978 12166 3988
rect 12128 3954 12130 3978
rect 12092 3944 12130 3954
rect 12164 3954 12166 3978
rect 12200 3954 12201 3988
rect 12164 3944 12201 3954
rect 12021 3914 12201 3944
rect 12021 3880 12022 3914
rect 12056 3910 12094 3914
rect 12056 3880 12058 3910
rect 12021 3876 12058 3880
rect 12092 3880 12094 3910
rect 12128 3910 12166 3914
rect 12128 3880 12130 3910
rect 12092 3876 12130 3880
rect 12164 3880 12166 3910
rect 12200 3880 12201 3914
rect 12164 3876 12201 3880
rect 12021 3842 12201 3876
rect 12021 3840 12058 3842
rect 12021 3806 12022 3840
rect 12056 3808 12058 3840
rect 12092 3840 12130 3842
rect 12092 3808 12094 3840
rect 12056 3806 12094 3808
rect 12128 3808 12130 3840
rect 12164 3840 12201 3842
rect 12164 3808 12166 3840
rect 12128 3806 12166 3808
rect 12200 3806 12201 3840
rect 12021 3774 12201 3806
rect 12021 3766 12058 3774
rect 12021 3732 12022 3766
rect 12056 3740 12058 3766
rect 12092 3766 12130 3774
rect 12092 3740 12094 3766
rect 12056 3732 12094 3740
rect 12128 3740 12130 3766
rect 12164 3766 12201 3774
rect 12164 3740 12166 3766
rect 12128 3732 12166 3740
rect 12200 3732 12201 3766
rect 12021 3706 12201 3732
rect 12021 3692 12058 3706
rect 12021 3658 12022 3692
rect 12056 3672 12058 3692
rect 12092 3692 12130 3706
rect 12092 3672 12094 3692
rect 12056 3658 12094 3672
rect 12128 3672 12130 3692
rect 12164 3692 12201 3706
rect 12164 3672 12166 3692
rect 12128 3658 12166 3672
rect 12200 3658 12201 3692
rect 12021 3638 12201 3658
rect 12021 3618 12058 3638
rect 12021 3584 12022 3618
rect 12056 3604 12058 3618
rect 12092 3618 12130 3638
rect 12092 3604 12094 3618
rect 12056 3584 12094 3604
rect 12128 3604 12130 3618
rect 12164 3618 12201 3638
rect 12164 3604 12166 3618
rect 12128 3584 12166 3604
rect 12200 3584 12201 3618
rect 12021 3570 12201 3584
rect 12021 3544 12058 3570
rect 12021 3510 12022 3544
rect 12056 3536 12058 3544
rect 12092 3544 12130 3570
rect 12092 3536 12094 3544
rect 12056 3510 12094 3536
rect 12128 3536 12130 3544
rect 12164 3544 12201 3570
rect 12164 3536 12166 3544
rect 12128 3510 12166 3536
rect 12200 3510 12201 3544
rect 12021 3502 12201 3510
rect 12021 3470 12058 3502
rect 12021 3436 12022 3470
rect 12056 3468 12058 3470
rect 12092 3470 12130 3502
rect 12092 3468 12094 3470
rect 12056 3436 12094 3468
rect 12128 3468 12130 3470
rect 12164 3470 12201 3502
rect 12164 3468 12166 3470
rect 12128 3436 12166 3468
rect 12200 3436 12201 3470
rect 12021 3434 12201 3436
rect 12021 3400 12058 3434
rect 12092 3400 12130 3434
rect 12164 3400 12201 3434
rect 12021 3396 12201 3400
rect 12021 3362 12022 3396
rect 12056 3366 12094 3396
rect 12056 3362 12058 3366
rect 12021 3332 12058 3362
rect 12092 3362 12094 3366
rect 12128 3366 12166 3396
rect 12128 3362 12130 3366
rect 12092 3332 12130 3362
rect 12164 3362 12166 3366
rect 12200 3362 12201 3396
rect 12164 3332 12201 3362
rect 12021 3322 12201 3332
rect 12021 3288 12022 3322
rect 12056 3298 12094 3322
rect 12056 3288 12058 3298
rect 12021 3264 12058 3288
rect 12092 3288 12094 3298
rect 12128 3298 12166 3322
rect 12128 3288 12130 3298
rect 12092 3264 12130 3288
rect 12164 3288 12166 3298
rect 12200 3288 12201 3322
rect 12164 3264 12201 3288
rect 12021 3248 12201 3264
rect 12021 3214 12022 3248
rect 12056 3230 12094 3248
rect 12056 3214 12058 3230
rect 12021 3196 12058 3214
rect 12092 3214 12094 3230
rect 12128 3230 12166 3248
rect 12128 3214 12130 3230
rect 12092 3196 12130 3214
rect 12164 3214 12166 3230
rect 12200 3214 12201 3248
rect 12164 3196 12201 3214
rect 12021 3174 12201 3196
rect 12021 3140 12022 3174
rect 12056 3162 12094 3174
rect 12056 3140 12058 3162
rect 12021 3128 12058 3140
rect 12092 3140 12094 3162
rect 12128 3162 12166 3174
rect 12128 3140 12130 3162
rect 12092 3128 12130 3140
rect 12164 3140 12166 3162
rect 12200 3140 12201 3174
rect 12164 3128 12201 3140
rect 12021 3100 12201 3128
rect 12021 3066 12022 3100
rect 12056 3066 12094 3100
rect 12128 3066 12166 3100
rect 12200 3066 12201 3100
rect 12021 3026 12201 3066
rect 12021 2992 12022 3026
rect 12056 2992 12094 3026
rect 12128 2992 12166 3026
rect 12200 2992 12201 3026
rect 12021 2952 12201 2992
rect 12021 2918 12022 2952
rect 12056 2918 12094 2952
rect 12128 2918 12166 2952
rect 12200 2918 12201 2952
rect 12021 2878 12201 2918
rect 12021 2844 12022 2878
rect 12056 2844 12094 2878
rect 12128 2844 12166 2878
rect 12200 2844 12201 2878
rect 12021 2804 12201 2844
rect 12021 2770 12022 2804
rect 12056 2770 12094 2804
rect 12128 2770 12166 2804
rect 12200 2770 12201 2804
rect 12021 2730 12201 2770
rect 12021 2696 12022 2730
rect 12056 2696 12094 2730
rect 12128 2696 12166 2730
rect 12200 2696 12201 2730
rect 12021 2656 12201 2696
rect 12021 2622 12022 2656
rect 12056 2622 12094 2656
rect 12128 2622 12166 2656
rect 12200 2622 12201 2656
rect 12021 2582 12201 2622
rect 12021 2548 12022 2582
rect 12056 2548 12094 2582
rect 12128 2548 12166 2582
rect 12200 2548 12201 2582
rect 12021 2508 12201 2548
rect 12021 2474 12022 2508
rect 12056 2474 12094 2508
rect 12128 2474 12166 2508
rect 12200 2474 12201 2508
rect 12021 2445 12201 2474
rect 12021 2434 12058 2445
rect 12021 2400 12022 2434
rect 12056 2411 12058 2434
rect 12092 2434 12130 2445
rect 12092 2411 12094 2434
rect 12056 2400 12094 2411
rect 12128 2411 12130 2434
rect 12164 2434 12201 2445
rect 12164 2411 12166 2434
rect 12128 2400 12166 2411
rect 12200 2400 12201 2434
rect 12021 2377 12201 2400
rect 12021 2360 12058 2377
rect 12021 2326 12022 2360
rect 12056 2343 12058 2360
rect 12092 2360 12130 2377
rect 12092 2343 12094 2360
rect 12056 2326 12094 2343
rect 12128 2343 12130 2360
rect 12164 2360 12201 2377
rect 12164 2343 12166 2360
rect 12128 2326 12166 2343
rect 12200 2326 12201 2360
rect 12021 2309 12201 2326
rect 12021 2286 12058 2309
rect 12021 2252 12022 2286
rect 12056 2275 12058 2286
rect 12092 2286 12130 2309
rect 12092 2275 12094 2286
rect 12056 2252 12094 2275
rect 12128 2275 12130 2286
rect 12164 2286 12201 2309
rect 12164 2275 12166 2286
rect 12128 2252 12166 2275
rect 12200 2252 12201 2286
rect 12021 2241 12201 2252
rect 12021 2212 12058 2241
rect 12021 2178 12022 2212
rect 12056 2207 12058 2212
rect 12092 2212 12130 2241
rect 12092 2207 12094 2212
rect 12056 2178 12094 2207
rect 12128 2207 12130 2212
rect 12164 2212 12201 2241
rect 12164 2207 12166 2212
rect 12128 2178 12166 2207
rect 12200 2178 12201 2212
rect 12021 2173 12201 2178
rect 12021 2139 12058 2173
rect 12092 2139 12130 2173
rect 12164 2139 12201 2173
rect 12021 2138 12201 2139
rect 12021 2104 12022 2138
rect 12056 2105 12094 2138
rect 12056 2104 12058 2105
rect 12021 2071 12058 2104
rect 12092 2104 12094 2105
rect 12128 2105 12166 2138
rect 12128 2104 12130 2105
rect 12092 2071 12130 2104
rect 12164 2104 12166 2105
rect 12200 2104 12201 2138
rect 12164 2071 12201 2104
rect 12021 2064 12201 2071
rect 12021 2030 12022 2064
rect 12056 2037 12094 2064
rect 12056 2030 12058 2037
rect 12021 2003 12058 2030
rect 12092 2030 12094 2037
rect 12128 2037 12166 2064
rect 12128 2030 12130 2037
rect 12092 2003 12130 2030
rect 12164 2030 12166 2037
rect 12200 2030 12201 2064
rect 12164 2003 12201 2030
rect 12021 1990 12201 2003
rect 12021 1956 12022 1990
rect 12056 1969 12094 1990
rect 12056 1956 12058 1969
rect 12021 1935 12058 1956
rect 12092 1956 12094 1969
rect 12128 1969 12166 1990
rect 12128 1956 12130 1969
rect 12092 1935 12130 1956
rect 12164 1956 12166 1969
rect 12200 1956 12201 1990
rect 12164 1935 12201 1956
rect 12021 1916 12201 1935
rect 12021 1882 12022 1916
rect 12056 1901 12094 1916
rect 12056 1882 12058 1901
rect 12021 1867 12058 1882
rect 12092 1882 12094 1901
rect 12128 1901 12166 1916
rect 12128 1882 12130 1901
rect 12092 1867 12130 1882
rect 12164 1882 12166 1901
rect 12200 1882 12201 1916
rect 12164 1867 12201 1882
rect 12021 1842 12201 1867
rect 12021 1808 12022 1842
rect 12056 1833 12094 1842
rect 12056 1808 12058 1833
rect 12021 1799 12058 1808
rect 12092 1808 12094 1833
rect 12128 1833 12166 1842
rect 12128 1808 12130 1833
rect 12092 1799 12130 1808
rect 12164 1808 12166 1833
rect 12200 1808 12201 1842
rect 12164 1799 12201 1808
rect 12021 1768 12201 1799
rect 12021 1734 12022 1768
rect 12056 1765 12094 1768
rect 12056 1734 12058 1765
rect 12021 1731 12058 1734
rect 12092 1734 12094 1765
rect 12128 1765 12166 1768
rect 12128 1734 12130 1765
rect 12092 1731 12130 1734
rect 12164 1734 12166 1765
rect 12200 1734 12201 1768
rect 12164 1731 12201 1734
rect 12021 1697 12201 1731
rect 12021 1694 12058 1697
rect 12021 1660 12022 1694
rect 12056 1663 12058 1694
rect 12092 1694 12130 1697
rect 12092 1663 12094 1694
rect 12056 1660 12094 1663
rect 12128 1663 12130 1694
rect 12164 1694 12201 1697
rect 12164 1663 12166 1694
rect 12128 1660 12166 1663
rect 12200 1660 12201 1694
rect 12021 1629 12201 1660
rect 12021 1620 12058 1629
rect 12021 1586 12022 1620
rect 12056 1595 12058 1620
rect 12092 1620 12130 1629
rect 12092 1595 12094 1620
rect 12056 1586 12094 1595
rect 12128 1595 12130 1620
rect 12164 1620 12201 1629
rect 12164 1595 12166 1620
rect 12128 1586 12166 1595
rect 12200 1586 12201 1620
rect 12021 1561 12201 1586
rect 12021 1545 12058 1561
rect 12021 1511 12022 1545
rect 12056 1527 12058 1545
rect 12092 1545 12130 1561
rect 12092 1527 12094 1545
rect 12056 1511 12094 1527
rect 12128 1527 12130 1545
rect 12164 1545 12201 1561
rect 12164 1527 12166 1545
rect 12128 1511 12166 1527
rect 12200 1511 12201 1545
rect 12266 3010 12386 4106
rect 12828 4388 12835 4494
rect 12941 4388 12948 4494
rect 12828 4214 12948 4388
rect 12828 4180 12871 4214
rect 12905 4180 12948 4214
rect 12828 4140 12948 4180
rect 12828 4106 12871 4140
rect 12905 4106 12948 4140
rect 12266 2976 12309 3010
rect 12343 2976 12386 3010
rect 12266 2932 12386 2976
rect 12266 2898 12309 2932
rect 12343 2898 12386 2932
rect 12266 2854 12386 2898
rect 12266 2820 12309 2854
rect 12343 2820 12386 2854
rect 12266 2776 12386 2820
rect 12266 2742 12309 2776
rect 12343 2742 12386 2776
rect 12266 2697 12386 2742
rect 12266 2663 12309 2697
rect 12343 2663 12386 2697
rect 12266 2618 12386 2663
rect 12266 2584 12309 2618
rect 12343 2584 12386 2618
rect 12266 2539 12386 2584
rect 12266 2505 12309 2539
rect 12343 2505 12386 2539
rect 12058 1491 12164 1511
rect 11836 1375 11879 1409
rect 11913 1375 11956 1409
rect 11836 1335 11956 1375
rect 11836 1301 11879 1335
rect 11913 1301 11956 1335
rect 11836 1285 11956 1301
rect 12266 1409 12386 2505
rect 12488 4050 12590 4062
rect 12624 4050 12726 4062
rect 12488 4046 12518 4050
rect 12696 4046 12726 4050
rect 12488 3978 12518 4012
rect 12696 3978 12726 4012
rect 12488 3910 12518 3944
rect 12696 3910 12726 3944
rect 12488 3842 12518 3876
rect 12696 3842 12726 3876
rect 12488 3774 12518 3808
rect 12696 3774 12726 3808
rect 12488 3706 12518 3740
rect 12696 3706 12726 3740
rect 12488 3638 12518 3672
rect 12696 3638 12726 3672
rect 12488 3570 12518 3604
rect 12696 3570 12726 3604
rect 12488 3502 12518 3536
rect 12696 3502 12726 3536
rect 12488 3434 12518 3468
rect 12696 3434 12726 3468
rect 12488 3366 12518 3400
rect 12696 3366 12726 3400
rect 12488 3298 12518 3332
rect 12696 3298 12726 3332
rect 12488 3230 12518 3264
rect 12696 3230 12726 3264
rect 12488 3162 12518 3196
rect 12696 3162 12726 3196
rect 12488 3080 12518 3128
rect 12552 3080 12662 3092
rect 12696 3080 12726 3128
rect 12488 3038 12726 3080
rect 12488 3004 12518 3038
rect 12552 3004 12590 3038
rect 12624 3004 12662 3038
rect 12696 3004 12726 3038
rect 12488 2955 12726 3004
rect 12488 2921 12518 2955
rect 12552 2935 12590 2955
rect 12624 2935 12662 2955
rect 12552 2921 12557 2935
rect 12624 2921 12625 2935
rect 12488 2901 12557 2921
rect 12591 2901 12625 2921
rect 12659 2921 12662 2935
rect 12696 2921 12726 2955
rect 12659 2901 12726 2921
rect 12488 2871 12726 2901
rect 12488 2837 12518 2871
rect 12552 2855 12590 2871
rect 12624 2855 12662 2871
rect 12552 2837 12557 2855
rect 12624 2837 12625 2855
rect 12488 2821 12557 2837
rect 12591 2821 12625 2837
rect 12659 2837 12662 2855
rect 12696 2837 12726 2871
rect 12659 2821 12726 2837
rect 12488 2787 12726 2821
rect 12488 2753 12518 2787
rect 12552 2775 12590 2787
rect 12624 2775 12662 2787
rect 12552 2753 12557 2775
rect 12624 2753 12625 2775
rect 12488 2741 12557 2753
rect 12591 2741 12625 2753
rect 12659 2753 12662 2775
rect 12696 2753 12726 2787
rect 12659 2741 12726 2753
rect 12488 2703 12726 2741
rect 12488 2669 12518 2703
rect 12552 2695 12590 2703
rect 12624 2695 12662 2703
rect 12552 2669 12557 2695
rect 12624 2669 12625 2695
rect 12488 2661 12557 2669
rect 12591 2661 12625 2669
rect 12659 2669 12662 2695
rect 12696 2669 12726 2703
rect 12659 2661 12726 2669
rect 12488 2619 12726 2661
rect 12488 2585 12518 2619
rect 12552 2614 12590 2619
rect 12624 2614 12662 2619
rect 12552 2585 12557 2614
rect 12624 2585 12625 2614
rect 12488 2580 12557 2585
rect 12591 2580 12625 2585
rect 12659 2585 12662 2614
rect 12696 2585 12726 2619
rect 12659 2580 12726 2585
rect 12488 2535 12726 2580
rect 12488 2501 12518 2535
rect 12552 2501 12590 2535
rect 12624 2501 12662 2535
rect 12696 2501 12726 2535
rect 12488 2461 12726 2501
rect 12488 2449 12590 2461
rect 12624 2449 12726 2461
rect 12488 2445 12518 2449
rect 12696 2445 12726 2449
rect 12488 2377 12518 2411
rect 12696 2377 12726 2411
rect 12488 2309 12518 2343
rect 12696 2309 12726 2343
rect 12488 2241 12518 2275
rect 12696 2241 12726 2275
rect 12488 2173 12518 2207
rect 12696 2173 12726 2207
rect 12488 2105 12518 2139
rect 12696 2105 12726 2139
rect 12488 2037 12518 2071
rect 12696 2037 12726 2071
rect 12488 1969 12518 2003
rect 12696 1969 12726 2003
rect 12488 1901 12518 1935
rect 12696 1901 12726 1935
rect 12488 1833 12518 1867
rect 12696 1833 12726 1867
rect 12488 1765 12518 1799
rect 12696 1765 12726 1799
rect 12488 1697 12518 1731
rect 12696 1697 12726 1731
rect 12488 1629 12518 1663
rect 12696 1629 12726 1663
rect 12488 1561 12518 1595
rect 12696 1561 12726 1595
rect 12488 1479 12518 1527
rect 12552 1479 12662 1491
rect 12696 1479 12726 1527
rect 12488 1464 12726 1479
rect 12828 3010 12948 4106
rect 13258 4388 13265 4494
rect 13371 4388 13378 4494
rect 13258 4214 13378 4388
rect 13258 4180 13301 4214
rect 13335 4180 13378 4214
rect 13258 4140 13378 4180
rect 13258 4106 13301 4140
rect 13335 4106 13378 4140
rect 12828 2976 12871 3010
rect 12905 2976 12948 3010
rect 12828 2932 12948 2976
rect 12828 2898 12871 2932
rect 12905 2898 12948 2932
rect 12828 2854 12948 2898
rect 12828 2820 12871 2854
rect 12905 2820 12948 2854
rect 12828 2776 12948 2820
rect 12828 2742 12871 2776
rect 12905 2742 12948 2776
rect 12828 2697 12948 2742
rect 12828 2663 12871 2697
rect 12905 2663 12948 2697
rect 12828 2618 12948 2663
rect 12828 2584 12871 2618
rect 12905 2584 12948 2618
rect 12828 2539 12948 2584
rect 12828 2505 12871 2539
rect 12905 2505 12948 2539
rect 12266 1375 12309 1409
rect 12343 1375 12386 1409
rect 12266 1335 12386 1375
rect 12266 1301 12309 1335
rect 12343 1301 12386 1335
rect 12266 1285 12386 1301
rect 12828 1409 12948 2505
rect 13013 4028 13014 4062
rect 13048 4046 13086 4062
rect 13048 4028 13050 4046
rect 13013 4012 13050 4028
rect 13084 4028 13086 4046
rect 13120 4046 13158 4062
rect 13120 4028 13122 4046
rect 13084 4012 13122 4028
rect 13156 4028 13158 4046
rect 13192 4028 13193 4062
rect 13156 4012 13193 4028
rect 13013 3988 13193 4012
rect 13013 3954 13014 3988
rect 13048 3978 13086 3988
rect 13048 3954 13050 3978
rect 13013 3944 13050 3954
rect 13084 3954 13086 3978
rect 13120 3978 13158 3988
rect 13120 3954 13122 3978
rect 13084 3944 13122 3954
rect 13156 3954 13158 3978
rect 13192 3954 13193 3988
rect 13156 3944 13193 3954
rect 13013 3914 13193 3944
rect 13013 3880 13014 3914
rect 13048 3910 13086 3914
rect 13048 3880 13050 3910
rect 13013 3876 13050 3880
rect 13084 3880 13086 3910
rect 13120 3910 13158 3914
rect 13120 3880 13122 3910
rect 13084 3876 13122 3880
rect 13156 3880 13158 3910
rect 13192 3880 13193 3914
rect 13156 3876 13193 3880
rect 13013 3842 13193 3876
rect 13013 3840 13050 3842
rect 13013 3806 13014 3840
rect 13048 3808 13050 3840
rect 13084 3840 13122 3842
rect 13084 3808 13086 3840
rect 13048 3806 13086 3808
rect 13120 3808 13122 3840
rect 13156 3840 13193 3842
rect 13156 3808 13158 3840
rect 13120 3806 13158 3808
rect 13192 3806 13193 3840
rect 13013 3774 13193 3806
rect 13013 3766 13050 3774
rect 13013 3732 13014 3766
rect 13048 3740 13050 3766
rect 13084 3766 13122 3774
rect 13084 3740 13086 3766
rect 13048 3732 13086 3740
rect 13120 3740 13122 3766
rect 13156 3766 13193 3774
rect 13156 3740 13158 3766
rect 13120 3732 13158 3740
rect 13192 3732 13193 3766
rect 13013 3706 13193 3732
rect 13013 3692 13050 3706
rect 13013 3658 13014 3692
rect 13048 3672 13050 3692
rect 13084 3692 13122 3706
rect 13084 3672 13086 3692
rect 13048 3658 13086 3672
rect 13120 3672 13122 3692
rect 13156 3692 13193 3706
rect 13156 3672 13158 3692
rect 13120 3658 13158 3672
rect 13192 3658 13193 3692
rect 13013 3638 13193 3658
rect 13013 3618 13050 3638
rect 13013 3584 13014 3618
rect 13048 3604 13050 3618
rect 13084 3618 13122 3638
rect 13084 3604 13086 3618
rect 13048 3584 13086 3604
rect 13120 3604 13122 3618
rect 13156 3618 13193 3638
rect 13156 3604 13158 3618
rect 13120 3584 13158 3604
rect 13192 3584 13193 3618
rect 13013 3570 13193 3584
rect 13013 3544 13050 3570
rect 13013 3510 13014 3544
rect 13048 3536 13050 3544
rect 13084 3544 13122 3570
rect 13084 3536 13086 3544
rect 13048 3510 13086 3536
rect 13120 3536 13122 3544
rect 13156 3544 13193 3570
rect 13156 3536 13158 3544
rect 13120 3510 13158 3536
rect 13192 3510 13193 3544
rect 13013 3502 13193 3510
rect 13013 3470 13050 3502
rect 13013 3436 13014 3470
rect 13048 3468 13050 3470
rect 13084 3470 13122 3502
rect 13084 3468 13086 3470
rect 13048 3436 13086 3468
rect 13120 3468 13122 3470
rect 13156 3470 13193 3502
rect 13156 3468 13158 3470
rect 13120 3436 13158 3468
rect 13192 3436 13193 3470
rect 13013 3434 13193 3436
rect 13013 3400 13050 3434
rect 13084 3400 13122 3434
rect 13156 3400 13193 3434
rect 13013 3396 13193 3400
rect 13013 3362 13014 3396
rect 13048 3366 13086 3396
rect 13048 3362 13050 3366
rect 13013 3332 13050 3362
rect 13084 3362 13086 3366
rect 13120 3366 13158 3396
rect 13120 3362 13122 3366
rect 13084 3332 13122 3362
rect 13156 3362 13158 3366
rect 13192 3362 13193 3396
rect 13156 3332 13193 3362
rect 13013 3322 13193 3332
rect 13013 3288 13014 3322
rect 13048 3298 13086 3322
rect 13048 3288 13050 3298
rect 13013 3264 13050 3288
rect 13084 3288 13086 3298
rect 13120 3298 13158 3322
rect 13120 3288 13122 3298
rect 13084 3264 13122 3288
rect 13156 3288 13158 3298
rect 13192 3288 13193 3322
rect 13156 3264 13193 3288
rect 13013 3248 13193 3264
rect 13013 3214 13014 3248
rect 13048 3230 13086 3248
rect 13048 3214 13050 3230
rect 13013 3196 13050 3214
rect 13084 3214 13086 3230
rect 13120 3230 13158 3248
rect 13120 3214 13122 3230
rect 13084 3196 13122 3214
rect 13156 3214 13158 3230
rect 13192 3214 13193 3248
rect 13156 3196 13193 3214
rect 13013 3174 13193 3196
rect 13013 3140 13014 3174
rect 13048 3162 13086 3174
rect 13048 3140 13050 3162
rect 13013 3128 13050 3140
rect 13084 3140 13086 3162
rect 13120 3162 13158 3174
rect 13120 3140 13122 3162
rect 13084 3128 13122 3140
rect 13156 3140 13158 3162
rect 13192 3140 13193 3174
rect 13156 3128 13193 3140
rect 13013 3100 13193 3128
rect 13013 3066 13014 3100
rect 13048 3066 13086 3100
rect 13120 3066 13158 3100
rect 13192 3066 13193 3100
rect 13013 3026 13193 3066
rect 13013 2992 13014 3026
rect 13048 2992 13086 3026
rect 13120 2992 13158 3026
rect 13192 2992 13193 3026
rect 13013 2952 13193 2992
rect 13013 2918 13014 2952
rect 13048 2918 13086 2952
rect 13120 2918 13158 2952
rect 13192 2918 13193 2952
rect 13013 2878 13193 2918
rect 13013 2844 13014 2878
rect 13048 2844 13086 2878
rect 13120 2844 13158 2878
rect 13192 2844 13193 2878
rect 13013 2804 13193 2844
rect 13013 2770 13014 2804
rect 13048 2770 13086 2804
rect 13120 2770 13158 2804
rect 13192 2770 13193 2804
rect 13013 2730 13193 2770
rect 13013 2696 13014 2730
rect 13048 2696 13086 2730
rect 13120 2696 13158 2730
rect 13192 2696 13193 2730
rect 13013 2656 13193 2696
rect 13013 2622 13014 2656
rect 13048 2622 13086 2656
rect 13120 2622 13158 2656
rect 13192 2622 13193 2656
rect 13013 2582 13193 2622
rect 13013 2548 13014 2582
rect 13048 2548 13086 2582
rect 13120 2548 13158 2582
rect 13192 2548 13193 2582
rect 13013 2508 13193 2548
rect 13013 2474 13014 2508
rect 13048 2474 13086 2508
rect 13120 2474 13158 2508
rect 13192 2474 13193 2508
rect 13013 2445 13193 2474
rect 13013 2434 13050 2445
rect 13013 2400 13014 2434
rect 13048 2411 13050 2434
rect 13084 2434 13122 2445
rect 13084 2411 13086 2434
rect 13048 2400 13086 2411
rect 13120 2411 13122 2434
rect 13156 2434 13193 2445
rect 13156 2411 13158 2434
rect 13120 2400 13158 2411
rect 13192 2400 13193 2434
rect 13013 2377 13193 2400
rect 13013 2360 13050 2377
rect 13013 2326 13014 2360
rect 13048 2343 13050 2360
rect 13084 2360 13122 2377
rect 13084 2343 13086 2360
rect 13048 2326 13086 2343
rect 13120 2343 13122 2360
rect 13156 2360 13193 2377
rect 13156 2343 13158 2360
rect 13120 2326 13158 2343
rect 13192 2326 13193 2360
rect 13013 2309 13193 2326
rect 13013 2286 13050 2309
rect 13013 2252 13014 2286
rect 13048 2275 13050 2286
rect 13084 2286 13122 2309
rect 13084 2275 13086 2286
rect 13048 2252 13086 2275
rect 13120 2275 13122 2286
rect 13156 2286 13193 2309
rect 13156 2275 13158 2286
rect 13120 2252 13158 2275
rect 13192 2252 13193 2286
rect 13013 2241 13193 2252
rect 13013 2212 13050 2241
rect 13013 2178 13014 2212
rect 13048 2207 13050 2212
rect 13084 2212 13122 2241
rect 13084 2207 13086 2212
rect 13048 2178 13086 2207
rect 13120 2207 13122 2212
rect 13156 2212 13193 2241
rect 13156 2207 13158 2212
rect 13120 2178 13158 2207
rect 13192 2178 13193 2212
rect 13013 2173 13193 2178
rect 13013 2139 13050 2173
rect 13084 2139 13122 2173
rect 13156 2139 13193 2173
rect 13013 2138 13193 2139
rect 13013 2104 13014 2138
rect 13048 2105 13086 2138
rect 13048 2104 13050 2105
rect 13013 2071 13050 2104
rect 13084 2104 13086 2105
rect 13120 2105 13158 2138
rect 13120 2104 13122 2105
rect 13084 2071 13122 2104
rect 13156 2104 13158 2105
rect 13192 2104 13193 2138
rect 13156 2071 13193 2104
rect 13013 2064 13193 2071
rect 13013 2030 13014 2064
rect 13048 2037 13086 2064
rect 13048 2030 13050 2037
rect 13013 2003 13050 2030
rect 13084 2030 13086 2037
rect 13120 2037 13158 2064
rect 13120 2030 13122 2037
rect 13084 2003 13122 2030
rect 13156 2030 13158 2037
rect 13192 2030 13193 2064
rect 13156 2003 13193 2030
rect 13013 1990 13193 2003
rect 13013 1956 13014 1990
rect 13048 1969 13086 1990
rect 13048 1956 13050 1969
rect 13013 1935 13050 1956
rect 13084 1956 13086 1969
rect 13120 1969 13158 1990
rect 13120 1956 13122 1969
rect 13084 1935 13122 1956
rect 13156 1956 13158 1969
rect 13192 1956 13193 1990
rect 13156 1935 13193 1956
rect 13013 1916 13193 1935
rect 13013 1882 13014 1916
rect 13048 1901 13086 1916
rect 13048 1882 13050 1901
rect 13013 1867 13050 1882
rect 13084 1882 13086 1901
rect 13120 1901 13158 1916
rect 13120 1882 13122 1901
rect 13084 1867 13122 1882
rect 13156 1882 13158 1901
rect 13192 1882 13193 1916
rect 13156 1867 13193 1882
rect 13013 1842 13193 1867
rect 13013 1808 13014 1842
rect 13048 1833 13086 1842
rect 13048 1808 13050 1833
rect 13013 1799 13050 1808
rect 13084 1808 13086 1833
rect 13120 1833 13158 1842
rect 13120 1808 13122 1833
rect 13084 1799 13122 1808
rect 13156 1808 13158 1833
rect 13192 1808 13193 1842
rect 13156 1799 13193 1808
rect 13013 1768 13193 1799
rect 13013 1734 13014 1768
rect 13048 1765 13086 1768
rect 13048 1734 13050 1765
rect 13013 1731 13050 1734
rect 13084 1734 13086 1765
rect 13120 1765 13158 1768
rect 13120 1734 13122 1765
rect 13084 1731 13122 1734
rect 13156 1734 13158 1765
rect 13192 1734 13193 1768
rect 13156 1731 13193 1734
rect 13013 1697 13193 1731
rect 13013 1694 13050 1697
rect 13013 1660 13014 1694
rect 13048 1663 13050 1694
rect 13084 1694 13122 1697
rect 13084 1663 13086 1694
rect 13048 1660 13086 1663
rect 13120 1663 13122 1694
rect 13156 1694 13193 1697
rect 13156 1663 13158 1694
rect 13120 1660 13158 1663
rect 13192 1660 13193 1694
rect 13013 1629 13193 1660
rect 13013 1620 13050 1629
rect 13013 1586 13014 1620
rect 13048 1595 13050 1620
rect 13084 1620 13122 1629
rect 13084 1595 13086 1620
rect 13048 1586 13086 1595
rect 13120 1595 13122 1620
rect 13156 1620 13193 1629
rect 13156 1595 13158 1620
rect 13120 1586 13158 1595
rect 13192 1586 13193 1620
rect 13013 1561 13193 1586
rect 13013 1545 13050 1561
rect 13013 1511 13014 1545
rect 13048 1527 13050 1545
rect 13084 1545 13122 1561
rect 13084 1527 13086 1545
rect 13048 1511 13086 1527
rect 13120 1527 13122 1545
rect 13156 1545 13193 1561
rect 13156 1527 13158 1545
rect 13120 1511 13158 1527
rect 13192 1511 13193 1545
rect 13258 3010 13378 4106
rect 13820 4388 13827 4494
rect 13933 4388 13940 4494
rect 13820 4214 13940 4388
rect 13820 4180 13863 4214
rect 13897 4180 13940 4214
rect 13820 4140 13940 4180
rect 13820 4106 13863 4140
rect 13897 4106 13940 4140
rect 13258 2976 13301 3010
rect 13335 2976 13378 3010
rect 13258 2932 13378 2976
rect 13258 2898 13301 2932
rect 13335 2898 13378 2932
rect 13258 2854 13378 2898
rect 13258 2820 13301 2854
rect 13335 2820 13378 2854
rect 13258 2776 13378 2820
rect 13258 2742 13301 2776
rect 13335 2742 13378 2776
rect 13258 2697 13378 2742
rect 13258 2663 13301 2697
rect 13335 2663 13378 2697
rect 13258 2618 13378 2663
rect 13258 2584 13301 2618
rect 13335 2584 13378 2618
rect 13258 2539 13378 2584
rect 13258 2505 13301 2539
rect 13335 2505 13378 2539
rect 12828 1375 12871 1409
rect 12905 1375 12948 1409
rect 12828 1335 12948 1375
rect 12828 1301 12871 1335
rect 12905 1301 12948 1335
rect 12828 1285 12948 1301
rect 13258 1409 13378 2505
rect 13480 4050 13582 4062
rect 13616 4050 13718 4062
rect 13480 4046 13510 4050
rect 13688 4046 13718 4050
rect 13480 3978 13510 4012
rect 13688 3978 13718 4012
rect 13480 3910 13510 3944
rect 13688 3910 13718 3944
rect 13480 3842 13510 3876
rect 13688 3842 13718 3876
rect 13480 3774 13510 3808
rect 13688 3774 13718 3808
rect 13480 3706 13510 3740
rect 13688 3706 13718 3740
rect 13480 3638 13510 3672
rect 13688 3638 13718 3672
rect 13480 3570 13510 3604
rect 13688 3570 13718 3604
rect 13480 3502 13510 3536
rect 13688 3502 13718 3536
rect 13480 3434 13510 3468
rect 13688 3434 13718 3468
rect 13480 3366 13510 3400
rect 13688 3366 13718 3400
rect 13480 3298 13510 3332
rect 13688 3298 13718 3332
rect 13480 3230 13510 3264
rect 13688 3230 13718 3264
rect 13480 3162 13510 3196
rect 13688 3162 13718 3196
rect 13480 3080 13510 3128
rect 13544 3080 13654 3092
rect 13688 3080 13718 3128
rect 13480 3040 13718 3080
rect 13480 2574 13510 3040
rect 13688 2574 13718 3040
rect 13480 2535 13718 2574
rect 13480 2501 13510 2535
rect 13544 2501 13582 2535
rect 13616 2501 13654 2535
rect 13688 2501 13718 2535
rect 13480 2461 13718 2501
rect 13480 2449 13582 2461
rect 13616 2449 13718 2461
rect 13480 2445 13510 2449
rect 13688 2445 13718 2449
rect 13480 2377 13510 2411
rect 13688 2377 13718 2411
rect 13480 2309 13510 2343
rect 13688 2309 13718 2343
rect 13480 2241 13510 2275
rect 13688 2241 13718 2275
rect 13480 2173 13510 2207
rect 13688 2173 13718 2207
rect 13480 2105 13510 2139
rect 13688 2105 13718 2139
rect 13480 2037 13510 2071
rect 13688 2037 13718 2071
rect 13480 1969 13510 2003
rect 13688 1969 13718 2003
rect 13480 1901 13510 1935
rect 13688 1901 13718 1935
rect 13480 1833 13510 1867
rect 13688 1833 13718 1867
rect 13480 1765 13510 1799
rect 13688 1765 13718 1799
rect 13480 1697 13510 1731
rect 13688 1697 13718 1731
rect 13480 1629 13510 1663
rect 13688 1629 13718 1663
rect 13480 1561 13510 1595
rect 13688 1561 13718 1595
rect 13480 1479 13510 1527
rect 13544 1479 13654 1491
rect 13688 1479 13718 1527
rect 13480 1464 13718 1479
rect 13820 3010 13940 4106
rect 14178 4388 14185 4494
rect 14291 4388 14298 4494
rect 14178 4214 14298 4388
rect 14178 4180 14221 4214
rect 14255 4180 14298 4214
rect 14178 4140 14298 4180
rect 14178 4106 14221 4140
rect 14255 4106 14298 4140
rect 13820 2976 13863 3010
rect 13897 2976 13940 3010
rect 13820 2932 13940 2976
rect 13820 2898 13863 2932
rect 13897 2898 13940 2932
rect 13820 2854 13940 2898
rect 13820 2820 13863 2854
rect 13897 2820 13940 2854
rect 13820 2776 13940 2820
rect 13820 2742 13863 2776
rect 13897 2742 13940 2776
rect 13820 2697 13940 2742
rect 13820 2663 13863 2697
rect 13897 2663 13940 2697
rect 13820 2618 13940 2663
rect 13820 2584 13863 2618
rect 13897 2584 13940 2618
rect 13820 2539 13940 2584
rect 13820 2505 13863 2539
rect 13897 2505 13940 2539
rect 13258 1375 13301 1409
rect 13335 1375 13378 1409
rect 13258 1335 13378 1375
rect 13258 1301 13301 1335
rect 13335 1301 13378 1335
rect 13258 1285 13378 1301
rect 13820 1409 13940 2505
rect 14006 2693 14112 2732
rect 14040 2659 14078 2693
rect 14006 2620 14112 2659
rect 14040 2586 14078 2620
rect 14006 2547 14112 2586
rect 14040 2513 14078 2547
rect 14006 2474 14112 2513
rect 14040 2445 14078 2474
rect 14040 2440 14042 2445
rect 14006 2411 14042 2440
rect 14076 2440 14078 2445
rect 14076 2411 14112 2440
rect 14006 2401 14112 2411
rect 14040 2377 14078 2401
rect 14040 2367 14042 2377
rect 14006 2343 14042 2367
rect 14076 2367 14078 2377
rect 14076 2343 14112 2367
rect 14006 2328 14112 2343
rect 14040 2309 14078 2328
rect 14040 2294 14042 2309
rect 14006 2275 14042 2294
rect 14076 2294 14078 2309
rect 14076 2275 14112 2294
rect 14006 2255 14112 2275
rect 14040 2241 14078 2255
rect 14040 2221 14042 2241
rect 14006 2207 14042 2221
rect 14076 2221 14078 2241
rect 14076 2207 14112 2221
rect 14006 2182 14112 2207
rect 14040 2173 14078 2182
rect 14040 2148 14042 2173
rect 14006 2139 14042 2148
rect 14076 2148 14078 2173
rect 14076 2139 14112 2148
rect 14006 2109 14112 2139
rect 14040 2105 14078 2109
rect 14040 2075 14042 2105
rect 14006 2071 14042 2075
rect 14076 2075 14078 2105
rect 14076 2071 14112 2075
rect 14006 2037 14112 2071
rect 14006 2036 14042 2037
rect 14040 2003 14042 2036
rect 14076 2036 14112 2037
rect 14076 2003 14078 2036
rect 14040 2002 14078 2003
rect 14006 1969 14112 2002
rect 14006 1963 14042 1969
rect 14040 1935 14042 1963
rect 14076 1963 14112 1969
rect 14076 1935 14078 1963
rect 14040 1929 14078 1935
rect 14006 1901 14112 1929
rect 14006 1890 14042 1901
rect 14040 1867 14042 1890
rect 14076 1890 14112 1901
rect 14076 1867 14078 1890
rect 14040 1856 14078 1867
rect 14006 1833 14112 1856
rect 14006 1817 14042 1833
rect 14040 1799 14042 1817
rect 14076 1817 14112 1833
rect 14076 1799 14078 1817
rect 14040 1783 14078 1799
rect 14006 1765 14112 1783
rect 14006 1744 14042 1765
rect 14040 1731 14042 1744
rect 14076 1744 14112 1765
rect 14076 1731 14078 1744
rect 14040 1710 14078 1731
rect 14006 1697 14112 1710
rect 14006 1671 14042 1697
rect 14040 1663 14042 1671
rect 14076 1671 14112 1697
rect 14076 1663 14078 1671
rect 14040 1637 14078 1663
rect 14006 1629 14112 1637
rect 14006 1598 14042 1629
rect 14040 1595 14042 1598
rect 14076 1598 14112 1629
rect 14076 1595 14078 1598
rect 14040 1564 14078 1595
rect 14006 1561 14112 1564
rect 14006 1527 14042 1561
rect 14076 1527 14112 1561
rect 14006 1525 14112 1527
rect 14040 1491 14078 1525
rect 14178 3010 14298 4106
rect 14400 4490 14510 4506
rect 14544 4504 14565 4524
rect 14616 4518 14633 4524
rect 14544 4490 14582 4504
rect 14616 4490 14667 4518
rect 14400 4482 14667 4490
rect 14400 4448 14431 4482
rect 14465 4479 14667 4482
rect 14465 4470 14633 4479
rect 14465 4448 14497 4470
rect 14531 4468 14633 4470
rect 14531 4451 14565 4468
rect 14599 4451 14633 4468
rect 14400 4436 14497 4448
rect 14400 4417 14510 4436
rect 14544 4434 14565 4451
rect 14616 4445 14633 4451
rect 14544 4417 14582 4434
rect 14616 4417 14667 4445
rect 14400 4409 14667 4417
rect 14400 4375 14431 4409
rect 14465 4406 14667 4409
rect 14465 4399 14633 4406
rect 14465 4375 14497 4399
rect 14531 4398 14633 4399
rect 14531 4378 14565 4398
rect 14599 4378 14633 4398
rect 14400 4365 14497 4375
rect 14400 4344 14510 4365
rect 14544 4364 14565 4378
rect 14616 4372 14633 4378
rect 14544 4344 14582 4364
rect 14616 4344 14667 4372
rect 14400 4336 14667 4344
rect 14400 4302 14431 4336
rect 14465 4333 14667 4336
rect 14465 4328 14633 4333
rect 14465 4302 14497 4328
rect 14531 4305 14565 4328
rect 14599 4305 14633 4328
rect 14400 4294 14497 4302
rect 14544 4294 14565 4305
rect 14616 4299 14633 4305
rect 14400 4271 14510 4294
rect 14544 4271 14582 4294
rect 14616 4271 14667 4299
rect 14400 4263 14667 4271
rect 14400 4229 14431 4263
rect 14465 4260 14667 4263
rect 14465 4257 14633 4260
rect 14465 4229 14497 4257
rect 14531 4232 14565 4257
rect 14599 4232 14633 4257
rect 14400 4223 14497 4229
rect 14544 4223 14565 4232
rect 14616 4226 14633 4232
rect 14400 4198 14510 4223
rect 14544 4198 14582 4223
rect 14616 4198 14667 4226
rect 14400 4190 14667 4198
rect 14400 4156 14431 4190
rect 14465 4186 14667 4190
rect 14465 4156 14497 4186
rect 14531 4159 14565 4186
rect 14599 4159 14633 4186
rect 14400 4152 14497 4156
rect 14544 4152 14565 4159
rect 14616 4152 14633 4159
rect 14400 4125 14510 4152
rect 14544 4125 14582 4152
rect 14616 4125 14667 4152
rect 14400 4117 14667 4125
rect 14400 4083 14431 4117
rect 14465 4115 14667 4117
rect 14465 4086 14565 4115
rect 14599 4086 14633 4115
rect 14465 4083 14510 4086
rect 14400 4062 14510 4083
rect 14386 4052 14510 4062
rect 14544 4081 14565 4086
rect 14616 4081 14633 4086
rect 14544 4052 14582 4081
rect 14616 4052 14667 4081
rect 14386 4046 14667 4052
rect 14420 4044 14667 4046
rect 14420 4012 14431 4044
rect 14465 4041 14667 4044
rect 14465 4034 14565 4041
rect 14386 4010 14431 4012
rect 14488 4013 14565 4034
rect 14599 4013 14633 4041
rect 14386 4000 14454 4010
rect 14488 4000 14510 4013
rect 14386 3979 14510 4000
rect 14544 4007 14565 4013
rect 14616 4007 14633 4013
rect 14544 3979 14582 4007
rect 14616 3979 14667 4007
rect 14386 3978 14667 3979
rect 14420 3971 14667 3978
rect 14420 3944 14431 3971
rect 14465 3970 14667 3971
rect 14465 3966 14565 3970
rect 14386 3937 14431 3944
rect 14488 3940 14565 3966
rect 14599 3940 14633 3970
rect 14386 3932 14454 3937
rect 14488 3932 14510 3940
rect 14386 3910 14510 3932
rect 14420 3906 14510 3910
rect 14544 3936 14565 3940
rect 14616 3936 14633 3940
rect 14544 3906 14582 3936
rect 14616 3906 14667 3936
rect 14420 3898 14667 3906
rect 14420 3876 14431 3898
rect 14386 3864 14431 3876
rect 14488 3896 14667 3898
rect 14488 3867 14565 3896
rect 14599 3867 14633 3896
rect 14488 3864 14510 3867
rect 14386 3842 14510 3864
rect 14420 3833 14510 3842
rect 14544 3862 14565 3867
rect 14616 3862 14633 3867
rect 14544 3833 14582 3862
rect 14616 3833 14667 3862
rect 14420 3830 14667 3833
rect 14420 3825 14454 3830
rect 14488 3825 14667 3830
rect 14420 3808 14431 3825
rect 14386 3791 14431 3808
rect 14488 3796 14565 3825
rect 14465 3794 14565 3796
rect 14599 3794 14633 3825
rect 14465 3791 14510 3794
rect 14386 3774 14510 3791
rect 14420 3762 14510 3774
rect 14420 3752 14454 3762
rect 14488 3760 14510 3762
rect 14544 3791 14565 3794
rect 14616 3791 14633 3794
rect 14544 3760 14582 3791
rect 14616 3760 14667 3791
rect 14420 3740 14431 3752
rect 14386 3718 14431 3740
rect 14488 3751 14667 3760
rect 14488 3728 14565 3751
rect 14465 3721 14565 3728
rect 14599 3721 14633 3751
rect 14465 3718 14510 3721
rect 14386 3706 14510 3718
rect 14420 3694 14510 3706
rect 14420 3679 14454 3694
rect 14488 3687 14510 3694
rect 14544 3717 14565 3721
rect 14616 3717 14633 3721
rect 14544 3687 14582 3717
rect 14616 3687 14667 3717
rect 14488 3680 14667 3687
rect 14420 3672 14431 3679
rect 14386 3645 14431 3672
rect 14488 3660 14565 3680
rect 14465 3648 14565 3660
rect 14599 3648 14633 3680
rect 14465 3645 14510 3648
rect 14386 3638 14510 3645
rect 14420 3626 14510 3638
rect 14420 3606 14454 3626
rect 14488 3614 14510 3626
rect 14544 3646 14565 3648
rect 14616 3646 14633 3648
rect 14544 3614 14582 3646
rect 14616 3614 14667 3646
rect 14488 3606 14667 3614
rect 14420 3604 14431 3606
rect 14386 3572 14431 3604
rect 14488 3592 14565 3606
rect 14465 3575 14565 3592
rect 14599 3575 14633 3606
rect 14465 3572 14510 3575
rect 14386 3570 14510 3572
rect 14420 3558 14510 3570
rect 14420 3536 14454 3558
rect 14386 3533 14454 3536
rect 14488 3541 14510 3558
rect 14544 3572 14565 3575
rect 14616 3572 14633 3575
rect 14544 3541 14582 3572
rect 14616 3541 14667 3572
rect 14488 3535 14667 3541
rect 14386 3502 14431 3533
rect 14488 3524 14565 3535
rect 14420 3499 14431 3502
rect 14465 3502 14565 3524
rect 14599 3502 14633 3535
rect 14465 3499 14510 3502
rect 14420 3490 14510 3499
rect 14420 3468 14454 3490
rect 14386 3460 14454 3468
rect 14488 3468 14510 3490
rect 14544 3501 14565 3502
rect 14616 3501 14633 3502
rect 14544 3468 14582 3501
rect 14616 3468 14667 3501
rect 14488 3461 14667 3468
rect 14386 3434 14431 3460
rect 14488 3456 14565 3461
rect 14420 3426 14431 3434
rect 14465 3429 14565 3456
rect 14599 3429 14633 3461
rect 14465 3426 14510 3429
rect 14420 3422 14510 3426
rect 14420 3400 14454 3422
rect 14386 3388 14454 3400
rect 14488 3395 14510 3422
rect 14544 3427 14565 3429
rect 14616 3427 14633 3429
rect 14544 3395 14582 3427
rect 14616 3395 14667 3427
rect 14488 3390 14667 3395
rect 14488 3388 14565 3390
rect 14386 3387 14565 3388
rect 14386 3366 14431 3387
rect 14420 3353 14431 3366
rect 14465 3356 14565 3387
rect 14599 3356 14633 3390
rect 14465 3354 14510 3356
rect 14420 3332 14454 3353
rect 14386 3320 14454 3332
rect 14488 3322 14510 3354
rect 14544 3322 14582 3356
rect 14616 3322 14667 3356
rect 14488 3320 14667 3322
rect 14386 3316 14667 3320
rect 14386 3314 14565 3316
rect 14386 3298 14431 3314
rect 14420 3280 14431 3298
rect 14465 3286 14565 3314
rect 14488 3283 14565 3286
rect 14599 3283 14633 3316
rect 14420 3264 14454 3280
rect 14386 3252 14454 3264
rect 14488 3252 14510 3283
rect 14386 3249 14510 3252
rect 14544 3282 14565 3283
rect 14616 3282 14633 3283
rect 14544 3249 14582 3282
rect 14616 3249 14667 3282
rect 14386 3245 14667 3249
rect 14386 3241 14565 3245
rect 14386 3230 14431 3241
rect 14420 3207 14431 3230
rect 14465 3218 14565 3241
rect 14488 3211 14565 3218
rect 14599 3211 14633 3245
rect 14488 3210 14667 3211
rect 14420 3196 14454 3207
rect 14386 3184 14454 3196
rect 14488 3184 14510 3210
rect 14386 3176 14510 3184
rect 14544 3176 14582 3210
rect 14616 3176 14667 3210
rect 14386 3168 14667 3176
rect 14386 3162 14431 3168
rect 14420 3134 14431 3162
rect 14465 3151 14667 3168
rect 14465 3150 14565 3151
rect 14488 3137 14565 3150
rect 14599 3137 14633 3151
rect 14420 3128 14454 3134
rect 14386 3116 14454 3128
rect 14488 3116 14510 3137
rect 14386 3103 14510 3116
rect 14544 3117 14565 3137
rect 14616 3117 14633 3137
rect 14544 3103 14582 3117
rect 14616 3103 14667 3117
rect 14386 3100 14667 3103
rect 14178 2976 14221 3010
rect 14255 2976 14298 3010
rect 14178 2932 14298 2976
rect 14178 2898 14221 2932
rect 14255 2898 14298 2932
rect 14178 2854 14298 2898
rect 14178 2820 14221 2854
rect 14255 2820 14298 2854
rect 14178 2776 14298 2820
rect 14178 2742 14221 2776
rect 14255 2742 14298 2776
rect 14178 2697 14298 2742
rect 14178 2663 14221 2697
rect 14255 2663 14298 2697
rect 14178 2618 14298 2663
rect 14178 2584 14221 2618
rect 14255 2584 14298 2618
rect 14178 2539 14298 2584
rect 14178 2505 14221 2539
rect 14255 2505 14298 2539
rect 13820 1375 13863 1409
rect 13897 1375 13940 1409
rect 13820 1335 13940 1375
rect 13820 1301 13863 1335
rect 13897 1301 13940 1335
rect 13820 1285 13940 1301
rect 14178 1409 14298 2505
rect 14400 3095 14667 3100
rect 14400 3061 14431 3095
rect 14465 3066 14667 3095
rect 14465 3064 14565 3066
rect 14599 3064 14633 3066
rect 14465 3061 14510 3064
rect 14400 3030 14510 3061
rect 14544 3032 14565 3064
rect 14616 3032 14633 3064
rect 14544 3030 14582 3032
rect 14616 3030 14667 3032
rect 14400 3022 14667 3030
rect 14400 2988 14431 3022
rect 14465 2991 14667 3022
rect 14465 2988 14510 2991
rect 14400 2972 14510 2988
rect 14544 2972 14582 2991
rect 14616 2972 14667 2991
rect 14400 2949 14497 2972
rect 14400 2915 14431 2949
rect 14465 2915 14497 2949
rect 14400 2876 14497 2915
rect 14400 2842 14431 2876
rect 14465 2842 14497 2876
rect 14400 2803 14497 2842
rect 14400 2769 14431 2803
rect 14465 2769 14497 2803
rect 14400 2730 14497 2769
rect 14400 2696 14431 2730
rect 14465 2696 14497 2730
rect 14400 2657 14497 2696
rect 14400 2623 14431 2657
rect 14465 2623 14497 2657
rect 14400 2584 14497 2623
rect 14400 2550 14431 2584
rect 14465 2550 14497 2584
rect 14400 2530 14497 2550
rect 14400 2519 14510 2530
rect 14544 2519 14582 2530
rect 14616 2519 14667 2530
rect 14400 2511 14667 2519
rect 14400 2477 14431 2511
rect 14465 2485 14667 2511
rect 14465 2480 14565 2485
rect 14599 2480 14633 2485
rect 14465 2477 14510 2480
rect 14400 2461 14510 2477
rect 14386 2446 14510 2461
rect 14544 2451 14565 2480
rect 14616 2451 14633 2480
rect 14544 2446 14582 2451
rect 14616 2446 14667 2451
rect 14386 2445 14667 2446
rect 14420 2438 14667 2445
rect 14420 2411 14431 2438
rect 14465 2433 14667 2438
rect 14386 2404 14431 2411
rect 14488 2407 14667 2433
rect 14386 2399 14454 2404
rect 14488 2399 14510 2407
rect 14386 2377 14510 2399
rect 14420 2373 14510 2377
rect 14544 2403 14582 2407
rect 14616 2403 14667 2407
rect 14544 2373 14565 2403
rect 14616 2373 14633 2403
rect 14420 2369 14565 2373
rect 14599 2369 14633 2373
rect 14420 2365 14667 2369
rect 14420 2343 14431 2365
rect 14386 2331 14431 2343
rect 14488 2334 14667 2365
rect 14488 2331 14510 2334
rect 14386 2309 14510 2331
rect 14420 2300 14510 2309
rect 14544 2327 14582 2334
rect 14616 2327 14667 2334
rect 14544 2300 14565 2327
rect 14616 2300 14633 2327
rect 14420 2297 14565 2300
rect 14420 2292 14454 2297
rect 14488 2293 14565 2297
rect 14599 2293 14633 2300
rect 14420 2275 14431 2292
rect 14386 2258 14431 2275
rect 14488 2263 14667 2293
rect 14465 2260 14667 2263
rect 14465 2258 14510 2260
rect 14386 2241 14510 2258
rect 14420 2229 14510 2241
rect 14420 2219 14454 2229
rect 14488 2226 14510 2229
rect 14544 2250 14582 2260
rect 14616 2250 14667 2260
rect 14544 2226 14565 2250
rect 14616 2226 14633 2250
rect 14420 2207 14431 2219
rect 14386 2185 14431 2207
rect 14488 2216 14565 2226
rect 14599 2216 14633 2226
rect 14488 2195 14667 2216
rect 14465 2186 14667 2195
rect 14465 2185 14510 2186
rect 14386 2173 14510 2185
rect 14420 2161 14510 2173
rect 14420 2146 14454 2161
rect 14488 2152 14510 2161
rect 14544 2156 14582 2186
rect 14616 2156 14667 2186
rect 14544 2152 14565 2156
rect 14616 2152 14633 2156
rect 14420 2139 14431 2146
rect 14386 2112 14431 2139
rect 14488 2127 14565 2152
rect 14465 2122 14565 2127
rect 14599 2122 14633 2152
rect 14465 2112 14667 2122
rect 14386 2105 14510 2112
rect 14420 2093 14510 2105
rect 14420 2073 14454 2093
rect 14488 2078 14510 2093
rect 14544 2085 14582 2112
rect 14616 2085 14667 2112
rect 14544 2078 14565 2085
rect 14616 2078 14633 2085
rect 14420 2071 14431 2073
rect 14386 2039 14431 2071
rect 14488 2059 14565 2078
rect 14465 2051 14565 2059
rect 14599 2051 14633 2078
rect 14465 2039 14667 2051
rect 14386 2038 14667 2039
rect 14386 2037 14510 2038
rect 14420 2025 14510 2037
rect 14420 2003 14454 2025
rect 14386 2000 14454 2003
rect 14488 2004 14510 2025
rect 14544 2011 14582 2038
rect 14616 2011 14667 2038
rect 14544 2004 14565 2011
rect 14616 2004 14633 2011
rect 14386 1969 14431 2000
rect 14488 1991 14565 2004
rect 14420 1966 14431 1969
rect 14465 1977 14565 1991
rect 14599 1977 14633 2004
rect 14465 1966 14667 1977
rect 14420 1964 14667 1966
rect 14420 1957 14510 1964
rect 14420 1935 14454 1957
rect 14386 1927 14454 1935
rect 14488 1930 14510 1957
rect 14544 1940 14582 1964
rect 14616 1940 14667 1964
rect 14544 1930 14565 1940
rect 14616 1930 14633 1940
rect 14386 1901 14431 1927
rect 14488 1923 14565 1930
rect 14420 1893 14431 1901
rect 14465 1906 14565 1923
rect 14599 1906 14633 1930
rect 14465 1893 14667 1906
rect 14420 1890 14667 1893
rect 14420 1889 14510 1890
rect 14420 1867 14454 1889
rect 14386 1855 14454 1867
rect 14488 1856 14510 1889
rect 14544 1866 14582 1890
rect 14616 1866 14667 1890
rect 14544 1856 14565 1866
rect 14616 1856 14633 1866
rect 14488 1855 14565 1856
rect 14386 1854 14565 1855
rect 14386 1833 14431 1854
rect 14420 1820 14431 1833
rect 14465 1832 14565 1854
rect 14599 1832 14633 1856
rect 14465 1821 14667 1832
rect 14420 1799 14454 1820
rect 14386 1787 14454 1799
rect 14488 1816 14667 1821
rect 14488 1787 14510 1816
rect 14386 1782 14510 1787
rect 14544 1795 14582 1816
rect 14616 1795 14667 1816
rect 14544 1782 14565 1795
rect 14616 1782 14633 1795
rect 14386 1781 14565 1782
rect 14386 1765 14431 1781
rect 14420 1747 14431 1765
rect 14465 1761 14565 1781
rect 14599 1761 14633 1782
rect 14465 1753 14667 1761
rect 14420 1731 14454 1747
rect 14386 1719 14454 1731
rect 14488 1742 14667 1753
rect 14488 1719 14510 1742
rect 14386 1708 14510 1719
rect 14544 1721 14582 1742
rect 14616 1721 14667 1742
rect 14544 1708 14565 1721
rect 14616 1708 14633 1721
rect 14386 1697 14431 1708
rect 14420 1674 14431 1697
rect 14465 1687 14565 1708
rect 14599 1687 14633 1708
rect 14465 1685 14667 1687
rect 14420 1663 14454 1674
rect 14386 1651 14454 1663
rect 14488 1668 14667 1685
rect 14488 1651 14510 1668
rect 14386 1635 14510 1651
rect 14386 1629 14431 1635
rect 14420 1601 14431 1629
rect 14465 1634 14510 1635
rect 14544 1650 14582 1668
rect 14616 1650 14667 1668
rect 14544 1634 14565 1650
rect 14616 1634 14633 1650
rect 14465 1617 14565 1634
rect 14488 1616 14565 1617
rect 14599 1616 14633 1634
rect 14420 1595 14454 1601
rect 14386 1583 14454 1595
rect 14488 1594 14667 1616
rect 14488 1583 14510 1594
rect 14386 1562 14510 1583
rect 14386 1561 14431 1562
rect 14420 1528 14431 1561
rect 14465 1560 14510 1562
rect 14544 1576 14582 1594
rect 14616 1576 14667 1594
rect 14544 1560 14565 1576
rect 14616 1560 14633 1576
rect 14465 1549 14565 1560
rect 14488 1542 14565 1549
rect 14599 1542 14633 1560
rect 14420 1527 14454 1528
rect 14386 1515 14454 1527
rect 14488 1520 14667 1542
rect 14488 1515 14510 1520
rect 14386 1499 14510 1515
rect 14178 1375 14221 1409
rect 14255 1375 14298 1409
rect 14178 1335 14298 1375
rect 14178 1301 14221 1335
rect 14255 1301 14298 1335
rect 14178 1285 14298 1301
rect 14400 1489 14510 1499
rect 14400 1455 14431 1489
rect 14465 1486 14510 1489
rect 14544 1505 14582 1520
rect 14616 1505 14667 1520
rect 14544 1486 14565 1505
rect 14616 1486 14633 1505
rect 14465 1471 14565 1486
rect 14599 1471 14633 1486
rect 14465 1455 14667 1471
rect 14400 1446 14667 1455
rect 14400 1416 14510 1446
rect 14400 1382 14431 1416
rect 14465 1412 14510 1416
rect 14544 1412 14582 1446
rect 14616 1412 14667 1446
rect 14465 1387 14667 1412
rect 14465 1382 14497 1387
rect 14400 1353 14497 1382
rect 14531 1372 14565 1387
rect 14599 1372 14633 1387
rect 14544 1353 14565 1372
rect 14616 1353 14633 1372
rect 14400 1342 14510 1353
rect 14400 1308 14431 1342
rect 14465 1338 14510 1342
rect 14544 1338 14582 1353
rect 14616 1338 14667 1353
rect 14465 1319 14667 1338
rect 14465 1311 14633 1319
rect 14465 1308 14565 1311
rect 555 1241 733 1268
rect 555 1221 587 1241
rect 621 1221 659 1241
rect 621 1207 623 1221
rect 589 1187 623 1207
rect 657 1207 659 1221
rect 693 1234 733 1241
rect 767 1234 822 1268
rect 693 1219 822 1234
rect 657 1187 691 1207
rect 555 1185 691 1187
rect 725 1194 822 1219
rect 725 1185 733 1194
rect 555 1160 733 1185
rect 767 1160 822 1194
rect 555 1150 822 1160
rect 555 1140 623 1150
rect 589 1116 623 1140
rect 657 1148 822 1150
rect 14400 1274 14497 1308
rect 14531 1298 14565 1308
rect 14599 1298 14633 1311
rect 14544 1277 14565 1298
rect 14616 1285 14633 1298
rect 14400 1268 14510 1274
rect 14400 1234 14431 1268
rect 14465 1264 14510 1268
rect 14544 1264 14582 1277
rect 14616 1264 14667 1285
rect 14465 1251 14667 1264
rect 14465 1234 14633 1251
rect 14400 1228 14565 1234
rect 14400 1194 14497 1228
rect 14531 1224 14565 1228
rect 14599 1224 14633 1234
rect 14544 1200 14565 1224
rect 14616 1217 14633 1224
rect 14400 1160 14431 1194
rect 14465 1190 14510 1194
rect 14544 1190 14582 1200
rect 14616 1190 14667 1217
rect 14465 1183 14667 1190
rect 14465 1160 14633 1183
rect 14400 1157 14633 1160
rect 14400 1148 14565 1157
rect 657 1116 691 1148
rect 589 1114 691 1116
rect 725 1114 760 1148
rect 794 1116 829 1148
rect 14531 1123 14565 1148
rect 14599 1149 14633 1157
rect 14599 1123 14667 1149
rect 589 1106 767 1114
rect 555 1082 767 1106
rect 801 1082 829 1116
rect 555 1080 829 1082
rect 555 1046 623 1080
rect 657 1046 692 1080
rect 726 1046 761 1080
rect 555 1012 761 1046
rect 555 978 589 1012
rect 623 978 658 1012
rect 692 978 727 1012
rect 14531 1115 14667 1123
rect 14531 1081 14633 1115
rect 14531 1080 14667 1081
rect 14599 1046 14667 1080
rect 14565 1012 14633 1046
rect 14565 978 14667 1012
rect 14990 4955 15003 4993
rect 14990 4883 15003 4921
rect 14990 4811 15003 4849
rect 14990 4739 15003 4777
rect 14990 4667 15003 4705
rect 14990 4595 15003 4633
rect 14990 4523 15003 4561
rect 14990 4451 15003 4489
rect 14990 4379 15003 4417
rect 14990 4307 15003 4345
rect 14990 4235 15003 4273
rect 14990 4163 15003 4201
rect 14990 4091 15003 4129
rect 14990 4019 15003 4057
rect 14990 3947 15003 3985
rect 14990 3875 15003 3913
rect 14990 3803 15003 3841
rect 14990 3731 15003 3769
rect 14990 3659 15003 3697
rect 14990 3587 15003 3625
rect 14990 3515 15003 3553
rect 14990 3443 15003 3481
rect 14990 3371 15003 3409
rect 14990 3299 15003 3337
rect 14990 3227 15003 3265
rect 14990 3155 15003 3193
rect 14990 3082 15003 3121
rect 14990 3009 15003 3048
rect 14990 2936 15003 2975
rect 14990 2863 15003 2902
rect 14990 2790 15003 2829
rect 14990 2717 15003 2756
rect 14990 2644 15003 2683
rect 14990 2571 15003 2610
rect 14990 2498 15003 2537
rect 14990 2425 15003 2464
rect 14990 2352 15003 2391
rect 14990 2279 15003 2318
rect 14990 2206 15003 2245
rect 14990 2133 15003 2172
rect 14990 2060 15003 2099
rect 14990 1987 15003 2026
rect 14990 1914 15003 1953
rect 14990 1841 15003 1880
rect 14990 1768 15003 1807
rect 14990 1695 15003 1734
rect 14990 1622 15003 1661
rect 14990 1549 15003 1588
rect 14990 1476 15003 1515
rect 14990 1403 15003 1442
rect 14990 1330 15003 1369
rect 14990 1257 15003 1296
rect 14990 1184 15003 1223
rect 14990 1111 15003 1150
rect 14990 1038 15003 1077
rect 402 872 403 910
rect 212 762 232 800
rect 402 800 403 838
rect 14990 965 15003 1004
rect 14990 892 15003 931
rect 14990 819 15003 858
rect 334 749 402 764
rect 212 696 232 728
rect 334 715 348 749
rect 382 729 402 749
rect 334 696 368 715
rect 212 695 368 696
rect 212 684 402 695
rect 246 664 402 684
rect 14990 746 15003 785
rect 14990 696 15003 712
rect 14820 673 15003 696
rect 14820 664 14969 673
rect 246 661 348 664
rect 212 627 232 650
rect 266 627 300 661
rect 334 630 348 661
rect 382 660 421 664
rect 455 660 494 664
rect 528 660 567 664
rect 601 660 640 664
rect 674 660 713 664
rect 747 660 786 664
rect 820 660 859 664
rect 893 660 932 664
rect 966 660 1005 664
rect 1039 660 1078 664
rect 1112 660 1151 664
rect 1185 660 1224 664
rect 1258 660 1297 664
rect 1331 660 1369 664
rect 1403 660 1441 664
rect 1475 660 1513 664
rect 1547 660 1585 664
rect 1619 660 1657 664
rect 1691 660 1729 664
rect 1763 660 1801 664
rect 1835 660 1873 664
rect 1907 660 1945 664
rect 1979 660 2017 664
rect 2051 660 2089 664
rect 2123 660 2161 664
rect 2195 660 2233 664
rect 2267 660 2305 664
rect 2339 660 2377 664
rect 2411 660 2449 664
rect 2483 660 2521 664
rect 2555 660 2593 664
rect 2627 660 2665 664
rect 2699 660 2737 664
rect 2771 660 2809 664
rect 2843 660 2881 664
rect 2915 660 2953 664
rect 2987 660 3025 664
rect 3059 660 3097 664
rect 3131 660 3169 664
rect 3203 660 3241 664
rect 3275 660 3313 664
rect 3347 660 3385 664
rect 3419 660 3457 664
rect 3491 660 3529 664
rect 3563 660 3601 664
rect 3635 660 3673 664
rect 3707 660 3745 664
rect 3779 660 3817 664
rect 3851 660 3889 664
rect 3923 660 3961 664
rect 3995 660 4033 664
rect 4067 660 4105 664
rect 4139 660 4177 664
rect 4211 660 4249 664
rect 4283 660 4321 664
rect 4355 660 4393 664
rect 4427 660 4465 664
rect 4499 660 4537 664
rect 4571 660 4609 664
rect 4643 660 4681 664
rect 4715 660 4753 664
rect 4787 660 4825 664
rect 4859 660 4897 664
rect 4931 660 4969 664
rect 5003 660 5041 664
rect 5075 660 5113 664
rect 5147 660 5185 664
rect 5219 660 5257 664
rect 5291 660 5329 664
rect 5363 660 5401 664
rect 5435 660 5473 664
rect 5507 660 5545 664
rect 5579 660 5617 664
rect 5651 660 5689 664
rect 5723 660 5761 664
rect 5795 660 5833 664
rect 5867 660 5905 664
rect 5939 660 5977 664
rect 6011 660 6049 664
rect 6083 660 6121 664
rect 6155 660 6193 664
rect 6227 660 6265 664
rect 6299 660 6337 664
rect 6371 660 6409 664
rect 6443 660 6481 664
rect 6515 660 6553 664
rect 6587 660 6625 664
rect 6659 660 6697 664
rect 6731 660 6769 664
rect 6803 660 6841 664
rect 6875 660 6913 664
rect 6947 660 6985 664
rect 7019 660 7057 664
rect 7091 660 7129 664
rect 7163 660 7201 664
rect 7235 660 7273 664
rect 7307 660 7345 664
rect 7379 660 7417 664
rect 7451 660 7489 664
rect 7523 660 7561 664
rect 7595 660 7633 664
rect 7667 660 7705 664
rect 7739 660 7777 664
rect 7811 660 7849 664
rect 7883 660 7921 664
rect 7955 660 7993 664
rect 8027 660 8065 664
rect 8099 660 8137 664
rect 8171 660 8209 664
rect 8243 660 8281 664
rect 8315 660 8353 664
rect 8387 660 8425 664
rect 8459 660 8497 664
rect 8531 660 8569 664
rect 8603 660 8641 664
rect 8675 660 8713 664
rect 8747 660 8785 664
rect 8819 660 8857 664
rect 8891 660 8929 664
rect 8963 660 9001 664
rect 9035 660 9073 664
rect 9107 660 9145 664
rect 9179 660 9217 664
rect 9251 660 9289 664
rect 9323 660 9361 664
rect 9395 660 9433 664
rect 9467 660 9505 664
rect 9539 660 9577 664
rect 9611 660 9649 664
rect 9683 660 9721 664
rect 9755 660 9793 664
rect 9827 660 9865 664
rect 9899 660 9937 664
rect 9971 660 10009 664
rect 10043 660 10081 664
rect 10115 660 10153 664
rect 10187 660 10225 664
rect 10259 660 10297 664
rect 10331 660 10369 664
rect 10403 660 10441 664
rect 10475 660 10513 664
rect 10547 660 10585 664
rect 10619 660 10657 664
rect 10691 660 10729 664
rect 10763 660 10801 664
rect 10835 660 10873 664
rect 10907 660 10945 664
rect 10979 660 11017 664
rect 11051 660 11089 664
rect 11123 660 11161 664
rect 11195 660 11233 664
rect 11267 660 11305 664
rect 11339 660 11377 664
rect 11411 660 11449 664
rect 11483 660 11521 664
rect 11555 660 11593 664
rect 11627 660 11665 664
rect 11699 660 11737 664
rect 11771 660 11809 664
rect 11843 660 11881 664
rect 11915 660 11953 664
rect 11987 660 12025 664
rect 12059 660 12097 664
rect 12131 660 12169 664
rect 12203 660 12241 664
rect 12275 660 12313 664
rect 12347 660 12385 664
rect 12419 660 12457 664
rect 12491 660 12529 664
rect 12563 660 12601 664
rect 12635 660 12673 664
rect 12707 660 12745 664
rect 12779 660 12817 664
rect 12851 660 12889 664
rect 12923 660 12961 664
rect 12995 660 13033 664
rect 13067 660 13105 664
rect 13139 660 13177 664
rect 13211 660 13249 664
rect 13283 660 13321 664
rect 13355 660 13393 664
rect 13427 660 13465 664
rect 12995 630 13017 660
rect 13067 630 13086 660
rect 13139 630 13155 660
rect 13211 630 13224 660
rect 13283 630 13293 660
rect 13355 630 13362 660
rect 13427 630 13431 660
rect 334 627 368 630
rect 212 606 368 627
rect 246 592 368 606
rect 12982 626 13017 630
rect 13051 626 13086 630
rect 13120 626 13155 630
rect 13189 626 13224 630
rect 13258 626 13293 630
rect 13327 626 13362 630
rect 13396 626 13431 630
rect 13499 660 13537 664
rect 13571 660 13609 664
rect 13643 660 13681 664
rect 13715 660 13753 664
rect 13787 660 13825 664
rect 13859 660 13897 664
rect 13931 660 13969 664
rect 14003 660 14041 664
rect 14075 660 14113 664
rect 14147 660 14185 664
rect 14219 660 14257 664
rect 14291 660 14329 664
rect 14363 660 14401 664
rect 14435 660 14473 664
rect 14507 660 14545 664
rect 14579 660 14617 664
rect 14651 660 14689 664
rect 14723 660 14761 664
rect 14795 660 14833 664
rect 14867 660 14969 664
rect 13499 630 13500 660
rect 13465 626 13500 630
rect 13534 630 13537 660
rect 13603 630 13609 660
rect 13672 630 13681 660
rect 13741 630 13753 660
rect 13810 630 13825 660
rect 13879 630 13897 660
rect 13948 630 13969 660
rect 14017 630 14041 660
rect 14086 630 14113 660
rect 14155 630 14185 660
rect 14224 630 14257 660
rect 13534 626 13569 630
rect 13603 626 13638 630
rect 13672 626 13707 630
rect 13741 626 13776 630
rect 13810 626 13845 630
rect 13879 626 13914 630
rect 13948 626 13983 630
rect 14017 626 14052 630
rect 14086 626 14121 630
rect 14155 626 14190 630
rect 14224 626 14259 630
rect 14293 626 14328 660
rect 14363 630 14397 660
rect 14435 630 14466 660
rect 14507 630 14535 660
rect 14579 630 14604 660
rect 14651 630 14673 660
rect 14723 630 14742 660
rect 14795 630 14811 660
rect 14867 630 14880 660
rect 14362 626 14397 630
rect 14431 626 14466 630
rect 14500 626 14535 630
rect 14569 626 14604 630
rect 14638 626 14673 630
rect 14707 626 14742 630
rect 14776 626 14811 630
rect 14845 626 14880 630
rect 14914 639 14969 660
rect 14914 626 15003 639
rect 12982 600 15003 626
rect 12982 592 14969 600
rect 212 558 232 572
rect 266 558 300 592
rect 212 528 300 558
rect 12982 558 13017 592
rect 13051 558 13086 592
rect 13120 558 13155 592
rect 13189 558 13224 592
rect 13258 558 13293 592
rect 13327 558 13362 592
rect 13396 558 13431 592
rect 13465 558 13500 592
rect 13534 558 13569 592
rect 13603 558 13638 592
rect 13672 558 13707 592
rect 13741 558 13776 592
rect 13810 558 13845 592
rect 13879 558 13914 592
rect 13948 558 13983 592
rect 14017 558 14052 592
rect 14086 558 14121 592
rect 14155 558 14190 592
rect 14224 558 14259 592
rect 14293 558 14328 592
rect 14362 558 14397 592
rect 14431 558 14466 592
rect 14500 558 14535 592
rect 14569 558 14604 592
rect 14638 558 14673 592
rect 14707 558 14742 592
rect 14776 558 14811 592
rect 14845 558 14880 592
rect 14914 566 14969 592
rect 14914 558 15003 566
rect 12982 528 15003 558
rect 212 494 284 528
rect 12987 524 13025 528
rect 13059 524 13097 528
rect 13131 524 13169 528
rect 13203 524 13241 528
rect 13275 524 13313 528
rect 13347 524 13385 528
rect 13419 524 13457 528
rect 13491 524 13529 528
rect 13563 524 13601 528
rect 13635 524 13673 528
rect 12987 494 13017 524
rect 13059 494 13086 524
rect 13131 494 13155 524
rect 13203 494 13224 524
rect 13275 494 13293 524
rect 13347 494 13362 524
rect 13419 494 13431 524
rect 13491 494 13500 524
rect 13563 494 13569 524
rect 13635 494 13638 524
rect 232 490 300 494
rect 12982 490 13017 494
rect 13051 490 13086 494
rect 13120 490 13155 494
rect 13189 490 13224 494
rect 13258 490 13293 494
rect 13327 490 13362 494
rect 13396 490 13431 494
rect 13465 490 13500 494
rect 13534 490 13569 494
rect 13603 490 13638 494
rect 13672 494 13673 524
rect 13707 524 13745 528
rect 13779 524 13817 528
rect 13851 524 13889 528
rect 13923 524 13961 528
rect 13995 524 14033 528
rect 14067 524 14105 528
rect 14139 524 14177 528
rect 14211 524 14249 528
rect 14283 524 14321 528
rect 14355 524 14393 528
rect 14427 524 14465 528
rect 14499 524 14537 528
rect 14571 524 14609 528
rect 14643 524 14681 528
rect 14715 524 14753 528
rect 14787 524 14825 528
rect 14859 524 14897 528
rect 13672 490 13707 494
rect 13741 494 13745 524
rect 13810 494 13817 524
rect 13879 494 13889 524
rect 13948 494 13961 524
rect 14017 494 14033 524
rect 14086 494 14105 524
rect 14155 494 14177 524
rect 14224 494 14249 524
rect 14293 494 14321 524
rect 14362 494 14393 524
rect 14431 494 14465 524
rect 13741 490 13776 494
rect 13810 490 13845 494
rect 13879 490 13914 494
rect 13948 490 13983 494
rect 14017 490 14052 494
rect 14086 490 14121 494
rect 14155 490 14190 494
rect 14224 490 14259 494
rect 14293 490 14328 494
rect 14362 490 14397 494
rect 14431 490 14466 494
rect 14500 490 14535 524
rect 14571 494 14604 524
rect 14643 494 14673 524
rect 14715 494 14742 524
rect 14787 494 14811 524
rect 14859 494 14880 524
rect 14931 494 15003 528
rect 14569 490 14604 494
rect 14638 490 14673 494
rect 14707 490 14742 494
rect 14776 490 14811 494
rect 14845 490 14880 494
rect 14914 490 14948 494
<< viali >>
rect 305 5425 339 5459
rect 377 5425 411 5459
rect 449 5425 483 5459
rect 521 5425 555 5459
rect 593 5425 627 5459
rect 665 5425 699 5459
rect 737 5425 771 5459
rect 809 5425 843 5459
rect 881 5425 915 5459
rect 953 5425 987 5459
rect 1025 5425 1059 5459
rect 1097 5425 1131 5459
rect 1169 5425 1203 5459
rect 1241 5425 1275 5459
rect 1313 5425 1347 5459
rect 1385 5425 1419 5459
rect 1457 5425 1491 5459
rect 1529 5425 1563 5459
rect 1601 5425 1635 5459
rect 1673 5425 1707 5459
rect 1745 5425 1779 5459
rect 1817 5425 1851 5459
rect 1889 5425 1923 5459
rect 1961 5425 1995 5459
rect 2033 5425 2067 5459
rect 2105 5425 2139 5459
rect 2177 5425 2211 5459
rect 2249 5425 2283 5459
rect 2321 5425 2355 5459
rect 2393 5425 2427 5459
rect 2465 5425 2499 5459
rect 2537 5425 2571 5459
rect 2609 5425 2643 5459
rect 2681 5425 2715 5459
rect 2753 5425 2787 5459
rect 2825 5425 2859 5459
rect 2897 5425 2931 5459
rect 2969 5425 3003 5459
rect 3041 5425 3075 5459
rect 3113 5425 3147 5459
rect 3185 5425 3219 5459
rect 3257 5425 3291 5459
rect 3329 5425 3363 5459
rect 3401 5425 3435 5459
rect 3473 5425 3507 5459
rect 3545 5425 3579 5459
rect 3617 5425 3651 5459
rect 3689 5425 3723 5459
rect 3761 5425 3795 5459
rect 3833 5425 3867 5459
rect 3905 5425 3939 5459
rect 3977 5425 4011 5459
rect 4049 5425 4083 5459
rect 4121 5425 4155 5459
rect 4193 5425 4227 5459
rect 4265 5425 4299 5459
rect 4337 5425 4371 5459
rect 4409 5425 4443 5459
rect 4481 5425 4515 5459
rect 4553 5425 4587 5459
rect 4625 5425 4659 5459
rect 4697 5425 4731 5459
rect 4769 5425 4803 5459
rect 4841 5425 4875 5459
rect 4913 5425 4947 5459
rect 4985 5425 5019 5459
rect 5057 5425 5091 5459
rect 5129 5425 5163 5459
rect 5201 5425 5235 5459
rect 5273 5425 5307 5459
rect 5345 5425 5379 5459
rect 5417 5425 5451 5459
rect 5489 5425 5523 5459
rect 5561 5425 5595 5459
rect 5633 5425 5667 5459
rect 5705 5425 5739 5459
rect 5777 5425 5811 5459
rect 5849 5425 5883 5459
rect 5921 5425 5955 5459
rect 5993 5425 6027 5459
rect 6065 5425 6099 5459
rect 6137 5425 6171 5459
rect 6209 5425 6243 5459
rect 6281 5425 6315 5459
rect 6353 5425 6387 5459
rect 6425 5425 6459 5459
rect 6497 5425 6531 5459
rect 6569 5425 6603 5459
rect 6641 5425 6675 5459
rect 6713 5425 6747 5459
rect 6785 5425 6819 5459
rect 6857 5425 6891 5459
rect 6929 5425 6963 5459
rect 7001 5425 7035 5459
rect 7073 5425 7107 5459
rect 7145 5425 7179 5459
rect 7217 5425 7251 5459
rect 7289 5425 7323 5459
rect 7361 5425 7395 5459
rect 7433 5425 7467 5459
rect 7505 5425 7539 5459
rect 7577 5425 7611 5459
rect 7649 5425 7683 5459
rect 7721 5425 7755 5459
rect 7793 5425 7827 5459
rect 7865 5425 7899 5459
rect 7937 5425 7971 5459
rect 8009 5425 8043 5459
rect 8081 5425 8115 5459
rect 8153 5425 8187 5459
rect 8225 5425 8259 5459
rect 8297 5425 8331 5459
rect 8369 5425 8403 5459
rect 8441 5425 8475 5459
rect 8513 5425 8547 5459
rect 8585 5425 8619 5459
rect 8657 5425 8691 5459
rect 8729 5425 8763 5459
rect 8801 5425 8835 5459
rect 8873 5425 8907 5459
rect 8945 5425 8979 5459
rect 9017 5425 9051 5459
rect 9089 5425 9123 5459
rect 9161 5425 9195 5459
rect 9233 5425 9267 5459
rect 9305 5425 9339 5459
rect 9377 5425 9411 5459
rect 9449 5425 9483 5459
rect 9521 5425 9555 5459
rect 9593 5425 9627 5459
rect 9665 5425 9699 5459
rect 9737 5425 9771 5459
rect 9809 5425 9843 5459
rect 9881 5425 9915 5459
rect 9953 5425 9987 5459
rect 10025 5425 10059 5459
rect 10097 5425 10131 5459
rect 10169 5425 10203 5459
rect 10241 5425 10275 5459
rect 10313 5425 10347 5459
rect 10385 5425 10419 5459
rect 10457 5425 10491 5459
rect 10529 5425 10563 5459
rect 10601 5425 10635 5459
rect 10673 5425 10707 5459
rect 10745 5425 10779 5459
rect 10817 5425 10851 5459
rect 10889 5425 10923 5459
rect 10961 5425 10995 5459
rect 11033 5425 11067 5459
rect 11105 5425 11139 5459
rect 11177 5425 11211 5459
rect 11249 5425 11283 5459
rect 11321 5425 11355 5459
rect 11393 5425 11427 5459
rect 11466 5425 11500 5459
rect 11539 5425 11573 5459
rect 11612 5425 11646 5459
rect 11685 5425 11719 5459
rect 11758 5425 11792 5459
rect 11831 5425 11865 5459
rect 11904 5425 11938 5459
rect 11977 5425 12011 5459
rect 12050 5425 12084 5459
rect 12123 5425 12157 5459
rect 12196 5425 12230 5459
rect 12269 5425 12303 5459
rect 12342 5425 12376 5459
rect 12415 5425 12449 5459
rect 12488 5425 12522 5459
rect 12561 5425 12595 5459
rect 12634 5425 12668 5459
rect 12707 5425 12741 5459
rect 12780 5425 12814 5459
rect 12853 5425 12887 5459
rect 12926 5425 12960 5459
rect 12999 5425 13033 5459
rect 13072 5425 13106 5459
rect 13145 5425 13179 5459
rect 13218 5425 13252 5459
rect 13291 5425 13325 5459
rect 13364 5425 13398 5459
rect 13437 5425 13471 5459
rect 13510 5425 13544 5459
rect 13583 5425 13617 5459
rect 13656 5425 13690 5459
rect 13729 5425 13763 5459
rect 13802 5425 13836 5459
rect 13875 5425 13909 5459
rect 13948 5425 13982 5459
rect 14021 5425 14055 5459
rect 14094 5425 14128 5459
rect 14167 5425 14201 5459
rect 14240 5425 14274 5459
rect 14313 5425 14347 5459
rect 14386 5425 14420 5459
rect 14459 5425 14493 5459
rect 14532 5425 14566 5459
rect 14605 5425 14639 5459
rect 14678 5425 14712 5459
rect 14751 5425 14785 5459
rect 14824 5425 14858 5459
rect 14897 5425 14931 5459
rect 233 5354 267 5387
rect 233 5353 267 5354
rect 233 5280 267 5314
rect 369 5320 403 5323
rect 441 5320 472 5323
rect 472 5320 475 5323
rect 513 5320 541 5323
rect 541 5320 547 5323
rect 585 5320 610 5323
rect 610 5320 619 5323
rect 657 5320 679 5323
rect 679 5320 691 5323
rect 729 5320 748 5323
rect 748 5320 763 5323
rect 801 5320 817 5323
rect 817 5320 835 5323
rect 873 5320 886 5323
rect 886 5320 907 5323
rect 945 5320 955 5323
rect 955 5320 979 5323
rect 1017 5320 1024 5323
rect 1024 5320 1051 5323
rect 1089 5320 1093 5323
rect 1093 5320 1123 5323
rect 1161 5320 1162 5323
rect 1162 5320 1195 5323
rect 1233 5320 1266 5323
rect 1266 5320 1267 5323
rect 1305 5320 1335 5323
rect 1335 5320 1339 5323
rect 1377 5320 1404 5323
rect 1404 5320 1411 5323
rect 1449 5320 1473 5323
rect 1473 5320 1483 5323
rect 1521 5320 1542 5323
rect 1542 5320 1555 5323
rect 1593 5320 1611 5323
rect 1611 5320 1627 5323
rect 1665 5320 1680 5323
rect 1680 5320 1699 5323
rect 1737 5320 1749 5323
rect 1749 5320 1771 5323
rect 1809 5320 1818 5323
rect 1818 5320 1843 5323
rect 1881 5320 1887 5323
rect 1887 5320 1915 5323
rect 1953 5320 1956 5323
rect 1956 5320 1987 5323
rect 2025 5320 2059 5323
rect 14969 5353 15003 5387
rect 2097 5320 2128 5323
rect 2128 5320 2131 5323
rect 2169 5320 2197 5323
rect 2197 5320 2203 5323
rect 2241 5320 2275 5323
rect 369 5289 403 5320
rect 441 5289 475 5320
rect 513 5289 547 5320
rect 585 5289 619 5320
rect 657 5289 691 5320
rect 729 5289 763 5320
rect 801 5289 835 5320
rect 873 5289 907 5320
rect 945 5289 979 5320
rect 1017 5289 1051 5320
rect 1089 5289 1123 5320
rect 1161 5289 1195 5320
rect 1233 5289 1267 5320
rect 1305 5289 1339 5320
rect 1377 5289 1411 5320
rect 1449 5289 1483 5320
rect 1521 5289 1555 5320
rect 1593 5289 1627 5320
rect 1665 5289 1699 5320
rect 1737 5289 1771 5320
rect 1809 5289 1843 5320
rect 1881 5289 1915 5320
rect 1953 5289 1987 5320
rect 2025 5289 2059 5320
rect 2097 5289 2131 5320
rect 2169 5289 2203 5320
rect 2241 5289 2275 5320
rect 2313 5289 2347 5323
rect 2385 5289 2419 5323
rect 2457 5289 2491 5323
rect 2529 5289 2563 5323
rect 2601 5289 2635 5323
rect 2673 5289 2707 5323
rect 2745 5289 2779 5323
rect 2817 5289 2851 5323
rect 2889 5289 2923 5323
rect 2961 5289 2995 5323
rect 3033 5289 3067 5323
rect 3105 5289 3139 5323
rect 3177 5289 3211 5323
rect 3249 5289 3283 5323
rect 3321 5289 3355 5323
rect 3393 5289 3427 5323
rect 3465 5289 3499 5323
rect 3537 5289 3571 5323
rect 3609 5289 3643 5323
rect 3681 5289 3715 5323
rect 3753 5289 3787 5323
rect 3825 5289 3859 5323
rect 3897 5289 3931 5323
rect 3969 5289 4003 5323
rect 4041 5289 4075 5323
rect 4113 5289 4147 5323
rect 4185 5289 4219 5323
rect 4257 5289 4291 5323
rect 4329 5289 4363 5323
rect 4401 5289 4435 5323
rect 4473 5289 4507 5323
rect 4545 5289 4579 5323
rect 4617 5289 4651 5323
rect 4689 5289 4723 5323
rect 4761 5289 4795 5323
rect 4833 5289 4867 5323
rect 4905 5289 4939 5323
rect 4977 5289 5011 5323
rect 5049 5289 5083 5323
rect 5121 5289 5155 5323
rect 5193 5289 5227 5323
rect 5265 5289 5299 5323
rect 5337 5289 5371 5323
rect 5409 5289 5443 5323
rect 5481 5289 5515 5323
rect 5553 5289 5587 5323
rect 5625 5289 5659 5323
rect 5697 5289 5731 5323
rect 5769 5289 5803 5323
rect 5841 5289 5875 5323
rect 5913 5289 5947 5323
rect 5985 5289 6019 5323
rect 6057 5289 6091 5323
rect 6129 5289 6163 5323
rect 6201 5289 6235 5323
rect 6273 5289 6307 5323
rect 6345 5289 6379 5323
rect 6417 5289 6451 5323
rect 6489 5289 6523 5323
rect 6561 5289 6595 5323
rect 6633 5289 6667 5323
rect 6705 5289 6739 5323
rect 6777 5289 6811 5323
rect 6849 5289 6883 5323
rect 6921 5289 6955 5323
rect 6993 5289 7027 5323
rect 7065 5289 7099 5323
rect 7137 5289 7171 5323
rect 7209 5289 7243 5323
rect 7281 5289 7315 5323
rect 7353 5289 7387 5323
rect 7425 5289 7459 5323
rect 7497 5289 7531 5323
rect 7569 5289 7603 5323
rect 7641 5289 7675 5323
rect 7713 5289 7747 5323
rect 7785 5289 7819 5323
rect 7857 5289 7891 5323
rect 7929 5289 7963 5323
rect 8001 5289 8035 5323
rect 8073 5289 8107 5323
rect 8145 5289 8179 5323
rect 8217 5289 8251 5323
rect 8289 5289 8323 5323
rect 8361 5289 8395 5323
rect 8433 5289 8467 5323
rect 8505 5289 8539 5323
rect 8577 5289 8611 5323
rect 8649 5289 8683 5323
rect 8721 5289 8755 5323
rect 8793 5289 8827 5323
rect 8865 5289 8899 5323
rect 8937 5289 8971 5323
rect 9009 5289 9043 5323
rect 9081 5289 9115 5323
rect 9153 5289 9187 5323
rect 9225 5289 9259 5323
rect 9297 5289 9331 5323
rect 9369 5289 9403 5323
rect 9441 5289 9475 5323
rect 9513 5289 9547 5323
rect 9585 5289 9619 5323
rect 9657 5289 9691 5323
rect 9729 5289 9763 5323
rect 9801 5289 9835 5323
rect 9873 5289 9907 5323
rect 9945 5289 9979 5323
rect 10017 5289 10051 5323
rect 10089 5289 10123 5323
rect 10161 5289 10195 5323
rect 10234 5289 10268 5323
rect 10307 5289 10341 5323
rect 10380 5289 10414 5323
rect 10453 5289 10487 5323
rect 10526 5289 10560 5323
rect 10599 5289 10633 5323
rect 10672 5289 10706 5323
rect 10745 5289 10779 5323
rect 10818 5289 10852 5323
rect 10891 5289 10925 5323
rect 10964 5289 10998 5323
rect 11037 5289 11071 5323
rect 11110 5289 11144 5323
rect 11183 5289 11217 5323
rect 11256 5289 11290 5323
rect 11329 5289 11363 5323
rect 11402 5289 11436 5323
rect 11475 5289 11509 5323
rect 11548 5289 11582 5323
rect 11621 5289 11655 5323
rect 11694 5289 11728 5323
rect 11767 5289 11801 5323
rect 11840 5289 11874 5323
rect 11913 5289 11947 5323
rect 11986 5289 12020 5323
rect 12059 5289 12093 5323
rect 12132 5289 12166 5323
rect 12205 5289 12239 5323
rect 12278 5289 12312 5323
rect 12351 5289 12385 5323
rect 12424 5289 12458 5323
rect 12497 5289 12531 5323
rect 12570 5289 12604 5323
rect 12643 5289 12677 5323
rect 12716 5289 12750 5323
rect 12789 5289 12823 5323
rect 12862 5289 12896 5323
rect 12935 5289 12969 5323
rect 13008 5289 13042 5323
rect 13081 5289 13115 5323
rect 13154 5289 13188 5323
rect 13227 5289 13261 5323
rect 13300 5289 13334 5323
rect 13373 5289 13407 5323
rect 13446 5289 13480 5323
rect 13519 5289 13553 5323
rect 13592 5289 13626 5323
rect 13665 5289 13699 5323
rect 13738 5289 13772 5323
rect 13811 5289 13845 5323
rect 13884 5289 13918 5323
rect 13957 5289 13991 5323
rect 14030 5289 14064 5323
rect 14103 5289 14137 5323
rect 14176 5289 14210 5323
rect 14249 5289 14283 5323
rect 14322 5289 14356 5323
rect 14395 5289 14429 5323
rect 14468 5289 14502 5323
rect 14541 5289 14575 5323
rect 14614 5289 14648 5323
rect 14687 5289 14721 5323
rect 14760 5289 14794 5323
rect 14833 5289 14867 5323
rect 14969 5281 15003 5315
rect 233 5207 267 5241
rect 369 5216 402 5250
rect 402 5216 403 5250
rect 233 5134 267 5168
rect 369 5143 402 5177
rect 402 5143 403 5177
rect 233 5061 267 5095
rect 369 5070 402 5104
rect 402 5070 403 5104
rect 233 4988 267 5022
rect 369 4997 402 5031
rect 402 4997 403 5031
rect 233 4915 267 4949
rect 369 4924 402 4958
rect 402 4924 403 4958
rect 14833 5217 14867 5251
rect 14969 5218 15003 5243
rect 14969 5209 14990 5218
rect 14990 5209 15003 5218
rect 14833 5145 14867 5179
rect 14969 5137 14990 5171
rect 14990 5137 15003 5171
rect 14833 5073 14867 5107
rect 14969 5065 14990 5099
rect 14990 5065 15003 5099
rect 14833 5001 14867 5035
rect 14969 4993 14990 5027
rect 14990 4993 15003 5027
rect 233 4842 267 4876
rect 369 4851 402 4885
rect 402 4851 403 4885
rect 233 4769 267 4803
rect 369 4778 402 4812
rect 402 4778 403 4812
rect 233 4696 267 4730
rect 369 4705 402 4739
rect 402 4705 403 4739
rect 233 4623 267 4657
rect 369 4632 402 4666
rect 402 4632 403 4666
rect 233 4550 267 4584
rect 369 4559 402 4593
rect 402 4559 403 4593
rect 233 4477 267 4511
rect 369 4486 402 4520
rect 402 4486 403 4520
rect 233 4404 267 4438
rect 369 4413 402 4447
rect 402 4413 403 4447
rect 233 4331 267 4365
rect 369 4340 402 4374
rect 402 4340 403 4374
rect 233 4258 267 4292
rect 369 4267 402 4301
rect 402 4267 403 4301
rect 233 4185 267 4219
rect 369 4194 402 4228
rect 402 4194 403 4228
rect 233 4112 267 4146
rect 369 4121 402 4155
rect 402 4121 403 4155
rect 233 4039 267 4073
rect 369 4048 402 4082
rect 402 4048 403 4082
rect 233 3966 267 4000
rect 369 3975 402 4009
rect 402 3975 403 4009
rect 233 3893 267 3927
rect 369 3902 402 3936
rect 402 3902 403 3936
rect 233 3820 267 3854
rect 369 3829 402 3863
rect 402 3829 403 3863
rect 233 3747 267 3781
rect 369 3756 402 3790
rect 402 3756 403 3790
rect 233 3674 267 3708
rect 369 3683 402 3717
rect 402 3683 403 3717
rect 233 3601 267 3635
rect 369 3610 402 3644
rect 402 3610 403 3644
rect 233 3528 267 3562
rect 369 3537 402 3571
rect 402 3537 403 3571
rect 233 3455 267 3489
rect 369 3464 402 3498
rect 402 3464 403 3498
rect 233 3382 267 3416
rect 369 3391 402 3425
rect 402 3391 403 3425
rect 233 3309 267 3343
rect 369 3318 402 3352
rect 402 3318 403 3352
rect 233 3236 267 3270
rect 369 3245 402 3279
rect 402 3245 403 3279
rect 233 3163 267 3197
rect 369 3172 402 3206
rect 402 3172 403 3206
rect 233 3090 267 3124
rect 369 3099 402 3133
rect 402 3099 403 3133
rect 233 3017 267 3051
rect 369 3026 402 3060
rect 402 3026 403 3060
rect 233 2944 267 2978
rect 369 2953 402 2987
rect 402 2953 403 2987
rect 233 2871 267 2905
rect 369 2880 402 2914
rect 402 2880 403 2914
rect 233 2798 267 2832
rect 369 2807 402 2841
rect 402 2807 403 2841
rect 233 2725 267 2759
rect 369 2734 402 2768
rect 402 2734 403 2768
rect 233 2652 267 2686
rect 369 2661 402 2695
rect 402 2661 403 2695
rect 233 2579 267 2613
rect 369 2588 402 2622
rect 402 2588 403 2622
rect 233 2506 267 2540
rect 369 2515 402 2549
rect 402 2515 403 2549
rect 233 2433 267 2467
rect 369 2442 402 2476
rect 402 2442 403 2476
rect 233 2360 267 2394
rect 369 2369 402 2403
rect 402 2369 403 2403
rect 233 2287 267 2321
rect 369 2296 402 2330
rect 402 2296 403 2330
rect 233 2214 267 2248
rect 369 2223 402 2257
rect 402 2223 403 2257
rect 233 2141 267 2175
rect 369 2150 402 2184
rect 402 2150 403 2184
rect 233 2068 267 2102
rect 369 2077 402 2111
rect 402 2077 403 2111
rect 233 1995 267 2029
rect 369 2004 402 2038
rect 402 2004 403 2038
rect 233 1922 267 1956
rect 369 1931 402 1965
rect 402 1931 403 1965
rect 233 1849 267 1883
rect 369 1858 402 1892
rect 402 1858 403 1892
rect 233 1776 267 1810
rect 369 1785 402 1819
rect 402 1785 403 1819
rect 233 1703 267 1737
rect 369 1712 402 1746
rect 402 1712 403 1746
rect 233 1630 267 1664
rect 369 1639 402 1673
rect 402 1639 403 1673
rect 233 1558 267 1592
rect 369 1566 402 1600
rect 402 1566 403 1600
rect 233 1486 267 1520
rect 369 1493 402 1527
rect 402 1493 403 1527
rect 233 1414 267 1448
rect 369 1420 402 1454
rect 402 1420 403 1454
rect 233 1342 267 1376
rect 369 1347 402 1381
rect 402 1347 403 1381
rect 233 1270 267 1304
rect 369 1274 402 1308
rect 402 1274 403 1308
rect 233 1198 267 1232
rect 369 1201 402 1235
rect 402 1201 403 1235
rect 233 1126 267 1160
rect 369 1128 402 1162
rect 402 1128 403 1162
rect 233 1054 267 1088
rect 369 1055 402 1089
rect 402 1055 403 1089
rect 233 982 267 1016
rect 369 982 402 1016
rect 402 982 403 1016
rect 767 4818 12465 4924
rect 12504 4890 12538 4924
rect 12577 4890 12611 4924
rect 12650 4890 12684 4924
rect 12723 4890 12757 4924
rect 12796 4890 12830 4924
rect 12869 4890 12903 4924
rect 12942 4890 12976 4924
rect 13015 4890 13049 4924
rect 13088 4890 13122 4924
rect 13161 4890 13195 4924
rect 13234 4890 13268 4924
rect 13307 4890 13341 4924
rect 13380 4890 13414 4924
rect 13453 4890 13487 4924
rect 13526 4890 13560 4924
rect 13599 4890 13633 4924
rect 13672 4890 13706 4924
rect 13745 4890 13779 4924
rect 13818 4890 13852 4924
rect 13891 4890 13925 4924
rect 13964 4890 13998 4924
rect 14037 4890 14071 4924
rect 14110 4890 14144 4924
rect 14183 4890 14217 4924
rect 14256 4890 14290 4924
rect 14329 4890 14363 4924
rect 14402 4890 14436 4924
rect 12504 4818 12538 4852
rect 12577 4818 12611 4852
rect 12650 4818 12684 4852
rect 12723 4818 12757 4852
rect 12796 4818 12830 4852
rect 12869 4818 12903 4852
rect 12942 4818 12976 4852
rect 13015 4818 13049 4852
rect 13088 4818 13122 4852
rect 13161 4818 13195 4852
rect 13234 4818 13268 4852
rect 13307 4818 13341 4852
rect 13380 4818 13414 4852
rect 13453 4818 13487 4852
rect 13526 4818 13560 4852
rect 13599 4818 13633 4852
rect 13672 4818 13706 4852
rect 13745 4818 13779 4852
rect 13818 4818 13852 4852
rect 13891 4818 13925 4852
rect 13964 4818 13998 4852
rect 14037 4818 14071 4852
rect 14110 4818 14144 4852
rect 14183 4818 14217 4852
rect 14256 4818 14290 4852
rect 14329 4818 14363 4852
rect 14402 4820 14436 4852
rect 14402 4818 14428 4820
rect 14428 4818 14436 4820
rect 587 4710 621 4744
rect 659 4717 691 4744
rect 691 4717 693 4744
rect 733 4740 767 4774
rect 659 4710 693 4717
rect 587 4636 621 4670
rect 659 4648 691 4670
rect 691 4648 693 4670
rect 733 4667 767 4701
rect 659 4636 693 4648
rect 587 4563 621 4596
rect 587 4562 589 4563
rect 589 4562 621 4563
rect 659 4562 693 4596
rect 733 4594 767 4628
rect 587 4492 621 4522
rect 587 4488 589 4492
rect 589 4488 621 4492
rect 659 4488 693 4522
rect 733 4521 767 4555
rect 14431 4740 14465 4774
rect 14510 4716 14531 4743
rect 14531 4716 14544 4743
rect 14510 4709 14544 4716
rect 14582 4714 14599 4743
rect 14599 4714 14616 4743
rect 14582 4709 14616 4714
rect 14431 4667 14465 4701
rect 14510 4646 14531 4670
rect 14531 4646 14544 4670
rect 14510 4636 14544 4646
rect 14582 4644 14599 4670
rect 14599 4644 14616 4670
rect 14582 4636 14616 4644
rect 14431 4594 14465 4628
rect 14510 4576 14531 4597
rect 14531 4576 14544 4597
rect 14510 4563 14544 4576
rect 14582 4574 14599 4597
rect 14599 4574 14616 4597
rect 14582 4563 14616 4574
rect 14431 4521 14465 4555
rect 14510 4506 14531 4524
rect 14531 4506 14544 4524
rect 587 4421 621 4449
rect 587 4415 589 4421
rect 589 4415 621 4421
rect 659 4415 693 4449
rect 733 4448 767 4482
rect 587 4350 621 4376
rect 587 4342 589 4350
rect 589 4342 621 4350
rect 659 4342 693 4376
rect 733 4375 767 4409
rect 587 4279 621 4303
rect 587 4269 589 4279
rect 589 4269 621 4279
rect 659 4269 693 4303
rect 733 4302 767 4336
rect 587 4208 621 4230
rect 587 4196 589 4208
rect 589 4196 621 4208
rect 659 4196 693 4230
rect 733 4229 767 4263
rect 587 4137 621 4157
rect 587 4123 589 4137
rect 589 4123 621 4137
rect 659 4123 693 4157
rect 733 4156 767 4190
rect 587 4050 621 4084
rect 659 4050 693 4084
rect 733 4083 767 4117
rect 931 4388 1037 4494
rect 587 4007 589 4011
rect 589 4007 621 4011
rect 733 4034 767 4044
rect 587 3977 621 4007
rect 659 3977 693 4011
rect 733 4010 734 4034
rect 734 4010 767 4034
rect 587 3936 589 3938
rect 589 3936 621 3938
rect 733 3966 767 3971
rect 587 3904 621 3936
rect 659 3904 693 3938
rect 733 3937 734 3966
rect 734 3937 767 3966
rect 587 3862 589 3865
rect 589 3862 621 3865
rect 587 3831 621 3862
rect 659 3831 693 3865
rect 733 3864 734 3898
rect 734 3864 767 3898
rect 587 3791 589 3792
rect 589 3791 621 3792
rect 733 3796 734 3825
rect 734 3796 767 3825
rect 587 3758 621 3791
rect 659 3758 693 3792
rect 733 3791 767 3796
rect 587 3717 589 3719
rect 589 3717 621 3719
rect 733 3728 734 3752
rect 734 3728 767 3752
rect 587 3685 621 3717
rect 659 3685 693 3719
rect 733 3718 767 3728
rect 733 3660 734 3679
rect 734 3660 767 3679
rect 587 3612 621 3646
rect 659 3612 693 3646
rect 733 3645 767 3660
rect 587 3572 589 3573
rect 589 3572 621 3573
rect 733 3592 734 3606
rect 734 3592 767 3606
rect 587 3539 621 3572
rect 659 3539 693 3573
rect 733 3572 767 3592
rect 733 3524 734 3533
rect 734 3524 767 3533
rect 587 3466 621 3500
rect 659 3466 693 3500
rect 733 3499 767 3524
rect 733 3456 734 3460
rect 734 3456 767 3460
rect 587 3393 621 3427
rect 659 3393 693 3427
rect 733 3426 767 3456
rect 733 3354 767 3387
rect 587 3320 621 3354
rect 659 3320 693 3354
rect 733 3353 734 3354
rect 734 3353 767 3354
rect 733 3286 767 3314
rect 587 3247 621 3281
rect 659 3247 693 3281
rect 733 3280 734 3286
rect 734 3280 767 3286
rect 733 3218 767 3241
rect 587 3174 621 3208
rect 659 3174 693 3208
rect 733 3207 734 3218
rect 734 3207 767 3218
rect 587 3117 589 3135
rect 589 3117 621 3135
rect 733 3150 767 3168
rect 587 3101 621 3117
rect 659 3101 693 3135
rect 733 3134 734 3150
rect 734 3134 767 3150
rect 587 3028 621 3062
rect 659 3028 693 3062
rect 733 3061 767 3095
rect 587 2955 621 2989
rect 659 2955 693 2989
rect 733 2988 767 3022
rect 587 2882 621 2916
rect 659 2882 693 2916
rect 733 2915 767 2949
rect 587 2809 621 2843
rect 659 2809 693 2843
rect 733 2842 767 2876
rect 587 2736 621 2770
rect 659 2736 693 2770
rect 733 2769 767 2803
rect 587 2663 621 2697
rect 659 2663 693 2697
rect 733 2696 767 2730
rect 587 2590 621 2624
rect 659 2590 693 2624
rect 733 2623 767 2657
rect 587 2517 621 2551
rect 659 2517 693 2551
rect 733 2550 767 2584
rect 587 2444 621 2478
rect 659 2444 693 2478
rect 733 2477 767 2511
rect 1361 4388 1467 4494
rect 733 2433 767 2438
rect 587 2371 621 2405
rect 659 2371 693 2405
rect 733 2404 734 2433
rect 734 2404 767 2433
rect 587 2327 621 2332
rect 587 2298 589 2327
rect 589 2298 621 2327
rect 659 2298 693 2332
rect 733 2331 734 2365
rect 734 2331 767 2365
rect 733 2263 734 2292
rect 734 2263 767 2292
rect 587 2250 621 2259
rect 587 2225 589 2250
rect 589 2225 621 2250
rect 659 2225 693 2259
rect 733 2258 767 2263
rect 733 2195 734 2219
rect 734 2195 767 2219
rect 587 2156 621 2186
rect 587 2152 589 2156
rect 589 2152 621 2156
rect 659 2152 693 2186
rect 733 2185 767 2195
rect 733 2127 734 2146
rect 734 2127 767 2146
rect 587 2085 621 2113
rect 587 2079 589 2085
rect 589 2079 621 2085
rect 659 2079 693 2113
rect 733 2112 767 2127
rect 733 2059 734 2073
rect 734 2059 767 2073
rect 587 2011 621 2040
rect 587 2006 589 2011
rect 589 2006 621 2011
rect 659 2006 693 2040
rect 733 2039 767 2059
rect 733 1991 734 2000
rect 734 1991 767 2000
rect 587 1940 621 1967
rect 587 1933 589 1940
rect 589 1933 621 1940
rect 659 1933 693 1967
rect 733 1966 767 1991
rect 733 1923 734 1927
rect 734 1923 767 1927
rect 587 1866 621 1894
rect 587 1860 589 1866
rect 589 1860 621 1866
rect 659 1860 693 1894
rect 733 1893 767 1923
rect 733 1821 767 1854
rect 587 1795 621 1821
rect 587 1787 589 1795
rect 589 1787 621 1795
rect 659 1787 693 1821
rect 733 1820 734 1821
rect 734 1820 767 1821
rect 733 1753 767 1781
rect 587 1721 621 1748
rect 587 1714 589 1721
rect 589 1714 621 1721
rect 659 1714 693 1748
rect 733 1747 734 1753
rect 734 1747 767 1753
rect 733 1685 767 1708
rect 587 1650 621 1675
rect 587 1641 589 1650
rect 589 1641 621 1650
rect 659 1641 693 1675
rect 733 1674 734 1685
rect 734 1674 767 1685
rect 733 1617 767 1635
rect 587 1576 621 1602
rect 587 1568 589 1576
rect 589 1568 621 1576
rect 659 1568 693 1602
rect 733 1601 734 1617
rect 734 1601 767 1617
rect 733 1549 767 1562
rect 587 1505 621 1529
rect 587 1495 589 1505
rect 589 1495 621 1505
rect 659 1495 693 1529
rect 733 1528 734 1549
rect 734 1528 767 1549
rect 733 1455 767 1489
rect 587 1385 621 1419
rect 659 1385 693 1419
rect 733 1382 767 1416
rect 587 1296 621 1330
rect 659 1296 693 1330
rect 733 1308 767 1342
rect 1110 4028 1144 4062
rect 1182 4028 1216 4062
rect 1254 4028 1288 4062
rect 1110 3954 1144 3988
rect 1182 3954 1216 3988
rect 1254 3954 1288 3988
rect 1110 3880 1144 3914
rect 1182 3880 1216 3914
rect 1254 3880 1288 3914
rect 1110 3806 1144 3840
rect 1182 3806 1216 3840
rect 1254 3806 1288 3840
rect 1110 3732 1144 3766
rect 1182 3732 1216 3766
rect 1254 3732 1288 3766
rect 1110 3658 1144 3692
rect 1182 3658 1216 3692
rect 1254 3658 1288 3692
rect 1110 3584 1144 3618
rect 1182 3584 1216 3618
rect 1254 3584 1288 3618
rect 1110 3510 1144 3544
rect 1182 3510 1216 3544
rect 1254 3510 1288 3544
rect 1110 3436 1144 3470
rect 1182 3436 1216 3470
rect 1254 3436 1288 3470
rect 1110 3362 1144 3396
rect 1182 3362 1216 3396
rect 1254 3362 1288 3396
rect 1110 3288 1144 3322
rect 1182 3288 1216 3322
rect 1254 3288 1288 3322
rect 1110 3214 1144 3248
rect 1182 3214 1216 3248
rect 1254 3214 1288 3248
rect 1110 3140 1144 3174
rect 1182 3140 1216 3174
rect 1254 3140 1288 3174
rect 1110 3066 1144 3100
rect 1182 3066 1216 3100
rect 1254 3066 1288 3100
rect 1110 2992 1144 3026
rect 1182 2992 1216 3026
rect 1254 2992 1288 3026
rect 1110 2918 1144 2952
rect 1182 2918 1216 2952
rect 1254 2918 1288 2952
rect 1110 2844 1144 2878
rect 1182 2844 1216 2878
rect 1254 2844 1288 2878
rect 1110 2770 1144 2804
rect 1182 2770 1216 2804
rect 1254 2770 1288 2804
rect 1110 2696 1144 2730
rect 1182 2696 1216 2730
rect 1254 2696 1288 2730
rect 1110 2622 1144 2656
rect 1182 2622 1216 2656
rect 1254 2622 1288 2656
rect 1110 2548 1144 2582
rect 1182 2548 1216 2582
rect 1254 2548 1288 2582
rect 1110 2474 1144 2508
rect 1182 2474 1216 2508
rect 1254 2474 1288 2508
rect 1110 2400 1144 2434
rect 1182 2400 1216 2434
rect 1254 2400 1288 2434
rect 1110 2326 1144 2360
rect 1182 2326 1216 2360
rect 1254 2326 1288 2360
rect 1110 2252 1144 2286
rect 1182 2252 1216 2286
rect 1254 2252 1288 2286
rect 1110 2178 1144 2212
rect 1182 2178 1216 2212
rect 1254 2178 1288 2212
rect 1110 2104 1144 2138
rect 1182 2104 1216 2138
rect 1254 2104 1288 2138
rect 1110 2030 1144 2064
rect 1182 2030 1216 2064
rect 1254 2030 1288 2064
rect 1110 1956 1144 1990
rect 1182 1956 1216 1990
rect 1254 1956 1288 1990
rect 1110 1882 1144 1916
rect 1182 1882 1216 1916
rect 1254 1882 1288 1916
rect 1110 1808 1144 1842
rect 1182 1808 1216 1842
rect 1254 1808 1288 1842
rect 1110 1734 1144 1768
rect 1182 1734 1216 1768
rect 1254 1734 1288 1768
rect 1110 1660 1144 1694
rect 1182 1660 1216 1694
rect 1254 1660 1288 1694
rect 1110 1586 1144 1620
rect 1182 1586 1216 1620
rect 1254 1586 1288 1620
rect 1110 1511 1144 1545
rect 1182 1511 1216 1545
rect 1254 1511 1288 1545
rect 1923 4388 2029 4494
rect 1678 4050 1712 4062
rect 1606 4046 1784 4050
rect 1606 4012 1610 4046
rect 1610 4012 1678 4046
rect 1678 4012 1712 4046
rect 1712 4012 1780 4046
rect 1780 4012 1784 4046
rect 1606 3978 1784 4012
rect 1606 3944 1610 3978
rect 1610 3944 1678 3978
rect 1678 3944 1712 3978
rect 1712 3944 1780 3978
rect 1780 3944 1784 3978
rect 1606 3910 1784 3944
rect 1606 3876 1610 3910
rect 1610 3876 1678 3910
rect 1678 3876 1712 3910
rect 1712 3876 1780 3910
rect 1780 3876 1784 3910
rect 1606 3842 1784 3876
rect 1606 3808 1610 3842
rect 1610 3808 1678 3842
rect 1678 3808 1712 3842
rect 1712 3808 1780 3842
rect 1780 3808 1784 3842
rect 1606 3774 1784 3808
rect 1606 3740 1610 3774
rect 1610 3740 1678 3774
rect 1678 3740 1712 3774
rect 1712 3740 1780 3774
rect 1780 3740 1784 3774
rect 1606 3706 1784 3740
rect 1606 3672 1610 3706
rect 1610 3672 1678 3706
rect 1678 3672 1712 3706
rect 1712 3672 1780 3706
rect 1780 3672 1784 3706
rect 1606 3638 1784 3672
rect 1606 3604 1610 3638
rect 1610 3604 1678 3638
rect 1678 3604 1712 3638
rect 1712 3604 1780 3638
rect 1780 3604 1784 3638
rect 1606 3570 1784 3604
rect 1606 3536 1610 3570
rect 1610 3536 1678 3570
rect 1678 3536 1712 3570
rect 1712 3536 1780 3570
rect 1780 3536 1784 3570
rect 1606 3502 1784 3536
rect 1606 3468 1610 3502
rect 1610 3468 1678 3502
rect 1678 3468 1712 3502
rect 1712 3468 1780 3502
rect 1780 3468 1784 3502
rect 1606 3434 1784 3468
rect 1606 3400 1610 3434
rect 1610 3400 1678 3434
rect 1678 3400 1712 3434
rect 1712 3400 1780 3434
rect 1780 3400 1784 3434
rect 1606 3366 1784 3400
rect 1606 3332 1610 3366
rect 1610 3332 1678 3366
rect 1678 3332 1712 3366
rect 1712 3332 1780 3366
rect 1780 3332 1784 3366
rect 1606 3298 1784 3332
rect 1606 3264 1610 3298
rect 1610 3264 1678 3298
rect 1678 3264 1712 3298
rect 1712 3264 1780 3298
rect 1780 3264 1784 3298
rect 1606 3230 1784 3264
rect 1606 3196 1610 3230
rect 1610 3196 1678 3230
rect 1678 3196 1712 3230
rect 1712 3196 1780 3230
rect 1780 3196 1784 3230
rect 1606 3162 1784 3196
rect 1606 3128 1610 3162
rect 1610 3128 1678 3162
rect 1678 3128 1712 3162
rect 1712 3128 1780 3162
rect 1780 3128 1784 3162
rect 1606 3092 1784 3128
rect 1606 3080 1640 3092
rect 1750 3080 1784 3092
rect 1606 2935 1784 3040
rect 1606 2901 1645 2935
rect 1645 2901 1679 2935
rect 1679 2901 1713 2935
rect 1713 2901 1747 2935
rect 1747 2901 1784 2935
rect 1606 2855 1784 2901
rect 1606 2821 1645 2855
rect 1645 2821 1679 2855
rect 1679 2821 1713 2855
rect 1713 2821 1747 2855
rect 1747 2821 1784 2855
rect 1606 2775 1784 2821
rect 1606 2741 1645 2775
rect 1645 2741 1679 2775
rect 1679 2741 1713 2775
rect 1713 2741 1747 2775
rect 1747 2741 1784 2775
rect 1606 2695 1784 2741
rect 1606 2661 1645 2695
rect 1645 2661 1679 2695
rect 1679 2661 1713 2695
rect 1713 2661 1747 2695
rect 1747 2661 1784 2695
rect 1606 2614 1784 2661
rect 1606 2580 1645 2614
rect 1645 2580 1679 2614
rect 1679 2580 1713 2614
rect 1713 2580 1747 2614
rect 1747 2580 1784 2614
rect 1606 2574 1784 2580
rect 1606 2501 1640 2535
rect 1678 2501 1712 2535
rect 1750 2501 1784 2535
rect 1678 2449 1712 2461
rect 1606 2445 1784 2449
rect 1606 2411 1610 2445
rect 1610 2411 1678 2445
rect 1678 2411 1712 2445
rect 1712 2411 1780 2445
rect 1780 2411 1784 2445
rect 1606 2377 1784 2411
rect 1606 2343 1610 2377
rect 1610 2343 1678 2377
rect 1678 2343 1712 2377
rect 1712 2343 1780 2377
rect 1780 2343 1784 2377
rect 1606 2309 1784 2343
rect 1606 2275 1610 2309
rect 1610 2275 1678 2309
rect 1678 2275 1712 2309
rect 1712 2275 1780 2309
rect 1780 2275 1784 2309
rect 1606 2241 1784 2275
rect 1606 2207 1610 2241
rect 1610 2207 1678 2241
rect 1678 2207 1712 2241
rect 1712 2207 1780 2241
rect 1780 2207 1784 2241
rect 1606 2173 1784 2207
rect 1606 2139 1610 2173
rect 1610 2139 1678 2173
rect 1678 2139 1712 2173
rect 1712 2139 1780 2173
rect 1780 2139 1784 2173
rect 1606 2105 1784 2139
rect 1606 2071 1610 2105
rect 1610 2071 1678 2105
rect 1678 2071 1712 2105
rect 1712 2071 1780 2105
rect 1780 2071 1784 2105
rect 1606 2037 1784 2071
rect 1606 2003 1610 2037
rect 1610 2003 1678 2037
rect 1678 2003 1712 2037
rect 1712 2003 1780 2037
rect 1780 2003 1784 2037
rect 1606 1969 1784 2003
rect 1606 1935 1610 1969
rect 1610 1935 1678 1969
rect 1678 1935 1712 1969
rect 1712 1935 1780 1969
rect 1780 1935 1784 1969
rect 1606 1901 1784 1935
rect 1606 1867 1610 1901
rect 1610 1867 1678 1901
rect 1678 1867 1712 1901
rect 1712 1867 1780 1901
rect 1780 1867 1784 1901
rect 1606 1833 1784 1867
rect 1606 1799 1610 1833
rect 1610 1799 1678 1833
rect 1678 1799 1712 1833
rect 1712 1799 1780 1833
rect 1780 1799 1784 1833
rect 1606 1765 1784 1799
rect 1606 1731 1610 1765
rect 1610 1731 1678 1765
rect 1678 1731 1712 1765
rect 1712 1731 1780 1765
rect 1780 1731 1784 1765
rect 1606 1697 1784 1731
rect 1606 1663 1610 1697
rect 1610 1663 1678 1697
rect 1678 1663 1712 1697
rect 1712 1663 1780 1697
rect 1780 1663 1784 1697
rect 1606 1629 1784 1663
rect 1606 1595 1610 1629
rect 1610 1595 1678 1629
rect 1678 1595 1712 1629
rect 1712 1595 1780 1629
rect 1780 1595 1784 1629
rect 1606 1561 1784 1595
rect 1606 1527 1610 1561
rect 1610 1527 1678 1561
rect 1678 1527 1712 1561
rect 1712 1527 1780 1561
rect 1780 1527 1784 1561
rect 1606 1491 1784 1527
rect 1606 1479 1640 1491
rect 1750 1479 1784 1491
rect 2353 4388 2459 4494
rect 2102 4028 2136 4062
rect 2174 4028 2208 4062
rect 2246 4028 2280 4062
rect 2102 3954 2136 3988
rect 2174 3954 2208 3988
rect 2246 3954 2280 3988
rect 2102 3880 2136 3914
rect 2174 3880 2208 3914
rect 2246 3880 2280 3914
rect 2102 3806 2136 3840
rect 2174 3806 2208 3840
rect 2246 3806 2280 3840
rect 2102 3732 2136 3766
rect 2174 3732 2208 3766
rect 2246 3732 2280 3766
rect 2102 3658 2136 3692
rect 2174 3658 2208 3692
rect 2246 3658 2280 3692
rect 2102 3584 2136 3618
rect 2174 3584 2208 3618
rect 2246 3584 2280 3618
rect 2102 3510 2136 3544
rect 2174 3510 2208 3544
rect 2246 3510 2280 3544
rect 2102 3436 2136 3470
rect 2174 3436 2208 3470
rect 2246 3436 2280 3470
rect 2102 3362 2136 3396
rect 2174 3362 2208 3396
rect 2246 3362 2280 3396
rect 2102 3288 2136 3322
rect 2174 3288 2208 3322
rect 2246 3288 2280 3322
rect 2102 3214 2136 3248
rect 2174 3214 2208 3248
rect 2246 3214 2280 3248
rect 2102 3140 2136 3174
rect 2174 3140 2208 3174
rect 2246 3140 2280 3174
rect 2102 3066 2136 3100
rect 2174 3066 2208 3100
rect 2246 3066 2280 3100
rect 2102 2992 2136 3026
rect 2174 2992 2208 3026
rect 2246 2992 2280 3026
rect 2102 2918 2136 2952
rect 2174 2918 2208 2952
rect 2246 2918 2280 2952
rect 2102 2844 2136 2878
rect 2174 2844 2208 2878
rect 2246 2844 2280 2878
rect 2102 2770 2136 2804
rect 2174 2770 2208 2804
rect 2246 2770 2280 2804
rect 2102 2696 2136 2730
rect 2174 2696 2208 2730
rect 2246 2696 2280 2730
rect 2102 2622 2136 2656
rect 2174 2622 2208 2656
rect 2246 2622 2280 2656
rect 2102 2548 2136 2582
rect 2174 2548 2208 2582
rect 2246 2548 2280 2582
rect 2102 2474 2136 2508
rect 2174 2474 2208 2508
rect 2246 2474 2280 2508
rect 2102 2400 2136 2434
rect 2174 2400 2208 2434
rect 2246 2400 2280 2434
rect 2102 2326 2136 2360
rect 2174 2326 2208 2360
rect 2246 2326 2280 2360
rect 2102 2252 2136 2286
rect 2174 2252 2208 2286
rect 2246 2252 2280 2286
rect 2102 2178 2136 2212
rect 2174 2178 2208 2212
rect 2246 2178 2280 2212
rect 2102 2104 2136 2138
rect 2174 2104 2208 2138
rect 2246 2104 2280 2138
rect 2102 2030 2136 2064
rect 2174 2030 2208 2064
rect 2246 2030 2280 2064
rect 2102 1956 2136 1990
rect 2174 1956 2208 1990
rect 2246 1956 2280 1990
rect 2102 1882 2136 1916
rect 2174 1882 2208 1916
rect 2246 1882 2280 1916
rect 2102 1808 2136 1842
rect 2174 1808 2208 1842
rect 2246 1808 2280 1842
rect 2102 1734 2136 1768
rect 2174 1734 2208 1768
rect 2246 1734 2280 1768
rect 2102 1660 2136 1694
rect 2174 1660 2208 1694
rect 2246 1660 2280 1694
rect 2102 1586 2136 1620
rect 2174 1586 2208 1620
rect 2246 1586 2280 1620
rect 2102 1511 2136 1545
rect 2174 1511 2208 1545
rect 2246 1511 2280 1545
rect 2915 4388 3021 4494
rect 2670 4050 2704 4062
rect 2598 4046 2776 4050
rect 2598 4012 2602 4046
rect 2602 4012 2670 4046
rect 2670 4012 2704 4046
rect 2704 4012 2772 4046
rect 2772 4012 2776 4046
rect 2598 3978 2776 4012
rect 2598 3944 2602 3978
rect 2602 3944 2670 3978
rect 2670 3944 2704 3978
rect 2704 3944 2772 3978
rect 2772 3944 2776 3978
rect 2598 3910 2776 3944
rect 2598 3876 2602 3910
rect 2602 3876 2670 3910
rect 2670 3876 2704 3910
rect 2704 3876 2772 3910
rect 2772 3876 2776 3910
rect 2598 3842 2776 3876
rect 2598 3808 2602 3842
rect 2602 3808 2670 3842
rect 2670 3808 2704 3842
rect 2704 3808 2772 3842
rect 2772 3808 2776 3842
rect 2598 3774 2776 3808
rect 2598 3740 2602 3774
rect 2602 3740 2670 3774
rect 2670 3740 2704 3774
rect 2704 3740 2772 3774
rect 2772 3740 2776 3774
rect 2598 3706 2776 3740
rect 2598 3672 2602 3706
rect 2602 3672 2670 3706
rect 2670 3672 2704 3706
rect 2704 3672 2772 3706
rect 2772 3672 2776 3706
rect 2598 3638 2776 3672
rect 2598 3604 2602 3638
rect 2602 3604 2670 3638
rect 2670 3604 2704 3638
rect 2704 3604 2772 3638
rect 2772 3604 2776 3638
rect 2598 3570 2776 3604
rect 2598 3536 2602 3570
rect 2602 3536 2670 3570
rect 2670 3536 2704 3570
rect 2704 3536 2772 3570
rect 2772 3536 2776 3570
rect 2598 3502 2776 3536
rect 2598 3468 2602 3502
rect 2602 3468 2670 3502
rect 2670 3468 2704 3502
rect 2704 3468 2772 3502
rect 2772 3468 2776 3502
rect 2598 3434 2776 3468
rect 2598 3400 2602 3434
rect 2602 3400 2670 3434
rect 2670 3400 2704 3434
rect 2704 3400 2772 3434
rect 2772 3400 2776 3434
rect 2598 3366 2776 3400
rect 2598 3332 2602 3366
rect 2602 3332 2670 3366
rect 2670 3332 2704 3366
rect 2704 3332 2772 3366
rect 2772 3332 2776 3366
rect 2598 3298 2776 3332
rect 2598 3264 2602 3298
rect 2602 3264 2670 3298
rect 2670 3264 2704 3298
rect 2704 3264 2772 3298
rect 2772 3264 2776 3298
rect 2598 3230 2776 3264
rect 2598 3196 2602 3230
rect 2602 3196 2670 3230
rect 2670 3196 2704 3230
rect 2704 3196 2772 3230
rect 2772 3196 2776 3230
rect 2598 3162 2776 3196
rect 2598 3128 2602 3162
rect 2602 3128 2670 3162
rect 2670 3128 2704 3162
rect 2704 3128 2772 3162
rect 2772 3128 2776 3162
rect 2598 3092 2776 3128
rect 2598 3080 2632 3092
rect 2742 3080 2776 3092
rect 2598 2935 2776 3040
rect 2598 2901 2637 2935
rect 2637 2901 2671 2935
rect 2671 2901 2705 2935
rect 2705 2901 2739 2935
rect 2739 2901 2776 2935
rect 2598 2855 2776 2901
rect 2598 2821 2637 2855
rect 2637 2821 2671 2855
rect 2671 2821 2705 2855
rect 2705 2821 2739 2855
rect 2739 2821 2776 2855
rect 2598 2775 2776 2821
rect 2598 2741 2637 2775
rect 2637 2741 2671 2775
rect 2671 2741 2705 2775
rect 2705 2741 2739 2775
rect 2739 2741 2776 2775
rect 2598 2695 2776 2741
rect 2598 2661 2637 2695
rect 2637 2661 2671 2695
rect 2671 2661 2705 2695
rect 2705 2661 2739 2695
rect 2739 2661 2776 2695
rect 2598 2614 2776 2661
rect 2598 2580 2637 2614
rect 2637 2580 2671 2614
rect 2671 2580 2705 2614
rect 2705 2580 2739 2614
rect 2739 2580 2776 2614
rect 2598 2574 2776 2580
rect 2598 2501 2632 2535
rect 2670 2501 2704 2535
rect 2742 2501 2776 2535
rect 2670 2449 2704 2461
rect 2598 2445 2776 2449
rect 2598 2411 2602 2445
rect 2602 2411 2670 2445
rect 2670 2411 2704 2445
rect 2704 2411 2772 2445
rect 2772 2411 2776 2445
rect 2598 2377 2776 2411
rect 2598 2343 2602 2377
rect 2602 2343 2670 2377
rect 2670 2343 2704 2377
rect 2704 2343 2772 2377
rect 2772 2343 2776 2377
rect 2598 2309 2776 2343
rect 2598 2275 2602 2309
rect 2602 2275 2670 2309
rect 2670 2275 2704 2309
rect 2704 2275 2772 2309
rect 2772 2275 2776 2309
rect 2598 2241 2776 2275
rect 2598 2207 2602 2241
rect 2602 2207 2670 2241
rect 2670 2207 2704 2241
rect 2704 2207 2772 2241
rect 2772 2207 2776 2241
rect 2598 2173 2776 2207
rect 2598 2139 2602 2173
rect 2602 2139 2670 2173
rect 2670 2139 2704 2173
rect 2704 2139 2772 2173
rect 2772 2139 2776 2173
rect 2598 2105 2776 2139
rect 2598 2071 2602 2105
rect 2602 2071 2670 2105
rect 2670 2071 2704 2105
rect 2704 2071 2772 2105
rect 2772 2071 2776 2105
rect 2598 2037 2776 2071
rect 2598 2003 2602 2037
rect 2602 2003 2670 2037
rect 2670 2003 2704 2037
rect 2704 2003 2772 2037
rect 2772 2003 2776 2037
rect 2598 1969 2776 2003
rect 2598 1935 2602 1969
rect 2602 1935 2670 1969
rect 2670 1935 2704 1969
rect 2704 1935 2772 1969
rect 2772 1935 2776 1969
rect 2598 1901 2776 1935
rect 2598 1867 2602 1901
rect 2602 1867 2670 1901
rect 2670 1867 2704 1901
rect 2704 1867 2772 1901
rect 2772 1867 2776 1901
rect 2598 1833 2776 1867
rect 2598 1799 2602 1833
rect 2602 1799 2670 1833
rect 2670 1799 2704 1833
rect 2704 1799 2772 1833
rect 2772 1799 2776 1833
rect 2598 1765 2776 1799
rect 2598 1731 2602 1765
rect 2602 1731 2670 1765
rect 2670 1731 2704 1765
rect 2704 1731 2772 1765
rect 2772 1731 2776 1765
rect 2598 1697 2776 1731
rect 2598 1663 2602 1697
rect 2602 1663 2670 1697
rect 2670 1663 2704 1697
rect 2704 1663 2772 1697
rect 2772 1663 2776 1697
rect 2598 1629 2776 1663
rect 2598 1595 2602 1629
rect 2602 1595 2670 1629
rect 2670 1595 2704 1629
rect 2704 1595 2772 1629
rect 2772 1595 2776 1629
rect 2598 1561 2776 1595
rect 2598 1527 2602 1561
rect 2602 1527 2670 1561
rect 2670 1527 2704 1561
rect 2704 1527 2772 1561
rect 2772 1527 2776 1561
rect 2598 1491 2776 1527
rect 2598 1479 2632 1491
rect 2742 1479 2776 1491
rect 3345 4388 3451 4494
rect 3094 4028 3128 4062
rect 3166 4028 3200 4062
rect 3238 4028 3272 4062
rect 3094 3954 3128 3988
rect 3166 3954 3200 3988
rect 3238 3954 3272 3988
rect 3094 3880 3128 3914
rect 3166 3880 3200 3914
rect 3238 3880 3272 3914
rect 3094 3806 3128 3840
rect 3166 3806 3200 3840
rect 3238 3806 3272 3840
rect 3094 3732 3128 3766
rect 3166 3732 3200 3766
rect 3238 3732 3272 3766
rect 3094 3658 3128 3692
rect 3166 3658 3200 3692
rect 3238 3658 3272 3692
rect 3094 3584 3128 3618
rect 3166 3584 3200 3618
rect 3238 3584 3272 3618
rect 3094 3510 3128 3544
rect 3166 3510 3200 3544
rect 3238 3510 3272 3544
rect 3094 3436 3128 3470
rect 3166 3436 3200 3470
rect 3238 3436 3272 3470
rect 3094 3362 3128 3396
rect 3166 3362 3200 3396
rect 3238 3362 3272 3396
rect 3094 3288 3128 3322
rect 3166 3288 3200 3322
rect 3238 3288 3272 3322
rect 3094 3214 3128 3248
rect 3166 3214 3200 3248
rect 3238 3214 3272 3248
rect 3094 3140 3128 3174
rect 3166 3140 3200 3174
rect 3238 3140 3272 3174
rect 3094 3066 3128 3100
rect 3166 3066 3200 3100
rect 3238 3066 3272 3100
rect 3094 2992 3128 3026
rect 3166 2992 3200 3026
rect 3238 2992 3272 3026
rect 3094 2918 3128 2952
rect 3166 2918 3200 2952
rect 3238 2918 3272 2952
rect 3094 2844 3128 2878
rect 3166 2844 3200 2878
rect 3238 2844 3272 2878
rect 3094 2770 3128 2804
rect 3166 2770 3200 2804
rect 3238 2770 3272 2804
rect 3094 2696 3128 2730
rect 3166 2696 3200 2730
rect 3238 2696 3272 2730
rect 3094 2622 3128 2656
rect 3166 2622 3200 2656
rect 3238 2622 3272 2656
rect 3094 2548 3128 2582
rect 3166 2548 3200 2582
rect 3238 2548 3272 2582
rect 3094 2474 3128 2508
rect 3166 2474 3200 2508
rect 3238 2474 3272 2508
rect 3094 2400 3128 2434
rect 3166 2400 3200 2434
rect 3238 2400 3272 2434
rect 3094 2326 3128 2360
rect 3166 2326 3200 2360
rect 3238 2326 3272 2360
rect 3094 2252 3128 2286
rect 3166 2252 3200 2286
rect 3238 2252 3272 2286
rect 3094 2178 3128 2212
rect 3166 2178 3200 2212
rect 3238 2178 3272 2212
rect 3094 2104 3128 2138
rect 3166 2104 3200 2138
rect 3238 2104 3272 2138
rect 3094 2030 3128 2064
rect 3166 2030 3200 2064
rect 3238 2030 3272 2064
rect 3094 1956 3128 1990
rect 3166 1956 3200 1990
rect 3238 1956 3272 1990
rect 3094 1882 3128 1916
rect 3166 1882 3200 1916
rect 3238 1882 3272 1916
rect 3094 1808 3128 1842
rect 3166 1808 3200 1842
rect 3238 1808 3272 1842
rect 3094 1734 3128 1768
rect 3166 1734 3200 1768
rect 3238 1734 3272 1768
rect 3094 1660 3128 1694
rect 3166 1660 3200 1694
rect 3238 1660 3272 1694
rect 3094 1586 3128 1620
rect 3166 1586 3200 1620
rect 3238 1586 3272 1620
rect 3094 1511 3128 1545
rect 3166 1511 3200 1545
rect 3238 1511 3272 1545
rect 3907 4388 4013 4494
rect 3662 4050 3696 4062
rect 3590 4046 3768 4050
rect 3590 4012 3594 4046
rect 3594 4012 3662 4046
rect 3662 4012 3696 4046
rect 3696 4012 3764 4046
rect 3764 4012 3768 4046
rect 3590 3978 3768 4012
rect 3590 3944 3594 3978
rect 3594 3944 3662 3978
rect 3662 3944 3696 3978
rect 3696 3944 3764 3978
rect 3764 3944 3768 3978
rect 3590 3910 3768 3944
rect 3590 3876 3594 3910
rect 3594 3876 3662 3910
rect 3662 3876 3696 3910
rect 3696 3876 3764 3910
rect 3764 3876 3768 3910
rect 3590 3842 3768 3876
rect 3590 3808 3594 3842
rect 3594 3808 3662 3842
rect 3662 3808 3696 3842
rect 3696 3808 3764 3842
rect 3764 3808 3768 3842
rect 3590 3774 3768 3808
rect 3590 3740 3594 3774
rect 3594 3740 3662 3774
rect 3662 3740 3696 3774
rect 3696 3740 3764 3774
rect 3764 3740 3768 3774
rect 3590 3706 3768 3740
rect 3590 3672 3594 3706
rect 3594 3672 3662 3706
rect 3662 3672 3696 3706
rect 3696 3672 3764 3706
rect 3764 3672 3768 3706
rect 3590 3638 3768 3672
rect 3590 3604 3594 3638
rect 3594 3604 3662 3638
rect 3662 3604 3696 3638
rect 3696 3604 3764 3638
rect 3764 3604 3768 3638
rect 3590 3570 3768 3604
rect 3590 3536 3594 3570
rect 3594 3536 3662 3570
rect 3662 3536 3696 3570
rect 3696 3536 3764 3570
rect 3764 3536 3768 3570
rect 3590 3502 3768 3536
rect 3590 3468 3594 3502
rect 3594 3468 3662 3502
rect 3662 3468 3696 3502
rect 3696 3468 3764 3502
rect 3764 3468 3768 3502
rect 3590 3434 3768 3468
rect 3590 3400 3594 3434
rect 3594 3400 3662 3434
rect 3662 3400 3696 3434
rect 3696 3400 3764 3434
rect 3764 3400 3768 3434
rect 3590 3366 3768 3400
rect 3590 3332 3594 3366
rect 3594 3332 3662 3366
rect 3662 3332 3696 3366
rect 3696 3332 3764 3366
rect 3764 3332 3768 3366
rect 3590 3298 3768 3332
rect 3590 3264 3594 3298
rect 3594 3264 3662 3298
rect 3662 3264 3696 3298
rect 3696 3264 3764 3298
rect 3764 3264 3768 3298
rect 3590 3230 3768 3264
rect 3590 3196 3594 3230
rect 3594 3196 3662 3230
rect 3662 3196 3696 3230
rect 3696 3196 3764 3230
rect 3764 3196 3768 3230
rect 3590 3162 3768 3196
rect 3590 3128 3594 3162
rect 3594 3128 3662 3162
rect 3662 3128 3696 3162
rect 3696 3128 3764 3162
rect 3764 3128 3768 3162
rect 3590 3092 3768 3128
rect 3590 3080 3624 3092
rect 3734 3080 3768 3092
rect 3590 2935 3768 3040
rect 3590 2901 3629 2935
rect 3629 2901 3663 2935
rect 3663 2901 3697 2935
rect 3697 2901 3731 2935
rect 3731 2901 3768 2935
rect 3590 2855 3768 2901
rect 3590 2821 3629 2855
rect 3629 2821 3663 2855
rect 3663 2821 3697 2855
rect 3697 2821 3731 2855
rect 3731 2821 3768 2855
rect 3590 2775 3768 2821
rect 3590 2741 3629 2775
rect 3629 2741 3663 2775
rect 3663 2741 3697 2775
rect 3697 2741 3731 2775
rect 3731 2741 3768 2775
rect 3590 2695 3768 2741
rect 3590 2661 3629 2695
rect 3629 2661 3663 2695
rect 3663 2661 3697 2695
rect 3697 2661 3731 2695
rect 3731 2661 3768 2695
rect 3590 2614 3768 2661
rect 3590 2580 3629 2614
rect 3629 2580 3663 2614
rect 3663 2580 3697 2614
rect 3697 2580 3731 2614
rect 3731 2580 3768 2614
rect 3590 2574 3768 2580
rect 3590 2501 3624 2535
rect 3662 2501 3696 2535
rect 3734 2501 3768 2535
rect 3662 2449 3696 2461
rect 3590 2445 3768 2449
rect 3590 2411 3594 2445
rect 3594 2411 3662 2445
rect 3662 2411 3696 2445
rect 3696 2411 3764 2445
rect 3764 2411 3768 2445
rect 3590 2377 3768 2411
rect 3590 2343 3594 2377
rect 3594 2343 3662 2377
rect 3662 2343 3696 2377
rect 3696 2343 3764 2377
rect 3764 2343 3768 2377
rect 3590 2309 3768 2343
rect 3590 2275 3594 2309
rect 3594 2275 3662 2309
rect 3662 2275 3696 2309
rect 3696 2275 3764 2309
rect 3764 2275 3768 2309
rect 3590 2241 3768 2275
rect 3590 2207 3594 2241
rect 3594 2207 3662 2241
rect 3662 2207 3696 2241
rect 3696 2207 3764 2241
rect 3764 2207 3768 2241
rect 3590 2173 3768 2207
rect 3590 2139 3594 2173
rect 3594 2139 3662 2173
rect 3662 2139 3696 2173
rect 3696 2139 3764 2173
rect 3764 2139 3768 2173
rect 3590 2105 3768 2139
rect 3590 2071 3594 2105
rect 3594 2071 3662 2105
rect 3662 2071 3696 2105
rect 3696 2071 3764 2105
rect 3764 2071 3768 2105
rect 3590 2037 3768 2071
rect 3590 2003 3594 2037
rect 3594 2003 3662 2037
rect 3662 2003 3696 2037
rect 3696 2003 3764 2037
rect 3764 2003 3768 2037
rect 3590 1969 3768 2003
rect 3590 1935 3594 1969
rect 3594 1935 3662 1969
rect 3662 1935 3696 1969
rect 3696 1935 3764 1969
rect 3764 1935 3768 1969
rect 3590 1901 3768 1935
rect 3590 1867 3594 1901
rect 3594 1867 3662 1901
rect 3662 1867 3696 1901
rect 3696 1867 3764 1901
rect 3764 1867 3768 1901
rect 3590 1833 3768 1867
rect 3590 1799 3594 1833
rect 3594 1799 3662 1833
rect 3662 1799 3696 1833
rect 3696 1799 3764 1833
rect 3764 1799 3768 1833
rect 3590 1765 3768 1799
rect 3590 1731 3594 1765
rect 3594 1731 3662 1765
rect 3662 1731 3696 1765
rect 3696 1731 3764 1765
rect 3764 1731 3768 1765
rect 3590 1697 3768 1731
rect 3590 1663 3594 1697
rect 3594 1663 3662 1697
rect 3662 1663 3696 1697
rect 3696 1663 3764 1697
rect 3764 1663 3768 1697
rect 3590 1629 3768 1663
rect 3590 1595 3594 1629
rect 3594 1595 3662 1629
rect 3662 1595 3696 1629
rect 3696 1595 3764 1629
rect 3764 1595 3768 1629
rect 3590 1561 3768 1595
rect 3590 1527 3594 1561
rect 3594 1527 3662 1561
rect 3662 1527 3696 1561
rect 3696 1527 3764 1561
rect 3764 1527 3768 1561
rect 3590 1491 3768 1527
rect 3590 1479 3624 1491
rect 3734 1479 3768 1491
rect 4337 4388 4443 4494
rect 4086 4028 4120 4062
rect 4158 4028 4192 4062
rect 4230 4028 4264 4062
rect 4086 3954 4120 3988
rect 4158 3954 4192 3988
rect 4230 3954 4264 3988
rect 4086 3880 4120 3914
rect 4158 3880 4192 3914
rect 4230 3880 4264 3914
rect 4086 3806 4120 3840
rect 4158 3806 4192 3840
rect 4230 3806 4264 3840
rect 4086 3732 4120 3766
rect 4158 3732 4192 3766
rect 4230 3732 4264 3766
rect 4086 3658 4120 3692
rect 4158 3658 4192 3692
rect 4230 3658 4264 3692
rect 4086 3584 4120 3618
rect 4158 3584 4192 3618
rect 4230 3584 4264 3618
rect 4086 3510 4120 3544
rect 4158 3510 4192 3544
rect 4230 3510 4264 3544
rect 4086 3436 4120 3470
rect 4158 3436 4192 3470
rect 4230 3436 4264 3470
rect 4086 3362 4120 3396
rect 4158 3362 4192 3396
rect 4230 3362 4264 3396
rect 4086 3288 4120 3322
rect 4158 3288 4192 3322
rect 4230 3288 4264 3322
rect 4086 3214 4120 3248
rect 4158 3214 4192 3248
rect 4230 3214 4264 3248
rect 4086 3140 4120 3174
rect 4158 3140 4192 3174
rect 4230 3140 4264 3174
rect 4086 3066 4120 3100
rect 4158 3066 4192 3100
rect 4230 3066 4264 3100
rect 4086 2992 4120 3026
rect 4158 2992 4192 3026
rect 4230 2992 4264 3026
rect 4086 2918 4120 2952
rect 4158 2918 4192 2952
rect 4230 2918 4264 2952
rect 4086 2844 4120 2878
rect 4158 2844 4192 2878
rect 4230 2844 4264 2878
rect 4086 2770 4120 2804
rect 4158 2770 4192 2804
rect 4230 2770 4264 2804
rect 4086 2696 4120 2730
rect 4158 2696 4192 2730
rect 4230 2696 4264 2730
rect 4086 2622 4120 2656
rect 4158 2622 4192 2656
rect 4230 2622 4264 2656
rect 4086 2548 4120 2582
rect 4158 2548 4192 2582
rect 4230 2548 4264 2582
rect 4086 2474 4120 2508
rect 4158 2474 4192 2508
rect 4230 2474 4264 2508
rect 4086 2400 4120 2434
rect 4158 2400 4192 2434
rect 4230 2400 4264 2434
rect 4086 2326 4120 2360
rect 4158 2326 4192 2360
rect 4230 2326 4264 2360
rect 4086 2252 4120 2286
rect 4158 2252 4192 2286
rect 4230 2252 4264 2286
rect 4086 2178 4120 2212
rect 4158 2178 4192 2212
rect 4230 2178 4264 2212
rect 4086 2104 4120 2138
rect 4158 2104 4192 2138
rect 4230 2104 4264 2138
rect 4086 2030 4120 2064
rect 4158 2030 4192 2064
rect 4230 2030 4264 2064
rect 4086 1956 4120 1990
rect 4158 1956 4192 1990
rect 4230 1956 4264 1990
rect 4086 1882 4120 1916
rect 4158 1882 4192 1916
rect 4230 1882 4264 1916
rect 4086 1808 4120 1842
rect 4158 1808 4192 1842
rect 4230 1808 4264 1842
rect 4086 1734 4120 1768
rect 4158 1734 4192 1768
rect 4230 1734 4264 1768
rect 4086 1660 4120 1694
rect 4158 1660 4192 1694
rect 4230 1660 4264 1694
rect 4086 1586 4120 1620
rect 4158 1586 4192 1620
rect 4230 1586 4264 1620
rect 4086 1511 4120 1545
rect 4158 1511 4192 1545
rect 4230 1511 4264 1545
rect 4899 4388 5005 4494
rect 4654 4050 4688 4062
rect 4582 4046 4760 4050
rect 4582 4012 4586 4046
rect 4586 4012 4654 4046
rect 4654 4012 4688 4046
rect 4688 4012 4756 4046
rect 4756 4012 4760 4046
rect 4582 3978 4760 4012
rect 4582 3944 4586 3978
rect 4586 3944 4654 3978
rect 4654 3944 4688 3978
rect 4688 3944 4756 3978
rect 4756 3944 4760 3978
rect 4582 3910 4760 3944
rect 4582 3876 4586 3910
rect 4586 3876 4654 3910
rect 4654 3876 4688 3910
rect 4688 3876 4756 3910
rect 4756 3876 4760 3910
rect 4582 3842 4760 3876
rect 4582 3808 4586 3842
rect 4586 3808 4654 3842
rect 4654 3808 4688 3842
rect 4688 3808 4756 3842
rect 4756 3808 4760 3842
rect 4582 3774 4760 3808
rect 4582 3740 4586 3774
rect 4586 3740 4654 3774
rect 4654 3740 4688 3774
rect 4688 3740 4756 3774
rect 4756 3740 4760 3774
rect 4582 3706 4760 3740
rect 4582 3672 4586 3706
rect 4586 3672 4654 3706
rect 4654 3672 4688 3706
rect 4688 3672 4756 3706
rect 4756 3672 4760 3706
rect 4582 3638 4760 3672
rect 4582 3604 4586 3638
rect 4586 3604 4654 3638
rect 4654 3604 4688 3638
rect 4688 3604 4756 3638
rect 4756 3604 4760 3638
rect 4582 3570 4760 3604
rect 4582 3536 4586 3570
rect 4586 3536 4654 3570
rect 4654 3536 4688 3570
rect 4688 3536 4756 3570
rect 4756 3536 4760 3570
rect 4582 3502 4760 3536
rect 4582 3468 4586 3502
rect 4586 3468 4654 3502
rect 4654 3468 4688 3502
rect 4688 3468 4756 3502
rect 4756 3468 4760 3502
rect 4582 3434 4760 3468
rect 4582 3400 4586 3434
rect 4586 3400 4654 3434
rect 4654 3400 4688 3434
rect 4688 3400 4756 3434
rect 4756 3400 4760 3434
rect 4582 3366 4760 3400
rect 4582 3332 4586 3366
rect 4586 3332 4654 3366
rect 4654 3332 4688 3366
rect 4688 3332 4756 3366
rect 4756 3332 4760 3366
rect 4582 3298 4760 3332
rect 4582 3264 4586 3298
rect 4586 3264 4654 3298
rect 4654 3264 4688 3298
rect 4688 3264 4756 3298
rect 4756 3264 4760 3298
rect 4582 3230 4760 3264
rect 4582 3196 4586 3230
rect 4586 3196 4654 3230
rect 4654 3196 4688 3230
rect 4688 3196 4756 3230
rect 4756 3196 4760 3230
rect 4582 3162 4760 3196
rect 4582 3128 4586 3162
rect 4586 3128 4654 3162
rect 4654 3128 4688 3162
rect 4688 3128 4756 3162
rect 4756 3128 4760 3162
rect 4582 3092 4760 3128
rect 4582 3080 4616 3092
rect 4726 3080 4760 3092
rect 4582 2935 4760 3040
rect 4582 2901 4621 2935
rect 4621 2901 4655 2935
rect 4655 2901 4689 2935
rect 4689 2901 4723 2935
rect 4723 2901 4760 2935
rect 4582 2855 4760 2901
rect 4582 2821 4621 2855
rect 4621 2821 4655 2855
rect 4655 2821 4689 2855
rect 4689 2821 4723 2855
rect 4723 2821 4760 2855
rect 4582 2775 4760 2821
rect 4582 2741 4621 2775
rect 4621 2741 4655 2775
rect 4655 2741 4689 2775
rect 4689 2741 4723 2775
rect 4723 2741 4760 2775
rect 4582 2695 4760 2741
rect 4582 2661 4621 2695
rect 4621 2661 4655 2695
rect 4655 2661 4689 2695
rect 4689 2661 4723 2695
rect 4723 2661 4760 2695
rect 4582 2614 4760 2661
rect 4582 2580 4621 2614
rect 4621 2580 4655 2614
rect 4655 2580 4689 2614
rect 4689 2580 4723 2614
rect 4723 2580 4760 2614
rect 4582 2574 4760 2580
rect 4582 2501 4616 2535
rect 4654 2501 4688 2535
rect 4726 2501 4760 2535
rect 4654 2449 4688 2461
rect 4582 2445 4760 2449
rect 4582 2411 4586 2445
rect 4586 2411 4654 2445
rect 4654 2411 4688 2445
rect 4688 2411 4756 2445
rect 4756 2411 4760 2445
rect 4582 2377 4760 2411
rect 4582 2343 4586 2377
rect 4586 2343 4654 2377
rect 4654 2343 4688 2377
rect 4688 2343 4756 2377
rect 4756 2343 4760 2377
rect 4582 2309 4760 2343
rect 4582 2275 4586 2309
rect 4586 2275 4654 2309
rect 4654 2275 4688 2309
rect 4688 2275 4756 2309
rect 4756 2275 4760 2309
rect 4582 2241 4760 2275
rect 4582 2207 4586 2241
rect 4586 2207 4654 2241
rect 4654 2207 4688 2241
rect 4688 2207 4756 2241
rect 4756 2207 4760 2241
rect 4582 2173 4760 2207
rect 4582 2139 4586 2173
rect 4586 2139 4654 2173
rect 4654 2139 4688 2173
rect 4688 2139 4756 2173
rect 4756 2139 4760 2173
rect 4582 2105 4760 2139
rect 4582 2071 4586 2105
rect 4586 2071 4654 2105
rect 4654 2071 4688 2105
rect 4688 2071 4756 2105
rect 4756 2071 4760 2105
rect 4582 2037 4760 2071
rect 4582 2003 4586 2037
rect 4586 2003 4654 2037
rect 4654 2003 4688 2037
rect 4688 2003 4756 2037
rect 4756 2003 4760 2037
rect 4582 1969 4760 2003
rect 4582 1935 4586 1969
rect 4586 1935 4654 1969
rect 4654 1935 4688 1969
rect 4688 1935 4756 1969
rect 4756 1935 4760 1969
rect 4582 1901 4760 1935
rect 4582 1867 4586 1901
rect 4586 1867 4654 1901
rect 4654 1867 4688 1901
rect 4688 1867 4756 1901
rect 4756 1867 4760 1901
rect 4582 1833 4760 1867
rect 4582 1799 4586 1833
rect 4586 1799 4654 1833
rect 4654 1799 4688 1833
rect 4688 1799 4756 1833
rect 4756 1799 4760 1833
rect 4582 1765 4760 1799
rect 4582 1731 4586 1765
rect 4586 1731 4654 1765
rect 4654 1731 4688 1765
rect 4688 1731 4756 1765
rect 4756 1731 4760 1765
rect 4582 1697 4760 1731
rect 4582 1663 4586 1697
rect 4586 1663 4654 1697
rect 4654 1663 4688 1697
rect 4688 1663 4756 1697
rect 4756 1663 4760 1697
rect 4582 1629 4760 1663
rect 4582 1595 4586 1629
rect 4586 1595 4654 1629
rect 4654 1595 4688 1629
rect 4688 1595 4756 1629
rect 4756 1595 4760 1629
rect 4582 1561 4760 1595
rect 4582 1527 4586 1561
rect 4586 1527 4654 1561
rect 4654 1527 4688 1561
rect 4688 1527 4756 1561
rect 4756 1527 4760 1561
rect 4582 1491 4760 1527
rect 4582 1479 4616 1491
rect 4726 1479 4760 1491
rect 5329 4388 5435 4494
rect 5078 4028 5112 4062
rect 5150 4028 5184 4062
rect 5222 4028 5256 4062
rect 5078 3954 5112 3988
rect 5150 3954 5184 3988
rect 5222 3954 5256 3988
rect 5078 3880 5112 3914
rect 5150 3880 5184 3914
rect 5222 3880 5256 3914
rect 5078 3806 5112 3840
rect 5150 3806 5184 3840
rect 5222 3806 5256 3840
rect 5078 3732 5112 3766
rect 5150 3732 5184 3766
rect 5222 3732 5256 3766
rect 5078 3658 5112 3692
rect 5150 3658 5184 3692
rect 5222 3658 5256 3692
rect 5078 3584 5112 3618
rect 5150 3584 5184 3618
rect 5222 3584 5256 3618
rect 5078 3510 5112 3544
rect 5150 3510 5184 3544
rect 5222 3510 5256 3544
rect 5078 3436 5112 3470
rect 5150 3436 5184 3470
rect 5222 3436 5256 3470
rect 5078 3362 5112 3396
rect 5150 3362 5184 3396
rect 5222 3362 5256 3396
rect 5078 3288 5112 3322
rect 5150 3288 5184 3322
rect 5222 3288 5256 3322
rect 5078 3214 5112 3248
rect 5150 3214 5184 3248
rect 5222 3214 5256 3248
rect 5078 3140 5112 3174
rect 5150 3140 5184 3174
rect 5222 3140 5256 3174
rect 5078 3066 5112 3100
rect 5150 3066 5184 3100
rect 5222 3066 5256 3100
rect 5078 2992 5112 3026
rect 5150 2992 5184 3026
rect 5222 2992 5256 3026
rect 5078 2918 5112 2952
rect 5150 2918 5184 2952
rect 5222 2918 5256 2952
rect 5078 2844 5112 2878
rect 5150 2844 5184 2878
rect 5222 2844 5256 2878
rect 5078 2770 5112 2804
rect 5150 2770 5184 2804
rect 5222 2770 5256 2804
rect 5078 2696 5112 2730
rect 5150 2696 5184 2730
rect 5222 2696 5256 2730
rect 5078 2622 5112 2656
rect 5150 2622 5184 2656
rect 5222 2622 5256 2656
rect 5078 2548 5112 2582
rect 5150 2548 5184 2582
rect 5222 2548 5256 2582
rect 5078 2474 5112 2508
rect 5150 2474 5184 2508
rect 5222 2474 5256 2508
rect 5078 2400 5112 2434
rect 5150 2400 5184 2434
rect 5222 2400 5256 2434
rect 5078 2326 5112 2360
rect 5150 2326 5184 2360
rect 5222 2326 5256 2360
rect 5078 2252 5112 2286
rect 5150 2252 5184 2286
rect 5222 2252 5256 2286
rect 5078 2178 5112 2212
rect 5150 2178 5184 2212
rect 5222 2178 5256 2212
rect 5078 2104 5112 2138
rect 5150 2104 5184 2138
rect 5222 2104 5256 2138
rect 5078 2030 5112 2064
rect 5150 2030 5184 2064
rect 5222 2030 5256 2064
rect 5078 1956 5112 1990
rect 5150 1956 5184 1990
rect 5222 1956 5256 1990
rect 5078 1882 5112 1916
rect 5150 1882 5184 1916
rect 5222 1882 5256 1916
rect 5078 1808 5112 1842
rect 5150 1808 5184 1842
rect 5222 1808 5256 1842
rect 5078 1734 5112 1768
rect 5150 1734 5184 1768
rect 5222 1734 5256 1768
rect 5078 1660 5112 1694
rect 5150 1660 5184 1694
rect 5222 1660 5256 1694
rect 5078 1586 5112 1620
rect 5150 1586 5184 1620
rect 5222 1586 5256 1620
rect 5078 1511 5112 1545
rect 5150 1511 5184 1545
rect 5222 1511 5256 1545
rect 5891 4388 5997 4494
rect 5646 4050 5680 4062
rect 5574 4046 5752 4050
rect 5574 4012 5578 4046
rect 5578 4012 5646 4046
rect 5646 4012 5680 4046
rect 5680 4012 5748 4046
rect 5748 4012 5752 4046
rect 5574 3978 5752 4012
rect 5574 3944 5578 3978
rect 5578 3944 5646 3978
rect 5646 3944 5680 3978
rect 5680 3944 5748 3978
rect 5748 3944 5752 3978
rect 5574 3910 5752 3944
rect 5574 3876 5578 3910
rect 5578 3876 5646 3910
rect 5646 3876 5680 3910
rect 5680 3876 5748 3910
rect 5748 3876 5752 3910
rect 5574 3842 5752 3876
rect 5574 3808 5578 3842
rect 5578 3808 5646 3842
rect 5646 3808 5680 3842
rect 5680 3808 5748 3842
rect 5748 3808 5752 3842
rect 5574 3774 5752 3808
rect 5574 3740 5578 3774
rect 5578 3740 5646 3774
rect 5646 3740 5680 3774
rect 5680 3740 5748 3774
rect 5748 3740 5752 3774
rect 5574 3706 5752 3740
rect 5574 3672 5578 3706
rect 5578 3672 5646 3706
rect 5646 3672 5680 3706
rect 5680 3672 5748 3706
rect 5748 3672 5752 3706
rect 5574 3638 5752 3672
rect 5574 3604 5578 3638
rect 5578 3604 5646 3638
rect 5646 3604 5680 3638
rect 5680 3604 5748 3638
rect 5748 3604 5752 3638
rect 5574 3570 5752 3604
rect 5574 3536 5578 3570
rect 5578 3536 5646 3570
rect 5646 3536 5680 3570
rect 5680 3536 5748 3570
rect 5748 3536 5752 3570
rect 5574 3502 5752 3536
rect 5574 3468 5578 3502
rect 5578 3468 5646 3502
rect 5646 3468 5680 3502
rect 5680 3468 5748 3502
rect 5748 3468 5752 3502
rect 5574 3434 5752 3468
rect 5574 3400 5578 3434
rect 5578 3400 5646 3434
rect 5646 3400 5680 3434
rect 5680 3400 5748 3434
rect 5748 3400 5752 3434
rect 5574 3366 5752 3400
rect 5574 3332 5578 3366
rect 5578 3332 5646 3366
rect 5646 3332 5680 3366
rect 5680 3332 5748 3366
rect 5748 3332 5752 3366
rect 5574 3298 5752 3332
rect 5574 3264 5578 3298
rect 5578 3264 5646 3298
rect 5646 3264 5680 3298
rect 5680 3264 5748 3298
rect 5748 3264 5752 3298
rect 5574 3230 5752 3264
rect 5574 3196 5578 3230
rect 5578 3196 5646 3230
rect 5646 3196 5680 3230
rect 5680 3196 5748 3230
rect 5748 3196 5752 3230
rect 5574 3162 5752 3196
rect 5574 3128 5578 3162
rect 5578 3128 5646 3162
rect 5646 3128 5680 3162
rect 5680 3128 5748 3162
rect 5748 3128 5752 3162
rect 5574 3092 5752 3128
rect 5574 3080 5608 3092
rect 5718 3080 5752 3092
rect 5574 2935 5752 3040
rect 5574 2901 5613 2935
rect 5613 2901 5647 2935
rect 5647 2901 5681 2935
rect 5681 2901 5715 2935
rect 5715 2901 5752 2935
rect 5574 2855 5752 2901
rect 5574 2821 5613 2855
rect 5613 2821 5647 2855
rect 5647 2821 5681 2855
rect 5681 2821 5715 2855
rect 5715 2821 5752 2855
rect 5574 2775 5752 2821
rect 5574 2741 5613 2775
rect 5613 2741 5647 2775
rect 5647 2741 5681 2775
rect 5681 2741 5715 2775
rect 5715 2741 5752 2775
rect 5574 2695 5752 2741
rect 5574 2661 5613 2695
rect 5613 2661 5647 2695
rect 5647 2661 5681 2695
rect 5681 2661 5715 2695
rect 5715 2661 5752 2695
rect 5574 2614 5752 2661
rect 5574 2580 5613 2614
rect 5613 2580 5647 2614
rect 5647 2580 5681 2614
rect 5681 2580 5715 2614
rect 5715 2580 5752 2614
rect 5574 2574 5752 2580
rect 5574 2501 5608 2535
rect 5646 2501 5680 2535
rect 5718 2501 5752 2535
rect 5646 2449 5680 2461
rect 5574 2445 5752 2449
rect 5574 2411 5578 2445
rect 5578 2411 5646 2445
rect 5646 2411 5680 2445
rect 5680 2411 5748 2445
rect 5748 2411 5752 2445
rect 5574 2377 5752 2411
rect 5574 2343 5578 2377
rect 5578 2343 5646 2377
rect 5646 2343 5680 2377
rect 5680 2343 5748 2377
rect 5748 2343 5752 2377
rect 5574 2309 5752 2343
rect 5574 2275 5578 2309
rect 5578 2275 5646 2309
rect 5646 2275 5680 2309
rect 5680 2275 5748 2309
rect 5748 2275 5752 2309
rect 5574 2241 5752 2275
rect 5574 2207 5578 2241
rect 5578 2207 5646 2241
rect 5646 2207 5680 2241
rect 5680 2207 5748 2241
rect 5748 2207 5752 2241
rect 5574 2173 5752 2207
rect 5574 2139 5578 2173
rect 5578 2139 5646 2173
rect 5646 2139 5680 2173
rect 5680 2139 5748 2173
rect 5748 2139 5752 2173
rect 5574 2105 5752 2139
rect 5574 2071 5578 2105
rect 5578 2071 5646 2105
rect 5646 2071 5680 2105
rect 5680 2071 5748 2105
rect 5748 2071 5752 2105
rect 5574 2037 5752 2071
rect 5574 2003 5578 2037
rect 5578 2003 5646 2037
rect 5646 2003 5680 2037
rect 5680 2003 5748 2037
rect 5748 2003 5752 2037
rect 5574 1969 5752 2003
rect 5574 1935 5578 1969
rect 5578 1935 5646 1969
rect 5646 1935 5680 1969
rect 5680 1935 5748 1969
rect 5748 1935 5752 1969
rect 5574 1901 5752 1935
rect 5574 1867 5578 1901
rect 5578 1867 5646 1901
rect 5646 1867 5680 1901
rect 5680 1867 5748 1901
rect 5748 1867 5752 1901
rect 5574 1833 5752 1867
rect 5574 1799 5578 1833
rect 5578 1799 5646 1833
rect 5646 1799 5680 1833
rect 5680 1799 5748 1833
rect 5748 1799 5752 1833
rect 5574 1765 5752 1799
rect 5574 1731 5578 1765
rect 5578 1731 5646 1765
rect 5646 1731 5680 1765
rect 5680 1731 5748 1765
rect 5748 1731 5752 1765
rect 5574 1697 5752 1731
rect 5574 1663 5578 1697
rect 5578 1663 5646 1697
rect 5646 1663 5680 1697
rect 5680 1663 5748 1697
rect 5748 1663 5752 1697
rect 5574 1629 5752 1663
rect 5574 1595 5578 1629
rect 5578 1595 5646 1629
rect 5646 1595 5680 1629
rect 5680 1595 5748 1629
rect 5748 1595 5752 1629
rect 5574 1561 5752 1595
rect 5574 1527 5578 1561
rect 5578 1527 5646 1561
rect 5646 1527 5680 1561
rect 5680 1527 5748 1561
rect 5748 1527 5752 1561
rect 5574 1491 5752 1527
rect 5574 1479 5608 1491
rect 5718 1479 5752 1491
rect 6321 4388 6427 4494
rect 6868 4388 6974 4494
rect 6070 4028 6104 4062
rect 6142 4028 6176 4062
rect 6214 4028 6248 4062
rect 6070 3954 6104 3988
rect 6142 3954 6176 3988
rect 6214 3954 6248 3988
rect 6070 3880 6104 3914
rect 6142 3880 6176 3914
rect 6214 3880 6248 3914
rect 6070 3806 6104 3840
rect 6142 3806 6176 3840
rect 6214 3806 6248 3840
rect 6070 3732 6104 3766
rect 6142 3732 6176 3766
rect 6214 3732 6248 3766
rect 6070 3658 6104 3692
rect 6142 3658 6176 3692
rect 6214 3658 6248 3692
rect 6070 3584 6104 3618
rect 6142 3584 6176 3618
rect 6214 3584 6248 3618
rect 6070 3510 6104 3544
rect 6142 3510 6176 3544
rect 6214 3510 6248 3544
rect 6070 3436 6104 3470
rect 6142 3436 6176 3470
rect 6214 3436 6248 3470
rect 6070 3362 6104 3396
rect 6142 3362 6176 3396
rect 6214 3362 6248 3396
rect 6070 3288 6104 3322
rect 6142 3288 6176 3322
rect 6214 3288 6248 3322
rect 6070 3214 6104 3248
rect 6142 3214 6176 3248
rect 6214 3214 6248 3248
rect 6070 3140 6104 3174
rect 6142 3140 6176 3174
rect 6214 3140 6248 3174
rect 6070 3066 6104 3100
rect 6142 3066 6176 3100
rect 6214 3066 6248 3100
rect 6070 2992 6104 3026
rect 6142 2992 6176 3026
rect 6214 2992 6248 3026
rect 6070 2918 6104 2952
rect 6142 2918 6176 2952
rect 6214 2918 6248 2952
rect 6070 2844 6104 2878
rect 6142 2844 6176 2878
rect 6214 2844 6248 2878
rect 6070 2770 6104 2804
rect 6142 2770 6176 2804
rect 6214 2770 6248 2804
rect 6070 2696 6104 2730
rect 6142 2696 6176 2730
rect 6214 2696 6248 2730
rect 6070 2622 6104 2656
rect 6142 2622 6176 2656
rect 6214 2622 6248 2656
rect 6070 2548 6104 2582
rect 6142 2548 6176 2582
rect 6214 2548 6248 2582
rect 6070 2474 6104 2508
rect 6142 2474 6176 2508
rect 6214 2474 6248 2508
rect 6070 2400 6104 2434
rect 6142 2400 6176 2434
rect 6214 2400 6248 2434
rect 6070 2326 6104 2360
rect 6142 2326 6176 2360
rect 6214 2326 6248 2360
rect 6070 2252 6104 2286
rect 6142 2252 6176 2286
rect 6214 2252 6248 2286
rect 6070 2178 6104 2212
rect 6142 2178 6176 2212
rect 6214 2178 6248 2212
rect 6070 2104 6104 2138
rect 6142 2104 6176 2138
rect 6214 2104 6248 2138
rect 6070 2030 6104 2064
rect 6142 2030 6176 2064
rect 6214 2030 6248 2064
rect 6070 1956 6104 1990
rect 6142 1956 6176 1990
rect 6214 1956 6248 1990
rect 6070 1882 6104 1916
rect 6142 1882 6176 1916
rect 6214 1882 6248 1916
rect 6070 1808 6104 1842
rect 6142 1808 6176 1842
rect 6214 1808 6248 1842
rect 6070 1734 6104 1768
rect 6142 1734 6176 1768
rect 6214 1734 6248 1768
rect 6070 1660 6104 1694
rect 6142 1660 6176 1694
rect 6214 1660 6248 1694
rect 6070 1586 6104 1620
rect 6142 1586 6176 1620
rect 6214 1586 6248 1620
rect 6070 1511 6104 1545
rect 6142 1511 6176 1545
rect 6214 1511 6248 1545
rect 6638 4050 6672 4062
rect 6566 4046 6744 4050
rect 6566 4012 6570 4046
rect 6570 4012 6638 4046
rect 6638 4012 6672 4046
rect 6672 4012 6740 4046
rect 6740 4012 6744 4046
rect 6566 3978 6744 4012
rect 6566 3944 6570 3978
rect 6570 3944 6638 3978
rect 6638 3944 6672 3978
rect 6672 3944 6740 3978
rect 6740 3944 6744 3978
rect 6566 3910 6744 3944
rect 6566 3876 6570 3910
rect 6570 3876 6638 3910
rect 6638 3876 6672 3910
rect 6672 3876 6740 3910
rect 6740 3876 6744 3910
rect 6566 3842 6744 3876
rect 6566 3808 6570 3842
rect 6570 3808 6638 3842
rect 6638 3808 6672 3842
rect 6672 3808 6740 3842
rect 6740 3808 6744 3842
rect 6566 3774 6744 3808
rect 6566 3740 6570 3774
rect 6570 3740 6638 3774
rect 6638 3740 6672 3774
rect 6672 3740 6740 3774
rect 6740 3740 6744 3774
rect 6566 3706 6744 3740
rect 6566 3672 6570 3706
rect 6570 3672 6638 3706
rect 6638 3672 6672 3706
rect 6672 3672 6740 3706
rect 6740 3672 6744 3706
rect 6566 3638 6744 3672
rect 6566 3604 6570 3638
rect 6570 3604 6638 3638
rect 6638 3604 6672 3638
rect 6672 3604 6740 3638
rect 6740 3604 6744 3638
rect 6566 3570 6744 3604
rect 6566 3536 6570 3570
rect 6570 3536 6638 3570
rect 6638 3536 6672 3570
rect 6672 3536 6740 3570
rect 6740 3536 6744 3570
rect 6566 3502 6744 3536
rect 6566 3468 6570 3502
rect 6570 3468 6638 3502
rect 6638 3468 6672 3502
rect 6672 3468 6740 3502
rect 6740 3468 6744 3502
rect 6566 3434 6744 3468
rect 6566 3400 6570 3434
rect 6570 3400 6638 3434
rect 6638 3400 6672 3434
rect 6672 3400 6740 3434
rect 6740 3400 6744 3434
rect 6566 3366 6744 3400
rect 6566 3332 6570 3366
rect 6570 3332 6638 3366
rect 6638 3332 6672 3366
rect 6672 3332 6740 3366
rect 6740 3332 6744 3366
rect 6566 3298 6744 3332
rect 6566 3264 6570 3298
rect 6570 3264 6638 3298
rect 6638 3264 6672 3298
rect 6672 3264 6740 3298
rect 6740 3264 6744 3298
rect 6566 3230 6744 3264
rect 6566 3196 6570 3230
rect 6570 3196 6638 3230
rect 6638 3196 6672 3230
rect 6672 3196 6740 3230
rect 6740 3196 6744 3230
rect 6566 3162 6744 3196
rect 6566 3128 6570 3162
rect 6570 3128 6638 3162
rect 6638 3128 6672 3162
rect 6672 3128 6740 3162
rect 6740 3128 6744 3162
rect 6566 3092 6744 3128
rect 6566 3080 6600 3092
rect 6710 3080 6744 3092
rect 6566 2935 6744 3040
rect 6566 2901 6605 2935
rect 6605 2901 6639 2935
rect 6639 2901 6673 2935
rect 6673 2901 6707 2935
rect 6707 2901 6744 2935
rect 6566 2855 6744 2901
rect 6566 2821 6605 2855
rect 6605 2821 6639 2855
rect 6639 2821 6673 2855
rect 6673 2821 6707 2855
rect 6707 2821 6744 2855
rect 6566 2775 6744 2821
rect 6566 2741 6605 2775
rect 6605 2741 6639 2775
rect 6639 2741 6673 2775
rect 6673 2741 6707 2775
rect 6707 2741 6744 2775
rect 6566 2695 6744 2741
rect 6566 2661 6605 2695
rect 6605 2661 6639 2695
rect 6639 2661 6673 2695
rect 6673 2661 6707 2695
rect 6707 2661 6744 2695
rect 6566 2614 6744 2661
rect 6566 2580 6605 2614
rect 6605 2580 6639 2614
rect 6639 2580 6673 2614
rect 6673 2580 6707 2614
rect 6707 2580 6744 2614
rect 6566 2574 6744 2580
rect 6566 2501 6600 2535
rect 6638 2501 6672 2535
rect 6710 2501 6744 2535
rect 6638 2449 6672 2461
rect 6566 2445 6744 2449
rect 6566 2411 6570 2445
rect 6570 2411 6638 2445
rect 6638 2411 6672 2445
rect 6672 2411 6740 2445
rect 6740 2411 6744 2445
rect 6566 2377 6744 2411
rect 6566 2343 6570 2377
rect 6570 2343 6638 2377
rect 6638 2343 6672 2377
rect 6672 2343 6740 2377
rect 6740 2343 6744 2377
rect 6566 2309 6744 2343
rect 6566 2275 6570 2309
rect 6570 2275 6638 2309
rect 6638 2275 6672 2309
rect 6672 2275 6740 2309
rect 6740 2275 6744 2309
rect 6566 2241 6744 2275
rect 6566 2207 6570 2241
rect 6570 2207 6638 2241
rect 6638 2207 6672 2241
rect 6672 2207 6740 2241
rect 6740 2207 6744 2241
rect 6566 2173 6744 2207
rect 6566 2139 6570 2173
rect 6570 2139 6638 2173
rect 6638 2139 6672 2173
rect 6672 2139 6740 2173
rect 6740 2139 6744 2173
rect 6566 2105 6744 2139
rect 6566 2071 6570 2105
rect 6570 2071 6638 2105
rect 6638 2071 6672 2105
rect 6672 2071 6740 2105
rect 6740 2071 6744 2105
rect 6566 2037 6744 2071
rect 6566 2003 6570 2037
rect 6570 2003 6638 2037
rect 6638 2003 6672 2037
rect 6672 2003 6740 2037
rect 6740 2003 6744 2037
rect 6566 1969 6744 2003
rect 6566 1935 6570 1969
rect 6570 1935 6638 1969
rect 6638 1935 6672 1969
rect 6672 1935 6740 1969
rect 6740 1935 6744 1969
rect 6566 1901 6744 1935
rect 6566 1867 6570 1901
rect 6570 1867 6638 1901
rect 6638 1867 6672 1901
rect 6672 1867 6740 1901
rect 6740 1867 6744 1901
rect 6566 1833 6744 1867
rect 6566 1799 6570 1833
rect 6570 1799 6638 1833
rect 6638 1799 6672 1833
rect 6672 1799 6740 1833
rect 6740 1799 6744 1833
rect 6566 1765 6744 1799
rect 6566 1731 6570 1765
rect 6570 1731 6638 1765
rect 6638 1731 6672 1765
rect 6672 1731 6740 1765
rect 6740 1731 6744 1765
rect 6566 1697 6744 1731
rect 6566 1663 6570 1697
rect 6570 1663 6638 1697
rect 6638 1663 6672 1697
rect 6672 1663 6740 1697
rect 6740 1663 6744 1697
rect 6566 1629 6744 1663
rect 6566 1595 6570 1629
rect 6570 1595 6638 1629
rect 6638 1595 6672 1629
rect 6672 1595 6740 1629
rect 6740 1595 6744 1629
rect 6566 1561 6744 1595
rect 6566 1527 6570 1561
rect 6570 1527 6638 1561
rect 6638 1527 6672 1561
rect 6672 1527 6740 1561
rect 6740 1527 6744 1561
rect 6566 1491 6744 1527
rect 6566 1479 6600 1491
rect 6710 1479 6744 1491
rect 7313 4388 7419 4494
rect 7062 4028 7096 4062
rect 7134 4028 7168 4062
rect 7206 4028 7240 4062
rect 7062 3954 7096 3988
rect 7134 3954 7168 3988
rect 7206 3954 7240 3988
rect 7062 3880 7096 3914
rect 7134 3880 7168 3914
rect 7206 3880 7240 3914
rect 7062 3806 7096 3840
rect 7134 3806 7168 3840
rect 7206 3806 7240 3840
rect 7062 3732 7096 3766
rect 7134 3732 7168 3766
rect 7206 3732 7240 3766
rect 7062 3658 7096 3692
rect 7134 3658 7168 3692
rect 7206 3658 7240 3692
rect 7062 3584 7096 3618
rect 7134 3584 7168 3618
rect 7206 3584 7240 3618
rect 7062 3510 7096 3544
rect 7134 3510 7168 3544
rect 7206 3510 7240 3544
rect 7062 3436 7096 3470
rect 7134 3436 7168 3470
rect 7206 3436 7240 3470
rect 7062 3362 7096 3396
rect 7134 3362 7168 3396
rect 7206 3362 7240 3396
rect 7062 3288 7096 3322
rect 7134 3288 7168 3322
rect 7206 3288 7240 3322
rect 7062 3214 7096 3248
rect 7134 3214 7168 3248
rect 7206 3214 7240 3248
rect 7062 3140 7096 3174
rect 7134 3140 7168 3174
rect 7206 3140 7240 3174
rect 7062 3066 7096 3100
rect 7134 3066 7168 3100
rect 7206 3066 7240 3100
rect 7062 2992 7096 3026
rect 7134 2992 7168 3026
rect 7206 2992 7240 3026
rect 7062 2918 7096 2952
rect 7134 2918 7168 2952
rect 7206 2918 7240 2952
rect 7062 2844 7096 2878
rect 7134 2844 7168 2878
rect 7206 2844 7240 2878
rect 7062 2770 7096 2804
rect 7134 2770 7168 2804
rect 7206 2770 7240 2804
rect 7062 2696 7096 2730
rect 7134 2696 7168 2730
rect 7206 2696 7240 2730
rect 7062 2622 7096 2656
rect 7134 2622 7168 2656
rect 7206 2622 7240 2656
rect 7062 2548 7096 2582
rect 7134 2548 7168 2582
rect 7206 2548 7240 2582
rect 7062 2474 7096 2508
rect 7134 2474 7168 2508
rect 7206 2474 7240 2508
rect 7062 2400 7096 2434
rect 7134 2400 7168 2434
rect 7206 2400 7240 2434
rect 7062 2326 7096 2360
rect 7134 2326 7168 2360
rect 7206 2326 7240 2360
rect 7062 2252 7096 2286
rect 7134 2252 7168 2286
rect 7206 2252 7240 2286
rect 7062 2178 7096 2212
rect 7134 2178 7168 2212
rect 7206 2178 7240 2212
rect 7062 2104 7096 2138
rect 7134 2104 7168 2138
rect 7206 2104 7240 2138
rect 7062 2030 7096 2064
rect 7134 2030 7168 2064
rect 7206 2030 7240 2064
rect 7062 1956 7096 1990
rect 7134 1956 7168 1990
rect 7206 1956 7240 1990
rect 7062 1882 7096 1916
rect 7134 1882 7168 1916
rect 7206 1882 7240 1916
rect 7062 1808 7096 1842
rect 7134 1808 7168 1842
rect 7206 1808 7240 1842
rect 7062 1734 7096 1768
rect 7134 1734 7168 1768
rect 7206 1734 7240 1768
rect 7062 1660 7096 1694
rect 7134 1660 7168 1694
rect 7206 1660 7240 1694
rect 7062 1586 7096 1620
rect 7134 1586 7168 1620
rect 7206 1586 7240 1620
rect 7062 1511 7096 1545
rect 7134 1511 7168 1545
rect 7206 1511 7240 1545
rect 7875 4388 7981 4494
rect 7630 4050 7664 4062
rect 7558 4046 7736 4050
rect 7558 4012 7562 4046
rect 7562 4012 7630 4046
rect 7630 4012 7664 4046
rect 7664 4012 7732 4046
rect 7732 4012 7736 4046
rect 7558 3978 7736 4012
rect 7558 3944 7562 3978
rect 7562 3944 7630 3978
rect 7630 3944 7664 3978
rect 7664 3944 7732 3978
rect 7732 3944 7736 3978
rect 7558 3910 7736 3944
rect 7558 3876 7562 3910
rect 7562 3876 7630 3910
rect 7630 3876 7664 3910
rect 7664 3876 7732 3910
rect 7732 3876 7736 3910
rect 7558 3842 7736 3876
rect 7558 3808 7562 3842
rect 7562 3808 7630 3842
rect 7630 3808 7664 3842
rect 7664 3808 7732 3842
rect 7732 3808 7736 3842
rect 7558 3774 7736 3808
rect 7558 3740 7562 3774
rect 7562 3740 7630 3774
rect 7630 3740 7664 3774
rect 7664 3740 7732 3774
rect 7732 3740 7736 3774
rect 7558 3706 7736 3740
rect 7558 3672 7562 3706
rect 7562 3672 7630 3706
rect 7630 3672 7664 3706
rect 7664 3672 7732 3706
rect 7732 3672 7736 3706
rect 7558 3638 7736 3672
rect 7558 3604 7562 3638
rect 7562 3604 7630 3638
rect 7630 3604 7664 3638
rect 7664 3604 7732 3638
rect 7732 3604 7736 3638
rect 7558 3570 7736 3604
rect 7558 3536 7562 3570
rect 7562 3536 7630 3570
rect 7630 3536 7664 3570
rect 7664 3536 7732 3570
rect 7732 3536 7736 3570
rect 7558 3502 7736 3536
rect 7558 3468 7562 3502
rect 7562 3468 7630 3502
rect 7630 3468 7664 3502
rect 7664 3468 7732 3502
rect 7732 3468 7736 3502
rect 7558 3434 7736 3468
rect 7558 3400 7562 3434
rect 7562 3400 7630 3434
rect 7630 3400 7664 3434
rect 7664 3400 7732 3434
rect 7732 3400 7736 3434
rect 7558 3366 7736 3400
rect 7558 3332 7562 3366
rect 7562 3332 7630 3366
rect 7630 3332 7664 3366
rect 7664 3332 7732 3366
rect 7732 3332 7736 3366
rect 7558 3298 7736 3332
rect 7558 3264 7562 3298
rect 7562 3264 7630 3298
rect 7630 3264 7664 3298
rect 7664 3264 7732 3298
rect 7732 3264 7736 3298
rect 7558 3230 7736 3264
rect 7558 3196 7562 3230
rect 7562 3196 7630 3230
rect 7630 3196 7664 3230
rect 7664 3196 7732 3230
rect 7732 3196 7736 3230
rect 7558 3162 7736 3196
rect 7558 3128 7562 3162
rect 7562 3128 7630 3162
rect 7630 3128 7664 3162
rect 7664 3128 7732 3162
rect 7732 3128 7736 3162
rect 7558 3092 7736 3128
rect 7558 3080 7592 3092
rect 7702 3080 7736 3092
rect 7558 2935 7736 3040
rect 7558 2901 7597 2935
rect 7597 2901 7631 2935
rect 7631 2901 7665 2935
rect 7665 2901 7699 2935
rect 7699 2901 7736 2935
rect 7558 2855 7736 2901
rect 7558 2821 7597 2855
rect 7597 2821 7631 2855
rect 7631 2821 7665 2855
rect 7665 2821 7699 2855
rect 7699 2821 7736 2855
rect 7558 2775 7736 2821
rect 7558 2741 7597 2775
rect 7597 2741 7631 2775
rect 7631 2741 7665 2775
rect 7665 2741 7699 2775
rect 7699 2741 7736 2775
rect 7558 2695 7736 2741
rect 7558 2661 7597 2695
rect 7597 2661 7631 2695
rect 7631 2661 7665 2695
rect 7665 2661 7699 2695
rect 7699 2661 7736 2695
rect 7558 2614 7736 2661
rect 7558 2580 7597 2614
rect 7597 2580 7631 2614
rect 7631 2580 7665 2614
rect 7665 2580 7699 2614
rect 7699 2580 7736 2614
rect 7558 2574 7736 2580
rect 7558 2501 7592 2535
rect 7630 2501 7664 2535
rect 7702 2501 7736 2535
rect 7630 2449 7664 2461
rect 7558 2445 7736 2449
rect 7558 2411 7562 2445
rect 7562 2411 7630 2445
rect 7630 2411 7664 2445
rect 7664 2411 7732 2445
rect 7732 2411 7736 2445
rect 7558 2377 7736 2411
rect 7558 2343 7562 2377
rect 7562 2343 7630 2377
rect 7630 2343 7664 2377
rect 7664 2343 7732 2377
rect 7732 2343 7736 2377
rect 7558 2309 7736 2343
rect 7558 2275 7562 2309
rect 7562 2275 7630 2309
rect 7630 2275 7664 2309
rect 7664 2275 7732 2309
rect 7732 2275 7736 2309
rect 7558 2241 7736 2275
rect 7558 2207 7562 2241
rect 7562 2207 7630 2241
rect 7630 2207 7664 2241
rect 7664 2207 7732 2241
rect 7732 2207 7736 2241
rect 7558 2173 7736 2207
rect 7558 2139 7562 2173
rect 7562 2139 7630 2173
rect 7630 2139 7664 2173
rect 7664 2139 7732 2173
rect 7732 2139 7736 2173
rect 7558 2105 7736 2139
rect 7558 2071 7562 2105
rect 7562 2071 7630 2105
rect 7630 2071 7664 2105
rect 7664 2071 7732 2105
rect 7732 2071 7736 2105
rect 7558 2037 7736 2071
rect 7558 2003 7562 2037
rect 7562 2003 7630 2037
rect 7630 2003 7664 2037
rect 7664 2003 7732 2037
rect 7732 2003 7736 2037
rect 7558 1969 7736 2003
rect 7558 1935 7562 1969
rect 7562 1935 7630 1969
rect 7630 1935 7664 1969
rect 7664 1935 7732 1969
rect 7732 1935 7736 1969
rect 7558 1901 7736 1935
rect 7558 1867 7562 1901
rect 7562 1867 7630 1901
rect 7630 1867 7664 1901
rect 7664 1867 7732 1901
rect 7732 1867 7736 1901
rect 7558 1833 7736 1867
rect 7558 1799 7562 1833
rect 7562 1799 7630 1833
rect 7630 1799 7664 1833
rect 7664 1799 7732 1833
rect 7732 1799 7736 1833
rect 7558 1765 7736 1799
rect 7558 1731 7562 1765
rect 7562 1731 7630 1765
rect 7630 1731 7664 1765
rect 7664 1731 7732 1765
rect 7732 1731 7736 1765
rect 7558 1697 7736 1731
rect 7558 1663 7562 1697
rect 7562 1663 7630 1697
rect 7630 1663 7664 1697
rect 7664 1663 7732 1697
rect 7732 1663 7736 1697
rect 7558 1629 7736 1663
rect 7558 1595 7562 1629
rect 7562 1595 7630 1629
rect 7630 1595 7664 1629
rect 7664 1595 7732 1629
rect 7732 1595 7736 1629
rect 7558 1561 7736 1595
rect 7558 1527 7562 1561
rect 7562 1527 7630 1561
rect 7630 1527 7664 1561
rect 7664 1527 7732 1561
rect 7732 1527 7736 1561
rect 7558 1491 7736 1527
rect 7558 1479 7592 1491
rect 7702 1479 7736 1491
rect 8305 4388 8411 4494
rect 8054 4028 8088 4062
rect 8126 4028 8160 4062
rect 8198 4028 8232 4062
rect 8054 3954 8088 3988
rect 8126 3954 8160 3988
rect 8198 3954 8232 3988
rect 8054 3880 8088 3914
rect 8126 3880 8160 3914
rect 8198 3880 8232 3914
rect 8054 3806 8088 3840
rect 8126 3806 8160 3840
rect 8198 3806 8232 3840
rect 8054 3732 8088 3766
rect 8126 3732 8160 3766
rect 8198 3732 8232 3766
rect 8054 3658 8088 3692
rect 8126 3658 8160 3692
rect 8198 3658 8232 3692
rect 8054 3584 8088 3618
rect 8126 3584 8160 3618
rect 8198 3584 8232 3618
rect 8054 3510 8088 3544
rect 8126 3510 8160 3544
rect 8198 3510 8232 3544
rect 8054 3436 8088 3470
rect 8126 3436 8160 3470
rect 8198 3436 8232 3470
rect 8054 3362 8088 3396
rect 8126 3362 8160 3396
rect 8198 3362 8232 3396
rect 8054 3288 8088 3322
rect 8126 3288 8160 3322
rect 8198 3288 8232 3322
rect 8054 3214 8088 3248
rect 8126 3214 8160 3248
rect 8198 3214 8232 3248
rect 8054 3140 8088 3174
rect 8126 3140 8160 3174
rect 8198 3140 8232 3174
rect 8054 3066 8088 3100
rect 8126 3066 8160 3100
rect 8198 3066 8232 3100
rect 8054 2992 8088 3026
rect 8126 2992 8160 3026
rect 8198 2992 8232 3026
rect 8054 2918 8088 2952
rect 8126 2918 8160 2952
rect 8198 2918 8232 2952
rect 8054 2844 8088 2878
rect 8126 2844 8160 2878
rect 8198 2844 8232 2878
rect 8054 2770 8088 2804
rect 8126 2770 8160 2804
rect 8198 2770 8232 2804
rect 8054 2696 8088 2730
rect 8126 2696 8160 2730
rect 8198 2696 8232 2730
rect 8054 2622 8088 2656
rect 8126 2622 8160 2656
rect 8198 2622 8232 2656
rect 8054 2548 8088 2582
rect 8126 2548 8160 2582
rect 8198 2548 8232 2582
rect 8054 2474 8088 2508
rect 8126 2474 8160 2508
rect 8198 2474 8232 2508
rect 8054 2400 8088 2434
rect 8126 2400 8160 2434
rect 8198 2400 8232 2434
rect 8054 2326 8088 2360
rect 8126 2326 8160 2360
rect 8198 2326 8232 2360
rect 8054 2252 8088 2286
rect 8126 2252 8160 2286
rect 8198 2252 8232 2286
rect 8054 2178 8088 2212
rect 8126 2178 8160 2212
rect 8198 2178 8232 2212
rect 8054 2104 8088 2138
rect 8126 2104 8160 2138
rect 8198 2104 8232 2138
rect 8054 2030 8088 2064
rect 8126 2030 8160 2064
rect 8198 2030 8232 2064
rect 8054 1956 8088 1990
rect 8126 1956 8160 1990
rect 8198 1956 8232 1990
rect 8054 1882 8088 1916
rect 8126 1882 8160 1916
rect 8198 1882 8232 1916
rect 8054 1808 8088 1842
rect 8126 1808 8160 1842
rect 8198 1808 8232 1842
rect 8054 1734 8088 1768
rect 8126 1734 8160 1768
rect 8198 1734 8232 1768
rect 8054 1660 8088 1694
rect 8126 1660 8160 1694
rect 8198 1660 8232 1694
rect 8054 1586 8088 1620
rect 8126 1586 8160 1620
rect 8198 1586 8232 1620
rect 8054 1511 8088 1545
rect 8126 1511 8160 1545
rect 8198 1511 8232 1545
rect 8867 4388 8973 4494
rect 8622 4050 8656 4062
rect 8550 4046 8728 4050
rect 8550 4012 8554 4046
rect 8554 4012 8622 4046
rect 8622 4012 8656 4046
rect 8656 4012 8724 4046
rect 8724 4012 8728 4046
rect 8550 3978 8728 4012
rect 8550 3944 8554 3978
rect 8554 3944 8622 3978
rect 8622 3944 8656 3978
rect 8656 3944 8724 3978
rect 8724 3944 8728 3978
rect 8550 3910 8728 3944
rect 8550 3876 8554 3910
rect 8554 3876 8622 3910
rect 8622 3876 8656 3910
rect 8656 3876 8724 3910
rect 8724 3876 8728 3910
rect 8550 3842 8728 3876
rect 8550 3808 8554 3842
rect 8554 3808 8622 3842
rect 8622 3808 8656 3842
rect 8656 3808 8724 3842
rect 8724 3808 8728 3842
rect 8550 3774 8728 3808
rect 8550 3740 8554 3774
rect 8554 3740 8622 3774
rect 8622 3740 8656 3774
rect 8656 3740 8724 3774
rect 8724 3740 8728 3774
rect 8550 3706 8728 3740
rect 8550 3672 8554 3706
rect 8554 3672 8622 3706
rect 8622 3672 8656 3706
rect 8656 3672 8724 3706
rect 8724 3672 8728 3706
rect 8550 3638 8728 3672
rect 8550 3604 8554 3638
rect 8554 3604 8622 3638
rect 8622 3604 8656 3638
rect 8656 3604 8724 3638
rect 8724 3604 8728 3638
rect 8550 3570 8728 3604
rect 8550 3536 8554 3570
rect 8554 3536 8622 3570
rect 8622 3536 8656 3570
rect 8656 3536 8724 3570
rect 8724 3536 8728 3570
rect 8550 3502 8728 3536
rect 8550 3468 8554 3502
rect 8554 3468 8622 3502
rect 8622 3468 8656 3502
rect 8656 3468 8724 3502
rect 8724 3468 8728 3502
rect 8550 3434 8728 3468
rect 8550 3400 8554 3434
rect 8554 3400 8622 3434
rect 8622 3400 8656 3434
rect 8656 3400 8724 3434
rect 8724 3400 8728 3434
rect 8550 3366 8728 3400
rect 8550 3332 8554 3366
rect 8554 3332 8622 3366
rect 8622 3332 8656 3366
rect 8656 3332 8724 3366
rect 8724 3332 8728 3366
rect 8550 3298 8728 3332
rect 8550 3264 8554 3298
rect 8554 3264 8622 3298
rect 8622 3264 8656 3298
rect 8656 3264 8724 3298
rect 8724 3264 8728 3298
rect 8550 3230 8728 3264
rect 8550 3196 8554 3230
rect 8554 3196 8622 3230
rect 8622 3196 8656 3230
rect 8656 3196 8724 3230
rect 8724 3196 8728 3230
rect 8550 3162 8728 3196
rect 8550 3128 8554 3162
rect 8554 3128 8622 3162
rect 8622 3128 8656 3162
rect 8656 3128 8724 3162
rect 8724 3128 8728 3162
rect 8550 3092 8728 3128
rect 8550 3080 8584 3092
rect 8694 3080 8728 3092
rect 8550 2935 8728 3040
rect 8550 2901 8589 2935
rect 8589 2901 8623 2935
rect 8623 2901 8657 2935
rect 8657 2901 8691 2935
rect 8691 2901 8728 2935
rect 8550 2855 8728 2901
rect 8550 2821 8589 2855
rect 8589 2821 8623 2855
rect 8623 2821 8657 2855
rect 8657 2821 8691 2855
rect 8691 2821 8728 2855
rect 8550 2775 8728 2821
rect 8550 2741 8589 2775
rect 8589 2741 8623 2775
rect 8623 2741 8657 2775
rect 8657 2741 8691 2775
rect 8691 2741 8728 2775
rect 8550 2695 8728 2741
rect 8550 2661 8589 2695
rect 8589 2661 8623 2695
rect 8623 2661 8657 2695
rect 8657 2661 8691 2695
rect 8691 2661 8728 2695
rect 8550 2614 8728 2661
rect 8550 2580 8589 2614
rect 8589 2580 8623 2614
rect 8623 2580 8657 2614
rect 8657 2580 8691 2614
rect 8691 2580 8728 2614
rect 8550 2574 8728 2580
rect 8550 2501 8584 2535
rect 8622 2501 8656 2535
rect 8694 2501 8728 2535
rect 8622 2449 8656 2461
rect 8550 2445 8728 2449
rect 8550 2411 8554 2445
rect 8554 2411 8622 2445
rect 8622 2411 8656 2445
rect 8656 2411 8724 2445
rect 8724 2411 8728 2445
rect 8550 2377 8728 2411
rect 8550 2343 8554 2377
rect 8554 2343 8622 2377
rect 8622 2343 8656 2377
rect 8656 2343 8724 2377
rect 8724 2343 8728 2377
rect 8550 2309 8728 2343
rect 8550 2275 8554 2309
rect 8554 2275 8622 2309
rect 8622 2275 8656 2309
rect 8656 2275 8724 2309
rect 8724 2275 8728 2309
rect 8550 2241 8728 2275
rect 8550 2207 8554 2241
rect 8554 2207 8622 2241
rect 8622 2207 8656 2241
rect 8656 2207 8724 2241
rect 8724 2207 8728 2241
rect 8550 2173 8728 2207
rect 8550 2139 8554 2173
rect 8554 2139 8622 2173
rect 8622 2139 8656 2173
rect 8656 2139 8724 2173
rect 8724 2139 8728 2173
rect 8550 2105 8728 2139
rect 8550 2071 8554 2105
rect 8554 2071 8622 2105
rect 8622 2071 8656 2105
rect 8656 2071 8724 2105
rect 8724 2071 8728 2105
rect 8550 2037 8728 2071
rect 8550 2003 8554 2037
rect 8554 2003 8622 2037
rect 8622 2003 8656 2037
rect 8656 2003 8724 2037
rect 8724 2003 8728 2037
rect 8550 1969 8728 2003
rect 8550 1935 8554 1969
rect 8554 1935 8622 1969
rect 8622 1935 8656 1969
rect 8656 1935 8724 1969
rect 8724 1935 8728 1969
rect 8550 1901 8728 1935
rect 8550 1867 8554 1901
rect 8554 1867 8622 1901
rect 8622 1867 8656 1901
rect 8656 1867 8724 1901
rect 8724 1867 8728 1901
rect 8550 1833 8728 1867
rect 8550 1799 8554 1833
rect 8554 1799 8622 1833
rect 8622 1799 8656 1833
rect 8656 1799 8724 1833
rect 8724 1799 8728 1833
rect 8550 1765 8728 1799
rect 8550 1731 8554 1765
rect 8554 1731 8622 1765
rect 8622 1731 8656 1765
rect 8656 1731 8724 1765
rect 8724 1731 8728 1765
rect 8550 1697 8728 1731
rect 8550 1663 8554 1697
rect 8554 1663 8622 1697
rect 8622 1663 8656 1697
rect 8656 1663 8724 1697
rect 8724 1663 8728 1697
rect 8550 1629 8728 1663
rect 8550 1595 8554 1629
rect 8554 1595 8622 1629
rect 8622 1595 8656 1629
rect 8656 1595 8724 1629
rect 8724 1595 8728 1629
rect 8550 1561 8728 1595
rect 8550 1527 8554 1561
rect 8554 1527 8622 1561
rect 8622 1527 8656 1561
rect 8656 1527 8724 1561
rect 8724 1527 8728 1561
rect 8550 1491 8728 1527
rect 8550 1479 8584 1491
rect 8694 1479 8728 1491
rect 9297 4388 9403 4494
rect 9046 4028 9080 4062
rect 9118 4028 9152 4062
rect 9190 4028 9224 4062
rect 9046 3954 9080 3988
rect 9118 3954 9152 3988
rect 9190 3954 9224 3988
rect 9046 3880 9080 3914
rect 9118 3880 9152 3914
rect 9190 3880 9224 3914
rect 9046 3806 9080 3840
rect 9118 3806 9152 3840
rect 9190 3806 9224 3840
rect 9046 3732 9080 3766
rect 9118 3732 9152 3766
rect 9190 3732 9224 3766
rect 9046 3658 9080 3692
rect 9118 3658 9152 3692
rect 9190 3658 9224 3692
rect 9046 3584 9080 3618
rect 9118 3584 9152 3618
rect 9190 3584 9224 3618
rect 9046 3510 9080 3544
rect 9118 3510 9152 3544
rect 9190 3510 9224 3544
rect 9046 3436 9080 3470
rect 9118 3436 9152 3470
rect 9190 3436 9224 3470
rect 9046 3362 9080 3396
rect 9118 3362 9152 3396
rect 9190 3362 9224 3396
rect 9046 3288 9080 3322
rect 9118 3288 9152 3322
rect 9190 3288 9224 3322
rect 9046 3214 9080 3248
rect 9118 3214 9152 3248
rect 9190 3214 9224 3248
rect 9046 3140 9080 3174
rect 9118 3140 9152 3174
rect 9190 3140 9224 3174
rect 9046 3066 9080 3100
rect 9118 3066 9152 3100
rect 9190 3066 9224 3100
rect 9046 2992 9080 3026
rect 9118 2992 9152 3026
rect 9190 2992 9224 3026
rect 9046 2918 9080 2952
rect 9118 2918 9152 2952
rect 9190 2918 9224 2952
rect 9046 2844 9080 2878
rect 9118 2844 9152 2878
rect 9190 2844 9224 2878
rect 9046 2770 9080 2804
rect 9118 2770 9152 2804
rect 9190 2770 9224 2804
rect 9046 2696 9080 2730
rect 9118 2696 9152 2730
rect 9190 2696 9224 2730
rect 9046 2622 9080 2656
rect 9118 2622 9152 2656
rect 9190 2622 9224 2656
rect 9046 2548 9080 2582
rect 9118 2548 9152 2582
rect 9190 2548 9224 2582
rect 9046 2474 9080 2508
rect 9118 2474 9152 2508
rect 9190 2474 9224 2508
rect 9046 2400 9080 2434
rect 9118 2400 9152 2434
rect 9190 2400 9224 2434
rect 9046 2326 9080 2360
rect 9118 2326 9152 2360
rect 9190 2326 9224 2360
rect 9046 2252 9080 2286
rect 9118 2252 9152 2286
rect 9190 2252 9224 2286
rect 9046 2178 9080 2212
rect 9118 2178 9152 2212
rect 9190 2178 9224 2212
rect 9046 2104 9080 2138
rect 9118 2104 9152 2138
rect 9190 2104 9224 2138
rect 9046 2030 9080 2064
rect 9118 2030 9152 2064
rect 9190 2030 9224 2064
rect 9046 1956 9080 1990
rect 9118 1956 9152 1990
rect 9190 1956 9224 1990
rect 9046 1882 9080 1916
rect 9118 1882 9152 1916
rect 9190 1882 9224 1916
rect 9046 1808 9080 1842
rect 9118 1808 9152 1842
rect 9190 1808 9224 1842
rect 9046 1734 9080 1768
rect 9118 1734 9152 1768
rect 9190 1734 9224 1768
rect 9046 1660 9080 1694
rect 9118 1660 9152 1694
rect 9190 1660 9224 1694
rect 9046 1586 9080 1620
rect 9118 1586 9152 1620
rect 9190 1586 9224 1620
rect 9046 1511 9080 1545
rect 9118 1511 9152 1545
rect 9190 1511 9224 1545
rect 9859 4388 9965 4494
rect 9614 4050 9648 4062
rect 9542 4046 9720 4050
rect 9542 4012 9546 4046
rect 9546 4012 9614 4046
rect 9614 4012 9648 4046
rect 9648 4012 9716 4046
rect 9716 4012 9720 4046
rect 9542 3978 9720 4012
rect 9542 3944 9546 3978
rect 9546 3944 9614 3978
rect 9614 3944 9648 3978
rect 9648 3944 9716 3978
rect 9716 3944 9720 3978
rect 9542 3910 9720 3944
rect 9542 3876 9546 3910
rect 9546 3876 9614 3910
rect 9614 3876 9648 3910
rect 9648 3876 9716 3910
rect 9716 3876 9720 3910
rect 9542 3842 9720 3876
rect 9542 3808 9546 3842
rect 9546 3808 9614 3842
rect 9614 3808 9648 3842
rect 9648 3808 9716 3842
rect 9716 3808 9720 3842
rect 9542 3774 9720 3808
rect 9542 3740 9546 3774
rect 9546 3740 9614 3774
rect 9614 3740 9648 3774
rect 9648 3740 9716 3774
rect 9716 3740 9720 3774
rect 9542 3706 9720 3740
rect 9542 3672 9546 3706
rect 9546 3672 9614 3706
rect 9614 3672 9648 3706
rect 9648 3672 9716 3706
rect 9716 3672 9720 3706
rect 9542 3638 9720 3672
rect 9542 3604 9546 3638
rect 9546 3604 9614 3638
rect 9614 3604 9648 3638
rect 9648 3604 9716 3638
rect 9716 3604 9720 3638
rect 9542 3570 9720 3604
rect 9542 3536 9546 3570
rect 9546 3536 9614 3570
rect 9614 3536 9648 3570
rect 9648 3536 9716 3570
rect 9716 3536 9720 3570
rect 9542 3502 9720 3536
rect 9542 3468 9546 3502
rect 9546 3468 9614 3502
rect 9614 3468 9648 3502
rect 9648 3468 9716 3502
rect 9716 3468 9720 3502
rect 9542 3434 9720 3468
rect 9542 3400 9546 3434
rect 9546 3400 9614 3434
rect 9614 3400 9648 3434
rect 9648 3400 9716 3434
rect 9716 3400 9720 3434
rect 9542 3366 9720 3400
rect 9542 3332 9546 3366
rect 9546 3332 9614 3366
rect 9614 3332 9648 3366
rect 9648 3332 9716 3366
rect 9716 3332 9720 3366
rect 9542 3298 9720 3332
rect 9542 3264 9546 3298
rect 9546 3264 9614 3298
rect 9614 3264 9648 3298
rect 9648 3264 9716 3298
rect 9716 3264 9720 3298
rect 9542 3230 9720 3264
rect 9542 3196 9546 3230
rect 9546 3196 9614 3230
rect 9614 3196 9648 3230
rect 9648 3196 9716 3230
rect 9716 3196 9720 3230
rect 9542 3162 9720 3196
rect 9542 3128 9546 3162
rect 9546 3128 9614 3162
rect 9614 3128 9648 3162
rect 9648 3128 9716 3162
rect 9716 3128 9720 3162
rect 9542 3092 9720 3128
rect 9542 3080 9576 3092
rect 9686 3080 9720 3092
rect 9542 2935 9720 3040
rect 9542 2901 9581 2935
rect 9581 2901 9615 2935
rect 9615 2901 9649 2935
rect 9649 2901 9683 2935
rect 9683 2901 9720 2935
rect 9542 2855 9720 2901
rect 9542 2821 9581 2855
rect 9581 2821 9615 2855
rect 9615 2821 9649 2855
rect 9649 2821 9683 2855
rect 9683 2821 9720 2855
rect 9542 2775 9720 2821
rect 9542 2741 9581 2775
rect 9581 2741 9615 2775
rect 9615 2741 9649 2775
rect 9649 2741 9683 2775
rect 9683 2741 9720 2775
rect 9542 2695 9720 2741
rect 9542 2661 9581 2695
rect 9581 2661 9615 2695
rect 9615 2661 9649 2695
rect 9649 2661 9683 2695
rect 9683 2661 9720 2695
rect 9542 2614 9720 2661
rect 9542 2580 9581 2614
rect 9581 2580 9615 2614
rect 9615 2580 9649 2614
rect 9649 2580 9683 2614
rect 9683 2580 9720 2614
rect 9542 2574 9720 2580
rect 9542 2501 9576 2535
rect 9614 2501 9648 2535
rect 9686 2501 9720 2535
rect 9614 2449 9648 2461
rect 9542 2445 9720 2449
rect 9542 2411 9546 2445
rect 9546 2411 9614 2445
rect 9614 2411 9648 2445
rect 9648 2411 9716 2445
rect 9716 2411 9720 2445
rect 9542 2377 9720 2411
rect 9542 2343 9546 2377
rect 9546 2343 9614 2377
rect 9614 2343 9648 2377
rect 9648 2343 9716 2377
rect 9716 2343 9720 2377
rect 9542 2309 9720 2343
rect 9542 2275 9546 2309
rect 9546 2275 9614 2309
rect 9614 2275 9648 2309
rect 9648 2275 9716 2309
rect 9716 2275 9720 2309
rect 9542 2241 9720 2275
rect 9542 2207 9546 2241
rect 9546 2207 9614 2241
rect 9614 2207 9648 2241
rect 9648 2207 9716 2241
rect 9716 2207 9720 2241
rect 9542 2173 9720 2207
rect 9542 2139 9546 2173
rect 9546 2139 9614 2173
rect 9614 2139 9648 2173
rect 9648 2139 9716 2173
rect 9716 2139 9720 2173
rect 9542 2105 9720 2139
rect 9542 2071 9546 2105
rect 9546 2071 9614 2105
rect 9614 2071 9648 2105
rect 9648 2071 9716 2105
rect 9716 2071 9720 2105
rect 9542 2037 9720 2071
rect 9542 2003 9546 2037
rect 9546 2003 9614 2037
rect 9614 2003 9648 2037
rect 9648 2003 9716 2037
rect 9716 2003 9720 2037
rect 9542 1969 9720 2003
rect 9542 1935 9546 1969
rect 9546 1935 9614 1969
rect 9614 1935 9648 1969
rect 9648 1935 9716 1969
rect 9716 1935 9720 1969
rect 9542 1901 9720 1935
rect 9542 1867 9546 1901
rect 9546 1867 9614 1901
rect 9614 1867 9648 1901
rect 9648 1867 9716 1901
rect 9716 1867 9720 1901
rect 9542 1833 9720 1867
rect 9542 1799 9546 1833
rect 9546 1799 9614 1833
rect 9614 1799 9648 1833
rect 9648 1799 9716 1833
rect 9716 1799 9720 1833
rect 9542 1765 9720 1799
rect 9542 1731 9546 1765
rect 9546 1731 9614 1765
rect 9614 1731 9648 1765
rect 9648 1731 9716 1765
rect 9716 1731 9720 1765
rect 9542 1697 9720 1731
rect 9542 1663 9546 1697
rect 9546 1663 9614 1697
rect 9614 1663 9648 1697
rect 9648 1663 9716 1697
rect 9716 1663 9720 1697
rect 9542 1629 9720 1663
rect 9542 1595 9546 1629
rect 9546 1595 9614 1629
rect 9614 1595 9648 1629
rect 9648 1595 9716 1629
rect 9716 1595 9720 1629
rect 9542 1561 9720 1595
rect 9542 1527 9546 1561
rect 9546 1527 9614 1561
rect 9614 1527 9648 1561
rect 9648 1527 9716 1561
rect 9716 1527 9720 1561
rect 9542 1491 9720 1527
rect 9542 1479 9576 1491
rect 9686 1479 9720 1491
rect 10289 4388 10395 4494
rect 10038 4028 10072 4062
rect 10110 4028 10144 4062
rect 10182 4028 10216 4062
rect 10038 3954 10072 3988
rect 10110 3954 10144 3988
rect 10182 3954 10216 3988
rect 10038 3880 10072 3914
rect 10110 3880 10144 3914
rect 10182 3880 10216 3914
rect 10038 3806 10072 3840
rect 10110 3806 10144 3840
rect 10182 3806 10216 3840
rect 10038 3732 10072 3766
rect 10110 3732 10144 3766
rect 10182 3732 10216 3766
rect 10038 3658 10072 3692
rect 10110 3658 10144 3692
rect 10182 3658 10216 3692
rect 10038 3584 10072 3618
rect 10110 3584 10144 3618
rect 10182 3584 10216 3618
rect 10038 3510 10072 3544
rect 10110 3510 10144 3544
rect 10182 3510 10216 3544
rect 10038 3436 10072 3470
rect 10110 3436 10144 3470
rect 10182 3436 10216 3470
rect 10038 3362 10072 3396
rect 10110 3362 10144 3396
rect 10182 3362 10216 3396
rect 10038 3288 10072 3322
rect 10110 3288 10144 3322
rect 10182 3288 10216 3322
rect 10038 3214 10072 3248
rect 10110 3214 10144 3248
rect 10182 3214 10216 3248
rect 10038 3140 10072 3174
rect 10110 3140 10144 3174
rect 10182 3140 10216 3174
rect 10038 3066 10072 3100
rect 10110 3066 10144 3100
rect 10182 3066 10216 3100
rect 10038 2992 10072 3026
rect 10110 2992 10144 3026
rect 10182 2992 10216 3026
rect 10038 2918 10072 2952
rect 10110 2918 10144 2952
rect 10182 2918 10216 2952
rect 10038 2844 10072 2878
rect 10110 2844 10144 2878
rect 10182 2844 10216 2878
rect 10038 2770 10072 2804
rect 10110 2770 10144 2804
rect 10182 2770 10216 2804
rect 10038 2696 10072 2730
rect 10110 2696 10144 2730
rect 10182 2696 10216 2730
rect 10038 2622 10072 2656
rect 10110 2622 10144 2656
rect 10182 2622 10216 2656
rect 10038 2548 10072 2582
rect 10110 2548 10144 2582
rect 10182 2548 10216 2582
rect 10038 2474 10072 2508
rect 10110 2474 10144 2508
rect 10182 2474 10216 2508
rect 10038 2400 10072 2434
rect 10110 2400 10144 2434
rect 10182 2400 10216 2434
rect 10038 2326 10072 2360
rect 10110 2326 10144 2360
rect 10182 2326 10216 2360
rect 10038 2252 10072 2286
rect 10110 2252 10144 2286
rect 10182 2252 10216 2286
rect 10038 2178 10072 2212
rect 10110 2178 10144 2212
rect 10182 2178 10216 2212
rect 10038 2104 10072 2138
rect 10110 2104 10144 2138
rect 10182 2104 10216 2138
rect 10038 2030 10072 2064
rect 10110 2030 10144 2064
rect 10182 2030 10216 2064
rect 10038 1956 10072 1990
rect 10110 1956 10144 1990
rect 10182 1956 10216 1990
rect 10038 1882 10072 1916
rect 10110 1882 10144 1916
rect 10182 1882 10216 1916
rect 10038 1808 10072 1842
rect 10110 1808 10144 1842
rect 10182 1808 10216 1842
rect 10038 1734 10072 1768
rect 10110 1734 10144 1768
rect 10182 1734 10216 1768
rect 10038 1660 10072 1694
rect 10110 1660 10144 1694
rect 10182 1660 10216 1694
rect 10038 1586 10072 1620
rect 10110 1586 10144 1620
rect 10182 1586 10216 1620
rect 10038 1511 10072 1545
rect 10110 1511 10144 1545
rect 10182 1511 10216 1545
rect 10851 4388 10957 4494
rect 10606 4050 10640 4062
rect 10534 4046 10712 4050
rect 10534 4012 10538 4046
rect 10538 4012 10606 4046
rect 10606 4012 10640 4046
rect 10640 4012 10708 4046
rect 10708 4012 10712 4046
rect 10534 3978 10712 4012
rect 10534 3944 10538 3978
rect 10538 3944 10606 3978
rect 10606 3944 10640 3978
rect 10640 3944 10708 3978
rect 10708 3944 10712 3978
rect 10534 3910 10712 3944
rect 10534 3876 10538 3910
rect 10538 3876 10606 3910
rect 10606 3876 10640 3910
rect 10640 3876 10708 3910
rect 10708 3876 10712 3910
rect 10534 3842 10712 3876
rect 10534 3808 10538 3842
rect 10538 3808 10606 3842
rect 10606 3808 10640 3842
rect 10640 3808 10708 3842
rect 10708 3808 10712 3842
rect 10534 3774 10712 3808
rect 10534 3740 10538 3774
rect 10538 3740 10606 3774
rect 10606 3740 10640 3774
rect 10640 3740 10708 3774
rect 10708 3740 10712 3774
rect 10534 3706 10712 3740
rect 10534 3672 10538 3706
rect 10538 3672 10606 3706
rect 10606 3672 10640 3706
rect 10640 3672 10708 3706
rect 10708 3672 10712 3706
rect 10534 3638 10712 3672
rect 10534 3604 10538 3638
rect 10538 3604 10606 3638
rect 10606 3604 10640 3638
rect 10640 3604 10708 3638
rect 10708 3604 10712 3638
rect 10534 3570 10712 3604
rect 10534 3536 10538 3570
rect 10538 3536 10606 3570
rect 10606 3536 10640 3570
rect 10640 3536 10708 3570
rect 10708 3536 10712 3570
rect 10534 3502 10712 3536
rect 10534 3468 10538 3502
rect 10538 3468 10606 3502
rect 10606 3468 10640 3502
rect 10640 3468 10708 3502
rect 10708 3468 10712 3502
rect 10534 3434 10712 3468
rect 10534 3400 10538 3434
rect 10538 3400 10606 3434
rect 10606 3400 10640 3434
rect 10640 3400 10708 3434
rect 10708 3400 10712 3434
rect 10534 3366 10712 3400
rect 10534 3332 10538 3366
rect 10538 3332 10606 3366
rect 10606 3332 10640 3366
rect 10640 3332 10708 3366
rect 10708 3332 10712 3366
rect 10534 3298 10712 3332
rect 10534 3264 10538 3298
rect 10538 3264 10606 3298
rect 10606 3264 10640 3298
rect 10640 3264 10708 3298
rect 10708 3264 10712 3298
rect 10534 3230 10712 3264
rect 10534 3196 10538 3230
rect 10538 3196 10606 3230
rect 10606 3196 10640 3230
rect 10640 3196 10708 3230
rect 10708 3196 10712 3230
rect 10534 3162 10712 3196
rect 10534 3128 10538 3162
rect 10538 3128 10606 3162
rect 10606 3128 10640 3162
rect 10640 3128 10708 3162
rect 10708 3128 10712 3162
rect 10534 3092 10712 3128
rect 10534 3080 10568 3092
rect 10678 3080 10712 3092
rect 10534 3003 10568 3037
rect 10606 3003 10640 3037
rect 10678 3003 10712 3037
rect 10534 2920 10568 2954
rect 10606 2935 10640 2954
rect 10606 2920 10607 2935
rect 10607 2920 10640 2935
rect 10678 2920 10712 2954
rect 10534 2837 10568 2871
rect 10606 2855 10640 2871
rect 10606 2837 10607 2855
rect 10607 2837 10640 2855
rect 10678 2837 10712 2871
rect 10534 2753 10568 2787
rect 10606 2775 10640 2787
rect 10606 2753 10607 2775
rect 10607 2753 10640 2775
rect 10678 2753 10712 2787
rect 10534 2669 10568 2703
rect 10606 2695 10640 2703
rect 10606 2669 10607 2695
rect 10607 2669 10640 2695
rect 10678 2669 10712 2703
rect 10534 2585 10568 2619
rect 10606 2614 10640 2619
rect 10606 2585 10607 2614
rect 10607 2585 10640 2614
rect 10678 2585 10712 2619
rect 10534 2501 10568 2535
rect 10606 2501 10640 2535
rect 10678 2501 10712 2535
rect 10606 2449 10640 2461
rect 10534 2445 10712 2449
rect 10534 2411 10538 2445
rect 10538 2411 10606 2445
rect 10606 2411 10640 2445
rect 10640 2411 10708 2445
rect 10708 2411 10712 2445
rect 10534 2377 10712 2411
rect 10534 2343 10538 2377
rect 10538 2343 10606 2377
rect 10606 2343 10640 2377
rect 10640 2343 10708 2377
rect 10708 2343 10712 2377
rect 10534 2309 10712 2343
rect 10534 2275 10538 2309
rect 10538 2275 10606 2309
rect 10606 2275 10640 2309
rect 10640 2275 10708 2309
rect 10708 2275 10712 2309
rect 10534 2241 10712 2275
rect 10534 2207 10538 2241
rect 10538 2207 10606 2241
rect 10606 2207 10640 2241
rect 10640 2207 10708 2241
rect 10708 2207 10712 2241
rect 10534 2173 10712 2207
rect 10534 2139 10538 2173
rect 10538 2139 10606 2173
rect 10606 2139 10640 2173
rect 10640 2139 10708 2173
rect 10708 2139 10712 2173
rect 10534 2105 10712 2139
rect 10534 2071 10538 2105
rect 10538 2071 10606 2105
rect 10606 2071 10640 2105
rect 10640 2071 10708 2105
rect 10708 2071 10712 2105
rect 10534 2037 10712 2071
rect 10534 2003 10538 2037
rect 10538 2003 10606 2037
rect 10606 2003 10640 2037
rect 10640 2003 10708 2037
rect 10708 2003 10712 2037
rect 10534 1969 10712 2003
rect 10534 1935 10538 1969
rect 10538 1935 10606 1969
rect 10606 1935 10640 1969
rect 10640 1935 10708 1969
rect 10708 1935 10712 1969
rect 10534 1901 10712 1935
rect 10534 1867 10538 1901
rect 10538 1867 10606 1901
rect 10606 1867 10640 1901
rect 10640 1867 10708 1901
rect 10708 1867 10712 1901
rect 10534 1833 10712 1867
rect 10534 1799 10538 1833
rect 10538 1799 10606 1833
rect 10606 1799 10640 1833
rect 10640 1799 10708 1833
rect 10708 1799 10712 1833
rect 10534 1765 10712 1799
rect 10534 1731 10538 1765
rect 10538 1731 10606 1765
rect 10606 1731 10640 1765
rect 10640 1731 10708 1765
rect 10708 1731 10712 1765
rect 10534 1697 10712 1731
rect 10534 1663 10538 1697
rect 10538 1663 10606 1697
rect 10606 1663 10640 1697
rect 10640 1663 10708 1697
rect 10708 1663 10712 1697
rect 10534 1629 10712 1663
rect 10534 1595 10538 1629
rect 10538 1595 10606 1629
rect 10606 1595 10640 1629
rect 10640 1595 10708 1629
rect 10708 1595 10712 1629
rect 10534 1561 10712 1595
rect 10534 1527 10538 1561
rect 10538 1527 10606 1561
rect 10606 1527 10640 1561
rect 10640 1527 10708 1561
rect 10708 1527 10712 1561
rect 10534 1491 10712 1527
rect 10534 1479 10568 1491
rect 10678 1479 10712 1491
rect 11281 4388 11387 4494
rect 11030 4028 11064 4062
rect 11102 4028 11136 4062
rect 11174 4028 11208 4062
rect 11030 3954 11064 3988
rect 11102 3954 11136 3988
rect 11174 3954 11208 3988
rect 11030 3880 11064 3914
rect 11102 3880 11136 3914
rect 11174 3880 11208 3914
rect 11030 3806 11064 3840
rect 11102 3806 11136 3840
rect 11174 3806 11208 3840
rect 11030 3732 11064 3766
rect 11102 3732 11136 3766
rect 11174 3732 11208 3766
rect 11030 3658 11064 3692
rect 11102 3658 11136 3692
rect 11174 3658 11208 3692
rect 11030 3584 11064 3618
rect 11102 3584 11136 3618
rect 11174 3584 11208 3618
rect 11030 3510 11064 3544
rect 11102 3510 11136 3544
rect 11174 3510 11208 3544
rect 11030 3436 11064 3470
rect 11102 3436 11136 3470
rect 11174 3436 11208 3470
rect 11030 3362 11064 3396
rect 11102 3362 11136 3396
rect 11174 3362 11208 3396
rect 11030 3288 11064 3322
rect 11102 3288 11136 3322
rect 11174 3288 11208 3322
rect 11030 3214 11064 3248
rect 11102 3214 11136 3248
rect 11174 3214 11208 3248
rect 11030 3140 11064 3174
rect 11102 3140 11136 3174
rect 11174 3140 11208 3174
rect 11030 3066 11064 3100
rect 11102 3066 11136 3100
rect 11174 3066 11208 3100
rect 11030 2992 11064 3026
rect 11102 2992 11136 3026
rect 11174 2992 11208 3026
rect 11030 2918 11064 2952
rect 11102 2918 11136 2952
rect 11174 2918 11208 2952
rect 11030 2844 11064 2878
rect 11102 2844 11136 2878
rect 11174 2844 11208 2878
rect 11030 2770 11064 2804
rect 11102 2770 11136 2804
rect 11174 2770 11208 2804
rect 11030 2696 11064 2730
rect 11102 2696 11136 2730
rect 11174 2696 11208 2730
rect 11030 2622 11064 2656
rect 11102 2622 11136 2656
rect 11174 2622 11208 2656
rect 11030 2548 11064 2582
rect 11102 2548 11136 2582
rect 11174 2548 11208 2582
rect 11030 2474 11064 2508
rect 11102 2474 11136 2508
rect 11174 2474 11208 2508
rect 11030 2400 11064 2434
rect 11102 2400 11136 2434
rect 11174 2400 11208 2434
rect 11030 2326 11064 2360
rect 11102 2326 11136 2360
rect 11174 2326 11208 2360
rect 11030 2252 11064 2286
rect 11102 2252 11136 2286
rect 11174 2252 11208 2286
rect 11030 2178 11064 2212
rect 11102 2178 11136 2212
rect 11174 2178 11208 2212
rect 11030 2104 11064 2138
rect 11102 2104 11136 2138
rect 11174 2104 11208 2138
rect 11030 2030 11064 2064
rect 11102 2030 11136 2064
rect 11174 2030 11208 2064
rect 11030 1956 11064 1990
rect 11102 1956 11136 1990
rect 11174 1956 11208 1990
rect 11030 1882 11064 1916
rect 11102 1882 11136 1916
rect 11174 1882 11208 1916
rect 11030 1808 11064 1842
rect 11102 1808 11136 1842
rect 11174 1808 11208 1842
rect 11030 1734 11064 1768
rect 11102 1734 11136 1768
rect 11174 1734 11208 1768
rect 11030 1660 11064 1694
rect 11102 1660 11136 1694
rect 11174 1660 11208 1694
rect 11030 1586 11064 1620
rect 11102 1586 11136 1620
rect 11174 1586 11208 1620
rect 11030 1511 11064 1545
rect 11102 1511 11136 1545
rect 11174 1511 11208 1545
rect 11843 4388 11949 4494
rect 11598 4050 11632 4062
rect 11526 4046 11704 4050
rect 11526 4012 11530 4046
rect 11530 4012 11598 4046
rect 11598 4012 11632 4046
rect 11632 4012 11700 4046
rect 11700 4012 11704 4046
rect 11526 3978 11704 4012
rect 11526 3944 11530 3978
rect 11530 3944 11598 3978
rect 11598 3944 11632 3978
rect 11632 3944 11700 3978
rect 11700 3944 11704 3978
rect 11526 3910 11704 3944
rect 11526 3876 11530 3910
rect 11530 3876 11598 3910
rect 11598 3876 11632 3910
rect 11632 3876 11700 3910
rect 11700 3876 11704 3910
rect 11526 3842 11704 3876
rect 11526 3808 11530 3842
rect 11530 3808 11598 3842
rect 11598 3808 11632 3842
rect 11632 3808 11700 3842
rect 11700 3808 11704 3842
rect 11526 3774 11704 3808
rect 11526 3740 11530 3774
rect 11530 3740 11598 3774
rect 11598 3740 11632 3774
rect 11632 3740 11700 3774
rect 11700 3740 11704 3774
rect 11526 3706 11704 3740
rect 11526 3672 11530 3706
rect 11530 3672 11598 3706
rect 11598 3672 11632 3706
rect 11632 3672 11700 3706
rect 11700 3672 11704 3706
rect 11526 3638 11704 3672
rect 11526 3604 11530 3638
rect 11530 3604 11598 3638
rect 11598 3604 11632 3638
rect 11632 3604 11700 3638
rect 11700 3604 11704 3638
rect 11526 3570 11704 3604
rect 11526 3536 11530 3570
rect 11530 3536 11598 3570
rect 11598 3536 11632 3570
rect 11632 3536 11700 3570
rect 11700 3536 11704 3570
rect 11526 3502 11704 3536
rect 11526 3468 11530 3502
rect 11530 3468 11598 3502
rect 11598 3468 11632 3502
rect 11632 3468 11700 3502
rect 11700 3468 11704 3502
rect 11526 3434 11704 3468
rect 11526 3400 11530 3434
rect 11530 3400 11598 3434
rect 11598 3400 11632 3434
rect 11632 3400 11700 3434
rect 11700 3400 11704 3434
rect 11526 3366 11704 3400
rect 11526 3332 11530 3366
rect 11530 3332 11598 3366
rect 11598 3332 11632 3366
rect 11632 3332 11700 3366
rect 11700 3332 11704 3366
rect 11526 3298 11704 3332
rect 11526 3264 11530 3298
rect 11530 3264 11598 3298
rect 11598 3264 11632 3298
rect 11632 3264 11700 3298
rect 11700 3264 11704 3298
rect 11526 3230 11704 3264
rect 11526 3196 11530 3230
rect 11530 3196 11598 3230
rect 11598 3196 11632 3230
rect 11632 3196 11700 3230
rect 11700 3196 11704 3230
rect 11526 3162 11704 3196
rect 11526 3128 11530 3162
rect 11530 3128 11598 3162
rect 11598 3128 11632 3162
rect 11632 3128 11700 3162
rect 11700 3128 11704 3162
rect 11526 3092 11704 3128
rect 11526 3080 11560 3092
rect 11670 3080 11704 3092
rect 11526 3003 11560 3037
rect 11598 3003 11632 3037
rect 11670 3003 11704 3037
rect 11526 2920 11560 2954
rect 11598 2935 11632 2954
rect 11598 2920 11599 2935
rect 11599 2920 11632 2935
rect 11670 2920 11704 2954
rect 11526 2837 11560 2871
rect 11598 2855 11632 2871
rect 11598 2837 11599 2855
rect 11599 2837 11632 2855
rect 11670 2837 11704 2871
rect 11526 2753 11560 2787
rect 11598 2775 11632 2787
rect 11598 2753 11599 2775
rect 11599 2753 11632 2775
rect 11670 2753 11704 2787
rect 11526 2669 11560 2703
rect 11598 2695 11632 2703
rect 11598 2669 11599 2695
rect 11599 2669 11632 2695
rect 11670 2669 11704 2703
rect 11526 2585 11560 2619
rect 11598 2614 11632 2619
rect 11598 2585 11599 2614
rect 11599 2585 11632 2614
rect 11670 2585 11704 2619
rect 11526 2501 11560 2535
rect 11598 2501 11632 2535
rect 11670 2501 11704 2535
rect 11598 2449 11632 2461
rect 11526 2445 11704 2449
rect 11526 2411 11530 2445
rect 11530 2411 11598 2445
rect 11598 2411 11632 2445
rect 11632 2411 11700 2445
rect 11700 2411 11704 2445
rect 11526 2377 11704 2411
rect 11526 2343 11530 2377
rect 11530 2343 11598 2377
rect 11598 2343 11632 2377
rect 11632 2343 11700 2377
rect 11700 2343 11704 2377
rect 11526 2309 11704 2343
rect 11526 2275 11530 2309
rect 11530 2275 11598 2309
rect 11598 2275 11632 2309
rect 11632 2275 11700 2309
rect 11700 2275 11704 2309
rect 11526 2241 11704 2275
rect 11526 2207 11530 2241
rect 11530 2207 11598 2241
rect 11598 2207 11632 2241
rect 11632 2207 11700 2241
rect 11700 2207 11704 2241
rect 11526 2173 11704 2207
rect 11526 2139 11530 2173
rect 11530 2139 11598 2173
rect 11598 2139 11632 2173
rect 11632 2139 11700 2173
rect 11700 2139 11704 2173
rect 11526 2105 11704 2139
rect 11526 2071 11530 2105
rect 11530 2071 11598 2105
rect 11598 2071 11632 2105
rect 11632 2071 11700 2105
rect 11700 2071 11704 2105
rect 11526 2037 11704 2071
rect 11526 2003 11530 2037
rect 11530 2003 11598 2037
rect 11598 2003 11632 2037
rect 11632 2003 11700 2037
rect 11700 2003 11704 2037
rect 11526 1969 11704 2003
rect 11526 1935 11530 1969
rect 11530 1935 11598 1969
rect 11598 1935 11632 1969
rect 11632 1935 11700 1969
rect 11700 1935 11704 1969
rect 11526 1901 11704 1935
rect 11526 1867 11530 1901
rect 11530 1867 11598 1901
rect 11598 1867 11632 1901
rect 11632 1867 11700 1901
rect 11700 1867 11704 1901
rect 11526 1833 11704 1867
rect 11526 1799 11530 1833
rect 11530 1799 11598 1833
rect 11598 1799 11632 1833
rect 11632 1799 11700 1833
rect 11700 1799 11704 1833
rect 11526 1765 11704 1799
rect 11526 1731 11530 1765
rect 11530 1731 11598 1765
rect 11598 1731 11632 1765
rect 11632 1731 11700 1765
rect 11700 1731 11704 1765
rect 11526 1697 11704 1731
rect 11526 1663 11530 1697
rect 11530 1663 11598 1697
rect 11598 1663 11632 1697
rect 11632 1663 11700 1697
rect 11700 1663 11704 1697
rect 11526 1629 11704 1663
rect 11526 1595 11530 1629
rect 11530 1595 11598 1629
rect 11598 1595 11632 1629
rect 11632 1595 11700 1629
rect 11700 1595 11704 1629
rect 11526 1561 11704 1595
rect 11526 1527 11530 1561
rect 11530 1527 11598 1561
rect 11598 1527 11632 1561
rect 11632 1527 11700 1561
rect 11700 1527 11704 1561
rect 11526 1491 11704 1527
rect 11526 1479 11560 1491
rect 11670 1479 11704 1491
rect 12273 4388 12379 4494
rect 12022 4028 12056 4062
rect 12094 4028 12128 4062
rect 12166 4028 12200 4062
rect 12022 3954 12056 3988
rect 12094 3954 12128 3988
rect 12166 3954 12200 3988
rect 12022 3880 12056 3914
rect 12094 3880 12128 3914
rect 12166 3880 12200 3914
rect 12022 3806 12056 3840
rect 12094 3806 12128 3840
rect 12166 3806 12200 3840
rect 12022 3732 12056 3766
rect 12094 3732 12128 3766
rect 12166 3732 12200 3766
rect 12022 3658 12056 3692
rect 12094 3658 12128 3692
rect 12166 3658 12200 3692
rect 12022 3584 12056 3618
rect 12094 3584 12128 3618
rect 12166 3584 12200 3618
rect 12022 3510 12056 3544
rect 12094 3510 12128 3544
rect 12166 3510 12200 3544
rect 12022 3436 12056 3470
rect 12094 3436 12128 3470
rect 12166 3436 12200 3470
rect 12022 3362 12056 3396
rect 12094 3362 12128 3396
rect 12166 3362 12200 3396
rect 12022 3288 12056 3322
rect 12094 3288 12128 3322
rect 12166 3288 12200 3322
rect 12022 3214 12056 3248
rect 12094 3214 12128 3248
rect 12166 3214 12200 3248
rect 12022 3140 12056 3174
rect 12094 3140 12128 3174
rect 12166 3140 12200 3174
rect 12022 3066 12056 3100
rect 12094 3066 12128 3100
rect 12166 3066 12200 3100
rect 12022 2992 12056 3026
rect 12094 2992 12128 3026
rect 12166 2992 12200 3026
rect 12022 2918 12056 2952
rect 12094 2918 12128 2952
rect 12166 2918 12200 2952
rect 12022 2844 12056 2878
rect 12094 2844 12128 2878
rect 12166 2844 12200 2878
rect 12022 2770 12056 2804
rect 12094 2770 12128 2804
rect 12166 2770 12200 2804
rect 12022 2696 12056 2730
rect 12094 2696 12128 2730
rect 12166 2696 12200 2730
rect 12022 2622 12056 2656
rect 12094 2622 12128 2656
rect 12166 2622 12200 2656
rect 12022 2548 12056 2582
rect 12094 2548 12128 2582
rect 12166 2548 12200 2582
rect 12022 2474 12056 2508
rect 12094 2474 12128 2508
rect 12166 2474 12200 2508
rect 12022 2400 12056 2434
rect 12094 2400 12128 2434
rect 12166 2400 12200 2434
rect 12022 2326 12056 2360
rect 12094 2326 12128 2360
rect 12166 2326 12200 2360
rect 12022 2252 12056 2286
rect 12094 2252 12128 2286
rect 12166 2252 12200 2286
rect 12022 2178 12056 2212
rect 12094 2178 12128 2212
rect 12166 2178 12200 2212
rect 12022 2104 12056 2138
rect 12094 2104 12128 2138
rect 12166 2104 12200 2138
rect 12022 2030 12056 2064
rect 12094 2030 12128 2064
rect 12166 2030 12200 2064
rect 12022 1956 12056 1990
rect 12094 1956 12128 1990
rect 12166 1956 12200 1990
rect 12022 1882 12056 1916
rect 12094 1882 12128 1916
rect 12166 1882 12200 1916
rect 12022 1808 12056 1842
rect 12094 1808 12128 1842
rect 12166 1808 12200 1842
rect 12022 1734 12056 1768
rect 12094 1734 12128 1768
rect 12166 1734 12200 1768
rect 12022 1660 12056 1694
rect 12094 1660 12128 1694
rect 12166 1660 12200 1694
rect 12022 1586 12056 1620
rect 12094 1586 12128 1620
rect 12166 1586 12200 1620
rect 12022 1511 12056 1545
rect 12094 1511 12128 1545
rect 12166 1511 12200 1545
rect 12835 4388 12941 4494
rect 12590 4050 12624 4062
rect 12518 4046 12696 4050
rect 12518 4012 12522 4046
rect 12522 4012 12590 4046
rect 12590 4012 12624 4046
rect 12624 4012 12692 4046
rect 12692 4012 12696 4046
rect 12518 3978 12696 4012
rect 12518 3944 12522 3978
rect 12522 3944 12590 3978
rect 12590 3944 12624 3978
rect 12624 3944 12692 3978
rect 12692 3944 12696 3978
rect 12518 3910 12696 3944
rect 12518 3876 12522 3910
rect 12522 3876 12590 3910
rect 12590 3876 12624 3910
rect 12624 3876 12692 3910
rect 12692 3876 12696 3910
rect 12518 3842 12696 3876
rect 12518 3808 12522 3842
rect 12522 3808 12590 3842
rect 12590 3808 12624 3842
rect 12624 3808 12692 3842
rect 12692 3808 12696 3842
rect 12518 3774 12696 3808
rect 12518 3740 12522 3774
rect 12522 3740 12590 3774
rect 12590 3740 12624 3774
rect 12624 3740 12692 3774
rect 12692 3740 12696 3774
rect 12518 3706 12696 3740
rect 12518 3672 12522 3706
rect 12522 3672 12590 3706
rect 12590 3672 12624 3706
rect 12624 3672 12692 3706
rect 12692 3672 12696 3706
rect 12518 3638 12696 3672
rect 12518 3604 12522 3638
rect 12522 3604 12590 3638
rect 12590 3604 12624 3638
rect 12624 3604 12692 3638
rect 12692 3604 12696 3638
rect 12518 3570 12696 3604
rect 12518 3536 12522 3570
rect 12522 3536 12590 3570
rect 12590 3536 12624 3570
rect 12624 3536 12692 3570
rect 12692 3536 12696 3570
rect 12518 3502 12696 3536
rect 12518 3468 12522 3502
rect 12522 3468 12590 3502
rect 12590 3468 12624 3502
rect 12624 3468 12692 3502
rect 12692 3468 12696 3502
rect 12518 3434 12696 3468
rect 12518 3400 12522 3434
rect 12522 3400 12590 3434
rect 12590 3400 12624 3434
rect 12624 3400 12692 3434
rect 12692 3400 12696 3434
rect 12518 3366 12696 3400
rect 12518 3332 12522 3366
rect 12522 3332 12590 3366
rect 12590 3332 12624 3366
rect 12624 3332 12692 3366
rect 12692 3332 12696 3366
rect 12518 3298 12696 3332
rect 12518 3264 12522 3298
rect 12522 3264 12590 3298
rect 12590 3264 12624 3298
rect 12624 3264 12692 3298
rect 12692 3264 12696 3298
rect 12518 3230 12696 3264
rect 12518 3196 12522 3230
rect 12522 3196 12590 3230
rect 12590 3196 12624 3230
rect 12624 3196 12692 3230
rect 12692 3196 12696 3230
rect 12518 3162 12696 3196
rect 12518 3128 12522 3162
rect 12522 3128 12590 3162
rect 12590 3128 12624 3162
rect 12624 3128 12692 3162
rect 12692 3128 12696 3162
rect 12518 3092 12696 3128
rect 12518 3080 12552 3092
rect 12662 3080 12696 3092
rect 12518 3004 12552 3038
rect 12590 3004 12624 3038
rect 12662 3004 12696 3038
rect 12518 2921 12552 2955
rect 12590 2935 12624 2955
rect 12590 2921 12591 2935
rect 12591 2921 12624 2935
rect 12662 2921 12696 2955
rect 12518 2837 12552 2871
rect 12590 2855 12624 2871
rect 12590 2837 12591 2855
rect 12591 2837 12624 2855
rect 12662 2837 12696 2871
rect 12518 2753 12552 2787
rect 12590 2775 12624 2787
rect 12590 2753 12591 2775
rect 12591 2753 12624 2775
rect 12662 2753 12696 2787
rect 12518 2669 12552 2703
rect 12590 2695 12624 2703
rect 12590 2669 12591 2695
rect 12591 2669 12624 2695
rect 12662 2669 12696 2703
rect 12518 2585 12552 2619
rect 12590 2614 12624 2619
rect 12590 2585 12591 2614
rect 12591 2585 12624 2614
rect 12662 2585 12696 2619
rect 12518 2501 12552 2535
rect 12590 2501 12624 2535
rect 12662 2501 12696 2535
rect 12590 2449 12624 2461
rect 12518 2445 12696 2449
rect 12518 2411 12522 2445
rect 12522 2411 12590 2445
rect 12590 2411 12624 2445
rect 12624 2411 12692 2445
rect 12692 2411 12696 2445
rect 12518 2377 12696 2411
rect 12518 2343 12522 2377
rect 12522 2343 12590 2377
rect 12590 2343 12624 2377
rect 12624 2343 12692 2377
rect 12692 2343 12696 2377
rect 12518 2309 12696 2343
rect 12518 2275 12522 2309
rect 12522 2275 12590 2309
rect 12590 2275 12624 2309
rect 12624 2275 12692 2309
rect 12692 2275 12696 2309
rect 12518 2241 12696 2275
rect 12518 2207 12522 2241
rect 12522 2207 12590 2241
rect 12590 2207 12624 2241
rect 12624 2207 12692 2241
rect 12692 2207 12696 2241
rect 12518 2173 12696 2207
rect 12518 2139 12522 2173
rect 12522 2139 12590 2173
rect 12590 2139 12624 2173
rect 12624 2139 12692 2173
rect 12692 2139 12696 2173
rect 12518 2105 12696 2139
rect 12518 2071 12522 2105
rect 12522 2071 12590 2105
rect 12590 2071 12624 2105
rect 12624 2071 12692 2105
rect 12692 2071 12696 2105
rect 12518 2037 12696 2071
rect 12518 2003 12522 2037
rect 12522 2003 12590 2037
rect 12590 2003 12624 2037
rect 12624 2003 12692 2037
rect 12692 2003 12696 2037
rect 12518 1969 12696 2003
rect 12518 1935 12522 1969
rect 12522 1935 12590 1969
rect 12590 1935 12624 1969
rect 12624 1935 12692 1969
rect 12692 1935 12696 1969
rect 12518 1901 12696 1935
rect 12518 1867 12522 1901
rect 12522 1867 12590 1901
rect 12590 1867 12624 1901
rect 12624 1867 12692 1901
rect 12692 1867 12696 1901
rect 12518 1833 12696 1867
rect 12518 1799 12522 1833
rect 12522 1799 12590 1833
rect 12590 1799 12624 1833
rect 12624 1799 12692 1833
rect 12692 1799 12696 1833
rect 12518 1765 12696 1799
rect 12518 1731 12522 1765
rect 12522 1731 12590 1765
rect 12590 1731 12624 1765
rect 12624 1731 12692 1765
rect 12692 1731 12696 1765
rect 12518 1697 12696 1731
rect 12518 1663 12522 1697
rect 12522 1663 12590 1697
rect 12590 1663 12624 1697
rect 12624 1663 12692 1697
rect 12692 1663 12696 1697
rect 12518 1629 12696 1663
rect 12518 1595 12522 1629
rect 12522 1595 12590 1629
rect 12590 1595 12624 1629
rect 12624 1595 12692 1629
rect 12692 1595 12696 1629
rect 12518 1561 12696 1595
rect 12518 1527 12522 1561
rect 12522 1527 12590 1561
rect 12590 1527 12624 1561
rect 12624 1527 12692 1561
rect 12692 1527 12696 1561
rect 12518 1491 12696 1527
rect 12518 1479 12552 1491
rect 12662 1479 12696 1491
rect 13265 4388 13371 4494
rect 13014 4028 13048 4062
rect 13086 4028 13120 4062
rect 13158 4028 13192 4062
rect 13014 3954 13048 3988
rect 13086 3954 13120 3988
rect 13158 3954 13192 3988
rect 13014 3880 13048 3914
rect 13086 3880 13120 3914
rect 13158 3880 13192 3914
rect 13014 3806 13048 3840
rect 13086 3806 13120 3840
rect 13158 3806 13192 3840
rect 13014 3732 13048 3766
rect 13086 3732 13120 3766
rect 13158 3732 13192 3766
rect 13014 3658 13048 3692
rect 13086 3658 13120 3692
rect 13158 3658 13192 3692
rect 13014 3584 13048 3618
rect 13086 3584 13120 3618
rect 13158 3584 13192 3618
rect 13014 3510 13048 3544
rect 13086 3510 13120 3544
rect 13158 3510 13192 3544
rect 13014 3436 13048 3470
rect 13086 3436 13120 3470
rect 13158 3436 13192 3470
rect 13014 3362 13048 3396
rect 13086 3362 13120 3396
rect 13158 3362 13192 3396
rect 13014 3288 13048 3322
rect 13086 3288 13120 3322
rect 13158 3288 13192 3322
rect 13014 3214 13048 3248
rect 13086 3214 13120 3248
rect 13158 3214 13192 3248
rect 13014 3140 13048 3174
rect 13086 3140 13120 3174
rect 13158 3140 13192 3174
rect 13014 3066 13048 3100
rect 13086 3066 13120 3100
rect 13158 3066 13192 3100
rect 13014 2992 13048 3026
rect 13086 2992 13120 3026
rect 13158 2992 13192 3026
rect 13014 2918 13048 2952
rect 13086 2918 13120 2952
rect 13158 2918 13192 2952
rect 13014 2844 13048 2878
rect 13086 2844 13120 2878
rect 13158 2844 13192 2878
rect 13014 2770 13048 2804
rect 13086 2770 13120 2804
rect 13158 2770 13192 2804
rect 13014 2696 13048 2730
rect 13086 2696 13120 2730
rect 13158 2696 13192 2730
rect 13014 2622 13048 2656
rect 13086 2622 13120 2656
rect 13158 2622 13192 2656
rect 13014 2548 13048 2582
rect 13086 2548 13120 2582
rect 13158 2548 13192 2582
rect 13014 2474 13048 2508
rect 13086 2474 13120 2508
rect 13158 2474 13192 2508
rect 13014 2400 13048 2434
rect 13086 2400 13120 2434
rect 13158 2400 13192 2434
rect 13014 2326 13048 2360
rect 13086 2326 13120 2360
rect 13158 2326 13192 2360
rect 13014 2252 13048 2286
rect 13086 2252 13120 2286
rect 13158 2252 13192 2286
rect 13014 2178 13048 2212
rect 13086 2178 13120 2212
rect 13158 2178 13192 2212
rect 13014 2104 13048 2138
rect 13086 2104 13120 2138
rect 13158 2104 13192 2138
rect 13014 2030 13048 2064
rect 13086 2030 13120 2064
rect 13158 2030 13192 2064
rect 13014 1956 13048 1990
rect 13086 1956 13120 1990
rect 13158 1956 13192 1990
rect 13014 1882 13048 1916
rect 13086 1882 13120 1916
rect 13158 1882 13192 1916
rect 13014 1808 13048 1842
rect 13086 1808 13120 1842
rect 13158 1808 13192 1842
rect 13014 1734 13048 1768
rect 13086 1734 13120 1768
rect 13158 1734 13192 1768
rect 13014 1660 13048 1694
rect 13086 1660 13120 1694
rect 13158 1660 13192 1694
rect 13014 1586 13048 1620
rect 13086 1586 13120 1620
rect 13158 1586 13192 1620
rect 13014 1511 13048 1545
rect 13086 1511 13120 1545
rect 13158 1511 13192 1545
rect 13827 4388 13933 4494
rect 13582 4050 13616 4062
rect 13510 4046 13688 4050
rect 13510 4012 13514 4046
rect 13514 4012 13582 4046
rect 13582 4012 13616 4046
rect 13616 4012 13684 4046
rect 13684 4012 13688 4046
rect 13510 3978 13688 4012
rect 13510 3944 13514 3978
rect 13514 3944 13582 3978
rect 13582 3944 13616 3978
rect 13616 3944 13684 3978
rect 13684 3944 13688 3978
rect 13510 3910 13688 3944
rect 13510 3876 13514 3910
rect 13514 3876 13582 3910
rect 13582 3876 13616 3910
rect 13616 3876 13684 3910
rect 13684 3876 13688 3910
rect 13510 3842 13688 3876
rect 13510 3808 13514 3842
rect 13514 3808 13582 3842
rect 13582 3808 13616 3842
rect 13616 3808 13684 3842
rect 13684 3808 13688 3842
rect 13510 3774 13688 3808
rect 13510 3740 13514 3774
rect 13514 3740 13582 3774
rect 13582 3740 13616 3774
rect 13616 3740 13684 3774
rect 13684 3740 13688 3774
rect 13510 3706 13688 3740
rect 13510 3672 13514 3706
rect 13514 3672 13582 3706
rect 13582 3672 13616 3706
rect 13616 3672 13684 3706
rect 13684 3672 13688 3706
rect 13510 3638 13688 3672
rect 13510 3604 13514 3638
rect 13514 3604 13582 3638
rect 13582 3604 13616 3638
rect 13616 3604 13684 3638
rect 13684 3604 13688 3638
rect 13510 3570 13688 3604
rect 13510 3536 13514 3570
rect 13514 3536 13582 3570
rect 13582 3536 13616 3570
rect 13616 3536 13684 3570
rect 13684 3536 13688 3570
rect 13510 3502 13688 3536
rect 13510 3468 13514 3502
rect 13514 3468 13582 3502
rect 13582 3468 13616 3502
rect 13616 3468 13684 3502
rect 13684 3468 13688 3502
rect 13510 3434 13688 3468
rect 13510 3400 13514 3434
rect 13514 3400 13582 3434
rect 13582 3400 13616 3434
rect 13616 3400 13684 3434
rect 13684 3400 13688 3434
rect 13510 3366 13688 3400
rect 13510 3332 13514 3366
rect 13514 3332 13582 3366
rect 13582 3332 13616 3366
rect 13616 3332 13684 3366
rect 13684 3332 13688 3366
rect 13510 3298 13688 3332
rect 13510 3264 13514 3298
rect 13514 3264 13582 3298
rect 13582 3264 13616 3298
rect 13616 3264 13684 3298
rect 13684 3264 13688 3298
rect 13510 3230 13688 3264
rect 13510 3196 13514 3230
rect 13514 3196 13582 3230
rect 13582 3196 13616 3230
rect 13616 3196 13684 3230
rect 13684 3196 13688 3230
rect 13510 3162 13688 3196
rect 13510 3128 13514 3162
rect 13514 3128 13582 3162
rect 13582 3128 13616 3162
rect 13616 3128 13684 3162
rect 13684 3128 13688 3162
rect 13510 3092 13688 3128
rect 13510 3080 13544 3092
rect 13654 3080 13688 3092
rect 13510 2935 13688 3040
rect 13510 2901 13549 2935
rect 13549 2901 13583 2935
rect 13583 2901 13617 2935
rect 13617 2901 13651 2935
rect 13651 2901 13688 2935
rect 13510 2855 13688 2901
rect 13510 2821 13549 2855
rect 13549 2821 13583 2855
rect 13583 2821 13617 2855
rect 13617 2821 13651 2855
rect 13651 2821 13688 2855
rect 13510 2775 13688 2821
rect 13510 2741 13549 2775
rect 13549 2741 13583 2775
rect 13583 2741 13617 2775
rect 13617 2741 13651 2775
rect 13651 2741 13688 2775
rect 13510 2695 13688 2741
rect 13510 2661 13549 2695
rect 13549 2661 13583 2695
rect 13583 2661 13617 2695
rect 13617 2661 13651 2695
rect 13651 2661 13688 2695
rect 13510 2614 13688 2661
rect 13510 2580 13549 2614
rect 13549 2580 13583 2614
rect 13583 2580 13617 2614
rect 13617 2580 13651 2614
rect 13651 2580 13688 2614
rect 13510 2574 13688 2580
rect 13510 2501 13544 2535
rect 13582 2501 13616 2535
rect 13654 2501 13688 2535
rect 13582 2449 13616 2461
rect 13510 2445 13688 2449
rect 13510 2411 13514 2445
rect 13514 2411 13582 2445
rect 13582 2411 13616 2445
rect 13616 2411 13684 2445
rect 13684 2411 13688 2445
rect 13510 2377 13688 2411
rect 13510 2343 13514 2377
rect 13514 2343 13582 2377
rect 13582 2343 13616 2377
rect 13616 2343 13684 2377
rect 13684 2343 13688 2377
rect 13510 2309 13688 2343
rect 13510 2275 13514 2309
rect 13514 2275 13582 2309
rect 13582 2275 13616 2309
rect 13616 2275 13684 2309
rect 13684 2275 13688 2309
rect 13510 2241 13688 2275
rect 13510 2207 13514 2241
rect 13514 2207 13582 2241
rect 13582 2207 13616 2241
rect 13616 2207 13684 2241
rect 13684 2207 13688 2241
rect 13510 2173 13688 2207
rect 13510 2139 13514 2173
rect 13514 2139 13582 2173
rect 13582 2139 13616 2173
rect 13616 2139 13684 2173
rect 13684 2139 13688 2173
rect 13510 2105 13688 2139
rect 13510 2071 13514 2105
rect 13514 2071 13582 2105
rect 13582 2071 13616 2105
rect 13616 2071 13684 2105
rect 13684 2071 13688 2105
rect 13510 2037 13688 2071
rect 13510 2003 13514 2037
rect 13514 2003 13582 2037
rect 13582 2003 13616 2037
rect 13616 2003 13684 2037
rect 13684 2003 13688 2037
rect 13510 1969 13688 2003
rect 13510 1935 13514 1969
rect 13514 1935 13582 1969
rect 13582 1935 13616 1969
rect 13616 1935 13684 1969
rect 13684 1935 13688 1969
rect 13510 1901 13688 1935
rect 13510 1867 13514 1901
rect 13514 1867 13582 1901
rect 13582 1867 13616 1901
rect 13616 1867 13684 1901
rect 13684 1867 13688 1901
rect 13510 1833 13688 1867
rect 13510 1799 13514 1833
rect 13514 1799 13582 1833
rect 13582 1799 13616 1833
rect 13616 1799 13684 1833
rect 13684 1799 13688 1833
rect 13510 1765 13688 1799
rect 13510 1731 13514 1765
rect 13514 1731 13582 1765
rect 13582 1731 13616 1765
rect 13616 1731 13684 1765
rect 13684 1731 13688 1765
rect 13510 1697 13688 1731
rect 13510 1663 13514 1697
rect 13514 1663 13582 1697
rect 13582 1663 13616 1697
rect 13616 1663 13684 1697
rect 13684 1663 13688 1697
rect 13510 1629 13688 1663
rect 13510 1595 13514 1629
rect 13514 1595 13582 1629
rect 13582 1595 13616 1629
rect 13616 1595 13684 1629
rect 13684 1595 13688 1629
rect 13510 1561 13688 1595
rect 13510 1527 13514 1561
rect 13514 1527 13582 1561
rect 13582 1527 13616 1561
rect 13616 1527 13684 1561
rect 13684 1527 13688 1561
rect 13510 1491 13688 1527
rect 13510 1479 13544 1491
rect 13654 1479 13688 1491
rect 14185 4388 14291 4494
rect 14006 4046 14112 4062
rect 14006 4012 14042 4046
rect 14042 4012 14076 4046
rect 14076 4012 14112 4046
rect 14006 3978 14112 4012
rect 14006 3944 14042 3978
rect 14042 3944 14076 3978
rect 14076 3944 14112 3978
rect 14006 3910 14112 3944
rect 14006 3876 14042 3910
rect 14042 3876 14076 3910
rect 14076 3876 14112 3910
rect 14006 3842 14112 3876
rect 14006 3808 14042 3842
rect 14042 3808 14076 3842
rect 14076 3808 14112 3842
rect 14006 3774 14112 3808
rect 14006 3740 14042 3774
rect 14042 3740 14076 3774
rect 14076 3740 14112 3774
rect 14006 3706 14112 3740
rect 14006 3672 14042 3706
rect 14042 3672 14076 3706
rect 14076 3672 14112 3706
rect 14006 3638 14112 3672
rect 14006 3604 14042 3638
rect 14042 3604 14076 3638
rect 14076 3604 14112 3638
rect 14006 3570 14112 3604
rect 14006 3536 14042 3570
rect 14042 3536 14076 3570
rect 14076 3536 14112 3570
rect 14006 3502 14112 3536
rect 14006 3468 14042 3502
rect 14042 3468 14076 3502
rect 14076 3468 14112 3502
rect 14006 3434 14112 3468
rect 14006 3400 14042 3434
rect 14042 3400 14076 3434
rect 14076 3400 14112 3434
rect 14006 3366 14112 3400
rect 14006 3332 14042 3366
rect 14042 3332 14076 3366
rect 14076 3332 14112 3366
rect 14006 3298 14112 3332
rect 14006 3264 14042 3298
rect 14042 3264 14076 3298
rect 14076 3264 14112 3298
rect 14006 3230 14112 3264
rect 14006 3196 14042 3230
rect 14042 3196 14076 3230
rect 14076 3196 14112 3230
rect 14006 3162 14112 3196
rect 14006 3128 14042 3162
rect 14042 3128 14076 3162
rect 14076 3128 14112 3162
rect 14006 2732 14112 3128
rect 14006 2659 14040 2693
rect 14078 2659 14112 2693
rect 14006 2586 14040 2620
rect 14078 2586 14112 2620
rect 14006 2513 14040 2547
rect 14078 2513 14112 2547
rect 14006 2440 14040 2474
rect 14078 2440 14112 2474
rect 14006 2367 14040 2401
rect 14078 2367 14112 2401
rect 14006 2294 14040 2328
rect 14078 2294 14112 2328
rect 14006 2221 14040 2255
rect 14078 2221 14112 2255
rect 14006 2148 14040 2182
rect 14078 2148 14112 2182
rect 14006 2075 14040 2109
rect 14078 2075 14112 2109
rect 14006 2002 14040 2036
rect 14078 2002 14112 2036
rect 14006 1929 14040 1963
rect 14078 1929 14112 1963
rect 14006 1856 14040 1890
rect 14078 1856 14112 1890
rect 14006 1783 14040 1817
rect 14078 1783 14112 1817
rect 14006 1710 14040 1744
rect 14078 1710 14112 1744
rect 14006 1637 14040 1671
rect 14078 1637 14112 1671
rect 14006 1564 14040 1598
rect 14078 1564 14112 1598
rect 14006 1491 14040 1525
rect 14078 1491 14112 1525
rect 14510 4490 14544 4506
rect 14582 4504 14599 4524
rect 14599 4504 14616 4524
rect 14582 4490 14616 4504
rect 14431 4448 14465 4482
rect 14510 4436 14531 4451
rect 14531 4436 14544 4451
rect 14510 4417 14544 4436
rect 14582 4434 14599 4451
rect 14599 4434 14616 4451
rect 14582 4417 14616 4434
rect 14431 4375 14465 4409
rect 14510 4365 14531 4378
rect 14531 4365 14544 4378
rect 14510 4344 14544 4365
rect 14582 4364 14599 4378
rect 14599 4364 14616 4378
rect 14582 4344 14616 4364
rect 14431 4302 14465 4336
rect 14510 4294 14531 4305
rect 14531 4294 14544 4305
rect 14582 4294 14599 4305
rect 14599 4294 14616 4305
rect 14510 4271 14544 4294
rect 14582 4271 14616 4294
rect 14431 4229 14465 4263
rect 14510 4223 14531 4232
rect 14531 4223 14544 4232
rect 14582 4223 14599 4232
rect 14599 4223 14616 4232
rect 14510 4198 14544 4223
rect 14582 4198 14616 4223
rect 14431 4156 14465 4190
rect 14510 4152 14531 4159
rect 14531 4152 14544 4159
rect 14582 4152 14599 4159
rect 14599 4152 14616 4159
rect 14510 4125 14544 4152
rect 14582 4125 14616 4152
rect 14431 4083 14465 4117
rect 14510 4052 14544 4086
rect 14582 4081 14599 4086
rect 14599 4081 14616 4086
rect 14582 4052 14616 4081
rect 14431 4034 14465 4044
rect 14431 4010 14454 4034
rect 14454 4010 14465 4034
rect 14510 3979 14544 4013
rect 14582 4007 14599 4013
rect 14599 4007 14616 4013
rect 14582 3979 14616 4007
rect 14431 3966 14465 3971
rect 14431 3937 14454 3966
rect 14454 3937 14465 3966
rect 14510 3906 14544 3940
rect 14582 3936 14599 3940
rect 14599 3936 14616 3940
rect 14582 3906 14616 3936
rect 14431 3864 14454 3898
rect 14454 3864 14465 3898
rect 14510 3833 14544 3867
rect 14582 3862 14599 3867
rect 14599 3862 14616 3867
rect 14582 3833 14616 3862
rect 14431 3796 14454 3825
rect 14454 3796 14465 3825
rect 14431 3791 14465 3796
rect 14510 3760 14544 3794
rect 14582 3791 14599 3794
rect 14599 3791 14616 3794
rect 14582 3760 14616 3791
rect 14431 3728 14454 3752
rect 14454 3728 14465 3752
rect 14431 3718 14465 3728
rect 14510 3687 14544 3721
rect 14582 3717 14599 3721
rect 14599 3717 14616 3721
rect 14582 3687 14616 3717
rect 14431 3660 14454 3679
rect 14454 3660 14465 3679
rect 14431 3645 14465 3660
rect 14510 3614 14544 3648
rect 14582 3646 14599 3648
rect 14599 3646 14616 3648
rect 14582 3614 14616 3646
rect 14431 3592 14454 3606
rect 14454 3592 14465 3606
rect 14431 3572 14465 3592
rect 14510 3541 14544 3575
rect 14582 3572 14599 3575
rect 14599 3572 14616 3575
rect 14582 3541 14616 3572
rect 14431 3524 14454 3533
rect 14454 3524 14465 3533
rect 14431 3499 14465 3524
rect 14510 3468 14544 3502
rect 14582 3501 14599 3502
rect 14599 3501 14616 3502
rect 14582 3468 14616 3501
rect 14431 3456 14454 3460
rect 14454 3456 14465 3460
rect 14431 3426 14465 3456
rect 14510 3395 14544 3429
rect 14582 3427 14599 3429
rect 14599 3427 14616 3429
rect 14582 3395 14616 3427
rect 14431 3354 14465 3387
rect 14431 3353 14454 3354
rect 14454 3353 14465 3354
rect 14510 3322 14544 3356
rect 14582 3322 14616 3356
rect 14431 3286 14465 3314
rect 14431 3280 14454 3286
rect 14454 3280 14465 3286
rect 14510 3249 14544 3283
rect 14582 3282 14599 3283
rect 14599 3282 14616 3283
rect 14582 3249 14616 3282
rect 14431 3218 14465 3241
rect 14431 3207 14454 3218
rect 14454 3207 14465 3218
rect 14510 3176 14544 3210
rect 14582 3176 14616 3210
rect 14431 3150 14465 3168
rect 14431 3134 14454 3150
rect 14454 3134 14465 3150
rect 14510 3103 14544 3137
rect 14582 3117 14599 3137
rect 14599 3117 14616 3137
rect 14582 3103 14616 3117
rect 14431 3061 14465 3095
rect 14510 3030 14544 3064
rect 14582 3032 14599 3064
rect 14599 3032 14616 3064
rect 14582 3030 14616 3032
rect 14431 2988 14465 3022
rect 14510 2972 14544 2991
rect 14582 2972 14616 2991
rect 14510 2957 14544 2972
rect 14582 2957 14616 2972
rect 14431 2915 14465 2949
rect 14510 2884 14544 2918
rect 14582 2884 14616 2918
rect 14431 2842 14465 2876
rect 14510 2811 14544 2845
rect 14582 2811 14616 2845
rect 14431 2769 14465 2803
rect 14510 2738 14544 2772
rect 14582 2738 14616 2772
rect 14431 2696 14465 2730
rect 14510 2665 14544 2699
rect 14582 2665 14616 2699
rect 14431 2623 14465 2657
rect 14510 2592 14544 2626
rect 14582 2592 14616 2626
rect 14431 2550 14465 2584
rect 14510 2530 14544 2553
rect 14582 2530 14616 2553
rect 14510 2519 14544 2530
rect 14582 2519 14616 2530
rect 14431 2477 14465 2511
rect 14510 2446 14544 2480
rect 14582 2451 14599 2480
rect 14599 2451 14616 2480
rect 14582 2446 14616 2451
rect 14431 2433 14465 2438
rect 14431 2404 14454 2433
rect 14454 2404 14465 2433
rect 14510 2373 14544 2407
rect 14582 2403 14616 2407
rect 14582 2373 14599 2403
rect 14599 2373 14616 2403
rect 14431 2331 14454 2365
rect 14454 2331 14465 2365
rect 14510 2300 14544 2334
rect 14582 2327 14616 2334
rect 14582 2300 14599 2327
rect 14599 2300 14616 2327
rect 14431 2263 14454 2292
rect 14454 2263 14465 2292
rect 14431 2258 14465 2263
rect 14510 2226 14544 2260
rect 14582 2250 14616 2260
rect 14582 2226 14599 2250
rect 14599 2226 14616 2250
rect 14431 2195 14454 2219
rect 14454 2195 14465 2219
rect 14431 2185 14465 2195
rect 14510 2152 14544 2186
rect 14582 2156 14616 2186
rect 14582 2152 14599 2156
rect 14599 2152 14616 2156
rect 14431 2127 14454 2146
rect 14454 2127 14465 2146
rect 14431 2112 14465 2127
rect 14510 2078 14544 2112
rect 14582 2085 14616 2112
rect 14582 2078 14599 2085
rect 14599 2078 14616 2085
rect 14431 2059 14454 2073
rect 14454 2059 14465 2073
rect 14431 2039 14465 2059
rect 14510 2004 14544 2038
rect 14582 2011 14616 2038
rect 14582 2004 14599 2011
rect 14599 2004 14616 2011
rect 14431 1991 14454 2000
rect 14454 1991 14465 2000
rect 14431 1966 14465 1991
rect 14510 1930 14544 1964
rect 14582 1940 14616 1964
rect 14582 1930 14599 1940
rect 14599 1930 14616 1940
rect 14431 1923 14454 1927
rect 14454 1923 14465 1927
rect 14431 1893 14465 1923
rect 14510 1856 14544 1890
rect 14582 1866 14616 1890
rect 14582 1856 14599 1866
rect 14599 1856 14616 1866
rect 14431 1821 14465 1854
rect 14431 1820 14454 1821
rect 14454 1820 14465 1821
rect 14510 1782 14544 1816
rect 14582 1795 14616 1816
rect 14582 1782 14599 1795
rect 14599 1782 14616 1795
rect 14431 1753 14465 1781
rect 14431 1747 14454 1753
rect 14454 1747 14465 1753
rect 14510 1708 14544 1742
rect 14582 1721 14616 1742
rect 14582 1708 14599 1721
rect 14599 1708 14616 1721
rect 14431 1685 14465 1708
rect 14431 1674 14454 1685
rect 14454 1674 14465 1685
rect 14431 1617 14465 1635
rect 14510 1634 14544 1668
rect 14582 1650 14616 1668
rect 14582 1634 14599 1650
rect 14599 1634 14616 1650
rect 14431 1601 14454 1617
rect 14454 1601 14465 1617
rect 14431 1549 14465 1562
rect 14510 1560 14544 1594
rect 14582 1576 14616 1594
rect 14582 1560 14599 1576
rect 14599 1560 14616 1576
rect 14431 1528 14454 1549
rect 14454 1528 14465 1549
rect 14431 1455 14465 1489
rect 14510 1486 14544 1520
rect 14582 1505 14616 1520
rect 14582 1486 14599 1505
rect 14599 1486 14616 1505
rect 14431 1382 14465 1416
rect 14510 1412 14544 1446
rect 14582 1412 14616 1446
rect 14510 1353 14531 1372
rect 14531 1353 14544 1372
rect 14582 1353 14599 1372
rect 14599 1353 14616 1372
rect 14431 1308 14465 1342
rect 14510 1338 14544 1353
rect 14582 1338 14616 1353
rect 587 1221 621 1241
rect 587 1207 589 1221
rect 589 1207 621 1221
rect 659 1219 693 1241
rect 733 1234 767 1268
rect 659 1207 691 1219
rect 691 1207 693 1219
rect 733 1160 767 1194
rect 14510 1274 14531 1298
rect 14531 1274 14544 1298
rect 14582 1277 14599 1298
rect 14599 1277 14616 1298
rect 14431 1234 14465 1268
rect 14510 1264 14544 1274
rect 14582 1264 14616 1277
rect 14510 1194 14531 1224
rect 14531 1194 14544 1224
rect 14582 1200 14599 1224
rect 14599 1200 14616 1224
rect 14431 1160 14465 1194
rect 14510 1190 14544 1194
rect 14582 1190 14616 1200
rect 767 1114 794 1116
rect 794 1114 801 1116
rect 767 1082 801 1114
rect 840 1082 874 1116
rect 913 1082 947 1116
rect 986 1082 1020 1116
rect 1059 1082 1093 1116
rect 1132 1082 1166 1116
rect 1205 1082 1239 1116
rect 1278 1082 1312 1116
rect 1351 1082 1385 1116
rect 1424 1082 1458 1116
rect 1497 1082 1531 1116
rect 1570 1082 1604 1116
rect 1643 1082 1677 1116
rect 1716 1082 1750 1116
rect 1789 1082 1823 1116
rect 1862 1082 1896 1116
rect 1935 1082 1969 1116
rect 2008 1082 2042 1116
rect 2081 1082 2115 1116
rect 2154 1082 2188 1116
rect 2227 1082 2261 1116
rect 2300 1082 2334 1116
rect 2373 1082 2407 1116
rect 2446 1082 2480 1116
rect 2519 1082 2553 1116
rect 2592 1082 2626 1116
rect 2665 1082 2699 1116
rect 767 1010 801 1044
rect 840 1010 874 1044
rect 913 1010 947 1044
rect 986 1010 1020 1044
rect 1059 1010 1093 1044
rect 1132 1010 1166 1044
rect 1205 1010 1239 1044
rect 1278 1010 1312 1044
rect 1351 1010 1385 1044
rect 1424 1010 1458 1044
rect 1497 1010 1531 1044
rect 1570 1010 1604 1044
rect 1643 1010 1677 1044
rect 1716 1010 1750 1044
rect 1789 1010 1823 1044
rect 1862 1010 1896 1044
rect 1935 1010 1969 1044
rect 2008 1010 2042 1044
rect 2081 1010 2115 1044
rect 2154 1010 2188 1044
rect 2227 1010 2261 1044
rect 2300 1010 2334 1044
rect 2373 1010 2407 1044
rect 2446 1010 2480 1044
rect 2519 1010 2553 1044
rect 2592 1010 2626 1044
rect 2665 1010 2699 1044
rect 2738 1010 14436 1116
rect 14833 4929 14867 4963
rect 14969 4921 14990 4955
rect 14990 4921 15003 4955
rect 14833 4857 14867 4891
rect 14969 4849 14990 4883
rect 14990 4849 15003 4883
rect 14833 4785 14867 4819
rect 14969 4777 14990 4811
rect 14990 4777 15003 4811
rect 14833 4713 14867 4747
rect 14969 4705 14990 4739
rect 14990 4705 15003 4739
rect 14833 4641 14867 4675
rect 14969 4633 14990 4667
rect 14990 4633 15003 4667
rect 14833 4569 14867 4603
rect 14969 4561 14990 4595
rect 14990 4561 15003 4595
rect 14833 4497 14867 4531
rect 14969 4489 14990 4523
rect 14990 4489 15003 4523
rect 14833 4425 14867 4459
rect 14969 4417 14990 4451
rect 14990 4417 15003 4451
rect 14833 4353 14867 4387
rect 14969 4345 14990 4379
rect 14990 4345 15003 4379
rect 14833 4280 14867 4314
rect 14969 4273 14990 4307
rect 14990 4273 15003 4307
rect 14833 4207 14867 4241
rect 14969 4201 14990 4235
rect 14990 4201 15003 4235
rect 14833 4134 14867 4168
rect 14969 4129 14990 4163
rect 14990 4129 15003 4163
rect 14833 4061 14867 4095
rect 14969 4057 14990 4091
rect 14990 4057 15003 4091
rect 14833 3988 14867 4022
rect 14969 3985 14990 4019
rect 14990 3985 15003 4019
rect 14833 3915 14867 3949
rect 14969 3913 14990 3947
rect 14990 3913 15003 3947
rect 14833 3842 14867 3876
rect 14969 3841 14990 3875
rect 14990 3841 15003 3875
rect 14833 3769 14867 3803
rect 14969 3769 14990 3803
rect 14990 3769 15003 3803
rect 14833 3696 14867 3730
rect 14969 3697 14990 3731
rect 14990 3697 15003 3731
rect 14833 3623 14867 3657
rect 14969 3625 14990 3659
rect 14990 3625 15003 3659
rect 14833 3550 14867 3584
rect 14969 3553 14990 3587
rect 14990 3553 15003 3587
rect 14833 3477 14867 3511
rect 14969 3481 14990 3515
rect 14990 3481 15003 3515
rect 14833 3404 14867 3438
rect 14969 3409 14990 3443
rect 14990 3409 15003 3443
rect 14833 3331 14867 3365
rect 14969 3337 14990 3371
rect 14990 3337 15003 3371
rect 14833 3258 14867 3292
rect 14969 3265 14990 3299
rect 14990 3265 15003 3299
rect 14833 3185 14867 3219
rect 14969 3193 14990 3227
rect 14990 3193 15003 3227
rect 14833 3112 14867 3146
rect 14969 3121 14990 3155
rect 14990 3121 15003 3155
rect 14833 3039 14867 3073
rect 14969 3048 14990 3082
rect 14990 3048 15003 3082
rect 14833 2966 14867 3000
rect 14969 2975 14990 3009
rect 14990 2975 15003 3009
rect 14833 2893 14867 2927
rect 14969 2902 14990 2936
rect 14990 2902 15003 2936
rect 14833 2820 14867 2854
rect 14969 2829 14990 2863
rect 14990 2829 15003 2863
rect 14833 2747 14867 2781
rect 14969 2756 14990 2790
rect 14990 2756 15003 2790
rect 14833 2674 14867 2708
rect 14969 2683 14990 2717
rect 14990 2683 15003 2717
rect 14833 2601 14867 2635
rect 14969 2610 14990 2644
rect 14990 2610 15003 2644
rect 14833 2528 14867 2562
rect 14969 2537 14990 2571
rect 14990 2537 15003 2571
rect 14833 2455 14867 2489
rect 14969 2464 14990 2498
rect 14990 2464 15003 2498
rect 14833 2382 14867 2416
rect 14969 2391 14990 2425
rect 14990 2391 15003 2425
rect 14833 2309 14867 2343
rect 14969 2318 14990 2352
rect 14990 2318 15003 2352
rect 14833 2236 14867 2270
rect 14969 2245 14990 2279
rect 14990 2245 15003 2279
rect 14833 2163 14867 2197
rect 14969 2172 14990 2206
rect 14990 2172 15003 2206
rect 14833 2090 14867 2124
rect 14969 2099 14990 2133
rect 14990 2099 15003 2133
rect 14833 2017 14867 2051
rect 14969 2026 14990 2060
rect 14990 2026 15003 2060
rect 14833 1944 14867 1978
rect 14969 1953 14990 1987
rect 14990 1953 15003 1987
rect 14833 1871 14867 1905
rect 14969 1880 14990 1914
rect 14990 1880 15003 1914
rect 14833 1798 14867 1832
rect 14969 1807 14990 1841
rect 14990 1807 15003 1841
rect 14833 1725 14867 1759
rect 14969 1734 14990 1768
rect 14990 1734 15003 1768
rect 14833 1652 14867 1686
rect 14969 1661 14990 1695
rect 14990 1661 15003 1695
rect 14833 1579 14867 1613
rect 14969 1588 14990 1622
rect 14990 1588 15003 1622
rect 14833 1506 14867 1540
rect 14969 1515 14990 1549
rect 14990 1515 15003 1549
rect 14833 1433 14867 1467
rect 14969 1442 14990 1476
rect 14990 1442 15003 1476
rect 14833 1360 14867 1394
rect 14969 1369 14990 1403
rect 14990 1369 15003 1403
rect 14833 1287 14867 1321
rect 14969 1296 14990 1330
rect 14990 1296 15003 1330
rect 14833 1214 14867 1248
rect 14969 1223 14990 1257
rect 14990 1223 15003 1257
rect 14833 1141 14867 1175
rect 14969 1150 14990 1184
rect 14990 1150 15003 1184
rect 14833 1068 14867 1102
rect 14969 1077 14990 1111
rect 14990 1077 15003 1111
rect 14833 995 14867 1029
rect 14969 1004 14990 1038
rect 14990 1004 15003 1038
rect 233 910 267 944
rect 369 910 402 944
rect 402 910 403 944
rect 233 838 267 872
rect 369 838 402 872
rect 402 838 403 872
rect 14833 922 14867 956
rect 14969 931 14990 965
rect 14990 931 15003 965
rect 14833 849 14867 883
rect 14969 858 14990 892
rect 14990 858 15003 892
rect 212 728 232 762
rect 232 728 246 762
rect 348 729 382 749
rect 348 715 368 729
rect 368 715 382 729
rect 212 661 246 684
rect 14833 776 14867 810
rect 14969 785 14990 819
rect 14990 785 15003 819
rect 14833 703 14867 737
rect 14969 712 14990 746
rect 14990 712 15003 746
rect 212 650 232 661
rect 232 650 246 661
rect 348 660 382 664
rect 421 660 455 664
rect 494 660 528 664
rect 567 660 601 664
rect 640 660 674 664
rect 713 660 747 664
rect 786 660 820 664
rect 859 660 893 664
rect 932 660 966 664
rect 1005 660 1039 664
rect 1078 660 1112 664
rect 1151 660 1185 664
rect 1224 660 1258 664
rect 1297 660 1331 664
rect 1369 660 1403 664
rect 1441 660 1475 664
rect 1513 660 1547 664
rect 1585 660 1619 664
rect 1657 660 1691 664
rect 1729 660 1763 664
rect 1801 660 1835 664
rect 1873 660 1907 664
rect 1945 660 1979 664
rect 2017 660 2051 664
rect 2089 660 2123 664
rect 2161 660 2195 664
rect 2233 660 2267 664
rect 2305 660 2339 664
rect 2377 660 2411 664
rect 2449 660 2483 664
rect 2521 660 2555 664
rect 2593 660 2627 664
rect 2665 660 2699 664
rect 2737 660 2771 664
rect 2809 660 2843 664
rect 2881 660 2915 664
rect 2953 660 2987 664
rect 3025 660 3059 664
rect 3097 660 3131 664
rect 3169 660 3203 664
rect 3241 660 3275 664
rect 3313 660 3347 664
rect 3385 660 3419 664
rect 3457 660 3491 664
rect 3529 660 3563 664
rect 3601 660 3635 664
rect 3673 660 3707 664
rect 3745 660 3779 664
rect 3817 660 3851 664
rect 3889 660 3923 664
rect 3961 660 3995 664
rect 4033 660 4067 664
rect 4105 660 4139 664
rect 4177 660 4211 664
rect 4249 660 4283 664
rect 4321 660 4355 664
rect 4393 660 4427 664
rect 4465 660 4499 664
rect 4537 660 4571 664
rect 4609 660 4643 664
rect 4681 660 4715 664
rect 4753 660 4787 664
rect 4825 660 4859 664
rect 4897 660 4931 664
rect 4969 660 5003 664
rect 5041 660 5075 664
rect 5113 660 5147 664
rect 5185 660 5219 664
rect 5257 660 5291 664
rect 5329 660 5363 664
rect 5401 660 5435 664
rect 5473 660 5507 664
rect 5545 660 5579 664
rect 5617 660 5651 664
rect 5689 660 5723 664
rect 5761 660 5795 664
rect 5833 660 5867 664
rect 5905 660 5939 664
rect 5977 660 6011 664
rect 6049 660 6083 664
rect 6121 660 6155 664
rect 6193 660 6227 664
rect 6265 660 6299 664
rect 6337 660 6371 664
rect 6409 660 6443 664
rect 6481 660 6515 664
rect 6553 660 6587 664
rect 6625 660 6659 664
rect 6697 660 6731 664
rect 6769 660 6803 664
rect 6841 660 6875 664
rect 6913 660 6947 664
rect 6985 660 7019 664
rect 7057 660 7091 664
rect 7129 660 7163 664
rect 7201 660 7235 664
rect 7273 660 7307 664
rect 7345 660 7379 664
rect 7417 660 7451 664
rect 7489 660 7523 664
rect 7561 660 7595 664
rect 7633 660 7667 664
rect 7705 660 7739 664
rect 7777 660 7811 664
rect 7849 660 7883 664
rect 7921 660 7955 664
rect 7993 660 8027 664
rect 8065 660 8099 664
rect 8137 660 8171 664
rect 8209 660 8243 664
rect 8281 660 8315 664
rect 8353 660 8387 664
rect 8425 660 8459 664
rect 8497 660 8531 664
rect 8569 660 8603 664
rect 8641 660 8675 664
rect 8713 660 8747 664
rect 8785 660 8819 664
rect 8857 660 8891 664
rect 8929 660 8963 664
rect 9001 660 9035 664
rect 9073 660 9107 664
rect 9145 660 9179 664
rect 9217 660 9251 664
rect 9289 660 9323 664
rect 9361 660 9395 664
rect 9433 660 9467 664
rect 9505 660 9539 664
rect 9577 660 9611 664
rect 9649 660 9683 664
rect 9721 660 9755 664
rect 9793 660 9827 664
rect 9865 660 9899 664
rect 9937 660 9971 664
rect 10009 660 10043 664
rect 10081 660 10115 664
rect 10153 660 10187 664
rect 10225 660 10259 664
rect 10297 660 10331 664
rect 10369 660 10403 664
rect 10441 660 10475 664
rect 10513 660 10547 664
rect 10585 660 10619 664
rect 10657 660 10691 664
rect 10729 660 10763 664
rect 10801 660 10835 664
rect 10873 660 10907 664
rect 10945 660 10979 664
rect 11017 660 11051 664
rect 11089 660 11123 664
rect 11161 660 11195 664
rect 11233 660 11267 664
rect 11305 660 11339 664
rect 11377 660 11411 664
rect 11449 660 11483 664
rect 11521 660 11555 664
rect 11593 660 11627 664
rect 11665 660 11699 664
rect 11737 660 11771 664
rect 11809 660 11843 664
rect 11881 660 11915 664
rect 11953 660 11987 664
rect 12025 660 12059 664
rect 12097 660 12131 664
rect 12169 660 12203 664
rect 12241 660 12275 664
rect 12313 660 12347 664
rect 12385 660 12419 664
rect 12457 660 12491 664
rect 12529 660 12563 664
rect 12601 660 12635 664
rect 12673 660 12707 664
rect 12745 660 12779 664
rect 12817 660 12851 664
rect 12889 660 12923 664
rect 12961 660 12995 664
rect 13033 660 13067 664
rect 13105 660 13139 664
rect 13177 660 13211 664
rect 13249 660 13283 664
rect 13321 660 13355 664
rect 13393 660 13427 664
rect 348 630 368 660
rect 368 630 382 660
rect 421 630 455 660
rect 494 630 528 660
rect 567 630 601 660
rect 640 630 674 660
rect 713 630 747 660
rect 786 630 820 660
rect 859 630 893 660
rect 932 630 966 660
rect 1005 630 1039 660
rect 1078 630 1112 660
rect 1151 630 1185 660
rect 1224 630 1258 660
rect 1297 630 1331 660
rect 1369 630 1403 660
rect 1441 630 1475 660
rect 1513 630 1547 660
rect 1585 630 1619 660
rect 1657 630 1691 660
rect 1729 630 1763 660
rect 1801 630 1835 660
rect 1873 630 1907 660
rect 1945 630 1979 660
rect 2017 630 2051 660
rect 2089 630 2123 660
rect 2161 630 2195 660
rect 2233 630 2267 660
rect 2305 630 2339 660
rect 2377 630 2411 660
rect 2449 630 2483 660
rect 2521 630 2555 660
rect 2593 630 2627 660
rect 2665 630 2699 660
rect 2737 630 2771 660
rect 2809 630 2843 660
rect 2881 630 2915 660
rect 2953 630 2987 660
rect 3025 630 3059 660
rect 3097 630 3131 660
rect 3169 630 3203 660
rect 3241 630 3275 660
rect 3313 630 3347 660
rect 3385 630 3419 660
rect 3457 630 3491 660
rect 3529 630 3563 660
rect 3601 630 3635 660
rect 3673 630 3707 660
rect 3745 630 3779 660
rect 3817 630 3851 660
rect 3889 630 3923 660
rect 3961 630 3995 660
rect 4033 630 4067 660
rect 4105 630 4139 660
rect 4177 630 4211 660
rect 4249 630 4283 660
rect 4321 630 4355 660
rect 4393 630 4427 660
rect 4465 630 4499 660
rect 4537 630 4571 660
rect 4609 630 4643 660
rect 4681 630 4715 660
rect 4753 630 4787 660
rect 4825 630 4859 660
rect 4897 630 4931 660
rect 4969 630 5003 660
rect 5041 630 5075 660
rect 5113 630 5147 660
rect 5185 630 5219 660
rect 5257 630 5291 660
rect 5329 630 5363 660
rect 5401 630 5435 660
rect 5473 630 5507 660
rect 5545 630 5579 660
rect 5617 630 5651 660
rect 5689 630 5723 660
rect 5761 630 5795 660
rect 5833 630 5867 660
rect 5905 630 5939 660
rect 5977 630 6011 660
rect 6049 630 6083 660
rect 6121 630 6155 660
rect 6193 630 6227 660
rect 6265 630 6299 660
rect 6337 630 6371 660
rect 6409 630 6443 660
rect 6481 630 6515 660
rect 6553 630 6587 660
rect 6625 630 6659 660
rect 6697 630 6731 660
rect 6769 630 6803 660
rect 6841 630 6875 660
rect 6913 630 6947 660
rect 6985 630 7019 660
rect 7057 630 7091 660
rect 7129 630 7163 660
rect 7201 630 7235 660
rect 7273 630 7307 660
rect 7345 630 7379 660
rect 7417 630 7451 660
rect 7489 630 7523 660
rect 7561 630 7595 660
rect 7633 630 7667 660
rect 7705 630 7739 660
rect 7777 630 7811 660
rect 7849 630 7883 660
rect 7921 630 7955 660
rect 7993 630 8027 660
rect 8065 630 8099 660
rect 8137 630 8171 660
rect 8209 630 8243 660
rect 8281 630 8315 660
rect 8353 630 8387 660
rect 8425 630 8459 660
rect 8497 630 8531 660
rect 8569 630 8603 660
rect 8641 630 8675 660
rect 8713 630 8747 660
rect 8785 630 8819 660
rect 8857 630 8891 660
rect 8929 630 8963 660
rect 9001 630 9035 660
rect 9073 630 9107 660
rect 9145 630 9179 660
rect 9217 630 9251 660
rect 9289 630 9323 660
rect 9361 630 9395 660
rect 9433 630 9467 660
rect 9505 630 9539 660
rect 9577 630 9611 660
rect 9649 630 9683 660
rect 9721 630 9755 660
rect 9793 630 9827 660
rect 9865 630 9899 660
rect 9937 630 9971 660
rect 10009 630 10043 660
rect 10081 630 10115 660
rect 10153 630 10187 660
rect 10225 630 10259 660
rect 10297 630 10331 660
rect 10369 630 10403 660
rect 10441 630 10475 660
rect 10513 630 10547 660
rect 10585 630 10619 660
rect 10657 630 10691 660
rect 10729 630 10763 660
rect 10801 630 10835 660
rect 10873 630 10907 660
rect 10945 630 10979 660
rect 11017 630 11051 660
rect 11089 630 11123 660
rect 11161 630 11195 660
rect 11233 630 11267 660
rect 11305 630 11339 660
rect 11377 630 11411 660
rect 11449 630 11483 660
rect 11521 630 11555 660
rect 11593 630 11627 660
rect 11665 630 11699 660
rect 11737 630 11771 660
rect 11809 630 11843 660
rect 11881 630 11915 660
rect 11953 630 11987 660
rect 12025 630 12059 660
rect 12097 630 12131 660
rect 12169 630 12203 660
rect 12241 630 12275 660
rect 12313 630 12347 660
rect 12385 630 12419 660
rect 12457 630 12491 660
rect 12529 630 12563 660
rect 12601 630 12635 660
rect 12673 630 12707 660
rect 12745 630 12779 660
rect 12817 630 12851 660
rect 12889 630 12923 660
rect 12961 630 12982 660
rect 12982 630 12995 660
rect 13033 630 13051 660
rect 13051 630 13067 660
rect 13105 630 13120 660
rect 13120 630 13139 660
rect 13177 630 13189 660
rect 13189 630 13211 660
rect 13249 630 13258 660
rect 13258 630 13283 660
rect 13321 630 13327 660
rect 13327 630 13355 660
rect 13393 630 13396 660
rect 13396 630 13427 660
rect 212 592 246 606
rect 13465 630 13499 664
rect 13537 660 13571 664
rect 13609 660 13643 664
rect 13681 660 13715 664
rect 13753 660 13787 664
rect 13825 660 13859 664
rect 13897 660 13931 664
rect 13969 660 14003 664
rect 14041 660 14075 664
rect 14113 660 14147 664
rect 14185 660 14219 664
rect 14257 660 14291 664
rect 14329 660 14363 664
rect 14401 660 14435 664
rect 14473 660 14507 664
rect 14545 660 14579 664
rect 14617 660 14651 664
rect 14689 660 14723 664
rect 14761 660 14795 664
rect 14833 660 14867 664
rect 13537 630 13569 660
rect 13569 630 13571 660
rect 13609 630 13638 660
rect 13638 630 13643 660
rect 13681 630 13707 660
rect 13707 630 13715 660
rect 13753 630 13776 660
rect 13776 630 13787 660
rect 13825 630 13845 660
rect 13845 630 13859 660
rect 13897 630 13914 660
rect 13914 630 13931 660
rect 13969 630 13983 660
rect 13983 630 14003 660
rect 14041 630 14052 660
rect 14052 630 14075 660
rect 14113 630 14121 660
rect 14121 630 14147 660
rect 14185 630 14190 660
rect 14190 630 14219 660
rect 14257 630 14259 660
rect 14259 630 14291 660
rect 14329 630 14362 660
rect 14362 630 14363 660
rect 14401 630 14431 660
rect 14431 630 14435 660
rect 14473 630 14500 660
rect 14500 630 14507 660
rect 14545 630 14569 660
rect 14569 630 14579 660
rect 14617 630 14638 660
rect 14638 630 14651 660
rect 14689 630 14707 660
rect 14707 630 14723 660
rect 14761 630 14776 660
rect 14776 630 14795 660
rect 14833 630 14845 660
rect 14845 630 14867 660
rect 14969 639 15003 673
rect 212 572 232 592
rect 232 572 246 592
rect 14969 566 15003 600
rect 284 494 300 528
rect 300 494 318 528
rect 357 494 391 528
rect 430 494 464 528
rect 503 494 537 528
rect 576 494 610 528
rect 649 494 683 528
rect 722 494 756 528
rect 795 494 829 528
rect 868 494 902 528
rect 941 494 975 528
rect 1014 494 1048 528
rect 1087 494 1121 528
rect 1160 494 1194 528
rect 1233 494 1267 528
rect 1306 494 1340 528
rect 1379 494 1413 528
rect 1452 494 1486 528
rect 1525 494 1559 528
rect 1598 494 1632 528
rect 1671 494 1705 528
rect 1744 494 1778 528
rect 1817 494 1851 528
rect 1890 494 1924 528
rect 1963 494 1997 528
rect 2036 494 2070 528
rect 2109 494 2143 528
rect 2182 494 2216 528
rect 2255 494 2289 528
rect 2328 494 2362 528
rect 2401 494 2435 528
rect 2474 494 2508 528
rect 2547 494 2581 528
rect 2620 494 2654 528
rect 2693 494 2727 528
rect 2766 494 2800 528
rect 2839 494 2873 528
rect 2912 494 2946 528
rect 2985 494 3019 528
rect 3058 494 3092 528
rect 3131 494 3165 528
rect 3204 494 3238 528
rect 3277 494 3311 528
rect 3350 494 3384 528
rect 3423 494 3457 528
rect 3496 494 3530 528
rect 3569 494 3603 528
rect 3642 494 3676 528
rect 3715 494 3749 528
rect 3788 494 3822 528
rect 3861 494 3895 528
rect 3934 494 3968 528
rect 4007 494 4041 528
rect 4080 494 4114 528
rect 4153 494 4187 528
rect 4226 494 4260 528
rect 4299 494 4333 528
rect 4372 494 4406 528
rect 4445 494 4479 528
rect 4518 494 4552 528
rect 4591 494 4625 528
rect 4664 494 4698 528
rect 4737 494 4771 528
rect 4810 494 4844 528
rect 4883 494 4917 528
rect 4956 494 4990 528
rect 5029 494 5063 528
rect 5102 494 5136 528
rect 5175 494 5209 528
rect 5248 494 5282 528
rect 5321 494 5355 528
rect 5393 494 5427 528
rect 5465 494 5499 528
rect 5537 494 5571 528
rect 5609 494 5643 528
rect 5681 494 5715 528
rect 5753 494 5787 528
rect 5825 494 5859 528
rect 5897 494 5931 528
rect 5969 494 6003 528
rect 6041 494 6075 528
rect 6113 494 6147 528
rect 6185 494 6219 528
rect 6257 494 6291 528
rect 6329 494 6363 528
rect 6401 494 6435 528
rect 6473 494 6507 528
rect 6545 494 6579 528
rect 6617 494 6651 528
rect 6689 494 6723 528
rect 6761 494 6795 528
rect 6833 494 6867 528
rect 6905 494 6939 528
rect 6977 494 7011 528
rect 7049 494 7083 528
rect 7121 494 7155 528
rect 7193 494 7227 528
rect 7265 494 7299 528
rect 7337 494 7371 528
rect 7409 494 7443 528
rect 7481 494 7515 528
rect 7553 494 7587 528
rect 7625 494 7659 528
rect 7697 494 7731 528
rect 7769 494 7803 528
rect 7841 494 7875 528
rect 7913 494 7947 528
rect 7985 494 8019 528
rect 8057 494 8091 528
rect 8129 494 8163 528
rect 8201 494 8235 528
rect 8273 494 8307 528
rect 8345 494 8379 528
rect 8417 494 8451 528
rect 8489 494 8523 528
rect 8561 494 8595 528
rect 8633 494 8667 528
rect 8705 494 8739 528
rect 8777 494 8811 528
rect 8849 494 8883 528
rect 8921 494 8955 528
rect 8993 494 9027 528
rect 9065 494 9099 528
rect 9137 494 9171 528
rect 9209 494 9243 528
rect 9281 494 9315 528
rect 9353 494 9387 528
rect 9425 494 9459 528
rect 9497 494 9531 528
rect 9569 494 9603 528
rect 9641 494 9675 528
rect 9713 494 9747 528
rect 9785 494 9819 528
rect 9857 494 9891 528
rect 9929 494 9963 528
rect 10001 494 10035 528
rect 10073 494 10107 528
rect 10145 494 10179 528
rect 10217 494 10251 528
rect 10289 494 10323 528
rect 10361 494 10395 528
rect 10433 494 10467 528
rect 10505 494 10539 528
rect 10577 494 10611 528
rect 10649 494 10683 528
rect 10721 494 10755 528
rect 10793 494 10827 528
rect 10865 494 10899 528
rect 10937 494 10971 528
rect 11009 494 11043 528
rect 11081 494 11115 528
rect 11153 494 11187 528
rect 11225 494 11259 528
rect 11297 494 11331 528
rect 11369 494 11403 528
rect 11441 494 11475 528
rect 11513 494 11547 528
rect 11585 494 11619 528
rect 11657 494 11691 528
rect 11729 494 11763 528
rect 11801 494 11835 528
rect 11873 494 11907 528
rect 11945 494 11979 528
rect 12017 494 12051 528
rect 12089 494 12123 528
rect 12161 494 12195 528
rect 12233 494 12267 528
rect 12305 494 12339 528
rect 12377 494 12411 528
rect 12449 494 12483 528
rect 12521 494 12555 528
rect 12593 494 12627 528
rect 12665 494 12699 528
rect 12737 494 12771 528
rect 12809 494 12843 528
rect 12881 494 12915 528
rect 12953 494 12982 528
rect 12982 494 12987 528
rect 13025 524 13059 528
rect 13097 524 13131 528
rect 13169 524 13203 528
rect 13241 524 13275 528
rect 13313 524 13347 528
rect 13385 524 13419 528
rect 13457 524 13491 528
rect 13529 524 13563 528
rect 13601 524 13635 528
rect 13025 494 13051 524
rect 13051 494 13059 524
rect 13097 494 13120 524
rect 13120 494 13131 524
rect 13169 494 13189 524
rect 13189 494 13203 524
rect 13241 494 13258 524
rect 13258 494 13275 524
rect 13313 494 13327 524
rect 13327 494 13347 524
rect 13385 494 13396 524
rect 13396 494 13419 524
rect 13457 494 13465 524
rect 13465 494 13491 524
rect 13529 494 13534 524
rect 13534 494 13563 524
rect 13601 494 13603 524
rect 13603 494 13635 524
rect 13673 494 13707 528
rect 13745 524 13779 528
rect 13817 524 13851 528
rect 13889 524 13923 528
rect 13961 524 13995 528
rect 14033 524 14067 528
rect 14105 524 14139 528
rect 14177 524 14211 528
rect 14249 524 14283 528
rect 14321 524 14355 528
rect 14393 524 14427 528
rect 14465 524 14499 528
rect 14537 524 14571 528
rect 14609 524 14643 528
rect 14681 524 14715 528
rect 14753 524 14787 528
rect 14825 524 14859 528
rect 14897 524 14931 528
rect 13745 494 13776 524
rect 13776 494 13779 524
rect 13817 494 13845 524
rect 13845 494 13851 524
rect 13889 494 13914 524
rect 13914 494 13923 524
rect 13961 494 13983 524
rect 13983 494 13995 524
rect 14033 494 14052 524
rect 14052 494 14067 524
rect 14105 494 14121 524
rect 14121 494 14139 524
rect 14177 494 14190 524
rect 14190 494 14211 524
rect 14249 494 14259 524
rect 14259 494 14283 524
rect 14321 494 14328 524
rect 14328 494 14355 524
rect 14393 494 14397 524
rect 14397 494 14427 524
rect 14465 494 14466 524
rect 14466 494 14499 524
rect 14537 494 14569 524
rect 14569 494 14571 524
rect 14609 494 14638 524
rect 14638 494 14643 524
rect 14681 494 14707 524
rect 14707 494 14715 524
rect 14753 494 14776 524
rect 14776 494 14787 524
rect 14825 494 14845 524
rect 14845 494 14859 524
rect 14897 494 14914 524
rect 14914 494 14931 524
<< metal1 >>
rect 59 5459 15117 5465
rect 59 5425 305 5459
rect 339 5425 377 5459
rect 411 5425 449 5459
rect 483 5425 521 5459
rect 555 5425 593 5459
rect 627 5425 665 5459
rect 699 5425 737 5459
rect 771 5425 809 5459
rect 843 5425 881 5459
rect 915 5425 953 5459
rect 987 5425 1025 5459
rect 1059 5425 1097 5459
rect 1131 5425 1169 5459
rect 1203 5425 1241 5459
rect 1275 5425 1313 5459
rect 1347 5425 1385 5459
rect 1419 5425 1457 5459
rect 1491 5425 1529 5459
rect 1563 5425 1601 5459
rect 1635 5425 1673 5459
rect 1707 5425 1745 5459
rect 1779 5425 1817 5459
rect 1851 5425 1889 5459
rect 1923 5425 1961 5459
rect 1995 5425 2033 5459
rect 2067 5425 2105 5459
rect 2139 5425 2177 5459
rect 2211 5425 2249 5459
rect 2283 5425 2321 5459
rect 2355 5425 2393 5459
rect 2427 5425 2465 5459
rect 2499 5425 2537 5459
rect 2571 5425 2609 5459
rect 2643 5425 2681 5459
rect 2715 5425 2753 5459
rect 2787 5425 2825 5459
rect 2859 5425 2897 5459
rect 2931 5425 2969 5459
rect 3003 5425 3041 5459
rect 3075 5425 3113 5459
rect 3147 5425 3185 5459
rect 3219 5425 3257 5459
rect 3291 5425 3329 5459
rect 3363 5425 3401 5459
rect 3435 5425 3473 5459
rect 3507 5425 3545 5459
rect 3579 5425 3617 5459
rect 3651 5425 3689 5459
rect 3723 5425 3761 5459
rect 3795 5425 3833 5459
rect 3867 5425 3905 5459
rect 3939 5425 3977 5459
rect 4011 5425 4049 5459
rect 4083 5425 4121 5459
rect 4155 5425 4193 5459
rect 4227 5425 4265 5459
rect 4299 5425 4337 5459
rect 4371 5425 4409 5459
rect 4443 5425 4481 5459
rect 4515 5425 4553 5459
rect 4587 5425 4625 5459
rect 4659 5425 4697 5459
rect 4731 5425 4769 5459
rect 4803 5425 4841 5459
rect 4875 5425 4913 5459
rect 4947 5425 4985 5459
rect 5019 5425 5057 5459
rect 5091 5425 5129 5459
rect 5163 5425 5201 5459
rect 5235 5425 5273 5459
rect 5307 5425 5345 5459
rect 5379 5425 5417 5459
rect 5451 5425 5489 5459
rect 5523 5425 5561 5459
rect 5595 5425 5633 5459
rect 5667 5425 5705 5459
rect 5739 5425 5777 5459
rect 5811 5425 5849 5459
rect 5883 5425 5921 5459
rect 5955 5425 5993 5459
rect 6027 5425 6065 5459
rect 6099 5425 6137 5459
rect 6171 5425 6209 5459
rect 6243 5425 6281 5459
rect 6315 5425 6353 5459
rect 6387 5425 6425 5459
rect 6459 5425 6497 5459
rect 6531 5425 6569 5459
rect 6603 5425 6641 5459
rect 6675 5425 6713 5459
rect 6747 5425 6785 5459
rect 6819 5425 6857 5459
rect 6891 5425 6929 5459
rect 6963 5425 7001 5459
rect 7035 5425 7073 5459
rect 7107 5425 7145 5459
rect 7179 5425 7217 5459
rect 7251 5425 7289 5459
rect 7323 5425 7361 5459
rect 7395 5425 7433 5459
rect 7467 5425 7505 5459
rect 7539 5425 7577 5459
rect 7611 5425 7649 5459
rect 7683 5425 7721 5459
rect 7755 5425 7793 5459
rect 7827 5425 7865 5459
rect 7899 5425 7937 5459
rect 7971 5425 8009 5459
rect 8043 5425 8081 5459
rect 8115 5425 8153 5459
rect 8187 5425 8225 5459
rect 8259 5425 8297 5459
rect 8331 5425 8369 5459
rect 8403 5425 8441 5459
rect 8475 5425 8513 5459
rect 8547 5425 8585 5459
rect 8619 5425 8657 5459
rect 8691 5425 8729 5459
rect 8763 5425 8801 5459
rect 8835 5425 8873 5459
rect 8907 5425 8945 5459
rect 8979 5425 9017 5459
rect 9051 5425 9089 5459
rect 9123 5425 9161 5459
rect 9195 5425 9233 5459
rect 9267 5425 9305 5459
rect 9339 5425 9377 5459
rect 9411 5425 9449 5459
rect 9483 5425 9521 5459
rect 9555 5425 9593 5459
rect 9627 5425 9665 5459
rect 9699 5425 9737 5459
rect 9771 5425 9809 5459
rect 9843 5425 9881 5459
rect 9915 5425 9953 5459
rect 9987 5425 10025 5459
rect 10059 5425 10097 5459
rect 10131 5425 10169 5459
rect 10203 5425 10241 5459
rect 10275 5425 10313 5459
rect 10347 5425 10385 5459
rect 10419 5425 10457 5459
rect 10491 5425 10529 5459
rect 10563 5425 10601 5459
rect 10635 5425 10673 5459
rect 10707 5425 10745 5459
rect 10779 5425 10817 5459
rect 10851 5425 10889 5459
rect 10923 5425 10961 5459
rect 10995 5425 11033 5459
rect 11067 5425 11105 5459
rect 11139 5425 11177 5459
rect 11211 5425 11249 5459
rect 11283 5425 11321 5459
rect 11355 5425 11393 5459
rect 11427 5425 11466 5459
rect 11500 5425 11539 5459
rect 11573 5425 11612 5459
rect 11646 5425 11685 5459
rect 11719 5425 11758 5459
rect 11792 5425 11831 5459
rect 11865 5425 11904 5459
rect 11938 5425 11977 5459
rect 12011 5425 12050 5459
rect 12084 5425 12123 5459
rect 12157 5425 12196 5459
rect 12230 5425 12269 5459
rect 12303 5425 12342 5459
rect 12376 5425 12415 5459
rect 12449 5425 12488 5459
rect 12522 5425 12561 5459
rect 12595 5425 12634 5459
rect 12668 5425 12707 5459
rect 12741 5425 12780 5459
rect 12814 5425 12853 5459
rect 12887 5425 12926 5459
rect 12960 5425 12999 5459
rect 13033 5425 13072 5459
rect 13106 5425 13145 5459
rect 13179 5425 13218 5459
rect 13252 5425 13291 5459
rect 13325 5425 13364 5459
rect 13398 5425 13437 5459
rect 13471 5425 13510 5459
rect 13544 5425 13583 5459
rect 13617 5425 13656 5459
rect 13690 5425 13729 5459
rect 13763 5425 13802 5459
rect 13836 5425 13875 5459
rect 13909 5425 13948 5459
rect 13982 5425 14021 5459
rect 14055 5425 14094 5459
rect 14128 5425 14167 5459
rect 14201 5425 14240 5459
rect 14274 5425 14313 5459
rect 14347 5425 14386 5459
rect 14420 5425 14459 5459
rect 14493 5425 14532 5459
rect 14566 5425 14605 5459
rect 14639 5425 14678 5459
rect 14712 5425 14751 5459
rect 14785 5425 14824 5459
rect 14858 5425 14897 5459
rect 14931 5425 15117 5459
rect 59 5387 15117 5425
rect 59 5353 233 5387
rect 267 5353 14969 5387
rect 15003 5353 15117 5387
rect 59 5323 15117 5353
rect 59 5314 369 5323
rect 59 5280 233 5314
rect 267 5289 369 5314
rect 403 5289 441 5323
rect 475 5289 513 5323
rect 547 5289 585 5323
rect 619 5289 657 5323
rect 691 5289 729 5323
rect 763 5289 801 5323
rect 835 5289 873 5323
rect 907 5289 945 5323
rect 979 5289 1017 5323
rect 1051 5289 1089 5323
rect 1123 5289 1161 5323
rect 1195 5289 1233 5323
rect 1267 5289 1305 5323
rect 1339 5289 1377 5323
rect 1411 5289 1449 5323
rect 1483 5289 1521 5323
rect 1555 5289 1593 5323
rect 1627 5289 1665 5323
rect 1699 5289 1737 5323
rect 1771 5289 1809 5323
rect 1843 5289 1881 5323
rect 1915 5289 1953 5323
rect 1987 5289 2025 5323
rect 2059 5289 2097 5323
rect 2131 5289 2169 5323
rect 2203 5289 2241 5323
rect 2275 5289 2313 5323
rect 2347 5289 2385 5323
rect 2419 5289 2457 5323
rect 2491 5289 2529 5323
rect 2563 5289 2601 5323
rect 2635 5289 2673 5323
rect 2707 5289 2745 5323
rect 2779 5289 2817 5323
rect 2851 5289 2889 5323
rect 2923 5289 2961 5323
rect 2995 5289 3033 5323
rect 3067 5289 3105 5323
rect 3139 5289 3177 5323
rect 3211 5289 3249 5323
rect 3283 5289 3321 5323
rect 3355 5289 3393 5323
rect 3427 5289 3465 5323
rect 3499 5289 3537 5323
rect 3571 5289 3609 5323
rect 3643 5289 3681 5323
rect 3715 5289 3753 5323
rect 3787 5289 3825 5323
rect 3859 5289 3897 5323
rect 3931 5289 3969 5323
rect 4003 5289 4041 5323
rect 4075 5289 4113 5323
rect 4147 5289 4185 5323
rect 4219 5289 4257 5323
rect 4291 5289 4329 5323
rect 4363 5289 4401 5323
rect 4435 5289 4473 5323
rect 4507 5289 4545 5323
rect 4579 5289 4617 5323
rect 4651 5289 4689 5323
rect 4723 5289 4761 5323
rect 4795 5289 4833 5323
rect 4867 5289 4905 5323
rect 4939 5289 4977 5323
rect 5011 5289 5049 5323
rect 5083 5289 5121 5323
rect 5155 5289 5193 5323
rect 5227 5289 5265 5323
rect 5299 5289 5337 5323
rect 5371 5289 5409 5323
rect 5443 5289 5481 5323
rect 5515 5289 5553 5323
rect 5587 5289 5625 5323
rect 5659 5289 5697 5323
rect 5731 5289 5769 5323
rect 5803 5289 5841 5323
rect 5875 5289 5913 5323
rect 5947 5289 5985 5323
rect 6019 5289 6057 5323
rect 6091 5289 6129 5323
rect 6163 5289 6201 5323
rect 6235 5289 6273 5323
rect 6307 5289 6345 5323
rect 6379 5289 6417 5323
rect 6451 5289 6489 5323
rect 6523 5289 6561 5323
rect 6595 5289 6633 5323
rect 6667 5289 6705 5323
rect 6739 5289 6777 5323
rect 6811 5289 6849 5323
rect 6883 5289 6921 5323
rect 6955 5289 6993 5323
rect 7027 5289 7065 5323
rect 7099 5289 7137 5323
rect 7171 5289 7209 5323
rect 7243 5289 7281 5323
rect 7315 5289 7353 5323
rect 7387 5289 7425 5323
rect 7459 5289 7497 5323
rect 7531 5289 7569 5323
rect 7603 5289 7641 5323
rect 7675 5289 7713 5323
rect 7747 5289 7785 5323
rect 7819 5289 7857 5323
rect 7891 5289 7929 5323
rect 7963 5289 8001 5323
rect 8035 5289 8073 5323
rect 8107 5289 8145 5323
rect 8179 5289 8217 5323
rect 8251 5289 8289 5323
rect 8323 5289 8361 5323
rect 8395 5289 8433 5323
rect 8467 5289 8505 5323
rect 8539 5289 8577 5323
rect 8611 5289 8649 5323
rect 8683 5289 8721 5323
rect 8755 5289 8793 5323
rect 8827 5289 8865 5323
rect 8899 5289 8937 5323
rect 8971 5289 9009 5323
rect 9043 5289 9081 5323
rect 9115 5289 9153 5323
rect 9187 5289 9225 5323
rect 9259 5289 9297 5323
rect 9331 5289 9369 5323
rect 9403 5289 9441 5323
rect 9475 5289 9513 5323
rect 9547 5289 9585 5323
rect 9619 5289 9657 5323
rect 9691 5289 9729 5323
rect 9763 5289 9801 5323
rect 9835 5289 9873 5323
rect 9907 5289 9945 5323
rect 9979 5289 10017 5323
rect 10051 5289 10089 5323
rect 10123 5289 10161 5323
rect 10195 5289 10234 5323
rect 10268 5289 10307 5323
rect 10341 5289 10380 5323
rect 10414 5289 10453 5323
rect 10487 5289 10526 5323
rect 10560 5289 10599 5323
rect 10633 5289 10672 5323
rect 10706 5289 10745 5323
rect 10779 5289 10818 5323
rect 10852 5289 10891 5323
rect 10925 5289 10964 5323
rect 10998 5289 11037 5323
rect 11071 5289 11110 5323
rect 11144 5289 11183 5323
rect 11217 5289 11256 5323
rect 11290 5289 11329 5323
rect 11363 5289 11402 5323
rect 11436 5289 11475 5323
rect 11509 5289 11548 5323
rect 11582 5289 11621 5323
rect 11655 5289 11694 5323
rect 11728 5289 11767 5323
rect 11801 5289 11840 5323
rect 11874 5289 11913 5323
rect 11947 5289 11986 5323
rect 12020 5289 12059 5323
rect 12093 5289 12132 5323
rect 12166 5289 12205 5323
rect 12239 5289 12278 5323
rect 12312 5289 12351 5323
rect 12385 5289 12424 5323
rect 12458 5289 12497 5323
rect 12531 5289 12570 5323
rect 12604 5289 12643 5323
rect 12677 5289 12716 5323
rect 12750 5289 12789 5323
rect 12823 5289 12862 5323
rect 12896 5289 12935 5323
rect 12969 5289 13008 5323
rect 13042 5289 13081 5323
rect 13115 5289 13154 5323
rect 13188 5289 13227 5323
rect 13261 5289 13300 5323
rect 13334 5289 13373 5323
rect 13407 5289 13446 5323
rect 13480 5289 13519 5323
rect 13553 5289 13592 5323
rect 13626 5289 13665 5323
rect 13699 5289 13738 5323
rect 13772 5289 13811 5323
rect 13845 5289 13884 5323
rect 13918 5289 13957 5323
rect 13991 5289 14030 5323
rect 14064 5289 14103 5323
rect 14137 5289 14176 5323
rect 14210 5289 14249 5323
rect 14283 5289 14322 5323
rect 14356 5289 14395 5323
rect 14429 5289 14468 5323
rect 14502 5289 14541 5323
rect 14575 5289 14614 5323
rect 14648 5289 14687 5323
rect 14721 5289 14760 5323
rect 14794 5289 14833 5323
rect 14867 5315 15117 5323
rect 14867 5289 14969 5315
rect 267 5281 14969 5289
rect 15003 5281 15117 5315
rect 267 5280 15117 5281
rect 59 5255 15117 5280
rect 59 5251 552 5255
tri 552 5251 556 5255 nw
tri 14619 5251 14623 5255 ne
rect 14623 5251 15117 5255
rect 59 5250 518 5251
rect 59 5241 369 5250
rect 59 5207 233 5241
rect 267 5216 369 5241
rect 403 5217 518 5250
tri 518 5217 552 5251 nw
tri 14623 5217 14657 5251 ne
rect 14657 5217 14833 5251
rect 14867 5243 15117 5251
rect 14867 5217 14969 5243
rect 403 5216 510 5217
rect 267 5209 510 5216
tri 510 5209 518 5217 nw
tri 14657 5209 14665 5217 ne
rect 14665 5209 14969 5217
rect 15003 5209 15117 5243
rect 267 5207 480 5209
rect 59 5179 480 5207
tri 480 5179 510 5209 nw
tri 14665 5179 14695 5209 ne
rect 14695 5179 15117 5209
rect 59 5177 446 5179
rect 59 5168 369 5177
rect 59 5134 233 5168
rect 267 5143 369 5168
rect 403 5145 446 5177
tri 446 5145 480 5179 nw
tri 14695 5145 14729 5179 ne
rect 14729 5145 14833 5179
rect 14867 5171 15117 5179
rect 14867 5145 14969 5171
rect 403 5143 438 5145
rect 267 5137 438 5143
tri 438 5137 446 5145 nw
tri 14729 5137 14737 5145 ne
rect 14737 5137 14969 5145
rect 15003 5137 15117 5171
rect 267 5134 409 5137
rect 59 5104 409 5134
tri 409 5108 438 5137 nw
tri 14737 5108 14766 5137 ne
rect 14766 5108 15117 5137
tri 14766 5107 14767 5108 ne
rect 14767 5107 15117 5108
rect 59 5095 369 5104
rect 59 5061 233 5095
rect 267 5070 369 5095
rect 403 5070 409 5104
tri 14767 5073 14801 5107 ne
rect 14801 5073 14833 5107
rect 14867 5099 15117 5107
rect 14867 5073 14969 5099
rect 267 5061 409 5070
tri 14801 5065 14809 5073 ne
rect 14809 5065 14969 5073
rect 15003 5065 15117 5099
rect 59 5031 409 5061
tri 14809 5056 14818 5065 ne
rect 59 5022 369 5031
rect 59 4988 233 5022
rect 267 4997 369 5022
rect 403 4997 409 5031
rect 267 4988 409 4997
rect 59 4958 409 4988
rect 59 4949 369 4958
rect 59 4915 233 4949
rect 267 4924 369 4949
rect 403 4924 409 4958
rect 14818 5035 15117 5065
rect 14818 5001 14833 5035
rect 14867 5027 15117 5035
rect 14867 5001 14969 5027
rect 14818 4993 14969 5001
rect 15003 4993 15117 5027
rect 14818 4963 15117 4993
tri 684 4929 691 4936 se
rect 691 4929 14512 4936
tri 14512 4929 14519 4936 sw
rect 14818 4929 14833 4963
rect 14867 4955 15117 4963
rect 14867 4929 14969 4955
tri 679 4924 684 4929 se
rect 684 4924 14519 4929
rect 267 4915 409 4924
rect 59 4885 409 4915
rect 59 4876 369 4885
rect 59 4842 233 4876
rect 267 4851 369 4876
rect 403 4851 409 4885
rect 267 4842 409 4851
rect 59 4812 409 4842
rect 59 4803 369 4812
rect 59 4769 233 4803
rect 267 4778 369 4803
rect 403 4778 409 4812
rect 267 4769 409 4778
rect 59 4739 409 4769
rect 59 4730 369 4739
rect 59 4696 233 4730
rect 267 4705 369 4730
rect 403 4705 409 4739
rect 267 4696 409 4705
rect 59 4666 409 4696
rect 59 4657 369 4666
rect 59 4623 233 4657
rect 267 4632 369 4657
rect 403 4632 409 4666
rect 267 4623 409 4632
rect 59 4593 409 4623
rect 59 4584 369 4593
rect 59 4550 233 4584
rect 267 4559 369 4584
rect 403 4559 409 4593
rect 267 4550 409 4559
rect 59 4520 409 4550
rect 59 4511 369 4520
rect 59 4477 233 4511
rect 267 4486 369 4511
rect 403 4486 409 4520
rect 267 4477 409 4486
rect 59 4447 409 4477
rect 59 4438 369 4447
rect 59 4404 233 4438
rect 267 4413 369 4438
rect 403 4413 409 4447
rect 267 4404 409 4413
rect 59 4374 409 4404
rect 59 4365 369 4374
rect 59 4331 233 4365
rect 267 4340 369 4365
rect 403 4340 409 4374
rect 267 4331 409 4340
rect 59 4301 409 4331
rect 59 4292 369 4301
rect 59 4258 233 4292
rect 267 4267 369 4292
rect 403 4267 409 4301
rect 267 4258 409 4267
rect 59 4228 409 4258
rect 59 4219 369 4228
rect 59 4185 233 4219
rect 267 4194 369 4219
rect 403 4194 409 4228
rect 267 4185 409 4194
rect 59 4155 409 4185
rect 59 4146 369 4155
rect 59 4112 233 4146
rect 267 4121 369 4146
rect 403 4121 409 4155
rect 267 4112 409 4121
rect 59 4082 409 4112
rect 59 4073 369 4082
rect 59 4039 233 4073
rect 267 4048 369 4073
rect 403 4048 409 4082
rect 267 4039 409 4048
rect 59 4009 409 4039
rect 59 4000 369 4009
rect 59 3966 233 4000
rect 267 3975 369 4000
rect 403 3975 409 4009
rect 267 3966 409 3975
rect 59 3936 409 3966
rect 59 3927 369 3936
rect 59 3893 233 3927
rect 267 3902 369 3927
rect 403 3902 409 3936
rect 267 3893 409 3902
rect 59 3863 409 3893
rect 59 3854 369 3863
rect 59 3820 233 3854
rect 267 3829 369 3854
rect 403 3829 409 3863
rect 267 3820 409 3829
rect 59 3790 409 3820
rect 59 3781 369 3790
rect 59 3747 233 3781
rect 267 3756 369 3781
rect 403 3756 409 3790
rect 267 3747 409 3756
rect 59 3717 409 3747
rect 59 3708 369 3717
rect 59 3674 233 3708
rect 267 3683 369 3708
rect 403 3683 409 3717
rect 267 3674 409 3683
rect 59 3644 409 3674
rect 59 3635 369 3644
rect 59 3601 233 3635
rect 267 3610 369 3635
rect 403 3610 409 3644
rect 267 3601 409 3610
rect 59 3571 409 3601
rect 59 3562 369 3571
rect 59 3528 233 3562
rect 267 3537 369 3562
rect 403 3537 409 3571
rect 267 3528 409 3537
rect 59 3498 409 3528
rect 59 3489 369 3498
rect 59 3455 233 3489
rect 267 3464 369 3489
rect 403 3464 409 3498
rect 267 3455 409 3464
rect 59 3425 409 3455
rect 59 3416 369 3425
rect 59 3382 233 3416
rect 267 3391 369 3416
rect 403 3391 409 3425
rect 267 3382 409 3391
rect 59 3352 409 3382
rect 59 3343 369 3352
rect 59 3309 233 3343
rect 267 3318 369 3343
rect 403 3318 409 3352
rect 267 3309 409 3318
rect 59 3279 409 3309
rect 59 3270 369 3279
rect 59 3236 233 3270
rect 267 3245 369 3270
rect 403 3245 409 3279
rect 267 3236 409 3245
rect 59 3206 409 3236
rect 59 3197 369 3206
rect 59 3163 233 3197
rect 267 3172 369 3197
rect 403 3172 409 3206
rect 267 3163 409 3172
rect 59 3133 409 3163
rect 59 3124 369 3133
rect 59 3090 233 3124
rect 267 3099 369 3124
rect 403 3099 409 3133
rect 267 3090 409 3099
rect 59 3060 409 3090
rect 59 3051 369 3060
rect 59 3017 233 3051
rect 267 3026 369 3051
rect 403 3026 409 3060
rect 267 3017 409 3026
rect 59 2987 409 3017
rect 59 2978 369 2987
rect 59 2944 233 2978
rect 267 2953 369 2978
rect 403 2953 409 2987
rect 267 2944 409 2953
rect 59 2914 409 2944
rect 59 2905 369 2914
rect 59 2871 233 2905
rect 267 2880 369 2905
rect 403 2880 409 2914
rect 267 2871 409 2880
rect 59 2841 409 2871
rect 59 2832 369 2841
rect 59 2798 233 2832
rect 267 2807 369 2832
rect 403 2807 409 2841
rect 267 2798 409 2807
rect 59 2768 409 2798
rect 59 2759 369 2768
rect 59 2725 233 2759
rect 267 2734 369 2759
rect 403 2734 409 2768
rect 267 2725 409 2734
rect 59 2695 409 2725
rect 59 2686 369 2695
rect 59 2652 233 2686
rect 267 2661 369 2686
rect 403 2661 409 2695
rect 267 2652 409 2661
rect 59 2622 409 2652
rect 59 2613 369 2622
rect 59 2579 233 2613
rect 267 2588 369 2613
rect 403 2588 409 2622
rect 267 2579 409 2588
rect 59 2549 409 2579
rect 59 2540 369 2549
rect 59 2506 233 2540
rect 267 2515 369 2540
rect 403 2515 409 2549
rect 267 2506 409 2515
rect 59 2476 409 2506
rect 59 2467 369 2476
rect 59 2433 233 2467
rect 267 2442 369 2467
rect 403 2442 409 2476
rect 267 2433 409 2442
rect 59 2403 409 2433
rect 59 2394 369 2403
rect 59 2360 233 2394
rect 267 2369 369 2394
rect 403 2369 409 2403
rect 267 2360 409 2369
rect 59 2330 409 2360
rect 59 2321 369 2330
rect 59 2287 233 2321
rect 267 2296 369 2321
rect 403 2296 409 2330
rect 267 2287 409 2296
rect 59 2257 409 2287
rect 59 2248 369 2257
rect 59 2214 233 2248
rect 267 2223 369 2248
rect 403 2223 409 2257
rect 267 2214 409 2223
rect 59 2184 409 2214
rect 59 2175 369 2184
rect 59 2141 233 2175
rect 267 2150 369 2175
rect 403 2150 409 2184
rect 267 2141 409 2150
rect 59 2111 409 2141
rect 59 2102 369 2111
rect 59 2068 233 2102
rect 267 2077 369 2102
rect 403 2077 409 2111
rect 267 2068 409 2077
rect 59 2038 409 2068
rect 59 2029 369 2038
rect 59 1995 233 2029
rect 267 2004 369 2029
rect 403 2004 409 2038
rect 267 1995 409 2004
rect 59 1965 409 1995
rect 59 1956 369 1965
rect 59 1922 233 1956
rect 267 1931 369 1956
rect 403 1931 409 1965
rect 267 1922 409 1931
rect 59 1892 409 1922
rect 59 1883 369 1892
rect 59 1849 233 1883
rect 267 1858 369 1883
rect 403 1858 409 1892
rect 267 1849 409 1858
rect 59 1819 409 1849
rect 59 1810 369 1819
rect 59 1776 233 1810
rect 267 1785 369 1810
rect 403 1785 409 1819
rect 267 1776 409 1785
rect 59 1746 409 1776
rect 59 1737 369 1746
rect 59 1703 233 1737
rect 267 1712 369 1737
rect 403 1712 409 1746
rect 267 1703 409 1712
rect 59 1673 409 1703
rect 59 1664 369 1673
rect 59 1630 233 1664
rect 267 1639 369 1664
rect 403 1639 409 1673
rect 267 1630 409 1639
rect 59 1600 409 1630
rect 59 1592 369 1600
rect 59 1558 233 1592
rect 267 1566 369 1592
rect 403 1566 409 1600
rect 267 1558 409 1566
rect 59 1527 409 1558
rect 59 1520 369 1527
rect 59 1486 233 1520
rect 267 1493 369 1520
rect 403 1493 409 1527
rect 267 1486 409 1493
rect 59 1454 409 1486
rect 59 1448 369 1454
rect 59 1414 233 1448
rect 267 1420 369 1448
rect 403 1420 409 1454
rect 267 1414 409 1420
rect 59 1381 409 1414
rect 59 1376 369 1381
rect 59 1342 233 1376
rect 267 1347 369 1376
rect 403 1347 409 1381
rect 267 1342 409 1347
rect 59 1308 409 1342
rect 59 1304 369 1308
rect 59 1270 233 1304
rect 267 1274 369 1304
rect 403 1274 409 1308
rect 267 1270 409 1274
rect 59 1235 409 1270
rect 59 1232 369 1235
rect 59 1198 233 1232
rect 267 1201 369 1232
rect 403 1201 409 1235
rect 267 1198 409 1201
rect 59 1162 409 1198
rect 59 1160 369 1162
rect 59 1126 233 1160
rect 267 1128 369 1160
rect 403 1128 409 1162
rect 267 1126 409 1128
rect 59 1089 409 1126
rect 59 1088 369 1089
rect 59 1054 233 1088
rect 267 1055 369 1088
rect 403 1055 409 1089
tri 575 4820 679 4924 se
rect 679 4820 767 4924
rect 575 4818 767 4820
rect 12465 4890 12504 4924
rect 12538 4890 12577 4924
rect 12611 4890 12650 4924
rect 12684 4890 12723 4924
rect 12757 4890 12796 4924
rect 12830 4890 12869 4924
rect 12903 4890 12942 4924
rect 12976 4890 13015 4924
rect 13049 4890 13088 4924
rect 13122 4890 13161 4924
rect 13195 4890 13234 4924
rect 13268 4890 13307 4924
rect 13341 4890 13380 4924
rect 13414 4890 13453 4924
rect 13487 4890 13526 4924
rect 13560 4890 13599 4924
rect 13633 4890 13672 4924
rect 13706 4890 13745 4924
rect 13779 4890 13818 4924
rect 13852 4890 13891 4924
rect 13925 4890 13964 4924
rect 13998 4890 14037 4924
rect 14071 4890 14110 4924
rect 14144 4890 14183 4924
rect 14217 4890 14256 4924
rect 14290 4890 14329 4924
rect 14363 4890 14402 4924
rect 14436 4921 14519 4924
tri 14519 4921 14527 4929 sw
rect 14818 4921 14969 4929
rect 15003 4921 15117 4955
rect 14436 4891 14527 4921
tri 14527 4891 14557 4921 sw
rect 14818 4891 15117 4921
rect 14436 4890 14557 4891
rect 12465 4857 14557 4890
tri 14557 4857 14591 4891 sw
rect 14818 4857 14833 4891
rect 14867 4883 15117 4891
rect 14867 4857 14969 4883
rect 12465 4852 14591 4857
rect 12465 4818 12504 4852
rect 12538 4818 12577 4852
rect 12611 4818 12650 4852
rect 12684 4818 12723 4852
rect 12757 4818 12796 4852
rect 12830 4818 12869 4852
rect 12903 4818 12942 4852
rect 12976 4818 13015 4852
rect 13049 4818 13088 4852
rect 13122 4818 13161 4852
rect 13195 4818 13234 4852
rect 13268 4818 13307 4852
rect 13341 4818 13380 4852
rect 13414 4818 13453 4852
rect 13487 4818 13526 4852
rect 13560 4818 13599 4852
rect 13633 4818 13672 4852
rect 13706 4818 13745 4852
rect 13779 4818 13818 4852
rect 13852 4818 13891 4852
rect 13925 4818 13964 4852
rect 13998 4818 14037 4852
rect 14071 4818 14110 4852
rect 14144 4818 14183 4852
rect 14217 4818 14256 4852
rect 14290 4818 14329 4852
rect 14363 4818 14402 4852
rect 14436 4849 14591 4852
tri 14591 4849 14599 4857 sw
rect 14818 4849 14969 4857
rect 15003 4849 15117 4883
rect 14436 4820 14599 4849
tri 14599 4820 14628 4849 sw
rect 14436 4818 14628 4820
rect 575 4806 14628 4818
rect 575 4785 991 4806
tri 991 4785 1012 4806 nw
tri 14210 4786 14230 4806 ne
rect 14230 4786 14628 4806
tri 14230 4785 14231 4786 ne
rect 14231 4785 14628 4786
rect 575 4777 983 4785
tri 983 4777 991 4785 nw
tri 14231 4777 14239 4785 ne
rect 14239 4777 14628 4785
rect 575 4774 980 4777
tri 980 4774 983 4777 nw
tri 14239 4774 14242 4777 ne
rect 14242 4774 14628 4777
rect 575 4744 733 4774
rect 575 4710 587 4744
rect 621 4710 659 4744
rect 693 4740 733 4744
rect 767 4740 946 4774
tri 946 4740 980 4774 nw
tri 14242 4740 14276 4774 ne
rect 14276 4740 14431 4774
rect 14465 4743 14628 4774
rect 14465 4740 14510 4743
rect 693 4710 915 4740
rect 575 4709 915 4710
tri 915 4709 946 4740 nw
tri 14276 4709 14307 4740 ne
rect 14307 4709 14510 4740
rect 14544 4709 14582 4743
rect 14616 4709 14628 4743
rect 575 4705 911 4709
tri 911 4705 915 4709 nw
tri 14307 4705 14311 4709 ne
rect 14311 4705 14628 4709
rect 575 4701 907 4705
tri 907 4701 911 4705 nw
tri 14311 4701 14315 4705 ne
rect 14315 4701 14628 4705
rect 575 4670 733 4701
rect 575 4636 587 4670
rect 621 4636 659 4670
rect 693 4667 733 4670
rect 767 4667 873 4701
tri 873 4667 907 4701 nw
tri 14315 4667 14349 4701 ne
rect 14349 4667 14431 4701
rect 14465 4670 14628 4701
rect 14465 4667 14510 4670
rect 693 4636 842 4667
tri 842 4636 873 4667 nw
tri 14349 4636 14380 4667 ne
rect 14380 4636 14510 4667
rect 14544 4636 14582 4670
rect 14616 4636 14628 4670
rect 575 4633 839 4636
tri 839 4633 842 4636 nw
tri 14380 4633 14383 4636 ne
rect 14383 4633 14628 4636
rect 575 4628 834 4633
tri 834 4628 839 4633 nw
tri 14383 4628 14388 4633 ne
rect 14388 4628 14628 4633
rect 575 4596 733 4628
rect 575 4562 587 4596
rect 621 4562 659 4596
rect 693 4594 733 4596
rect 767 4594 803 4628
tri 803 4597 834 4628 nw
tri 14388 4616 14400 4628 ne
rect 693 4562 803 4594
rect 575 4555 803 4562
rect 575 4522 733 4555
rect 575 4488 587 4522
rect 621 4488 659 4522
rect 693 4521 733 4522
rect 767 4521 803 4555
rect 693 4488 803 4521
rect 14400 4594 14431 4628
rect 14465 4597 14628 4628
rect 14465 4594 14510 4597
rect 14400 4563 14510 4594
rect 14544 4563 14582 4597
rect 14616 4563 14628 4597
rect 14400 4555 14628 4563
rect 14400 4521 14431 4555
rect 14465 4524 14628 4555
rect 14465 4521 14510 4524
rect 575 4482 803 4488
rect 575 4449 733 4482
rect 575 4415 587 4449
rect 621 4415 659 4449
rect 693 4448 733 4449
rect 767 4448 803 4482
rect 693 4415 803 4448
rect 575 4409 803 4415
rect 575 4376 733 4409
rect 575 4342 587 4376
rect 621 4342 659 4376
rect 693 4375 733 4376
rect 767 4375 803 4409
rect 919 4494 1049 4506
rect 919 4388 931 4494
rect 1037 4388 1049 4494
rect 919 4376 1049 4388
rect 1349 4494 1479 4506
rect 1349 4388 1361 4494
rect 1467 4388 1479 4494
rect 1349 4376 1479 4388
rect 1911 4494 2041 4506
rect 1911 4388 1923 4494
rect 2029 4388 2041 4494
rect 1911 4376 2041 4388
rect 2341 4494 2471 4506
rect 2341 4388 2353 4494
rect 2459 4388 2471 4494
rect 2341 4376 2471 4388
rect 2903 4494 3033 4506
rect 2903 4388 2915 4494
rect 3021 4388 3033 4494
rect 2903 4376 3033 4388
rect 3333 4494 3463 4506
rect 3333 4388 3345 4494
rect 3451 4388 3463 4494
rect 3333 4376 3463 4388
rect 3895 4494 4025 4506
rect 3895 4388 3907 4494
rect 4013 4388 4025 4494
rect 3895 4376 4025 4388
rect 4325 4494 4455 4506
rect 4325 4388 4337 4494
rect 4443 4388 4455 4494
rect 4325 4376 4455 4388
rect 4887 4494 5017 4506
rect 4887 4388 4899 4494
rect 5005 4388 5017 4494
rect 4887 4376 5017 4388
rect 5317 4494 5447 4506
rect 5317 4388 5329 4494
rect 5435 4388 5447 4494
rect 5317 4376 5447 4388
rect 5879 4494 6009 4506
rect 5879 4388 5891 4494
rect 5997 4388 6009 4494
rect 5879 4376 6009 4388
rect 6309 4494 6439 4506
rect 6309 4388 6321 4494
rect 6427 4388 6439 4494
rect 6309 4376 6439 4388
rect 6856 4494 6986 4506
rect 6856 4388 6868 4494
rect 6974 4388 6986 4494
rect 6856 4376 6986 4388
rect 7301 4494 7431 4506
rect 7301 4388 7313 4494
rect 7419 4388 7431 4494
rect 7301 4376 7431 4388
rect 7863 4494 7993 4506
rect 7863 4388 7875 4494
rect 7981 4388 7993 4494
rect 7863 4376 7993 4388
rect 8293 4494 8423 4506
rect 8293 4388 8305 4494
rect 8411 4388 8423 4494
rect 8293 4376 8423 4388
rect 8855 4494 8985 4506
rect 8855 4388 8867 4494
rect 8973 4388 8985 4494
rect 8855 4376 8985 4388
rect 9285 4494 9415 4506
rect 9285 4388 9297 4494
rect 9403 4388 9415 4494
rect 9285 4376 9415 4388
rect 9847 4494 9977 4506
rect 9847 4388 9859 4494
rect 9965 4388 9977 4494
rect 9847 4376 9977 4388
rect 10277 4494 10407 4506
rect 10277 4388 10289 4494
rect 10395 4388 10407 4494
rect 10277 4376 10407 4388
rect 10839 4494 10969 4506
rect 10839 4388 10851 4494
rect 10957 4388 10969 4494
rect 10839 4376 10969 4388
rect 11269 4494 11399 4506
rect 11269 4388 11281 4494
rect 11387 4388 11399 4494
rect 11269 4376 11399 4388
rect 11831 4494 11961 4506
rect 11831 4388 11843 4494
rect 11949 4388 11961 4494
rect 11831 4376 11961 4388
rect 12261 4494 12391 4506
rect 12261 4388 12273 4494
rect 12379 4388 12391 4494
rect 12261 4376 12391 4388
rect 12823 4494 12953 4506
rect 12823 4388 12835 4494
rect 12941 4388 12953 4494
rect 12823 4376 12953 4388
rect 13253 4494 13383 4506
rect 13253 4388 13265 4494
rect 13371 4388 13383 4494
rect 13253 4376 13383 4388
rect 13815 4494 13945 4506
rect 13815 4388 13827 4494
rect 13933 4388 13945 4494
rect 13815 4376 13945 4388
rect 14173 4494 14303 4506
rect 14173 4388 14185 4494
rect 14291 4388 14303 4494
rect 14173 4376 14303 4388
rect 14400 4490 14510 4521
rect 14544 4490 14582 4524
rect 14616 4490 14628 4524
rect 14400 4482 14628 4490
rect 14400 4448 14431 4482
rect 14465 4451 14628 4482
rect 14465 4448 14510 4451
rect 14400 4417 14510 4448
rect 14544 4417 14582 4451
rect 14616 4417 14628 4451
rect 14400 4409 14628 4417
rect 693 4342 803 4375
rect 575 4336 803 4342
rect 575 4303 733 4336
rect 575 4269 587 4303
rect 621 4269 659 4303
rect 693 4302 733 4303
rect 767 4302 803 4336
rect 693 4269 803 4302
rect 575 4263 803 4269
rect 575 4230 733 4263
rect 575 4196 587 4230
rect 621 4196 659 4230
rect 693 4229 733 4230
rect 767 4229 803 4263
rect 693 4196 803 4229
rect 575 4190 803 4196
rect 575 4157 733 4190
rect 575 4123 587 4157
rect 621 4123 659 4157
rect 693 4156 733 4157
rect 767 4156 803 4190
rect 693 4123 803 4156
rect 575 4117 803 4123
rect 575 4084 733 4117
rect 575 4068 587 4084
rect 621 4068 659 4084
rect 693 4083 733 4084
rect 767 4083 803 4117
rect 693 4068 803 4083
rect 14400 4375 14431 4409
rect 14465 4378 14628 4409
rect 14465 4375 14510 4378
rect 14400 4344 14510 4375
rect 14544 4344 14582 4378
rect 14616 4344 14628 4378
rect 14400 4336 14628 4344
rect 14400 4302 14431 4336
rect 14465 4305 14628 4336
rect 14465 4302 14510 4305
rect 14400 4271 14510 4302
rect 14544 4271 14582 4305
rect 14616 4271 14628 4305
rect 14400 4263 14628 4271
rect 14400 4229 14431 4263
rect 14465 4232 14628 4263
rect 14465 4229 14510 4232
rect 14400 4198 14510 4229
rect 14544 4198 14582 4232
rect 14616 4198 14628 4232
rect 14400 4190 14628 4198
rect 14400 4156 14431 4190
rect 14465 4159 14628 4190
rect 14465 4156 14510 4159
rect 14400 4125 14510 4156
rect 14544 4125 14582 4159
rect 14616 4125 14628 4159
rect 14400 4117 14628 4125
rect 14400 4083 14431 4117
rect 14465 4086 14628 4117
rect 14465 4083 14510 4086
rect 627 4050 659 4068
rect 627 4016 663 4050
rect 715 4044 751 4068
rect 715 4016 733 4044
rect 575 4011 733 4016
rect 575 4003 587 4011
rect 621 4003 659 4011
rect 693 4010 733 4011
rect 767 4010 803 4016
rect 693 4003 803 4010
rect 627 3977 659 4003
rect 627 3951 663 3977
rect 715 3971 751 4003
rect 715 3951 733 3971
rect 575 3938 733 3951
rect 767 3938 803 3951
rect 627 3904 659 3938
rect 715 3937 733 3938
rect 627 3886 663 3904
rect 715 3898 751 3937
rect 715 3886 733 3898
rect 575 3873 733 3886
rect 767 3873 803 3886
rect 627 3865 663 3873
rect 627 3831 659 3865
rect 715 3864 733 3873
rect 627 3821 663 3831
rect 715 3825 751 3864
rect 715 3821 733 3825
rect 575 3808 733 3821
rect 767 3808 803 3821
rect 627 3792 663 3808
rect 627 3758 659 3792
rect 715 3791 733 3808
rect 627 3756 663 3758
rect 715 3756 751 3791
rect 575 3752 803 3756
rect 575 3743 733 3752
rect 767 3743 803 3752
rect 627 3719 663 3743
rect 627 3691 659 3719
rect 715 3718 733 3743
rect 715 3691 751 3718
rect 575 3685 587 3691
rect 621 3685 659 3691
rect 693 3685 803 3691
rect 575 3679 803 3685
rect 575 3678 733 3679
rect 767 3678 803 3679
rect 627 3646 663 3678
rect 627 3626 659 3646
rect 715 3645 733 3678
rect 715 3626 751 3645
rect 575 3613 587 3626
rect 621 3613 659 3626
rect 693 3613 803 3626
rect 627 3612 659 3613
rect 627 3573 663 3612
rect 715 3606 751 3613
rect 627 3561 659 3573
rect 715 3572 733 3606
rect 715 3561 751 3572
rect 575 3548 587 3561
rect 621 3548 659 3561
rect 693 3548 803 3561
rect 627 3539 659 3548
rect 627 3500 663 3539
rect 715 3533 751 3548
rect 627 3496 659 3500
rect 715 3499 733 3533
rect 715 3496 751 3499
rect 575 3483 587 3496
rect 621 3483 659 3496
rect 693 3483 803 3496
rect 627 3466 659 3483
rect 627 3431 663 3466
rect 715 3460 751 3483
rect 715 3431 733 3460
rect 575 3427 733 3431
rect 575 3418 587 3427
rect 621 3418 659 3427
rect 693 3426 733 3427
rect 767 3426 803 3431
rect 693 3418 803 3426
rect 627 3393 659 3418
rect 627 3366 663 3393
rect 715 3387 751 3418
rect 715 3366 733 3387
rect 575 3354 733 3366
rect 575 3353 587 3354
rect 621 3353 659 3354
rect 693 3353 733 3354
rect 767 3353 803 3366
rect 627 3320 659 3353
rect 627 3301 663 3320
rect 715 3314 751 3353
rect 715 3301 733 3314
rect 575 3288 733 3301
rect 767 3288 803 3301
rect 627 3281 663 3288
rect 627 3247 659 3281
rect 715 3280 733 3288
rect 627 3236 663 3247
rect 715 3241 751 3280
rect 715 3236 733 3241
rect 575 3223 733 3236
rect 767 3223 803 3236
rect 627 3208 663 3223
rect 627 3174 659 3208
rect 715 3207 733 3223
rect 627 3171 663 3174
rect 715 3171 751 3207
rect 575 3168 803 3171
rect 575 3158 733 3168
rect 767 3158 803 3168
rect 627 3135 663 3158
rect 627 3106 659 3135
rect 715 3134 733 3158
rect 715 3106 751 3134
rect 575 3101 587 3106
rect 621 3101 659 3106
rect 693 3101 803 3106
rect 575 3095 803 3101
rect 575 3093 733 3095
rect 767 3093 803 3095
rect 627 3062 663 3093
rect 627 3041 659 3062
rect 715 3061 733 3093
rect 715 3041 751 3061
rect 575 3028 587 3041
rect 621 3028 659 3041
rect 693 3028 803 3041
rect 627 2989 663 3028
rect 715 3022 751 3028
rect 627 2976 659 2989
rect 715 2988 733 3022
rect 715 2976 751 2988
rect 575 2963 587 2976
rect 621 2963 659 2976
rect 693 2963 803 2976
rect 627 2955 659 2963
rect 627 2916 663 2955
rect 715 2949 751 2963
rect 627 2911 659 2916
rect 715 2915 733 2949
rect 715 2911 751 2915
rect 575 2898 587 2911
rect 621 2898 659 2911
rect 693 2898 803 2911
rect 627 2882 659 2898
rect 627 2846 663 2882
rect 715 2876 751 2898
rect 715 2846 733 2876
rect 575 2843 733 2846
rect 575 2833 587 2843
rect 621 2833 659 2843
rect 693 2842 733 2843
rect 767 2842 803 2846
rect 693 2833 803 2842
rect 627 2809 659 2833
rect 627 2781 663 2809
rect 715 2803 751 2833
rect 715 2781 733 2803
rect 575 2770 733 2781
rect 575 2768 587 2770
rect 621 2768 659 2770
rect 693 2769 733 2770
rect 767 2769 803 2781
rect 693 2768 803 2769
rect 627 2736 659 2768
rect 627 2716 663 2736
rect 715 2730 751 2768
rect 715 2716 733 2730
rect 575 2703 733 2716
rect 767 2703 803 2716
rect 627 2697 663 2703
rect 627 2663 659 2697
rect 715 2696 733 2703
rect 627 2651 663 2663
rect 715 2657 751 2696
rect 715 2651 733 2657
rect 575 2638 733 2651
rect 767 2638 803 2651
rect 627 2624 663 2638
rect 627 2590 659 2624
rect 715 2623 733 2638
rect 627 2586 663 2590
rect 715 2586 751 2623
rect 575 2584 803 2586
rect 575 2573 733 2584
rect 767 2573 803 2584
rect 627 2551 663 2573
rect 627 2521 659 2551
rect 715 2550 733 2573
rect 715 2521 751 2550
rect 575 2517 587 2521
rect 621 2517 659 2521
rect 693 2517 803 2521
rect 575 2511 803 2517
rect 575 2508 733 2511
rect 767 2508 803 2511
rect 627 2478 663 2508
rect 627 2456 659 2478
rect 715 2477 733 2508
rect 715 2456 751 2477
rect 575 2444 587 2456
rect 621 2444 659 2456
rect 693 2444 803 2456
rect 575 2443 803 2444
rect 627 2405 663 2443
rect 715 2438 751 2443
rect 627 2391 659 2405
rect 715 2404 733 2438
rect 715 2391 751 2404
rect 575 2378 587 2391
rect 621 2378 659 2391
rect 693 2378 803 2391
rect 627 2371 659 2378
rect 627 2332 663 2371
rect 715 2365 751 2378
rect 627 2326 659 2332
rect 715 2331 733 2365
rect 715 2326 751 2331
rect 575 2313 587 2326
rect 621 2313 659 2326
rect 693 2313 803 2326
rect 627 2298 659 2313
rect 627 2261 663 2298
rect 715 2292 751 2313
rect 715 2261 733 2292
rect 575 2259 733 2261
rect 575 2248 587 2259
rect 621 2248 659 2259
rect 693 2258 733 2259
rect 767 2258 803 2261
rect 693 2248 803 2258
rect 627 2225 659 2248
rect 627 2196 663 2225
rect 715 2219 751 2248
rect 715 2196 733 2219
rect 575 2186 733 2196
rect 575 2183 587 2186
rect 621 2183 659 2186
rect 693 2185 733 2186
rect 767 2185 803 2196
rect 693 2183 803 2185
rect 627 2152 659 2183
rect 627 2131 663 2152
rect 715 2146 751 2183
rect 715 2131 733 2146
rect 575 2118 733 2131
rect 767 2118 803 2131
rect 627 2113 663 2118
rect 627 2079 659 2113
rect 715 2112 733 2118
rect 627 2066 663 2079
rect 715 2073 751 2112
rect 715 2066 733 2073
rect 575 2053 733 2066
rect 767 2053 803 2066
rect 627 2040 663 2053
rect 627 2006 659 2040
rect 715 2039 733 2053
rect 627 2001 663 2006
rect 715 2001 751 2039
rect 575 2000 803 2001
rect 575 1987 733 2000
rect 767 1987 803 2000
rect 627 1967 663 1987
rect 627 1935 659 1967
rect 715 1966 733 1987
rect 715 1935 751 1966
rect 575 1933 587 1935
rect 621 1933 659 1935
rect 693 1933 803 1935
rect 575 1927 803 1933
rect 575 1921 733 1927
rect 767 1921 803 1927
rect 627 1894 663 1921
rect 627 1869 659 1894
rect 715 1893 733 1921
rect 715 1869 751 1893
rect 575 1860 587 1869
rect 621 1860 659 1869
rect 693 1860 803 1869
rect 575 1855 803 1860
rect 627 1821 663 1855
rect 715 1854 751 1855
rect 627 1803 659 1821
rect 715 1820 733 1854
rect 715 1803 751 1820
rect 575 1789 587 1803
rect 621 1789 659 1803
rect 693 1789 803 1803
rect 627 1787 659 1789
rect 627 1748 663 1787
rect 715 1781 751 1789
rect 627 1737 659 1748
rect 715 1747 733 1781
rect 715 1737 751 1747
rect 575 1723 587 1737
rect 621 1723 659 1737
rect 693 1723 803 1737
rect 627 1714 659 1723
rect 627 1675 663 1714
rect 715 1708 751 1723
rect 627 1671 659 1675
rect 715 1674 733 1708
rect 715 1671 751 1674
rect 575 1657 587 1671
rect 621 1657 659 1671
rect 693 1657 803 1671
rect 627 1641 659 1657
rect 627 1605 663 1641
rect 715 1635 751 1657
rect 715 1605 733 1635
rect 575 1602 733 1605
rect 575 1591 587 1602
rect 621 1591 659 1602
rect 693 1601 733 1602
rect 767 1601 803 1605
rect 693 1591 803 1601
rect 627 1568 659 1591
rect 627 1539 663 1568
rect 715 1562 751 1591
rect 715 1539 733 1562
rect 575 1529 733 1539
rect 575 1525 587 1529
rect 621 1525 659 1529
rect 693 1528 733 1529
rect 767 1528 803 1539
rect 693 1525 803 1528
rect 627 1495 659 1525
rect 627 1473 663 1495
rect 715 1489 751 1525
rect 715 1473 733 1489
rect 575 1455 733 1473
rect 767 1455 803 1473
rect 1103 4068 1295 4074
rect 1103 4016 1109 4068
rect 1161 4016 1173 4068
rect 1225 4016 1237 4068
rect 1289 4016 1295 4068
rect 1103 4003 1295 4016
rect 1103 3951 1109 4003
rect 1161 3951 1173 4003
rect 1225 3951 1237 4003
rect 1289 3951 1295 4003
rect 1103 3938 1295 3951
rect 1103 3886 1109 3938
rect 1161 3886 1173 3938
rect 1225 3886 1237 3938
rect 1289 3886 1295 3938
rect 1103 3880 1110 3886
rect 1144 3880 1182 3886
rect 1216 3880 1254 3886
rect 1288 3880 1295 3886
rect 1103 3873 1295 3880
rect 1103 3821 1109 3873
rect 1161 3821 1173 3873
rect 1225 3821 1237 3873
rect 1289 3821 1295 3873
rect 1103 3808 1110 3821
rect 1144 3808 1182 3821
rect 1216 3808 1254 3821
rect 1288 3808 1295 3821
rect 1103 3756 1109 3808
rect 1161 3756 1173 3808
rect 1225 3756 1237 3808
rect 1289 3756 1295 3808
rect 1103 3743 1110 3756
rect 1144 3743 1182 3756
rect 1216 3743 1254 3756
rect 1288 3743 1295 3756
rect 1103 3691 1109 3743
rect 1161 3691 1173 3743
rect 1225 3691 1237 3743
rect 1289 3691 1295 3743
rect 1103 3678 1110 3691
rect 1144 3678 1182 3691
rect 1216 3678 1254 3691
rect 1288 3678 1295 3691
rect 1103 3626 1109 3678
rect 1161 3626 1173 3678
rect 1225 3626 1237 3678
rect 1289 3626 1295 3678
rect 1103 3618 1295 3626
rect 1103 3613 1110 3618
rect 1144 3613 1182 3618
rect 1216 3613 1254 3618
rect 1288 3613 1295 3618
rect 1103 3561 1109 3613
rect 1161 3561 1173 3613
rect 1225 3561 1237 3613
rect 1289 3561 1295 3613
rect 1103 3548 1295 3561
rect 1103 3496 1109 3548
rect 1161 3496 1173 3548
rect 1225 3496 1237 3548
rect 1289 3496 1295 3548
rect 1103 3483 1295 3496
rect 1103 3431 1109 3483
rect 1161 3431 1173 3483
rect 1225 3431 1237 3483
rect 1289 3431 1295 3483
rect 1103 3418 1295 3431
rect 1103 3366 1109 3418
rect 1161 3366 1173 3418
rect 1225 3366 1237 3418
rect 1289 3366 1295 3418
rect 1103 3362 1110 3366
rect 1144 3362 1182 3366
rect 1216 3362 1254 3366
rect 1288 3362 1295 3366
rect 1103 3353 1295 3362
rect 1103 3301 1109 3353
rect 1161 3301 1173 3353
rect 1225 3301 1237 3353
rect 1289 3301 1295 3353
rect 1103 3288 1110 3301
rect 1144 3288 1182 3301
rect 1216 3288 1254 3301
rect 1288 3288 1295 3301
rect 1103 3236 1109 3288
rect 1161 3236 1173 3288
rect 1225 3236 1237 3288
rect 1289 3236 1295 3288
rect 1103 3223 1110 3236
rect 1144 3223 1182 3236
rect 1216 3223 1254 3236
rect 1288 3223 1295 3236
rect 1103 3171 1109 3223
rect 1161 3171 1173 3223
rect 1225 3171 1237 3223
rect 1289 3171 1295 3223
rect 1103 3158 1110 3171
rect 1144 3158 1182 3171
rect 1216 3158 1254 3171
rect 1288 3158 1295 3171
rect 1103 3106 1109 3158
rect 1161 3106 1173 3158
rect 1225 3106 1237 3158
rect 1289 3106 1295 3158
rect 1103 3100 1295 3106
rect 1103 3093 1110 3100
rect 1144 3093 1182 3100
rect 1216 3093 1254 3100
rect 1288 3093 1295 3100
rect 1103 3041 1109 3093
rect 1161 3041 1173 3093
rect 1225 3041 1237 3093
rect 1289 3041 1295 3093
rect 1103 3028 1295 3041
rect 1103 2976 1109 3028
rect 1161 2976 1173 3028
rect 1225 2976 1237 3028
rect 1289 2976 1295 3028
rect 1103 2963 1295 2976
rect 1103 2911 1109 2963
rect 1161 2911 1173 2963
rect 1225 2911 1237 2963
rect 1289 2911 1295 2963
rect 1103 2898 1295 2911
rect 1103 2846 1109 2898
rect 1161 2846 1173 2898
rect 1225 2846 1237 2898
rect 1289 2846 1295 2898
rect 1103 2844 1110 2846
rect 1144 2844 1182 2846
rect 1216 2844 1254 2846
rect 1288 2844 1295 2846
rect 1103 2833 1295 2844
rect 1103 2781 1109 2833
rect 1161 2781 1173 2833
rect 1225 2781 1237 2833
rect 1289 2781 1295 2833
rect 1103 2770 1110 2781
rect 1144 2770 1182 2781
rect 1216 2770 1254 2781
rect 1288 2770 1295 2781
rect 1103 2768 1295 2770
rect 1103 2716 1109 2768
rect 1161 2716 1173 2768
rect 1225 2716 1237 2768
rect 1289 2716 1295 2768
rect 1103 2703 1110 2716
rect 1144 2703 1182 2716
rect 1216 2703 1254 2716
rect 1288 2703 1295 2716
rect 1103 2651 1109 2703
rect 1161 2651 1173 2703
rect 1225 2651 1237 2703
rect 1289 2651 1295 2703
rect 1103 2638 1110 2651
rect 1144 2638 1182 2651
rect 1216 2638 1254 2651
rect 1288 2638 1295 2651
rect 1103 2586 1109 2638
rect 1161 2586 1173 2638
rect 1225 2586 1237 2638
rect 1289 2586 1295 2638
rect 1103 2582 1295 2586
rect 1103 2573 1110 2582
rect 1144 2573 1182 2582
rect 1216 2573 1254 2582
rect 1288 2573 1295 2582
rect 1103 2521 1109 2573
rect 1161 2521 1173 2573
rect 1225 2521 1237 2573
rect 1289 2521 1295 2573
rect 1103 2508 1295 2521
rect 1103 2456 1109 2508
rect 1161 2456 1173 2508
rect 1225 2456 1237 2508
rect 1289 2456 1295 2508
rect 1103 2443 1295 2456
rect 1103 2391 1109 2443
rect 1161 2391 1173 2443
rect 1225 2391 1237 2443
rect 1289 2391 1295 2443
rect 1103 2378 1295 2391
rect 1103 2326 1109 2378
rect 1161 2326 1173 2378
rect 1225 2326 1237 2378
rect 1289 2326 1295 2378
rect 1103 2313 1295 2326
rect 1103 2261 1109 2313
rect 1161 2261 1173 2313
rect 1225 2261 1237 2313
rect 1289 2261 1295 2313
rect 1103 2252 1110 2261
rect 1144 2252 1182 2261
rect 1216 2252 1254 2261
rect 1288 2252 1295 2261
rect 1103 2248 1295 2252
rect 1103 2196 1109 2248
rect 1161 2196 1173 2248
rect 1225 2196 1237 2248
rect 1289 2196 1295 2248
rect 1103 2183 1110 2196
rect 1144 2183 1182 2196
rect 1216 2183 1254 2196
rect 1288 2183 1295 2196
rect 1103 2131 1109 2183
rect 1161 2131 1173 2183
rect 1225 2131 1237 2183
rect 1289 2131 1295 2183
rect 1103 2118 1110 2131
rect 1144 2118 1182 2131
rect 1216 2118 1254 2131
rect 1288 2118 1295 2131
rect 1103 2066 1109 2118
rect 1161 2066 1173 2118
rect 1225 2066 1237 2118
rect 1289 2066 1295 2118
rect 1103 2064 1295 2066
rect 1103 2053 1110 2064
rect 1144 2053 1182 2064
rect 1216 2053 1254 2064
rect 1288 2053 1295 2064
rect 1103 2001 1109 2053
rect 1161 2001 1173 2053
rect 1225 2001 1237 2053
rect 1289 2001 1295 2053
rect 1103 1990 1295 2001
rect 1103 1987 1110 1990
rect 1144 1987 1182 1990
rect 1216 1987 1254 1990
rect 1288 1987 1295 1990
rect 1103 1935 1109 1987
rect 1161 1935 1173 1987
rect 1225 1935 1237 1987
rect 1289 1935 1295 1987
rect 1103 1921 1295 1935
rect 1103 1869 1109 1921
rect 1161 1869 1173 1921
rect 1225 1869 1237 1921
rect 1289 1869 1295 1921
rect 1103 1855 1295 1869
rect 1103 1803 1109 1855
rect 1161 1803 1173 1855
rect 1225 1803 1237 1855
rect 1289 1803 1295 1855
rect 1103 1789 1295 1803
rect 1103 1737 1109 1789
rect 1161 1737 1173 1789
rect 1225 1737 1237 1789
rect 1289 1737 1295 1789
rect 1103 1734 1110 1737
rect 1144 1734 1182 1737
rect 1216 1734 1254 1737
rect 1288 1734 1295 1737
rect 1103 1723 1295 1734
rect 1103 1671 1109 1723
rect 1161 1671 1173 1723
rect 1225 1671 1237 1723
rect 1289 1671 1295 1723
rect 1103 1660 1110 1671
rect 1144 1660 1182 1671
rect 1216 1660 1254 1671
rect 1288 1660 1295 1671
rect 1103 1657 1295 1660
rect 1103 1605 1109 1657
rect 1161 1605 1173 1657
rect 1225 1605 1237 1657
rect 1289 1605 1295 1657
rect 1103 1591 1110 1605
rect 1144 1591 1182 1605
rect 1216 1591 1254 1605
rect 1288 1591 1295 1605
rect 1103 1539 1109 1591
rect 1161 1539 1173 1591
rect 1225 1539 1237 1591
rect 1289 1539 1295 1591
rect 1103 1525 1110 1539
rect 1144 1525 1182 1539
rect 1216 1525 1254 1539
rect 1288 1525 1295 1539
rect 1103 1473 1109 1525
rect 1161 1473 1173 1525
rect 1225 1473 1237 1525
rect 1289 1473 1295 1525
rect 1103 1467 1295 1473
rect 1599 4068 1791 4074
rect 1599 4016 1605 4068
rect 1657 4050 1669 4068
rect 1721 4050 1733 4068
rect 1785 4016 1791 4068
rect 1599 4003 1606 4016
rect 1784 4003 1791 4016
rect 1599 3951 1605 4003
rect 1785 3951 1791 4003
rect 1599 3938 1606 3951
rect 1784 3938 1791 3951
rect 1599 3886 1605 3938
rect 1785 3886 1791 3938
rect 1599 3873 1606 3886
rect 1784 3873 1791 3886
rect 1599 3821 1605 3873
rect 1785 3821 1791 3873
rect 1599 3808 1606 3821
rect 1784 3808 1791 3821
rect 1599 3756 1605 3808
rect 1785 3756 1791 3808
rect 1599 3743 1606 3756
rect 1784 3743 1791 3756
rect 1599 3691 1605 3743
rect 1785 3691 1791 3743
rect 1599 3678 1606 3691
rect 1784 3678 1791 3691
rect 1599 3626 1605 3678
rect 1785 3626 1791 3678
rect 1599 3613 1606 3626
rect 1784 3613 1791 3626
rect 1599 3561 1605 3613
rect 1785 3561 1791 3613
rect 1599 3548 1606 3561
rect 1784 3548 1791 3561
rect 1599 3496 1605 3548
rect 1785 3496 1791 3548
rect 1599 3483 1606 3496
rect 1784 3483 1791 3496
rect 1599 3431 1605 3483
rect 1785 3431 1791 3483
rect 1599 3418 1606 3431
rect 1784 3418 1791 3431
rect 1599 3366 1605 3418
rect 1785 3366 1791 3418
rect 1599 3353 1606 3366
rect 1784 3353 1791 3366
rect 1599 3301 1605 3353
rect 1785 3301 1791 3353
rect 1599 3288 1606 3301
rect 1784 3288 1791 3301
rect 1599 3236 1605 3288
rect 1785 3236 1791 3288
rect 1599 3223 1606 3236
rect 1784 3223 1791 3236
rect 1599 3171 1605 3223
rect 1785 3171 1791 3223
rect 1599 3158 1606 3171
rect 1784 3158 1791 3171
rect 1599 3106 1605 3158
rect 1785 3106 1791 3158
rect 1599 3093 1606 3106
rect 1784 3093 1791 3106
rect 1599 3041 1605 3093
rect 1657 3041 1669 3092
rect 1721 3041 1733 3092
rect 1785 3041 1791 3093
rect 1599 3040 1791 3041
rect 1599 3028 1606 3040
rect 1784 3028 1791 3040
rect 1599 2976 1605 3028
rect 1785 2976 1791 3028
rect 1599 2963 1606 2976
rect 1784 2963 1791 2976
rect 1599 2911 1605 2963
rect 1785 2911 1791 2963
rect 1599 2898 1606 2911
rect 1784 2898 1791 2911
rect 1599 2846 1605 2898
rect 1785 2846 1791 2898
rect 1599 2833 1606 2846
rect 1784 2833 1791 2846
rect 1599 2781 1605 2833
rect 1785 2781 1791 2833
rect 1599 2768 1606 2781
rect 1784 2768 1791 2781
rect 1599 2716 1605 2768
rect 1785 2716 1791 2768
rect 1599 2703 1606 2716
rect 1784 2703 1791 2716
rect 1599 2651 1605 2703
rect 1785 2651 1791 2703
rect 1599 2638 1606 2651
rect 1784 2638 1791 2651
rect 1599 2586 1605 2638
rect 1785 2586 1791 2638
rect 1599 2574 1606 2586
rect 1784 2574 1791 2586
rect 1599 2573 1791 2574
rect 1599 2521 1605 2573
rect 1657 2521 1669 2573
rect 1721 2521 1733 2573
rect 1785 2521 1791 2573
rect 1599 2508 1606 2521
rect 1640 2508 1678 2521
rect 1712 2508 1750 2521
rect 1784 2508 1791 2521
rect 1599 2456 1605 2508
rect 1657 2456 1669 2508
rect 1721 2456 1733 2508
rect 1785 2456 1791 2508
rect 1599 2449 1678 2456
rect 1712 2449 1791 2456
rect 1599 2443 1606 2449
rect 1784 2443 1791 2449
rect 1599 2391 1605 2443
rect 1785 2391 1791 2443
rect 1599 2378 1606 2391
rect 1784 2378 1791 2391
rect 1599 2326 1605 2378
rect 1785 2326 1791 2378
rect 1599 2313 1606 2326
rect 1784 2313 1791 2326
rect 1599 2261 1605 2313
rect 1785 2261 1791 2313
rect 1599 2248 1606 2261
rect 1784 2248 1791 2261
rect 1599 2196 1605 2248
rect 1785 2196 1791 2248
rect 1599 2183 1606 2196
rect 1784 2183 1791 2196
rect 1599 2131 1605 2183
rect 1785 2131 1791 2183
rect 1599 2118 1606 2131
rect 1784 2118 1791 2131
rect 1599 2066 1605 2118
rect 1785 2066 1791 2118
rect 1599 2053 1606 2066
rect 1784 2053 1791 2066
rect 1599 2001 1605 2053
rect 1785 2001 1791 2053
rect 1599 1987 1606 2001
rect 1784 1987 1791 2001
rect 1599 1935 1605 1987
rect 1785 1935 1791 1987
rect 1599 1921 1606 1935
rect 1784 1921 1791 1935
rect 1599 1869 1605 1921
rect 1785 1869 1791 1921
rect 1599 1855 1606 1869
rect 1784 1855 1791 1869
rect 1599 1803 1605 1855
rect 1785 1803 1791 1855
rect 1599 1789 1606 1803
rect 1784 1789 1791 1803
rect 1599 1737 1605 1789
rect 1785 1737 1791 1789
rect 1599 1723 1606 1737
rect 1784 1723 1791 1737
rect 1599 1671 1605 1723
rect 1785 1671 1791 1723
rect 1599 1657 1606 1671
rect 1784 1657 1791 1671
rect 1599 1605 1605 1657
rect 1785 1605 1791 1657
rect 1599 1591 1606 1605
rect 1784 1591 1791 1605
rect 1599 1539 1605 1591
rect 1785 1539 1791 1591
rect 1599 1525 1606 1539
rect 1784 1525 1791 1539
rect 1599 1473 1605 1525
rect 1657 1473 1669 1491
rect 1721 1473 1733 1491
rect 1785 1473 1791 1525
rect 1599 1467 1791 1473
rect 2095 4068 2287 4074
rect 2095 4016 2101 4068
rect 2153 4016 2165 4068
rect 2217 4016 2229 4068
rect 2281 4016 2287 4068
rect 2095 4003 2287 4016
rect 2095 3951 2101 4003
rect 2153 3951 2165 4003
rect 2217 3951 2229 4003
rect 2281 3951 2287 4003
rect 2095 3938 2287 3951
rect 2095 3886 2101 3938
rect 2153 3886 2165 3938
rect 2217 3886 2229 3938
rect 2281 3886 2287 3938
rect 2095 3880 2102 3886
rect 2136 3880 2174 3886
rect 2208 3880 2246 3886
rect 2280 3880 2287 3886
rect 2095 3873 2287 3880
rect 2095 3821 2101 3873
rect 2153 3821 2165 3873
rect 2217 3821 2229 3873
rect 2281 3821 2287 3873
rect 2095 3808 2102 3821
rect 2136 3808 2174 3821
rect 2208 3808 2246 3821
rect 2280 3808 2287 3821
rect 2095 3756 2101 3808
rect 2153 3756 2165 3808
rect 2217 3756 2229 3808
rect 2281 3756 2287 3808
rect 2095 3743 2102 3756
rect 2136 3743 2174 3756
rect 2208 3743 2246 3756
rect 2280 3743 2287 3756
rect 2095 3691 2101 3743
rect 2153 3691 2165 3743
rect 2217 3691 2229 3743
rect 2281 3691 2287 3743
rect 2095 3678 2102 3691
rect 2136 3678 2174 3691
rect 2208 3678 2246 3691
rect 2280 3678 2287 3691
rect 2095 3626 2101 3678
rect 2153 3626 2165 3678
rect 2217 3626 2229 3678
rect 2281 3626 2287 3678
rect 2095 3618 2287 3626
rect 2095 3613 2102 3618
rect 2136 3613 2174 3618
rect 2208 3613 2246 3618
rect 2280 3613 2287 3618
rect 2095 3561 2101 3613
rect 2153 3561 2165 3613
rect 2217 3561 2229 3613
rect 2281 3561 2287 3613
rect 2095 3548 2287 3561
rect 2095 3496 2101 3548
rect 2153 3496 2165 3548
rect 2217 3496 2229 3548
rect 2281 3496 2287 3548
rect 2095 3483 2287 3496
rect 2095 3431 2101 3483
rect 2153 3431 2165 3483
rect 2217 3431 2229 3483
rect 2281 3431 2287 3483
rect 2095 3418 2287 3431
rect 2095 3366 2101 3418
rect 2153 3366 2165 3418
rect 2217 3366 2229 3418
rect 2281 3366 2287 3418
rect 2095 3362 2102 3366
rect 2136 3362 2174 3366
rect 2208 3362 2246 3366
rect 2280 3362 2287 3366
rect 2095 3353 2287 3362
rect 2095 3301 2101 3353
rect 2153 3301 2165 3353
rect 2217 3301 2229 3353
rect 2281 3301 2287 3353
rect 2095 3288 2102 3301
rect 2136 3288 2174 3301
rect 2208 3288 2246 3301
rect 2280 3288 2287 3301
rect 2095 3236 2101 3288
rect 2153 3236 2165 3288
rect 2217 3236 2229 3288
rect 2281 3236 2287 3288
rect 2095 3223 2102 3236
rect 2136 3223 2174 3236
rect 2208 3223 2246 3236
rect 2280 3223 2287 3236
rect 2095 3171 2101 3223
rect 2153 3171 2165 3223
rect 2217 3171 2229 3223
rect 2281 3171 2287 3223
rect 2095 3158 2102 3171
rect 2136 3158 2174 3171
rect 2208 3158 2246 3171
rect 2280 3158 2287 3171
rect 2095 3106 2101 3158
rect 2153 3106 2165 3158
rect 2217 3106 2229 3158
rect 2281 3106 2287 3158
rect 2095 3100 2287 3106
rect 2095 3093 2102 3100
rect 2136 3093 2174 3100
rect 2208 3093 2246 3100
rect 2280 3093 2287 3100
rect 2095 3041 2101 3093
rect 2153 3041 2165 3093
rect 2217 3041 2229 3093
rect 2281 3041 2287 3093
rect 2095 3028 2287 3041
rect 2095 2976 2101 3028
rect 2153 2976 2165 3028
rect 2217 2976 2229 3028
rect 2281 2976 2287 3028
rect 2095 2963 2287 2976
rect 2095 2911 2101 2963
rect 2153 2911 2165 2963
rect 2217 2911 2229 2963
rect 2281 2911 2287 2963
rect 2095 2898 2287 2911
rect 2095 2846 2101 2898
rect 2153 2846 2165 2898
rect 2217 2846 2229 2898
rect 2281 2846 2287 2898
rect 2095 2844 2102 2846
rect 2136 2844 2174 2846
rect 2208 2844 2246 2846
rect 2280 2844 2287 2846
rect 2095 2833 2287 2844
rect 2095 2781 2101 2833
rect 2153 2781 2165 2833
rect 2217 2781 2229 2833
rect 2281 2781 2287 2833
rect 2095 2770 2102 2781
rect 2136 2770 2174 2781
rect 2208 2770 2246 2781
rect 2280 2770 2287 2781
rect 2095 2768 2287 2770
rect 2095 2716 2101 2768
rect 2153 2716 2165 2768
rect 2217 2716 2229 2768
rect 2281 2716 2287 2768
rect 2095 2703 2102 2716
rect 2136 2703 2174 2716
rect 2208 2703 2246 2716
rect 2280 2703 2287 2716
rect 2095 2651 2101 2703
rect 2153 2651 2165 2703
rect 2217 2651 2229 2703
rect 2281 2651 2287 2703
rect 2095 2638 2102 2651
rect 2136 2638 2174 2651
rect 2208 2638 2246 2651
rect 2280 2638 2287 2651
rect 2095 2586 2101 2638
rect 2153 2586 2165 2638
rect 2217 2586 2229 2638
rect 2281 2586 2287 2638
rect 2095 2582 2287 2586
rect 2095 2573 2102 2582
rect 2136 2573 2174 2582
rect 2208 2573 2246 2582
rect 2280 2573 2287 2582
rect 2095 2521 2101 2573
rect 2153 2521 2165 2573
rect 2217 2521 2229 2573
rect 2281 2521 2287 2573
rect 2095 2508 2287 2521
rect 2095 2456 2101 2508
rect 2153 2456 2165 2508
rect 2217 2456 2229 2508
rect 2281 2456 2287 2508
rect 2095 2443 2287 2456
rect 2095 2391 2101 2443
rect 2153 2391 2165 2443
rect 2217 2391 2229 2443
rect 2281 2391 2287 2443
rect 2095 2378 2287 2391
rect 2095 2326 2101 2378
rect 2153 2326 2165 2378
rect 2217 2326 2229 2378
rect 2281 2326 2287 2378
rect 2095 2313 2287 2326
rect 2095 2261 2101 2313
rect 2153 2261 2165 2313
rect 2217 2261 2229 2313
rect 2281 2261 2287 2313
rect 2095 2252 2102 2261
rect 2136 2252 2174 2261
rect 2208 2252 2246 2261
rect 2280 2252 2287 2261
rect 2095 2248 2287 2252
rect 2095 2196 2101 2248
rect 2153 2196 2165 2248
rect 2217 2196 2229 2248
rect 2281 2196 2287 2248
rect 2095 2183 2102 2196
rect 2136 2183 2174 2196
rect 2208 2183 2246 2196
rect 2280 2183 2287 2196
rect 2095 2131 2101 2183
rect 2153 2131 2165 2183
rect 2217 2131 2229 2183
rect 2281 2131 2287 2183
rect 2095 2118 2102 2131
rect 2136 2118 2174 2131
rect 2208 2118 2246 2131
rect 2280 2118 2287 2131
rect 2095 2066 2101 2118
rect 2153 2066 2165 2118
rect 2217 2066 2229 2118
rect 2281 2066 2287 2118
rect 2095 2064 2287 2066
rect 2095 2053 2102 2064
rect 2136 2053 2174 2064
rect 2208 2053 2246 2064
rect 2280 2053 2287 2064
rect 2095 2001 2101 2053
rect 2153 2001 2165 2053
rect 2217 2001 2229 2053
rect 2281 2001 2287 2053
rect 2095 1990 2287 2001
rect 2095 1987 2102 1990
rect 2136 1987 2174 1990
rect 2208 1987 2246 1990
rect 2280 1987 2287 1990
rect 2095 1935 2101 1987
rect 2153 1935 2165 1987
rect 2217 1935 2229 1987
rect 2281 1935 2287 1987
rect 2095 1921 2287 1935
rect 2095 1869 2101 1921
rect 2153 1869 2165 1921
rect 2217 1869 2229 1921
rect 2281 1869 2287 1921
rect 2095 1855 2287 1869
rect 2095 1803 2101 1855
rect 2153 1803 2165 1855
rect 2217 1803 2229 1855
rect 2281 1803 2287 1855
rect 2095 1789 2287 1803
rect 2095 1737 2101 1789
rect 2153 1737 2165 1789
rect 2217 1737 2229 1789
rect 2281 1737 2287 1789
rect 2095 1734 2102 1737
rect 2136 1734 2174 1737
rect 2208 1734 2246 1737
rect 2280 1734 2287 1737
rect 2095 1723 2287 1734
rect 2095 1671 2101 1723
rect 2153 1671 2165 1723
rect 2217 1671 2229 1723
rect 2281 1671 2287 1723
rect 2095 1660 2102 1671
rect 2136 1660 2174 1671
rect 2208 1660 2246 1671
rect 2280 1660 2287 1671
rect 2095 1657 2287 1660
rect 2095 1605 2101 1657
rect 2153 1605 2165 1657
rect 2217 1605 2229 1657
rect 2281 1605 2287 1657
rect 2095 1591 2102 1605
rect 2136 1591 2174 1605
rect 2208 1591 2246 1605
rect 2280 1591 2287 1605
rect 2095 1539 2101 1591
rect 2153 1539 2165 1591
rect 2217 1539 2229 1591
rect 2281 1539 2287 1591
rect 2095 1525 2102 1539
rect 2136 1525 2174 1539
rect 2208 1525 2246 1539
rect 2280 1525 2287 1539
rect 2095 1473 2101 1525
rect 2153 1473 2165 1525
rect 2217 1473 2229 1525
rect 2281 1473 2287 1525
rect 2095 1467 2287 1473
rect 2591 4068 2783 4074
rect 2591 4016 2597 4068
rect 2649 4050 2661 4068
rect 2713 4050 2725 4068
rect 2777 4016 2783 4068
rect 2591 4003 2598 4016
rect 2776 4003 2783 4016
rect 2591 3951 2597 4003
rect 2777 3951 2783 4003
rect 2591 3938 2598 3951
rect 2776 3938 2783 3951
rect 2591 3886 2597 3938
rect 2777 3886 2783 3938
rect 2591 3873 2598 3886
rect 2776 3873 2783 3886
rect 2591 3821 2597 3873
rect 2777 3821 2783 3873
rect 2591 3808 2598 3821
rect 2776 3808 2783 3821
rect 2591 3756 2597 3808
rect 2777 3756 2783 3808
rect 2591 3743 2598 3756
rect 2776 3743 2783 3756
rect 2591 3691 2597 3743
rect 2777 3691 2783 3743
rect 2591 3678 2598 3691
rect 2776 3678 2783 3691
rect 2591 3626 2597 3678
rect 2777 3626 2783 3678
rect 2591 3613 2598 3626
rect 2776 3613 2783 3626
rect 2591 3561 2597 3613
rect 2777 3561 2783 3613
rect 2591 3548 2598 3561
rect 2776 3548 2783 3561
rect 2591 3496 2597 3548
rect 2777 3496 2783 3548
rect 2591 3483 2598 3496
rect 2776 3483 2783 3496
rect 2591 3431 2597 3483
rect 2777 3431 2783 3483
rect 2591 3418 2598 3431
rect 2776 3418 2783 3431
rect 2591 3366 2597 3418
rect 2777 3366 2783 3418
rect 2591 3353 2598 3366
rect 2776 3353 2783 3366
rect 2591 3301 2597 3353
rect 2777 3301 2783 3353
rect 2591 3288 2598 3301
rect 2776 3288 2783 3301
rect 2591 3236 2597 3288
rect 2777 3236 2783 3288
rect 2591 3223 2598 3236
rect 2776 3223 2783 3236
rect 2591 3171 2597 3223
rect 2777 3171 2783 3223
rect 2591 3158 2598 3171
rect 2776 3158 2783 3171
rect 2591 3106 2597 3158
rect 2777 3106 2783 3158
rect 2591 3093 2598 3106
rect 2776 3093 2783 3106
rect 2591 3041 2597 3093
rect 2649 3041 2661 3092
rect 2713 3041 2725 3092
rect 2777 3041 2783 3093
rect 2591 3040 2783 3041
rect 2591 3028 2598 3040
rect 2776 3028 2783 3040
rect 2591 2976 2597 3028
rect 2777 2976 2783 3028
rect 2591 2963 2598 2976
rect 2776 2963 2783 2976
rect 2591 2911 2597 2963
rect 2777 2911 2783 2963
rect 2591 2898 2598 2911
rect 2776 2898 2783 2911
rect 2591 2846 2597 2898
rect 2777 2846 2783 2898
rect 2591 2833 2598 2846
rect 2776 2833 2783 2846
rect 2591 2781 2597 2833
rect 2777 2781 2783 2833
rect 2591 2768 2598 2781
rect 2776 2768 2783 2781
rect 2591 2716 2597 2768
rect 2777 2716 2783 2768
rect 2591 2703 2598 2716
rect 2776 2703 2783 2716
rect 2591 2651 2597 2703
rect 2777 2651 2783 2703
rect 2591 2638 2598 2651
rect 2776 2638 2783 2651
rect 2591 2586 2597 2638
rect 2777 2586 2783 2638
rect 2591 2574 2598 2586
rect 2776 2574 2783 2586
rect 2591 2573 2783 2574
rect 2591 2521 2597 2573
rect 2649 2521 2661 2573
rect 2713 2521 2725 2573
rect 2777 2521 2783 2573
rect 2591 2508 2598 2521
rect 2632 2508 2670 2521
rect 2704 2508 2742 2521
rect 2776 2508 2783 2521
rect 2591 2456 2597 2508
rect 2649 2456 2661 2508
rect 2713 2456 2725 2508
rect 2777 2456 2783 2508
rect 2591 2449 2670 2456
rect 2704 2449 2783 2456
rect 2591 2443 2598 2449
rect 2776 2443 2783 2449
rect 2591 2391 2597 2443
rect 2777 2391 2783 2443
rect 2591 2378 2598 2391
rect 2776 2378 2783 2391
rect 2591 2326 2597 2378
rect 2777 2326 2783 2378
rect 2591 2313 2598 2326
rect 2776 2313 2783 2326
rect 2591 2261 2597 2313
rect 2777 2261 2783 2313
rect 2591 2248 2598 2261
rect 2776 2248 2783 2261
rect 2591 2196 2597 2248
rect 2777 2196 2783 2248
rect 2591 2183 2598 2196
rect 2776 2183 2783 2196
rect 2591 2131 2597 2183
rect 2777 2131 2783 2183
rect 2591 2118 2598 2131
rect 2776 2118 2783 2131
rect 2591 2066 2597 2118
rect 2777 2066 2783 2118
rect 2591 2053 2598 2066
rect 2776 2053 2783 2066
rect 2591 2001 2597 2053
rect 2777 2001 2783 2053
rect 2591 1987 2598 2001
rect 2776 1987 2783 2001
rect 2591 1935 2597 1987
rect 2777 1935 2783 1987
rect 2591 1921 2598 1935
rect 2776 1921 2783 1935
rect 2591 1869 2597 1921
rect 2777 1869 2783 1921
rect 2591 1855 2598 1869
rect 2776 1855 2783 1869
rect 2591 1803 2597 1855
rect 2777 1803 2783 1855
rect 2591 1789 2598 1803
rect 2776 1789 2783 1803
rect 2591 1737 2597 1789
rect 2777 1737 2783 1789
rect 2591 1723 2598 1737
rect 2776 1723 2783 1737
rect 2591 1671 2597 1723
rect 2777 1671 2783 1723
rect 2591 1657 2598 1671
rect 2776 1657 2783 1671
rect 2591 1605 2597 1657
rect 2777 1605 2783 1657
rect 2591 1591 2598 1605
rect 2776 1591 2783 1605
rect 2591 1539 2597 1591
rect 2777 1539 2783 1591
rect 2591 1525 2598 1539
rect 2776 1525 2783 1539
rect 2591 1473 2597 1525
rect 2649 1473 2661 1491
rect 2713 1473 2725 1491
rect 2777 1473 2783 1525
rect 2591 1467 2783 1473
rect 3087 4068 3279 4074
rect 3087 4016 3093 4068
rect 3145 4016 3157 4068
rect 3209 4016 3221 4068
rect 3273 4016 3279 4068
rect 3087 4003 3279 4016
rect 3087 3951 3093 4003
rect 3145 3951 3157 4003
rect 3209 3951 3221 4003
rect 3273 3951 3279 4003
rect 3087 3938 3279 3951
rect 3087 3886 3093 3938
rect 3145 3886 3157 3938
rect 3209 3886 3221 3938
rect 3273 3886 3279 3938
rect 3087 3880 3094 3886
rect 3128 3880 3166 3886
rect 3200 3880 3238 3886
rect 3272 3880 3279 3886
rect 3087 3873 3279 3880
rect 3087 3821 3093 3873
rect 3145 3821 3157 3873
rect 3209 3821 3221 3873
rect 3273 3821 3279 3873
rect 3087 3808 3094 3821
rect 3128 3808 3166 3821
rect 3200 3808 3238 3821
rect 3272 3808 3279 3821
rect 3087 3756 3093 3808
rect 3145 3756 3157 3808
rect 3209 3756 3221 3808
rect 3273 3756 3279 3808
rect 3087 3743 3094 3756
rect 3128 3743 3166 3756
rect 3200 3743 3238 3756
rect 3272 3743 3279 3756
rect 3087 3691 3093 3743
rect 3145 3691 3157 3743
rect 3209 3691 3221 3743
rect 3273 3691 3279 3743
rect 3087 3678 3094 3691
rect 3128 3678 3166 3691
rect 3200 3678 3238 3691
rect 3272 3678 3279 3691
rect 3087 3626 3093 3678
rect 3145 3626 3157 3678
rect 3209 3626 3221 3678
rect 3273 3626 3279 3678
rect 3087 3618 3279 3626
rect 3087 3613 3094 3618
rect 3128 3613 3166 3618
rect 3200 3613 3238 3618
rect 3272 3613 3279 3618
rect 3087 3561 3093 3613
rect 3145 3561 3157 3613
rect 3209 3561 3221 3613
rect 3273 3561 3279 3613
rect 3087 3548 3279 3561
rect 3087 3496 3093 3548
rect 3145 3496 3157 3548
rect 3209 3496 3221 3548
rect 3273 3496 3279 3548
rect 3087 3483 3279 3496
rect 3087 3431 3093 3483
rect 3145 3431 3157 3483
rect 3209 3431 3221 3483
rect 3273 3431 3279 3483
rect 3087 3418 3279 3431
rect 3087 3366 3093 3418
rect 3145 3366 3157 3418
rect 3209 3366 3221 3418
rect 3273 3366 3279 3418
rect 3087 3362 3094 3366
rect 3128 3362 3166 3366
rect 3200 3362 3238 3366
rect 3272 3362 3279 3366
rect 3087 3353 3279 3362
rect 3087 3301 3093 3353
rect 3145 3301 3157 3353
rect 3209 3301 3221 3353
rect 3273 3301 3279 3353
rect 3087 3288 3094 3301
rect 3128 3288 3166 3301
rect 3200 3288 3238 3301
rect 3272 3288 3279 3301
rect 3087 3236 3093 3288
rect 3145 3236 3157 3288
rect 3209 3236 3221 3288
rect 3273 3236 3279 3288
rect 3087 3223 3094 3236
rect 3128 3223 3166 3236
rect 3200 3223 3238 3236
rect 3272 3223 3279 3236
rect 3087 3171 3093 3223
rect 3145 3171 3157 3223
rect 3209 3171 3221 3223
rect 3273 3171 3279 3223
rect 3087 3158 3094 3171
rect 3128 3158 3166 3171
rect 3200 3158 3238 3171
rect 3272 3158 3279 3171
rect 3087 3106 3093 3158
rect 3145 3106 3157 3158
rect 3209 3106 3221 3158
rect 3273 3106 3279 3158
rect 3087 3100 3279 3106
rect 3087 3093 3094 3100
rect 3128 3093 3166 3100
rect 3200 3093 3238 3100
rect 3272 3093 3279 3100
rect 3087 3041 3093 3093
rect 3145 3041 3157 3093
rect 3209 3041 3221 3093
rect 3273 3041 3279 3093
rect 3087 3028 3279 3041
rect 3087 2976 3093 3028
rect 3145 2976 3157 3028
rect 3209 2976 3221 3028
rect 3273 2976 3279 3028
rect 3087 2963 3279 2976
rect 3087 2911 3093 2963
rect 3145 2911 3157 2963
rect 3209 2911 3221 2963
rect 3273 2911 3279 2963
rect 3087 2898 3279 2911
rect 3087 2846 3093 2898
rect 3145 2846 3157 2898
rect 3209 2846 3221 2898
rect 3273 2846 3279 2898
rect 3087 2844 3094 2846
rect 3128 2844 3166 2846
rect 3200 2844 3238 2846
rect 3272 2844 3279 2846
rect 3087 2833 3279 2844
rect 3087 2781 3093 2833
rect 3145 2781 3157 2833
rect 3209 2781 3221 2833
rect 3273 2781 3279 2833
rect 3087 2770 3094 2781
rect 3128 2770 3166 2781
rect 3200 2770 3238 2781
rect 3272 2770 3279 2781
rect 3087 2768 3279 2770
rect 3087 2716 3093 2768
rect 3145 2716 3157 2768
rect 3209 2716 3221 2768
rect 3273 2716 3279 2768
rect 3087 2703 3094 2716
rect 3128 2703 3166 2716
rect 3200 2703 3238 2716
rect 3272 2703 3279 2716
rect 3087 2651 3093 2703
rect 3145 2651 3157 2703
rect 3209 2651 3221 2703
rect 3273 2651 3279 2703
rect 3087 2638 3094 2651
rect 3128 2638 3166 2651
rect 3200 2638 3238 2651
rect 3272 2638 3279 2651
rect 3087 2586 3093 2638
rect 3145 2586 3157 2638
rect 3209 2586 3221 2638
rect 3273 2586 3279 2638
rect 3087 2582 3279 2586
rect 3087 2573 3094 2582
rect 3128 2573 3166 2582
rect 3200 2573 3238 2582
rect 3272 2573 3279 2582
rect 3087 2521 3093 2573
rect 3145 2521 3157 2573
rect 3209 2521 3221 2573
rect 3273 2521 3279 2573
rect 3087 2508 3279 2521
rect 3087 2456 3093 2508
rect 3145 2456 3157 2508
rect 3209 2456 3221 2508
rect 3273 2456 3279 2508
rect 3087 2443 3279 2456
rect 3087 2391 3093 2443
rect 3145 2391 3157 2443
rect 3209 2391 3221 2443
rect 3273 2391 3279 2443
rect 3087 2378 3279 2391
rect 3087 2326 3093 2378
rect 3145 2326 3157 2378
rect 3209 2326 3221 2378
rect 3273 2326 3279 2378
rect 3087 2313 3279 2326
rect 3087 2261 3093 2313
rect 3145 2261 3157 2313
rect 3209 2261 3221 2313
rect 3273 2261 3279 2313
rect 3087 2252 3094 2261
rect 3128 2252 3166 2261
rect 3200 2252 3238 2261
rect 3272 2252 3279 2261
rect 3087 2248 3279 2252
rect 3087 2196 3093 2248
rect 3145 2196 3157 2248
rect 3209 2196 3221 2248
rect 3273 2196 3279 2248
rect 3087 2183 3094 2196
rect 3128 2183 3166 2196
rect 3200 2183 3238 2196
rect 3272 2183 3279 2196
rect 3087 2131 3093 2183
rect 3145 2131 3157 2183
rect 3209 2131 3221 2183
rect 3273 2131 3279 2183
rect 3087 2118 3094 2131
rect 3128 2118 3166 2131
rect 3200 2118 3238 2131
rect 3272 2118 3279 2131
rect 3087 2066 3093 2118
rect 3145 2066 3157 2118
rect 3209 2066 3221 2118
rect 3273 2066 3279 2118
rect 3087 2064 3279 2066
rect 3087 2053 3094 2064
rect 3128 2053 3166 2064
rect 3200 2053 3238 2064
rect 3272 2053 3279 2064
rect 3087 2001 3093 2053
rect 3145 2001 3157 2053
rect 3209 2001 3221 2053
rect 3273 2001 3279 2053
rect 3087 1990 3279 2001
rect 3087 1987 3094 1990
rect 3128 1987 3166 1990
rect 3200 1987 3238 1990
rect 3272 1987 3279 1990
rect 3087 1935 3093 1987
rect 3145 1935 3157 1987
rect 3209 1935 3221 1987
rect 3273 1935 3279 1987
rect 3087 1921 3279 1935
rect 3087 1869 3093 1921
rect 3145 1869 3157 1921
rect 3209 1869 3221 1921
rect 3273 1869 3279 1921
rect 3087 1855 3279 1869
rect 3087 1803 3093 1855
rect 3145 1803 3157 1855
rect 3209 1803 3221 1855
rect 3273 1803 3279 1855
rect 3087 1789 3279 1803
rect 3087 1737 3093 1789
rect 3145 1737 3157 1789
rect 3209 1737 3221 1789
rect 3273 1737 3279 1789
rect 3087 1734 3094 1737
rect 3128 1734 3166 1737
rect 3200 1734 3238 1737
rect 3272 1734 3279 1737
rect 3087 1723 3279 1734
rect 3087 1671 3093 1723
rect 3145 1671 3157 1723
rect 3209 1671 3221 1723
rect 3273 1671 3279 1723
rect 3087 1660 3094 1671
rect 3128 1660 3166 1671
rect 3200 1660 3238 1671
rect 3272 1660 3279 1671
rect 3087 1657 3279 1660
rect 3087 1605 3093 1657
rect 3145 1605 3157 1657
rect 3209 1605 3221 1657
rect 3273 1605 3279 1657
rect 3087 1591 3094 1605
rect 3128 1591 3166 1605
rect 3200 1591 3238 1605
rect 3272 1591 3279 1605
rect 3087 1539 3093 1591
rect 3145 1539 3157 1591
rect 3209 1539 3221 1591
rect 3273 1539 3279 1591
rect 3087 1525 3094 1539
rect 3128 1525 3166 1539
rect 3200 1525 3238 1539
rect 3272 1525 3279 1539
rect 3087 1473 3093 1525
rect 3145 1473 3157 1525
rect 3209 1473 3221 1525
rect 3273 1473 3279 1525
rect 3087 1467 3279 1473
rect 3583 4068 3775 4074
rect 3583 4016 3589 4068
rect 3641 4050 3653 4068
rect 3705 4050 3717 4068
rect 3769 4016 3775 4068
rect 3583 4003 3590 4016
rect 3768 4003 3775 4016
rect 3583 3951 3589 4003
rect 3769 3951 3775 4003
rect 3583 3938 3590 3951
rect 3768 3938 3775 3951
rect 3583 3886 3589 3938
rect 3769 3886 3775 3938
rect 3583 3873 3590 3886
rect 3768 3873 3775 3886
rect 3583 3821 3589 3873
rect 3769 3821 3775 3873
rect 3583 3808 3590 3821
rect 3768 3808 3775 3821
rect 3583 3756 3589 3808
rect 3769 3756 3775 3808
rect 3583 3743 3590 3756
rect 3768 3743 3775 3756
rect 3583 3691 3589 3743
rect 3769 3691 3775 3743
rect 3583 3678 3590 3691
rect 3768 3678 3775 3691
rect 3583 3626 3589 3678
rect 3769 3626 3775 3678
rect 3583 3613 3590 3626
rect 3768 3613 3775 3626
rect 3583 3561 3589 3613
rect 3769 3561 3775 3613
rect 3583 3548 3590 3561
rect 3768 3548 3775 3561
rect 3583 3496 3589 3548
rect 3769 3496 3775 3548
rect 3583 3483 3590 3496
rect 3768 3483 3775 3496
rect 3583 3431 3589 3483
rect 3769 3431 3775 3483
rect 3583 3418 3590 3431
rect 3768 3418 3775 3431
rect 3583 3366 3589 3418
rect 3769 3366 3775 3418
rect 3583 3353 3590 3366
rect 3768 3353 3775 3366
rect 3583 3301 3589 3353
rect 3769 3301 3775 3353
rect 3583 3288 3590 3301
rect 3768 3288 3775 3301
rect 3583 3236 3589 3288
rect 3769 3236 3775 3288
rect 3583 3223 3590 3236
rect 3768 3223 3775 3236
rect 3583 3171 3589 3223
rect 3769 3171 3775 3223
rect 3583 3158 3590 3171
rect 3768 3158 3775 3171
rect 3583 3106 3589 3158
rect 3769 3106 3775 3158
rect 3583 3093 3590 3106
rect 3768 3093 3775 3106
rect 3583 3041 3589 3093
rect 3641 3041 3653 3092
rect 3705 3041 3717 3092
rect 3769 3041 3775 3093
rect 3583 3040 3775 3041
rect 3583 3028 3590 3040
rect 3768 3028 3775 3040
rect 3583 2976 3589 3028
rect 3769 2976 3775 3028
rect 3583 2963 3590 2976
rect 3768 2963 3775 2976
rect 3583 2911 3589 2963
rect 3769 2911 3775 2963
rect 3583 2898 3590 2911
rect 3768 2898 3775 2911
rect 3583 2846 3589 2898
rect 3769 2846 3775 2898
rect 3583 2833 3590 2846
rect 3768 2833 3775 2846
rect 3583 2781 3589 2833
rect 3769 2781 3775 2833
rect 3583 2768 3590 2781
rect 3768 2768 3775 2781
rect 3583 2716 3589 2768
rect 3769 2716 3775 2768
rect 3583 2703 3590 2716
rect 3768 2703 3775 2716
rect 3583 2651 3589 2703
rect 3769 2651 3775 2703
rect 3583 2638 3590 2651
rect 3768 2638 3775 2651
rect 3583 2586 3589 2638
rect 3769 2586 3775 2638
rect 3583 2574 3590 2586
rect 3768 2574 3775 2586
rect 3583 2573 3775 2574
rect 3583 2521 3589 2573
rect 3641 2521 3653 2573
rect 3705 2521 3717 2573
rect 3769 2521 3775 2573
rect 3583 2508 3590 2521
rect 3624 2508 3662 2521
rect 3696 2508 3734 2521
rect 3768 2508 3775 2521
rect 3583 2456 3589 2508
rect 3641 2456 3653 2508
rect 3705 2456 3717 2508
rect 3769 2456 3775 2508
rect 3583 2449 3662 2456
rect 3696 2449 3775 2456
rect 3583 2443 3590 2449
rect 3768 2443 3775 2449
rect 3583 2391 3589 2443
rect 3769 2391 3775 2443
rect 3583 2378 3590 2391
rect 3768 2378 3775 2391
rect 3583 2326 3589 2378
rect 3769 2326 3775 2378
rect 3583 2313 3590 2326
rect 3768 2313 3775 2326
rect 3583 2261 3589 2313
rect 3769 2261 3775 2313
rect 3583 2248 3590 2261
rect 3768 2248 3775 2261
rect 3583 2196 3589 2248
rect 3769 2196 3775 2248
rect 3583 2183 3590 2196
rect 3768 2183 3775 2196
rect 3583 2131 3589 2183
rect 3769 2131 3775 2183
rect 3583 2118 3590 2131
rect 3768 2118 3775 2131
rect 3583 2066 3589 2118
rect 3769 2066 3775 2118
rect 3583 2053 3590 2066
rect 3768 2053 3775 2066
rect 3583 2001 3589 2053
rect 3769 2001 3775 2053
rect 3583 1987 3590 2001
rect 3768 1987 3775 2001
rect 3583 1935 3589 1987
rect 3769 1935 3775 1987
rect 3583 1921 3590 1935
rect 3768 1921 3775 1935
rect 3583 1869 3589 1921
rect 3769 1869 3775 1921
rect 3583 1855 3590 1869
rect 3768 1855 3775 1869
rect 3583 1803 3589 1855
rect 3769 1803 3775 1855
rect 3583 1789 3590 1803
rect 3768 1789 3775 1803
rect 3583 1737 3589 1789
rect 3769 1737 3775 1789
rect 3583 1723 3590 1737
rect 3768 1723 3775 1737
rect 3583 1671 3589 1723
rect 3769 1671 3775 1723
rect 3583 1657 3590 1671
rect 3768 1657 3775 1671
rect 3583 1605 3589 1657
rect 3769 1605 3775 1657
rect 3583 1591 3590 1605
rect 3768 1591 3775 1605
rect 3583 1539 3589 1591
rect 3769 1539 3775 1591
rect 3583 1525 3590 1539
rect 3768 1525 3775 1539
rect 3583 1473 3589 1525
rect 3641 1473 3653 1491
rect 3705 1473 3717 1491
rect 3769 1473 3775 1525
rect 3583 1467 3775 1473
rect 4079 4068 4271 4074
rect 4079 4016 4085 4068
rect 4137 4016 4149 4068
rect 4201 4016 4213 4068
rect 4265 4016 4271 4068
rect 4079 4003 4271 4016
rect 4079 3951 4085 4003
rect 4137 3951 4149 4003
rect 4201 3951 4213 4003
rect 4265 3951 4271 4003
rect 4079 3938 4271 3951
rect 4079 3886 4085 3938
rect 4137 3886 4149 3938
rect 4201 3886 4213 3938
rect 4265 3886 4271 3938
rect 4079 3880 4086 3886
rect 4120 3880 4158 3886
rect 4192 3880 4230 3886
rect 4264 3880 4271 3886
rect 4079 3873 4271 3880
rect 4079 3821 4085 3873
rect 4137 3821 4149 3873
rect 4201 3821 4213 3873
rect 4265 3821 4271 3873
rect 4079 3808 4086 3821
rect 4120 3808 4158 3821
rect 4192 3808 4230 3821
rect 4264 3808 4271 3821
rect 4079 3756 4085 3808
rect 4137 3756 4149 3808
rect 4201 3756 4213 3808
rect 4265 3756 4271 3808
rect 4079 3743 4086 3756
rect 4120 3743 4158 3756
rect 4192 3743 4230 3756
rect 4264 3743 4271 3756
rect 4079 3691 4085 3743
rect 4137 3691 4149 3743
rect 4201 3691 4213 3743
rect 4265 3691 4271 3743
rect 4079 3678 4086 3691
rect 4120 3678 4158 3691
rect 4192 3678 4230 3691
rect 4264 3678 4271 3691
rect 4079 3626 4085 3678
rect 4137 3626 4149 3678
rect 4201 3626 4213 3678
rect 4265 3626 4271 3678
rect 4079 3618 4271 3626
rect 4079 3613 4086 3618
rect 4120 3613 4158 3618
rect 4192 3613 4230 3618
rect 4264 3613 4271 3618
rect 4079 3561 4085 3613
rect 4137 3561 4149 3613
rect 4201 3561 4213 3613
rect 4265 3561 4271 3613
rect 4079 3548 4271 3561
rect 4079 3496 4085 3548
rect 4137 3496 4149 3548
rect 4201 3496 4213 3548
rect 4265 3496 4271 3548
rect 4079 3483 4271 3496
rect 4079 3431 4085 3483
rect 4137 3431 4149 3483
rect 4201 3431 4213 3483
rect 4265 3431 4271 3483
rect 4079 3418 4271 3431
rect 4079 3366 4085 3418
rect 4137 3366 4149 3418
rect 4201 3366 4213 3418
rect 4265 3366 4271 3418
rect 4079 3362 4086 3366
rect 4120 3362 4158 3366
rect 4192 3362 4230 3366
rect 4264 3362 4271 3366
rect 4079 3353 4271 3362
rect 4079 3301 4085 3353
rect 4137 3301 4149 3353
rect 4201 3301 4213 3353
rect 4265 3301 4271 3353
rect 4079 3288 4086 3301
rect 4120 3288 4158 3301
rect 4192 3288 4230 3301
rect 4264 3288 4271 3301
rect 4079 3236 4085 3288
rect 4137 3236 4149 3288
rect 4201 3236 4213 3288
rect 4265 3236 4271 3288
rect 4079 3223 4086 3236
rect 4120 3223 4158 3236
rect 4192 3223 4230 3236
rect 4264 3223 4271 3236
rect 4079 3171 4085 3223
rect 4137 3171 4149 3223
rect 4201 3171 4213 3223
rect 4265 3171 4271 3223
rect 4079 3158 4086 3171
rect 4120 3158 4158 3171
rect 4192 3158 4230 3171
rect 4264 3158 4271 3171
rect 4079 3106 4085 3158
rect 4137 3106 4149 3158
rect 4201 3106 4213 3158
rect 4265 3106 4271 3158
rect 4079 3100 4271 3106
rect 4079 3093 4086 3100
rect 4120 3093 4158 3100
rect 4192 3093 4230 3100
rect 4264 3093 4271 3100
rect 4079 3041 4085 3093
rect 4137 3041 4149 3093
rect 4201 3041 4213 3093
rect 4265 3041 4271 3093
rect 4079 3028 4271 3041
rect 4079 2976 4085 3028
rect 4137 2976 4149 3028
rect 4201 2976 4213 3028
rect 4265 2976 4271 3028
rect 4079 2963 4271 2976
rect 4079 2911 4085 2963
rect 4137 2911 4149 2963
rect 4201 2911 4213 2963
rect 4265 2911 4271 2963
rect 4079 2898 4271 2911
rect 4079 2846 4085 2898
rect 4137 2846 4149 2898
rect 4201 2846 4213 2898
rect 4265 2846 4271 2898
rect 4079 2844 4086 2846
rect 4120 2844 4158 2846
rect 4192 2844 4230 2846
rect 4264 2844 4271 2846
rect 4079 2833 4271 2844
rect 4079 2781 4085 2833
rect 4137 2781 4149 2833
rect 4201 2781 4213 2833
rect 4265 2781 4271 2833
rect 4079 2770 4086 2781
rect 4120 2770 4158 2781
rect 4192 2770 4230 2781
rect 4264 2770 4271 2781
rect 4079 2768 4271 2770
rect 4079 2716 4085 2768
rect 4137 2716 4149 2768
rect 4201 2716 4213 2768
rect 4265 2716 4271 2768
rect 4079 2703 4086 2716
rect 4120 2703 4158 2716
rect 4192 2703 4230 2716
rect 4264 2703 4271 2716
rect 4079 2651 4085 2703
rect 4137 2651 4149 2703
rect 4201 2651 4213 2703
rect 4265 2651 4271 2703
rect 4079 2638 4086 2651
rect 4120 2638 4158 2651
rect 4192 2638 4230 2651
rect 4264 2638 4271 2651
rect 4079 2586 4085 2638
rect 4137 2586 4149 2638
rect 4201 2586 4213 2638
rect 4265 2586 4271 2638
rect 4079 2582 4271 2586
rect 4079 2573 4086 2582
rect 4120 2573 4158 2582
rect 4192 2573 4230 2582
rect 4264 2573 4271 2582
rect 4079 2521 4085 2573
rect 4137 2521 4149 2573
rect 4201 2521 4213 2573
rect 4265 2521 4271 2573
rect 4079 2508 4271 2521
rect 4079 2456 4085 2508
rect 4137 2456 4149 2508
rect 4201 2456 4213 2508
rect 4265 2456 4271 2508
rect 4079 2443 4271 2456
rect 4079 2391 4085 2443
rect 4137 2391 4149 2443
rect 4201 2391 4213 2443
rect 4265 2391 4271 2443
rect 4079 2378 4271 2391
rect 4079 2326 4085 2378
rect 4137 2326 4149 2378
rect 4201 2326 4213 2378
rect 4265 2326 4271 2378
rect 4079 2313 4271 2326
rect 4079 2261 4085 2313
rect 4137 2261 4149 2313
rect 4201 2261 4213 2313
rect 4265 2261 4271 2313
rect 4079 2252 4086 2261
rect 4120 2252 4158 2261
rect 4192 2252 4230 2261
rect 4264 2252 4271 2261
rect 4079 2248 4271 2252
rect 4079 2196 4085 2248
rect 4137 2196 4149 2248
rect 4201 2196 4213 2248
rect 4265 2196 4271 2248
rect 4079 2183 4086 2196
rect 4120 2183 4158 2196
rect 4192 2183 4230 2196
rect 4264 2183 4271 2196
rect 4079 2131 4085 2183
rect 4137 2131 4149 2183
rect 4201 2131 4213 2183
rect 4265 2131 4271 2183
rect 4079 2118 4086 2131
rect 4120 2118 4158 2131
rect 4192 2118 4230 2131
rect 4264 2118 4271 2131
rect 4079 2066 4085 2118
rect 4137 2066 4149 2118
rect 4201 2066 4213 2118
rect 4265 2066 4271 2118
rect 4079 2064 4271 2066
rect 4079 2053 4086 2064
rect 4120 2053 4158 2064
rect 4192 2053 4230 2064
rect 4264 2053 4271 2064
rect 4079 2001 4085 2053
rect 4137 2001 4149 2053
rect 4201 2001 4213 2053
rect 4265 2001 4271 2053
rect 4079 1990 4271 2001
rect 4079 1987 4086 1990
rect 4120 1987 4158 1990
rect 4192 1987 4230 1990
rect 4264 1987 4271 1990
rect 4079 1935 4085 1987
rect 4137 1935 4149 1987
rect 4201 1935 4213 1987
rect 4265 1935 4271 1987
rect 4079 1921 4271 1935
rect 4079 1869 4085 1921
rect 4137 1869 4149 1921
rect 4201 1869 4213 1921
rect 4265 1869 4271 1921
rect 4079 1855 4271 1869
rect 4079 1803 4085 1855
rect 4137 1803 4149 1855
rect 4201 1803 4213 1855
rect 4265 1803 4271 1855
rect 4079 1789 4271 1803
rect 4079 1737 4085 1789
rect 4137 1737 4149 1789
rect 4201 1737 4213 1789
rect 4265 1737 4271 1789
rect 4079 1734 4086 1737
rect 4120 1734 4158 1737
rect 4192 1734 4230 1737
rect 4264 1734 4271 1737
rect 4079 1723 4271 1734
rect 4079 1671 4085 1723
rect 4137 1671 4149 1723
rect 4201 1671 4213 1723
rect 4265 1671 4271 1723
rect 4079 1660 4086 1671
rect 4120 1660 4158 1671
rect 4192 1660 4230 1671
rect 4264 1660 4271 1671
rect 4079 1657 4271 1660
rect 4079 1605 4085 1657
rect 4137 1605 4149 1657
rect 4201 1605 4213 1657
rect 4265 1605 4271 1657
rect 4079 1591 4086 1605
rect 4120 1591 4158 1605
rect 4192 1591 4230 1605
rect 4264 1591 4271 1605
rect 4079 1539 4085 1591
rect 4137 1539 4149 1591
rect 4201 1539 4213 1591
rect 4265 1539 4271 1591
rect 4079 1525 4086 1539
rect 4120 1525 4158 1539
rect 4192 1525 4230 1539
rect 4264 1525 4271 1539
rect 4079 1473 4085 1525
rect 4137 1473 4149 1525
rect 4201 1473 4213 1525
rect 4265 1473 4271 1525
rect 4079 1467 4271 1473
rect 4575 4068 4767 4074
rect 4575 4016 4581 4068
rect 4633 4050 4645 4068
rect 4697 4050 4709 4068
rect 4761 4016 4767 4068
rect 4575 4003 4582 4016
rect 4760 4003 4767 4016
rect 4575 3951 4581 4003
rect 4761 3951 4767 4003
rect 4575 3938 4582 3951
rect 4760 3938 4767 3951
rect 4575 3886 4581 3938
rect 4761 3886 4767 3938
rect 4575 3873 4582 3886
rect 4760 3873 4767 3886
rect 4575 3821 4581 3873
rect 4761 3821 4767 3873
rect 4575 3808 4582 3821
rect 4760 3808 4767 3821
rect 4575 3756 4581 3808
rect 4761 3756 4767 3808
rect 4575 3743 4582 3756
rect 4760 3743 4767 3756
rect 4575 3691 4581 3743
rect 4761 3691 4767 3743
rect 4575 3678 4582 3691
rect 4760 3678 4767 3691
rect 4575 3626 4581 3678
rect 4761 3626 4767 3678
rect 4575 3613 4582 3626
rect 4760 3613 4767 3626
rect 4575 3561 4581 3613
rect 4761 3561 4767 3613
rect 4575 3548 4582 3561
rect 4760 3548 4767 3561
rect 4575 3496 4581 3548
rect 4761 3496 4767 3548
rect 4575 3483 4582 3496
rect 4760 3483 4767 3496
rect 4575 3431 4581 3483
rect 4761 3431 4767 3483
rect 4575 3418 4582 3431
rect 4760 3418 4767 3431
rect 4575 3366 4581 3418
rect 4761 3366 4767 3418
rect 4575 3353 4582 3366
rect 4760 3353 4767 3366
rect 4575 3301 4581 3353
rect 4761 3301 4767 3353
rect 4575 3288 4582 3301
rect 4760 3288 4767 3301
rect 4575 3236 4581 3288
rect 4761 3236 4767 3288
rect 4575 3223 4582 3236
rect 4760 3223 4767 3236
rect 4575 3171 4581 3223
rect 4761 3171 4767 3223
rect 4575 3158 4582 3171
rect 4760 3158 4767 3171
rect 4575 3106 4581 3158
rect 4761 3106 4767 3158
rect 4575 3093 4582 3106
rect 4760 3093 4767 3106
rect 4575 3041 4581 3093
rect 4633 3041 4645 3092
rect 4697 3041 4709 3092
rect 4761 3041 4767 3093
rect 4575 3040 4767 3041
rect 4575 3028 4582 3040
rect 4760 3028 4767 3040
rect 4575 2976 4581 3028
rect 4761 2976 4767 3028
rect 4575 2963 4582 2976
rect 4760 2963 4767 2976
rect 4575 2911 4581 2963
rect 4761 2911 4767 2963
rect 4575 2898 4582 2911
rect 4760 2898 4767 2911
rect 4575 2846 4581 2898
rect 4761 2846 4767 2898
rect 4575 2833 4582 2846
rect 4760 2833 4767 2846
rect 4575 2781 4581 2833
rect 4761 2781 4767 2833
rect 4575 2768 4582 2781
rect 4760 2768 4767 2781
rect 4575 2716 4581 2768
rect 4761 2716 4767 2768
rect 4575 2703 4582 2716
rect 4760 2703 4767 2716
rect 4575 2651 4581 2703
rect 4761 2651 4767 2703
rect 4575 2638 4582 2651
rect 4760 2638 4767 2651
rect 4575 2586 4581 2638
rect 4761 2586 4767 2638
rect 4575 2574 4582 2586
rect 4760 2574 4767 2586
rect 4575 2573 4767 2574
rect 4575 2521 4581 2573
rect 4633 2521 4645 2573
rect 4697 2521 4709 2573
rect 4761 2521 4767 2573
rect 4575 2508 4582 2521
rect 4616 2508 4654 2521
rect 4688 2508 4726 2521
rect 4760 2508 4767 2521
rect 4575 2456 4581 2508
rect 4633 2456 4645 2508
rect 4697 2456 4709 2508
rect 4761 2456 4767 2508
rect 4575 2449 4654 2456
rect 4688 2449 4767 2456
rect 4575 2443 4582 2449
rect 4760 2443 4767 2449
rect 4575 2391 4581 2443
rect 4761 2391 4767 2443
rect 4575 2378 4582 2391
rect 4760 2378 4767 2391
rect 4575 2326 4581 2378
rect 4761 2326 4767 2378
rect 4575 2313 4582 2326
rect 4760 2313 4767 2326
rect 4575 2261 4581 2313
rect 4761 2261 4767 2313
rect 4575 2248 4582 2261
rect 4760 2248 4767 2261
rect 4575 2196 4581 2248
rect 4761 2196 4767 2248
rect 4575 2183 4582 2196
rect 4760 2183 4767 2196
rect 4575 2131 4581 2183
rect 4761 2131 4767 2183
rect 4575 2118 4582 2131
rect 4760 2118 4767 2131
rect 4575 2066 4581 2118
rect 4761 2066 4767 2118
rect 4575 2053 4582 2066
rect 4760 2053 4767 2066
rect 4575 2001 4581 2053
rect 4761 2001 4767 2053
rect 4575 1987 4582 2001
rect 4760 1987 4767 2001
rect 4575 1935 4581 1987
rect 4761 1935 4767 1987
rect 4575 1921 4582 1935
rect 4760 1921 4767 1935
rect 4575 1869 4581 1921
rect 4761 1869 4767 1921
rect 4575 1855 4582 1869
rect 4760 1855 4767 1869
rect 4575 1803 4581 1855
rect 4761 1803 4767 1855
rect 4575 1789 4582 1803
rect 4760 1789 4767 1803
rect 4575 1737 4581 1789
rect 4761 1737 4767 1789
rect 4575 1723 4582 1737
rect 4760 1723 4767 1737
rect 4575 1671 4581 1723
rect 4761 1671 4767 1723
rect 4575 1657 4582 1671
rect 4760 1657 4767 1671
rect 4575 1605 4581 1657
rect 4761 1605 4767 1657
rect 4575 1591 4582 1605
rect 4760 1591 4767 1605
rect 4575 1539 4581 1591
rect 4761 1539 4767 1591
rect 4575 1525 4582 1539
rect 4760 1525 4767 1539
rect 4575 1473 4581 1525
rect 4633 1473 4645 1491
rect 4697 1473 4709 1491
rect 4761 1473 4767 1525
rect 4575 1467 4767 1473
rect 5071 4068 5263 4074
rect 5071 4016 5077 4068
rect 5129 4016 5141 4068
rect 5193 4016 5205 4068
rect 5257 4016 5263 4068
rect 5071 4003 5263 4016
rect 5071 3951 5077 4003
rect 5129 3951 5141 4003
rect 5193 3951 5205 4003
rect 5257 3951 5263 4003
rect 5071 3938 5263 3951
rect 5071 3886 5077 3938
rect 5129 3886 5141 3938
rect 5193 3886 5205 3938
rect 5257 3886 5263 3938
rect 5071 3880 5078 3886
rect 5112 3880 5150 3886
rect 5184 3880 5222 3886
rect 5256 3880 5263 3886
rect 5071 3873 5263 3880
rect 5071 3821 5077 3873
rect 5129 3821 5141 3873
rect 5193 3821 5205 3873
rect 5257 3821 5263 3873
rect 5071 3808 5078 3821
rect 5112 3808 5150 3821
rect 5184 3808 5222 3821
rect 5256 3808 5263 3821
rect 5071 3756 5077 3808
rect 5129 3756 5141 3808
rect 5193 3756 5205 3808
rect 5257 3756 5263 3808
rect 5071 3743 5078 3756
rect 5112 3743 5150 3756
rect 5184 3743 5222 3756
rect 5256 3743 5263 3756
rect 5071 3691 5077 3743
rect 5129 3691 5141 3743
rect 5193 3691 5205 3743
rect 5257 3691 5263 3743
rect 5071 3678 5078 3691
rect 5112 3678 5150 3691
rect 5184 3678 5222 3691
rect 5256 3678 5263 3691
rect 5071 3626 5077 3678
rect 5129 3626 5141 3678
rect 5193 3626 5205 3678
rect 5257 3626 5263 3678
rect 5071 3618 5263 3626
rect 5071 3613 5078 3618
rect 5112 3613 5150 3618
rect 5184 3613 5222 3618
rect 5256 3613 5263 3618
rect 5071 3561 5077 3613
rect 5129 3561 5141 3613
rect 5193 3561 5205 3613
rect 5257 3561 5263 3613
rect 5071 3548 5263 3561
rect 5071 3496 5077 3548
rect 5129 3496 5141 3548
rect 5193 3496 5205 3548
rect 5257 3496 5263 3548
rect 5071 3483 5263 3496
rect 5071 3431 5077 3483
rect 5129 3431 5141 3483
rect 5193 3431 5205 3483
rect 5257 3431 5263 3483
rect 5071 3418 5263 3431
rect 5071 3366 5077 3418
rect 5129 3366 5141 3418
rect 5193 3366 5205 3418
rect 5257 3366 5263 3418
rect 5071 3362 5078 3366
rect 5112 3362 5150 3366
rect 5184 3362 5222 3366
rect 5256 3362 5263 3366
rect 5071 3353 5263 3362
rect 5071 3301 5077 3353
rect 5129 3301 5141 3353
rect 5193 3301 5205 3353
rect 5257 3301 5263 3353
rect 5071 3288 5078 3301
rect 5112 3288 5150 3301
rect 5184 3288 5222 3301
rect 5256 3288 5263 3301
rect 5071 3236 5077 3288
rect 5129 3236 5141 3288
rect 5193 3236 5205 3288
rect 5257 3236 5263 3288
rect 5071 3223 5078 3236
rect 5112 3223 5150 3236
rect 5184 3223 5222 3236
rect 5256 3223 5263 3236
rect 5071 3171 5077 3223
rect 5129 3171 5141 3223
rect 5193 3171 5205 3223
rect 5257 3171 5263 3223
rect 5071 3158 5078 3171
rect 5112 3158 5150 3171
rect 5184 3158 5222 3171
rect 5256 3158 5263 3171
rect 5071 3106 5077 3158
rect 5129 3106 5141 3158
rect 5193 3106 5205 3158
rect 5257 3106 5263 3158
rect 5071 3100 5263 3106
rect 5071 3093 5078 3100
rect 5112 3093 5150 3100
rect 5184 3093 5222 3100
rect 5256 3093 5263 3100
rect 5071 3041 5077 3093
rect 5129 3041 5141 3093
rect 5193 3041 5205 3093
rect 5257 3041 5263 3093
rect 5071 3028 5263 3041
rect 5071 2976 5077 3028
rect 5129 2976 5141 3028
rect 5193 2976 5205 3028
rect 5257 2976 5263 3028
rect 5071 2963 5263 2976
rect 5071 2911 5077 2963
rect 5129 2911 5141 2963
rect 5193 2911 5205 2963
rect 5257 2911 5263 2963
rect 5071 2898 5263 2911
rect 5071 2846 5077 2898
rect 5129 2846 5141 2898
rect 5193 2846 5205 2898
rect 5257 2846 5263 2898
rect 5071 2844 5078 2846
rect 5112 2844 5150 2846
rect 5184 2844 5222 2846
rect 5256 2844 5263 2846
rect 5071 2833 5263 2844
rect 5071 2781 5077 2833
rect 5129 2781 5141 2833
rect 5193 2781 5205 2833
rect 5257 2781 5263 2833
rect 5071 2770 5078 2781
rect 5112 2770 5150 2781
rect 5184 2770 5222 2781
rect 5256 2770 5263 2781
rect 5071 2768 5263 2770
rect 5071 2716 5077 2768
rect 5129 2716 5141 2768
rect 5193 2716 5205 2768
rect 5257 2716 5263 2768
rect 5071 2703 5078 2716
rect 5112 2703 5150 2716
rect 5184 2703 5222 2716
rect 5256 2703 5263 2716
rect 5071 2651 5077 2703
rect 5129 2651 5141 2703
rect 5193 2651 5205 2703
rect 5257 2651 5263 2703
rect 5071 2638 5078 2651
rect 5112 2638 5150 2651
rect 5184 2638 5222 2651
rect 5256 2638 5263 2651
rect 5071 2586 5077 2638
rect 5129 2586 5141 2638
rect 5193 2586 5205 2638
rect 5257 2586 5263 2638
rect 5071 2582 5263 2586
rect 5071 2573 5078 2582
rect 5112 2573 5150 2582
rect 5184 2573 5222 2582
rect 5256 2573 5263 2582
rect 5071 2521 5077 2573
rect 5129 2521 5141 2573
rect 5193 2521 5205 2573
rect 5257 2521 5263 2573
rect 5071 2508 5263 2521
rect 5071 2456 5077 2508
rect 5129 2456 5141 2508
rect 5193 2456 5205 2508
rect 5257 2456 5263 2508
rect 5071 2443 5263 2456
rect 5071 2391 5077 2443
rect 5129 2391 5141 2443
rect 5193 2391 5205 2443
rect 5257 2391 5263 2443
rect 5071 2378 5263 2391
rect 5071 2326 5077 2378
rect 5129 2326 5141 2378
rect 5193 2326 5205 2378
rect 5257 2326 5263 2378
rect 5071 2313 5263 2326
rect 5071 2261 5077 2313
rect 5129 2261 5141 2313
rect 5193 2261 5205 2313
rect 5257 2261 5263 2313
rect 5071 2252 5078 2261
rect 5112 2252 5150 2261
rect 5184 2252 5222 2261
rect 5256 2252 5263 2261
rect 5071 2248 5263 2252
rect 5071 2196 5077 2248
rect 5129 2196 5141 2248
rect 5193 2196 5205 2248
rect 5257 2196 5263 2248
rect 5071 2183 5078 2196
rect 5112 2183 5150 2196
rect 5184 2183 5222 2196
rect 5256 2183 5263 2196
rect 5071 2131 5077 2183
rect 5129 2131 5141 2183
rect 5193 2131 5205 2183
rect 5257 2131 5263 2183
rect 5071 2118 5078 2131
rect 5112 2118 5150 2131
rect 5184 2118 5222 2131
rect 5256 2118 5263 2131
rect 5071 2066 5077 2118
rect 5129 2066 5141 2118
rect 5193 2066 5205 2118
rect 5257 2066 5263 2118
rect 5071 2064 5263 2066
rect 5071 2053 5078 2064
rect 5112 2053 5150 2064
rect 5184 2053 5222 2064
rect 5256 2053 5263 2064
rect 5071 2001 5077 2053
rect 5129 2001 5141 2053
rect 5193 2001 5205 2053
rect 5257 2001 5263 2053
rect 5071 1990 5263 2001
rect 5071 1987 5078 1990
rect 5112 1987 5150 1990
rect 5184 1987 5222 1990
rect 5256 1987 5263 1990
rect 5071 1935 5077 1987
rect 5129 1935 5141 1987
rect 5193 1935 5205 1987
rect 5257 1935 5263 1987
rect 5071 1921 5263 1935
rect 5071 1869 5077 1921
rect 5129 1869 5141 1921
rect 5193 1869 5205 1921
rect 5257 1869 5263 1921
rect 5071 1855 5263 1869
rect 5071 1803 5077 1855
rect 5129 1803 5141 1855
rect 5193 1803 5205 1855
rect 5257 1803 5263 1855
rect 5071 1789 5263 1803
rect 5071 1737 5077 1789
rect 5129 1737 5141 1789
rect 5193 1737 5205 1789
rect 5257 1737 5263 1789
rect 5071 1734 5078 1737
rect 5112 1734 5150 1737
rect 5184 1734 5222 1737
rect 5256 1734 5263 1737
rect 5071 1723 5263 1734
rect 5071 1671 5077 1723
rect 5129 1671 5141 1723
rect 5193 1671 5205 1723
rect 5257 1671 5263 1723
rect 5071 1660 5078 1671
rect 5112 1660 5150 1671
rect 5184 1660 5222 1671
rect 5256 1660 5263 1671
rect 5071 1657 5263 1660
rect 5071 1605 5077 1657
rect 5129 1605 5141 1657
rect 5193 1605 5205 1657
rect 5257 1605 5263 1657
rect 5071 1591 5078 1605
rect 5112 1591 5150 1605
rect 5184 1591 5222 1605
rect 5256 1591 5263 1605
rect 5071 1539 5077 1591
rect 5129 1539 5141 1591
rect 5193 1539 5205 1591
rect 5257 1539 5263 1591
rect 5071 1525 5078 1539
rect 5112 1525 5150 1539
rect 5184 1525 5222 1539
rect 5256 1525 5263 1539
rect 5071 1473 5077 1525
rect 5129 1473 5141 1525
rect 5193 1473 5205 1525
rect 5257 1473 5263 1525
rect 5071 1467 5263 1473
rect 5567 4068 5759 4074
rect 5567 4016 5573 4068
rect 5625 4050 5637 4068
rect 5689 4050 5701 4068
rect 5753 4016 5759 4068
rect 5567 4003 5574 4016
rect 5752 4003 5759 4016
rect 5567 3951 5573 4003
rect 5753 3951 5759 4003
rect 5567 3938 5574 3951
rect 5752 3938 5759 3951
rect 5567 3886 5573 3938
rect 5753 3886 5759 3938
rect 5567 3873 5574 3886
rect 5752 3873 5759 3886
rect 5567 3821 5573 3873
rect 5753 3821 5759 3873
rect 5567 3808 5574 3821
rect 5752 3808 5759 3821
rect 5567 3756 5573 3808
rect 5753 3756 5759 3808
rect 5567 3743 5574 3756
rect 5752 3743 5759 3756
rect 5567 3691 5573 3743
rect 5753 3691 5759 3743
rect 5567 3678 5574 3691
rect 5752 3678 5759 3691
rect 5567 3626 5573 3678
rect 5753 3626 5759 3678
rect 5567 3613 5574 3626
rect 5752 3613 5759 3626
rect 5567 3561 5573 3613
rect 5753 3561 5759 3613
rect 5567 3548 5574 3561
rect 5752 3548 5759 3561
rect 5567 3496 5573 3548
rect 5753 3496 5759 3548
rect 5567 3483 5574 3496
rect 5752 3483 5759 3496
rect 5567 3431 5573 3483
rect 5753 3431 5759 3483
rect 5567 3418 5574 3431
rect 5752 3418 5759 3431
rect 5567 3366 5573 3418
rect 5753 3366 5759 3418
rect 5567 3353 5574 3366
rect 5752 3353 5759 3366
rect 5567 3301 5573 3353
rect 5753 3301 5759 3353
rect 5567 3288 5574 3301
rect 5752 3288 5759 3301
rect 5567 3236 5573 3288
rect 5753 3236 5759 3288
rect 5567 3223 5574 3236
rect 5752 3223 5759 3236
rect 5567 3171 5573 3223
rect 5753 3171 5759 3223
rect 5567 3158 5574 3171
rect 5752 3158 5759 3171
rect 5567 3106 5573 3158
rect 5753 3106 5759 3158
rect 5567 3093 5574 3106
rect 5752 3093 5759 3106
rect 5567 3041 5573 3093
rect 5625 3041 5637 3092
rect 5689 3041 5701 3092
rect 5753 3041 5759 3093
rect 5567 3040 5759 3041
rect 5567 3028 5574 3040
rect 5752 3028 5759 3040
rect 5567 2976 5573 3028
rect 5753 2976 5759 3028
rect 5567 2963 5574 2976
rect 5752 2963 5759 2976
rect 5567 2911 5573 2963
rect 5753 2911 5759 2963
rect 5567 2898 5574 2911
rect 5752 2898 5759 2911
rect 5567 2846 5573 2898
rect 5753 2846 5759 2898
rect 5567 2833 5574 2846
rect 5752 2833 5759 2846
rect 5567 2781 5573 2833
rect 5753 2781 5759 2833
rect 5567 2768 5574 2781
rect 5752 2768 5759 2781
rect 5567 2716 5573 2768
rect 5753 2716 5759 2768
rect 5567 2703 5574 2716
rect 5752 2703 5759 2716
rect 5567 2651 5573 2703
rect 5753 2651 5759 2703
rect 5567 2638 5574 2651
rect 5752 2638 5759 2651
rect 5567 2586 5573 2638
rect 5753 2586 5759 2638
rect 5567 2574 5574 2586
rect 5752 2574 5759 2586
rect 5567 2573 5759 2574
rect 5567 2521 5573 2573
rect 5625 2521 5637 2573
rect 5689 2521 5701 2573
rect 5753 2521 5759 2573
rect 5567 2508 5574 2521
rect 5608 2508 5646 2521
rect 5680 2508 5718 2521
rect 5752 2508 5759 2521
rect 5567 2456 5573 2508
rect 5625 2456 5637 2508
rect 5689 2456 5701 2508
rect 5753 2456 5759 2508
rect 5567 2449 5646 2456
rect 5680 2449 5759 2456
rect 5567 2443 5574 2449
rect 5752 2443 5759 2449
rect 5567 2391 5573 2443
rect 5753 2391 5759 2443
rect 5567 2378 5574 2391
rect 5752 2378 5759 2391
rect 5567 2326 5573 2378
rect 5753 2326 5759 2378
rect 5567 2313 5574 2326
rect 5752 2313 5759 2326
rect 5567 2261 5573 2313
rect 5753 2261 5759 2313
rect 5567 2248 5574 2261
rect 5752 2248 5759 2261
rect 5567 2196 5573 2248
rect 5753 2196 5759 2248
rect 5567 2183 5574 2196
rect 5752 2183 5759 2196
rect 5567 2131 5573 2183
rect 5753 2131 5759 2183
rect 5567 2118 5574 2131
rect 5752 2118 5759 2131
rect 5567 2066 5573 2118
rect 5753 2066 5759 2118
rect 5567 2053 5574 2066
rect 5752 2053 5759 2066
rect 5567 2001 5573 2053
rect 5753 2001 5759 2053
rect 5567 1987 5574 2001
rect 5752 1987 5759 2001
rect 5567 1935 5573 1987
rect 5753 1935 5759 1987
rect 5567 1921 5574 1935
rect 5752 1921 5759 1935
rect 5567 1869 5573 1921
rect 5753 1869 5759 1921
rect 5567 1855 5574 1869
rect 5752 1855 5759 1869
rect 5567 1803 5573 1855
rect 5753 1803 5759 1855
rect 5567 1789 5574 1803
rect 5752 1789 5759 1803
rect 5567 1737 5573 1789
rect 5753 1737 5759 1789
rect 5567 1723 5574 1737
rect 5752 1723 5759 1737
rect 5567 1671 5573 1723
rect 5753 1671 5759 1723
rect 5567 1657 5574 1671
rect 5752 1657 5759 1671
rect 5567 1605 5573 1657
rect 5753 1605 5759 1657
rect 5567 1591 5574 1605
rect 5752 1591 5759 1605
rect 5567 1539 5573 1591
rect 5753 1539 5759 1591
rect 5567 1525 5574 1539
rect 5752 1525 5759 1539
rect 5567 1473 5573 1525
rect 5625 1473 5637 1491
rect 5689 1473 5701 1491
rect 5753 1473 5759 1525
rect 5567 1467 5759 1473
rect 6063 4068 6255 4074
rect 6063 4016 6069 4068
rect 6121 4016 6133 4068
rect 6185 4016 6197 4068
rect 6249 4016 6255 4068
rect 6063 4003 6255 4016
rect 6063 3951 6069 4003
rect 6121 3951 6133 4003
rect 6185 3951 6197 4003
rect 6249 3951 6255 4003
rect 6063 3938 6255 3951
rect 6063 3886 6069 3938
rect 6121 3886 6133 3938
rect 6185 3886 6197 3938
rect 6249 3886 6255 3938
rect 6063 3880 6070 3886
rect 6104 3880 6142 3886
rect 6176 3880 6214 3886
rect 6248 3880 6255 3886
rect 6063 3873 6255 3880
rect 6063 3821 6069 3873
rect 6121 3821 6133 3873
rect 6185 3821 6197 3873
rect 6249 3821 6255 3873
rect 6063 3808 6070 3821
rect 6104 3808 6142 3821
rect 6176 3808 6214 3821
rect 6248 3808 6255 3821
rect 6063 3756 6069 3808
rect 6121 3756 6133 3808
rect 6185 3756 6197 3808
rect 6249 3756 6255 3808
rect 6063 3743 6070 3756
rect 6104 3743 6142 3756
rect 6176 3743 6214 3756
rect 6248 3743 6255 3756
rect 6063 3691 6069 3743
rect 6121 3691 6133 3743
rect 6185 3691 6197 3743
rect 6249 3691 6255 3743
rect 6063 3678 6070 3691
rect 6104 3678 6142 3691
rect 6176 3678 6214 3691
rect 6248 3678 6255 3691
rect 6063 3626 6069 3678
rect 6121 3626 6133 3678
rect 6185 3626 6197 3678
rect 6249 3626 6255 3678
rect 6063 3618 6255 3626
rect 6063 3613 6070 3618
rect 6104 3613 6142 3618
rect 6176 3613 6214 3618
rect 6248 3613 6255 3618
rect 6063 3561 6069 3613
rect 6121 3561 6133 3613
rect 6185 3561 6197 3613
rect 6249 3561 6255 3613
rect 6063 3548 6255 3561
rect 6063 3496 6069 3548
rect 6121 3496 6133 3548
rect 6185 3496 6197 3548
rect 6249 3496 6255 3548
rect 6063 3483 6255 3496
rect 6063 3431 6069 3483
rect 6121 3431 6133 3483
rect 6185 3431 6197 3483
rect 6249 3431 6255 3483
rect 6063 3418 6255 3431
rect 6063 3366 6069 3418
rect 6121 3366 6133 3418
rect 6185 3366 6197 3418
rect 6249 3366 6255 3418
rect 6063 3362 6070 3366
rect 6104 3362 6142 3366
rect 6176 3362 6214 3366
rect 6248 3362 6255 3366
rect 6063 3353 6255 3362
rect 6063 3301 6069 3353
rect 6121 3301 6133 3353
rect 6185 3301 6197 3353
rect 6249 3301 6255 3353
rect 6063 3288 6070 3301
rect 6104 3288 6142 3301
rect 6176 3288 6214 3301
rect 6248 3288 6255 3301
rect 6063 3236 6069 3288
rect 6121 3236 6133 3288
rect 6185 3236 6197 3288
rect 6249 3236 6255 3288
rect 6063 3223 6070 3236
rect 6104 3223 6142 3236
rect 6176 3223 6214 3236
rect 6248 3223 6255 3236
rect 6063 3171 6069 3223
rect 6121 3171 6133 3223
rect 6185 3171 6197 3223
rect 6249 3171 6255 3223
rect 6063 3158 6070 3171
rect 6104 3158 6142 3171
rect 6176 3158 6214 3171
rect 6248 3158 6255 3171
rect 6063 3106 6069 3158
rect 6121 3106 6133 3158
rect 6185 3106 6197 3158
rect 6249 3106 6255 3158
rect 6063 3100 6255 3106
rect 6063 3093 6070 3100
rect 6104 3093 6142 3100
rect 6176 3093 6214 3100
rect 6248 3093 6255 3100
rect 6063 3041 6069 3093
rect 6121 3041 6133 3093
rect 6185 3041 6197 3093
rect 6249 3041 6255 3093
rect 6063 3028 6255 3041
rect 6063 2976 6069 3028
rect 6121 2976 6133 3028
rect 6185 2976 6197 3028
rect 6249 2976 6255 3028
rect 6063 2963 6255 2976
rect 6063 2911 6069 2963
rect 6121 2911 6133 2963
rect 6185 2911 6197 2963
rect 6249 2911 6255 2963
rect 6063 2898 6255 2911
rect 6063 2846 6069 2898
rect 6121 2846 6133 2898
rect 6185 2846 6197 2898
rect 6249 2846 6255 2898
rect 6063 2844 6070 2846
rect 6104 2844 6142 2846
rect 6176 2844 6214 2846
rect 6248 2844 6255 2846
rect 6063 2833 6255 2844
rect 6063 2781 6069 2833
rect 6121 2781 6133 2833
rect 6185 2781 6197 2833
rect 6249 2781 6255 2833
rect 6063 2770 6070 2781
rect 6104 2770 6142 2781
rect 6176 2770 6214 2781
rect 6248 2770 6255 2781
rect 6063 2768 6255 2770
rect 6063 2716 6069 2768
rect 6121 2716 6133 2768
rect 6185 2716 6197 2768
rect 6249 2716 6255 2768
rect 6063 2703 6070 2716
rect 6104 2703 6142 2716
rect 6176 2703 6214 2716
rect 6248 2703 6255 2716
rect 6063 2651 6069 2703
rect 6121 2651 6133 2703
rect 6185 2651 6197 2703
rect 6249 2651 6255 2703
rect 6063 2638 6070 2651
rect 6104 2638 6142 2651
rect 6176 2638 6214 2651
rect 6248 2638 6255 2651
rect 6063 2586 6069 2638
rect 6121 2586 6133 2638
rect 6185 2586 6197 2638
rect 6249 2586 6255 2638
rect 6063 2582 6255 2586
rect 6063 2573 6070 2582
rect 6104 2573 6142 2582
rect 6176 2573 6214 2582
rect 6248 2573 6255 2582
rect 6063 2521 6069 2573
rect 6121 2521 6133 2573
rect 6185 2521 6197 2573
rect 6249 2521 6255 2573
rect 6063 2508 6255 2521
rect 6063 2456 6069 2508
rect 6121 2456 6133 2508
rect 6185 2456 6197 2508
rect 6249 2456 6255 2508
rect 6063 2443 6255 2456
rect 6063 2391 6069 2443
rect 6121 2391 6133 2443
rect 6185 2391 6197 2443
rect 6249 2391 6255 2443
rect 6063 2378 6255 2391
rect 6063 2326 6069 2378
rect 6121 2326 6133 2378
rect 6185 2326 6197 2378
rect 6249 2326 6255 2378
rect 6063 2313 6255 2326
rect 6063 2261 6069 2313
rect 6121 2261 6133 2313
rect 6185 2261 6197 2313
rect 6249 2261 6255 2313
rect 6063 2252 6070 2261
rect 6104 2252 6142 2261
rect 6176 2252 6214 2261
rect 6248 2252 6255 2261
rect 6063 2248 6255 2252
rect 6063 2196 6069 2248
rect 6121 2196 6133 2248
rect 6185 2196 6197 2248
rect 6249 2196 6255 2248
rect 6063 2183 6070 2196
rect 6104 2183 6142 2196
rect 6176 2183 6214 2196
rect 6248 2183 6255 2196
rect 6063 2131 6069 2183
rect 6121 2131 6133 2183
rect 6185 2131 6197 2183
rect 6249 2131 6255 2183
rect 6063 2118 6070 2131
rect 6104 2118 6142 2131
rect 6176 2118 6214 2131
rect 6248 2118 6255 2131
rect 6063 2066 6069 2118
rect 6121 2066 6133 2118
rect 6185 2066 6197 2118
rect 6249 2066 6255 2118
rect 6063 2064 6255 2066
rect 6063 2053 6070 2064
rect 6104 2053 6142 2064
rect 6176 2053 6214 2064
rect 6248 2053 6255 2064
rect 6063 2001 6069 2053
rect 6121 2001 6133 2053
rect 6185 2001 6197 2053
rect 6249 2001 6255 2053
rect 6063 1990 6255 2001
rect 6063 1987 6070 1990
rect 6104 1987 6142 1990
rect 6176 1987 6214 1990
rect 6248 1987 6255 1990
rect 6063 1935 6069 1987
rect 6121 1935 6133 1987
rect 6185 1935 6197 1987
rect 6249 1935 6255 1987
rect 6063 1921 6255 1935
rect 6063 1869 6069 1921
rect 6121 1869 6133 1921
rect 6185 1869 6197 1921
rect 6249 1869 6255 1921
rect 6063 1855 6255 1869
rect 6063 1803 6069 1855
rect 6121 1803 6133 1855
rect 6185 1803 6197 1855
rect 6249 1803 6255 1855
rect 6063 1789 6255 1803
rect 6063 1737 6069 1789
rect 6121 1737 6133 1789
rect 6185 1737 6197 1789
rect 6249 1737 6255 1789
rect 6063 1734 6070 1737
rect 6104 1734 6142 1737
rect 6176 1734 6214 1737
rect 6248 1734 6255 1737
rect 6063 1723 6255 1734
rect 6063 1671 6069 1723
rect 6121 1671 6133 1723
rect 6185 1671 6197 1723
rect 6249 1671 6255 1723
rect 6063 1660 6070 1671
rect 6104 1660 6142 1671
rect 6176 1660 6214 1671
rect 6248 1660 6255 1671
rect 6063 1657 6255 1660
rect 6063 1605 6069 1657
rect 6121 1605 6133 1657
rect 6185 1605 6197 1657
rect 6249 1605 6255 1657
rect 6063 1591 6070 1605
rect 6104 1591 6142 1605
rect 6176 1591 6214 1605
rect 6248 1591 6255 1605
rect 6063 1539 6069 1591
rect 6121 1539 6133 1591
rect 6185 1539 6197 1591
rect 6249 1539 6255 1591
rect 6063 1525 6070 1539
rect 6104 1525 6142 1539
rect 6176 1525 6214 1539
rect 6248 1525 6255 1539
rect 6063 1473 6069 1525
rect 6121 1473 6133 1525
rect 6185 1473 6197 1525
rect 6249 1473 6255 1525
rect 6063 1467 6255 1473
rect 6559 4068 6751 4074
rect 6559 4016 6565 4068
rect 6617 4050 6629 4068
rect 6681 4050 6693 4068
rect 6745 4016 6751 4068
rect 6559 4003 6566 4016
rect 6744 4003 6751 4016
rect 6559 3951 6565 4003
rect 6745 3951 6751 4003
rect 6559 3938 6566 3951
rect 6744 3938 6751 3951
rect 6559 3886 6565 3938
rect 6745 3886 6751 3938
rect 6559 3873 6566 3886
rect 6744 3873 6751 3886
rect 6559 3821 6565 3873
rect 6745 3821 6751 3873
rect 6559 3808 6566 3821
rect 6744 3808 6751 3821
rect 6559 3756 6565 3808
rect 6745 3756 6751 3808
rect 6559 3743 6566 3756
rect 6744 3743 6751 3756
rect 6559 3691 6565 3743
rect 6745 3691 6751 3743
rect 6559 3678 6566 3691
rect 6744 3678 6751 3691
rect 6559 3626 6565 3678
rect 6745 3626 6751 3678
rect 6559 3613 6566 3626
rect 6744 3613 6751 3626
rect 6559 3561 6565 3613
rect 6745 3561 6751 3613
rect 6559 3548 6566 3561
rect 6744 3548 6751 3561
rect 6559 3496 6565 3548
rect 6745 3496 6751 3548
rect 6559 3483 6566 3496
rect 6744 3483 6751 3496
rect 6559 3431 6565 3483
rect 6745 3431 6751 3483
rect 6559 3418 6566 3431
rect 6744 3418 6751 3431
rect 6559 3366 6565 3418
rect 6745 3366 6751 3418
rect 6559 3353 6566 3366
rect 6744 3353 6751 3366
rect 6559 3301 6565 3353
rect 6745 3301 6751 3353
rect 6559 3288 6566 3301
rect 6744 3288 6751 3301
rect 6559 3236 6565 3288
rect 6745 3236 6751 3288
rect 6559 3223 6566 3236
rect 6744 3223 6751 3236
rect 6559 3171 6565 3223
rect 6745 3171 6751 3223
rect 6559 3158 6566 3171
rect 6744 3158 6751 3171
rect 6559 3106 6565 3158
rect 6745 3106 6751 3158
rect 6559 3093 6566 3106
rect 6744 3093 6751 3106
rect 6559 3041 6565 3093
rect 6617 3041 6629 3092
rect 6681 3041 6693 3092
rect 6745 3041 6751 3093
rect 6559 3040 6751 3041
rect 6559 3028 6566 3040
rect 6744 3028 6751 3040
rect 6559 2976 6565 3028
rect 6745 2976 6751 3028
rect 6559 2963 6566 2976
rect 6744 2963 6751 2976
rect 6559 2911 6565 2963
rect 6745 2911 6751 2963
rect 6559 2898 6566 2911
rect 6744 2898 6751 2911
rect 6559 2846 6565 2898
rect 6745 2846 6751 2898
rect 6559 2833 6566 2846
rect 6744 2833 6751 2846
rect 6559 2781 6565 2833
rect 6745 2781 6751 2833
rect 6559 2768 6566 2781
rect 6744 2768 6751 2781
rect 6559 2716 6565 2768
rect 6745 2716 6751 2768
rect 6559 2703 6566 2716
rect 6744 2703 6751 2716
rect 6559 2651 6565 2703
rect 6745 2651 6751 2703
rect 6559 2638 6566 2651
rect 6744 2638 6751 2651
rect 6559 2586 6565 2638
rect 6745 2586 6751 2638
rect 6559 2574 6566 2586
rect 6744 2574 6751 2586
rect 6559 2573 6751 2574
rect 6559 2521 6565 2573
rect 6617 2521 6629 2573
rect 6681 2521 6693 2573
rect 6745 2521 6751 2573
rect 6559 2508 6566 2521
rect 6600 2508 6638 2521
rect 6672 2508 6710 2521
rect 6744 2508 6751 2521
rect 6559 2456 6565 2508
rect 6617 2456 6629 2508
rect 6681 2456 6693 2508
rect 6745 2456 6751 2508
rect 6559 2449 6638 2456
rect 6672 2449 6751 2456
rect 6559 2443 6566 2449
rect 6744 2443 6751 2449
rect 6559 2391 6565 2443
rect 6745 2391 6751 2443
rect 6559 2378 6566 2391
rect 6744 2378 6751 2391
rect 6559 2326 6565 2378
rect 6745 2326 6751 2378
rect 6559 2313 6566 2326
rect 6744 2313 6751 2326
rect 6559 2261 6565 2313
rect 6745 2261 6751 2313
rect 6559 2248 6566 2261
rect 6744 2248 6751 2261
rect 6559 2196 6565 2248
rect 6745 2196 6751 2248
rect 6559 2183 6566 2196
rect 6744 2183 6751 2196
rect 6559 2131 6565 2183
rect 6745 2131 6751 2183
rect 6559 2118 6566 2131
rect 6744 2118 6751 2131
rect 6559 2066 6565 2118
rect 6745 2066 6751 2118
rect 6559 2053 6566 2066
rect 6744 2053 6751 2066
rect 6559 2001 6565 2053
rect 6745 2001 6751 2053
rect 6559 1987 6566 2001
rect 6744 1987 6751 2001
rect 6559 1935 6565 1987
rect 6745 1935 6751 1987
rect 6559 1921 6566 1935
rect 6744 1921 6751 1935
rect 6559 1869 6565 1921
rect 6745 1869 6751 1921
rect 6559 1855 6566 1869
rect 6744 1855 6751 1869
rect 6559 1803 6565 1855
rect 6745 1803 6751 1855
rect 6559 1789 6566 1803
rect 6744 1789 6751 1803
rect 6559 1737 6565 1789
rect 6745 1737 6751 1789
rect 6559 1723 6566 1737
rect 6744 1723 6751 1737
rect 6559 1671 6565 1723
rect 6745 1671 6751 1723
rect 6559 1657 6566 1671
rect 6744 1657 6751 1671
rect 6559 1605 6565 1657
rect 6745 1605 6751 1657
rect 6559 1591 6566 1605
rect 6744 1591 6751 1605
rect 6559 1539 6565 1591
rect 6745 1539 6751 1591
rect 6559 1525 6566 1539
rect 6744 1525 6751 1539
rect 6559 1473 6565 1525
rect 6617 1473 6629 1491
rect 6681 1473 6693 1491
rect 6745 1473 6751 1525
rect 6559 1467 6751 1473
rect 7055 4068 7247 4074
rect 7055 4016 7061 4068
rect 7113 4016 7125 4068
rect 7177 4016 7189 4068
rect 7241 4016 7247 4068
rect 7055 4003 7247 4016
rect 7055 3951 7061 4003
rect 7113 3951 7125 4003
rect 7177 3951 7189 4003
rect 7241 3951 7247 4003
rect 7055 3938 7247 3951
rect 7055 3886 7061 3938
rect 7113 3886 7125 3938
rect 7177 3886 7189 3938
rect 7241 3886 7247 3938
rect 7055 3880 7062 3886
rect 7096 3880 7134 3886
rect 7168 3880 7206 3886
rect 7240 3880 7247 3886
rect 7055 3873 7247 3880
rect 7055 3821 7061 3873
rect 7113 3821 7125 3873
rect 7177 3821 7189 3873
rect 7241 3821 7247 3873
rect 7055 3808 7062 3821
rect 7096 3808 7134 3821
rect 7168 3808 7206 3821
rect 7240 3808 7247 3821
rect 7055 3756 7061 3808
rect 7113 3756 7125 3808
rect 7177 3756 7189 3808
rect 7241 3756 7247 3808
rect 7055 3743 7062 3756
rect 7096 3743 7134 3756
rect 7168 3743 7206 3756
rect 7240 3743 7247 3756
rect 7055 3691 7061 3743
rect 7113 3691 7125 3743
rect 7177 3691 7189 3743
rect 7241 3691 7247 3743
rect 7055 3678 7062 3691
rect 7096 3678 7134 3691
rect 7168 3678 7206 3691
rect 7240 3678 7247 3691
rect 7055 3626 7061 3678
rect 7113 3626 7125 3678
rect 7177 3626 7189 3678
rect 7241 3626 7247 3678
rect 7055 3618 7247 3626
rect 7055 3613 7062 3618
rect 7096 3613 7134 3618
rect 7168 3613 7206 3618
rect 7240 3613 7247 3618
rect 7055 3561 7061 3613
rect 7113 3561 7125 3613
rect 7177 3561 7189 3613
rect 7241 3561 7247 3613
rect 7055 3548 7247 3561
rect 7055 3496 7061 3548
rect 7113 3496 7125 3548
rect 7177 3496 7189 3548
rect 7241 3496 7247 3548
rect 7055 3483 7247 3496
rect 7055 3431 7061 3483
rect 7113 3431 7125 3483
rect 7177 3431 7189 3483
rect 7241 3431 7247 3483
rect 7055 3418 7247 3431
rect 7055 3366 7061 3418
rect 7113 3366 7125 3418
rect 7177 3366 7189 3418
rect 7241 3366 7247 3418
rect 7055 3362 7062 3366
rect 7096 3362 7134 3366
rect 7168 3362 7206 3366
rect 7240 3362 7247 3366
rect 7055 3353 7247 3362
rect 7055 3301 7061 3353
rect 7113 3301 7125 3353
rect 7177 3301 7189 3353
rect 7241 3301 7247 3353
rect 7055 3288 7062 3301
rect 7096 3288 7134 3301
rect 7168 3288 7206 3301
rect 7240 3288 7247 3301
rect 7055 3236 7061 3288
rect 7113 3236 7125 3288
rect 7177 3236 7189 3288
rect 7241 3236 7247 3288
rect 7055 3223 7062 3236
rect 7096 3223 7134 3236
rect 7168 3223 7206 3236
rect 7240 3223 7247 3236
rect 7055 3171 7061 3223
rect 7113 3171 7125 3223
rect 7177 3171 7189 3223
rect 7241 3171 7247 3223
rect 7055 3158 7062 3171
rect 7096 3158 7134 3171
rect 7168 3158 7206 3171
rect 7240 3158 7247 3171
rect 7055 3106 7061 3158
rect 7113 3106 7125 3158
rect 7177 3106 7189 3158
rect 7241 3106 7247 3158
rect 7055 3100 7247 3106
rect 7055 3093 7062 3100
rect 7096 3093 7134 3100
rect 7168 3093 7206 3100
rect 7240 3093 7247 3100
rect 7055 3041 7061 3093
rect 7113 3041 7125 3093
rect 7177 3041 7189 3093
rect 7241 3041 7247 3093
rect 7055 3028 7247 3041
rect 7055 2976 7061 3028
rect 7113 2976 7125 3028
rect 7177 2976 7189 3028
rect 7241 2976 7247 3028
rect 7055 2963 7247 2976
rect 7055 2911 7061 2963
rect 7113 2911 7125 2963
rect 7177 2911 7189 2963
rect 7241 2911 7247 2963
rect 7055 2898 7247 2911
rect 7055 2846 7061 2898
rect 7113 2846 7125 2898
rect 7177 2846 7189 2898
rect 7241 2846 7247 2898
rect 7055 2844 7062 2846
rect 7096 2844 7134 2846
rect 7168 2844 7206 2846
rect 7240 2844 7247 2846
rect 7055 2833 7247 2844
rect 7055 2781 7061 2833
rect 7113 2781 7125 2833
rect 7177 2781 7189 2833
rect 7241 2781 7247 2833
rect 7055 2770 7062 2781
rect 7096 2770 7134 2781
rect 7168 2770 7206 2781
rect 7240 2770 7247 2781
rect 7055 2768 7247 2770
rect 7055 2716 7061 2768
rect 7113 2716 7125 2768
rect 7177 2716 7189 2768
rect 7241 2716 7247 2768
rect 7055 2703 7062 2716
rect 7096 2703 7134 2716
rect 7168 2703 7206 2716
rect 7240 2703 7247 2716
rect 7055 2651 7061 2703
rect 7113 2651 7125 2703
rect 7177 2651 7189 2703
rect 7241 2651 7247 2703
rect 7055 2638 7062 2651
rect 7096 2638 7134 2651
rect 7168 2638 7206 2651
rect 7240 2638 7247 2651
rect 7055 2586 7061 2638
rect 7113 2586 7125 2638
rect 7177 2586 7189 2638
rect 7241 2586 7247 2638
rect 7055 2582 7247 2586
rect 7055 2573 7062 2582
rect 7096 2573 7134 2582
rect 7168 2573 7206 2582
rect 7240 2573 7247 2582
rect 7055 2521 7061 2573
rect 7113 2521 7125 2573
rect 7177 2521 7189 2573
rect 7241 2521 7247 2573
rect 7055 2508 7247 2521
rect 7055 2456 7061 2508
rect 7113 2456 7125 2508
rect 7177 2456 7189 2508
rect 7241 2456 7247 2508
rect 7055 2443 7247 2456
rect 7055 2391 7061 2443
rect 7113 2391 7125 2443
rect 7177 2391 7189 2443
rect 7241 2391 7247 2443
rect 7055 2378 7247 2391
rect 7055 2326 7061 2378
rect 7113 2326 7125 2378
rect 7177 2326 7189 2378
rect 7241 2326 7247 2378
rect 7055 2313 7247 2326
rect 7055 2261 7061 2313
rect 7113 2261 7125 2313
rect 7177 2261 7189 2313
rect 7241 2261 7247 2313
rect 7055 2252 7062 2261
rect 7096 2252 7134 2261
rect 7168 2252 7206 2261
rect 7240 2252 7247 2261
rect 7055 2248 7247 2252
rect 7055 2196 7061 2248
rect 7113 2196 7125 2248
rect 7177 2196 7189 2248
rect 7241 2196 7247 2248
rect 7055 2183 7062 2196
rect 7096 2183 7134 2196
rect 7168 2183 7206 2196
rect 7240 2183 7247 2196
rect 7055 2131 7061 2183
rect 7113 2131 7125 2183
rect 7177 2131 7189 2183
rect 7241 2131 7247 2183
rect 7055 2118 7062 2131
rect 7096 2118 7134 2131
rect 7168 2118 7206 2131
rect 7240 2118 7247 2131
rect 7055 2066 7061 2118
rect 7113 2066 7125 2118
rect 7177 2066 7189 2118
rect 7241 2066 7247 2118
rect 7055 2064 7247 2066
rect 7055 2053 7062 2064
rect 7096 2053 7134 2064
rect 7168 2053 7206 2064
rect 7240 2053 7247 2064
rect 7055 2001 7061 2053
rect 7113 2001 7125 2053
rect 7177 2001 7189 2053
rect 7241 2001 7247 2053
rect 7055 1990 7247 2001
rect 7055 1987 7062 1990
rect 7096 1987 7134 1990
rect 7168 1987 7206 1990
rect 7240 1987 7247 1990
rect 7055 1935 7061 1987
rect 7113 1935 7125 1987
rect 7177 1935 7189 1987
rect 7241 1935 7247 1987
rect 7055 1921 7247 1935
rect 7055 1869 7061 1921
rect 7113 1869 7125 1921
rect 7177 1869 7189 1921
rect 7241 1869 7247 1921
rect 7055 1855 7247 1869
rect 7055 1803 7061 1855
rect 7113 1803 7125 1855
rect 7177 1803 7189 1855
rect 7241 1803 7247 1855
rect 7055 1789 7247 1803
rect 7055 1737 7061 1789
rect 7113 1737 7125 1789
rect 7177 1737 7189 1789
rect 7241 1737 7247 1789
rect 7055 1734 7062 1737
rect 7096 1734 7134 1737
rect 7168 1734 7206 1737
rect 7240 1734 7247 1737
rect 7055 1723 7247 1734
rect 7055 1671 7061 1723
rect 7113 1671 7125 1723
rect 7177 1671 7189 1723
rect 7241 1671 7247 1723
rect 7055 1660 7062 1671
rect 7096 1660 7134 1671
rect 7168 1660 7206 1671
rect 7240 1660 7247 1671
rect 7055 1657 7247 1660
rect 7055 1605 7061 1657
rect 7113 1605 7125 1657
rect 7177 1605 7189 1657
rect 7241 1605 7247 1657
rect 7055 1591 7062 1605
rect 7096 1591 7134 1605
rect 7168 1591 7206 1605
rect 7240 1591 7247 1605
rect 7055 1539 7061 1591
rect 7113 1539 7125 1591
rect 7177 1539 7189 1591
rect 7241 1539 7247 1591
rect 7055 1525 7062 1539
rect 7096 1525 7134 1539
rect 7168 1525 7206 1539
rect 7240 1525 7247 1539
rect 7055 1473 7061 1525
rect 7113 1473 7125 1525
rect 7177 1473 7189 1525
rect 7241 1473 7247 1525
rect 7055 1467 7247 1473
rect 7551 4068 7743 4074
rect 7551 4016 7557 4068
rect 7609 4050 7621 4068
rect 7673 4050 7685 4068
rect 7737 4016 7743 4068
rect 7551 4003 7558 4016
rect 7736 4003 7743 4016
rect 7551 3951 7557 4003
rect 7737 3951 7743 4003
rect 7551 3938 7558 3951
rect 7736 3938 7743 3951
rect 7551 3886 7557 3938
rect 7737 3886 7743 3938
rect 7551 3873 7558 3886
rect 7736 3873 7743 3886
rect 7551 3821 7557 3873
rect 7737 3821 7743 3873
rect 7551 3808 7558 3821
rect 7736 3808 7743 3821
rect 7551 3756 7557 3808
rect 7737 3756 7743 3808
rect 7551 3743 7558 3756
rect 7736 3743 7743 3756
rect 7551 3691 7557 3743
rect 7737 3691 7743 3743
rect 7551 3678 7558 3691
rect 7736 3678 7743 3691
rect 7551 3626 7557 3678
rect 7737 3626 7743 3678
rect 7551 3613 7558 3626
rect 7736 3613 7743 3626
rect 7551 3561 7557 3613
rect 7737 3561 7743 3613
rect 7551 3548 7558 3561
rect 7736 3548 7743 3561
rect 7551 3496 7557 3548
rect 7737 3496 7743 3548
rect 7551 3483 7558 3496
rect 7736 3483 7743 3496
rect 7551 3431 7557 3483
rect 7737 3431 7743 3483
rect 7551 3418 7558 3431
rect 7736 3418 7743 3431
rect 7551 3366 7557 3418
rect 7737 3366 7743 3418
rect 7551 3353 7558 3366
rect 7736 3353 7743 3366
rect 7551 3301 7557 3353
rect 7737 3301 7743 3353
rect 7551 3288 7558 3301
rect 7736 3288 7743 3301
rect 7551 3236 7557 3288
rect 7737 3236 7743 3288
rect 7551 3223 7558 3236
rect 7736 3223 7743 3236
rect 7551 3171 7557 3223
rect 7737 3171 7743 3223
rect 7551 3158 7558 3171
rect 7736 3158 7743 3171
rect 7551 3106 7557 3158
rect 7737 3106 7743 3158
rect 7551 3093 7558 3106
rect 7736 3093 7743 3106
rect 7551 3041 7557 3093
rect 7609 3041 7621 3092
rect 7673 3041 7685 3092
rect 7737 3041 7743 3093
rect 7551 3040 7743 3041
rect 7551 3028 7558 3040
rect 7736 3028 7743 3040
rect 7551 2976 7557 3028
rect 7737 2976 7743 3028
rect 7551 2963 7558 2976
rect 7736 2963 7743 2976
rect 7551 2911 7557 2963
rect 7737 2911 7743 2963
rect 7551 2898 7558 2911
rect 7736 2898 7743 2911
rect 7551 2846 7557 2898
rect 7737 2846 7743 2898
rect 7551 2833 7558 2846
rect 7736 2833 7743 2846
rect 7551 2781 7557 2833
rect 7737 2781 7743 2833
rect 7551 2768 7558 2781
rect 7736 2768 7743 2781
rect 7551 2716 7557 2768
rect 7737 2716 7743 2768
rect 7551 2703 7558 2716
rect 7736 2703 7743 2716
rect 7551 2651 7557 2703
rect 7737 2651 7743 2703
rect 7551 2638 7558 2651
rect 7736 2638 7743 2651
rect 7551 2586 7557 2638
rect 7737 2586 7743 2638
rect 7551 2574 7558 2586
rect 7736 2574 7743 2586
rect 7551 2573 7743 2574
rect 7551 2521 7557 2573
rect 7609 2521 7621 2573
rect 7673 2521 7685 2573
rect 7737 2521 7743 2573
rect 7551 2508 7558 2521
rect 7592 2508 7630 2521
rect 7664 2508 7702 2521
rect 7736 2508 7743 2521
rect 7551 2456 7557 2508
rect 7609 2456 7621 2508
rect 7673 2456 7685 2508
rect 7737 2456 7743 2508
rect 7551 2449 7630 2456
rect 7664 2449 7743 2456
rect 7551 2443 7558 2449
rect 7736 2443 7743 2449
rect 7551 2391 7557 2443
rect 7737 2391 7743 2443
rect 7551 2378 7558 2391
rect 7736 2378 7743 2391
rect 7551 2326 7557 2378
rect 7737 2326 7743 2378
rect 7551 2313 7558 2326
rect 7736 2313 7743 2326
rect 7551 2261 7557 2313
rect 7737 2261 7743 2313
rect 7551 2248 7558 2261
rect 7736 2248 7743 2261
rect 7551 2196 7557 2248
rect 7737 2196 7743 2248
rect 7551 2183 7558 2196
rect 7736 2183 7743 2196
rect 7551 2131 7557 2183
rect 7737 2131 7743 2183
rect 7551 2118 7558 2131
rect 7736 2118 7743 2131
rect 7551 2066 7557 2118
rect 7737 2066 7743 2118
rect 7551 2053 7558 2066
rect 7736 2053 7743 2066
rect 7551 2001 7557 2053
rect 7737 2001 7743 2053
rect 7551 1987 7558 2001
rect 7736 1987 7743 2001
rect 7551 1935 7557 1987
rect 7737 1935 7743 1987
rect 7551 1921 7558 1935
rect 7736 1921 7743 1935
rect 7551 1869 7557 1921
rect 7737 1869 7743 1921
rect 7551 1855 7558 1869
rect 7736 1855 7743 1869
rect 7551 1803 7557 1855
rect 7737 1803 7743 1855
rect 7551 1789 7558 1803
rect 7736 1789 7743 1803
rect 7551 1737 7557 1789
rect 7737 1737 7743 1789
rect 7551 1723 7558 1737
rect 7736 1723 7743 1737
rect 7551 1671 7557 1723
rect 7737 1671 7743 1723
rect 7551 1657 7558 1671
rect 7736 1657 7743 1671
rect 7551 1605 7557 1657
rect 7737 1605 7743 1657
rect 7551 1591 7558 1605
rect 7736 1591 7743 1605
rect 7551 1539 7557 1591
rect 7737 1539 7743 1591
rect 7551 1525 7558 1539
rect 7736 1525 7743 1539
rect 7551 1473 7557 1525
rect 7609 1473 7621 1491
rect 7673 1473 7685 1491
rect 7737 1473 7743 1525
rect 7551 1467 7743 1473
rect 8047 4068 8239 4074
rect 8047 4016 8053 4068
rect 8105 4016 8117 4068
rect 8169 4016 8181 4068
rect 8233 4016 8239 4068
rect 8047 4003 8239 4016
rect 8047 3951 8053 4003
rect 8105 3951 8117 4003
rect 8169 3951 8181 4003
rect 8233 3951 8239 4003
rect 8047 3938 8239 3951
rect 8047 3886 8053 3938
rect 8105 3886 8117 3938
rect 8169 3886 8181 3938
rect 8233 3886 8239 3938
rect 8047 3880 8054 3886
rect 8088 3880 8126 3886
rect 8160 3880 8198 3886
rect 8232 3880 8239 3886
rect 8047 3873 8239 3880
rect 8047 3821 8053 3873
rect 8105 3821 8117 3873
rect 8169 3821 8181 3873
rect 8233 3821 8239 3873
rect 8047 3808 8054 3821
rect 8088 3808 8126 3821
rect 8160 3808 8198 3821
rect 8232 3808 8239 3821
rect 8047 3756 8053 3808
rect 8105 3756 8117 3808
rect 8169 3756 8181 3808
rect 8233 3756 8239 3808
rect 8047 3743 8054 3756
rect 8088 3743 8126 3756
rect 8160 3743 8198 3756
rect 8232 3743 8239 3756
rect 8047 3691 8053 3743
rect 8105 3691 8117 3743
rect 8169 3691 8181 3743
rect 8233 3691 8239 3743
rect 8047 3678 8054 3691
rect 8088 3678 8126 3691
rect 8160 3678 8198 3691
rect 8232 3678 8239 3691
rect 8047 3626 8053 3678
rect 8105 3626 8117 3678
rect 8169 3626 8181 3678
rect 8233 3626 8239 3678
rect 8047 3618 8239 3626
rect 8047 3613 8054 3618
rect 8088 3613 8126 3618
rect 8160 3613 8198 3618
rect 8232 3613 8239 3618
rect 8047 3561 8053 3613
rect 8105 3561 8117 3613
rect 8169 3561 8181 3613
rect 8233 3561 8239 3613
rect 8047 3548 8239 3561
rect 8047 3496 8053 3548
rect 8105 3496 8117 3548
rect 8169 3496 8181 3548
rect 8233 3496 8239 3548
rect 8047 3483 8239 3496
rect 8047 3431 8053 3483
rect 8105 3431 8117 3483
rect 8169 3431 8181 3483
rect 8233 3431 8239 3483
rect 8047 3418 8239 3431
rect 8047 3366 8053 3418
rect 8105 3366 8117 3418
rect 8169 3366 8181 3418
rect 8233 3366 8239 3418
rect 8047 3362 8054 3366
rect 8088 3362 8126 3366
rect 8160 3362 8198 3366
rect 8232 3362 8239 3366
rect 8047 3353 8239 3362
rect 8047 3301 8053 3353
rect 8105 3301 8117 3353
rect 8169 3301 8181 3353
rect 8233 3301 8239 3353
rect 8047 3288 8054 3301
rect 8088 3288 8126 3301
rect 8160 3288 8198 3301
rect 8232 3288 8239 3301
rect 8047 3236 8053 3288
rect 8105 3236 8117 3288
rect 8169 3236 8181 3288
rect 8233 3236 8239 3288
rect 8047 3223 8054 3236
rect 8088 3223 8126 3236
rect 8160 3223 8198 3236
rect 8232 3223 8239 3236
rect 8047 3171 8053 3223
rect 8105 3171 8117 3223
rect 8169 3171 8181 3223
rect 8233 3171 8239 3223
rect 8047 3158 8054 3171
rect 8088 3158 8126 3171
rect 8160 3158 8198 3171
rect 8232 3158 8239 3171
rect 8047 3106 8053 3158
rect 8105 3106 8117 3158
rect 8169 3106 8181 3158
rect 8233 3106 8239 3158
rect 8047 3100 8239 3106
rect 8047 3093 8054 3100
rect 8088 3093 8126 3100
rect 8160 3093 8198 3100
rect 8232 3093 8239 3100
rect 8047 3041 8053 3093
rect 8105 3041 8117 3093
rect 8169 3041 8181 3093
rect 8233 3041 8239 3093
rect 8047 3028 8239 3041
rect 8047 2976 8053 3028
rect 8105 2976 8117 3028
rect 8169 2976 8181 3028
rect 8233 2976 8239 3028
rect 8047 2963 8239 2976
rect 8047 2911 8053 2963
rect 8105 2911 8117 2963
rect 8169 2911 8181 2963
rect 8233 2911 8239 2963
rect 8047 2898 8239 2911
rect 8047 2846 8053 2898
rect 8105 2846 8117 2898
rect 8169 2846 8181 2898
rect 8233 2846 8239 2898
rect 8047 2844 8054 2846
rect 8088 2844 8126 2846
rect 8160 2844 8198 2846
rect 8232 2844 8239 2846
rect 8047 2833 8239 2844
rect 8047 2781 8053 2833
rect 8105 2781 8117 2833
rect 8169 2781 8181 2833
rect 8233 2781 8239 2833
rect 8047 2770 8054 2781
rect 8088 2770 8126 2781
rect 8160 2770 8198 2781
rect 8232 2770 8239 2781
rect 8047 2768 8239 2770
rect 8047 2716 8053 2768
rect 8105 2716 8117 2768
rect 8169 2716 8181 2768
rect 8233 2716 8239 2768
rect 8047 2703 8054 2716
rect 8088 2703 8126 2716
rect 8160 2703 8198 2716
rect 8232 2703 8239 2716
rect 8047 2651 8053 2703
rect 8105 2651 8117 2703
rect 8169 2651 8181 2703
rect 8233 2651 8239 2703
rect 8047 2638 8054 2651
rect 8088 2638 8126 2651
rect 8160 2638 8198 2651
rect 8232 2638 8239 2651
rect 8047 2586 8053 2638
rect 8105 2586 8117 2638
rect 8169 2586 8181 2638
rect 8233 2586 8239 2638
rect 8047 2582 8239 2586
rect 8047 2573 8054 2582
rect 8088 2573 8126 2582
rect 8160 2573 8198 2582
rect 8232 2573 8239 2582
rect 8047 2521 8053 2573
rect 8105 2521 8117 2573
rect 8169 2521 8181 2573
rect 8233 2521 8239 2573
rect 8047 2508 8239 2521
rect 8047 2456 8053 2508
rect 8105 2456 8117 2508
rect 8169 2456 8181 2508
rect 8233 2456 8239 2508
rect 8047 2443 8239 2456
rect 8047 2391 8053 2443
rect 8105 2391 8117 2443
rect 8169 2391 8181 2443
rect 8233 2391 8239 2443
rect 8047 2378 8239 2391
rect 8047 2326 8053 2378
rect 8105 2326 8117 2378
rect 8169 2326 8181 2378
rect 8233 2326 8239 2378
rect 8047 2313 8239 2326
rect 8047 2261 8053 2313
rect 8105 2261 8117 2313
rect 8169 2261 8181 2313
rect 8233 2261 8239 2313
rect 8047 2252 8054 2261
rect 8088 2252 8126 2261
rect 8160 2252 8198 2261
rect 8232 2252 8239 2261
rect 8047 2248 8239 2252
rect 8047 2196 8053 2248
rect 8105 2196 8117 2248
rect 8169 2196 8181 2248
rect 8233 2196 8239 2248
rect 8047 2183 8054 2196
rect 8088 2183 8126 2196
rect 8160 2183 8198 2196
rect 8232 2183 8239 2196
rect 8047 2131 8053 2183
rect 8105 2131 8117 2183
rect 8169 2131 8181 2183
rect 8233 2131 8239 2183
rect 8047 2118 8054 2131
rect 8088 2118 8126 2131
rect 8160 2118 8198 2131
rect 8232 2118 8239 2131
rect 8047 2066 8053 2118
rect 8105 2066 8117 2118
rect 8169 2066 8181 2118
rect 8233 2066 8239 2118
rect 8047 2064 8239 2066
rect 8047 2053 8054 2064
rect 8088 2053 8126 2064
rect 8160 2053 8198 2064
rect 8232 2053 8239 2064
rect 8047 2001 8053 2053
rect 8105 2001 8117 2053
rect 8169 2001 8181 2053
rect 8233 2001 8239 2053
rect 8047 1990 8239 2001
rect 8047 1987 8054 1990
rect 8088 1987 8126 1990
rect 8160 1987 8198 1990
rect 8232 1987 8239 1990
rect 8047 1935 8053 1987
rect 8105 1935 8117 1987
rect 8169 1935 8181 1987
rect 8233 1935 8239 1987
rect 8047 1921 8239 1935
rect 8047 1869 8053 1921
rect 8105 1869 8117 1921
rect 8169 1869 8181 1921
rect 8233 1869 8239 1921
rect 8047 1855 8239 1869
rect 8047 1803 8053 1855
rect 8105 1803 8117 1855
rect 8169 1803 8181 1855
rect 8233 1803 8239 1855
rect 8047 1789 8239 1803
rect 8047 1737 8053 1789
rect 8105 1737 8117 1789
rect 8169 1737 8181 1789
rect 8233 1737 8239 1789
rect 8047 1734 8054 1737
rect 8088 1734 8126 1737
rect 8160 1734 8198 1737
rect 8232 1734 8239 1737
rect 8047 1723 8239 1734
rect 8047 1671 8053 1723
rect 8105 1671 8117 1723
rect 8169 1671 8181 1723
rect 8233 1671 8239 1723
rect 8047 1660 8054 1671
rect 8088 1660 8126 1671
rect 8160 1660 8198 1671
rect 8232 1660 8239 1671
rect 8047 1657 8239 1660
rect 8047 1605 8053 1657
rect 8105 1605 8117 1657
rect 8169 1605 8181 1657
rect 8233 1605 8239 1657
rect 8047 1591 8054 1605
rect 8088 1591 8126 1605
rect 8160 1591 8198 1605
rect 8232 1591 8239 1605
rect 8047 1539 8053 1591
rect 8105 1539 8117 1591
rect 8169 1539 8181 1591
rect 8233 1539 8239 1591
rect 8047 1525 8054 1539
rect 8088 1525 8126 1539
rect 8160 1525 8198 1539
rect 8232 1525 8239 1539
rect 8047 1473 8053 1525
rect 8105 1473 8117 1525
rect 8169 1473 8181 1525
rect 8233 1473 8239 1525
rect 8047 1467 8239 1473
rect 8543 4068 8735 4074
rect 8543 4016 8549 4068
rect 8601 4050 8613 4068
rect 8665 4050 8677 4068
rect 8729 4016 8735 4068
rect 8543 4003 8550 4016
rect 8728 4003 8735 4016
rect 8543 3951 8549 4003
rect 8729 3951 8735 4003
rect 8543 3938 8550 3951
rect 8728 3938 8735 3951
rect 8543 3886 8549 3938
rect 8729 3886 8735 3938
rect 8543 3873 8550 3886
rect 8728 3873 8735 3886
rect 8543 3821 8549 3873
rect 8729 3821 8735 3873
rect 8543 3808 8550 3821
rect 8728 3808 8735 3821
rect 8543 3756 8549 3808
rect 8729 3756 8735 3808
rect 8543 3743 8550 3756
rect 8728 3743 8735 3756
rect 8543 3691 8549 3743
rect 8729 3691 8735 3743
rect 8543 3678 8550 3691
rect 8728 3678 8735 3691
rect 8543 3626 8549 3678
rect 8729 3626 8735 3678
rect 8543 3613 8550 3626
rect 8728 3613 8735 3626
rect 8543 3561 8549 3613
rect 8729 3561 8735 3613
rect 8543 3548 8550 3561
rect 8728 3548 8735 3561
rect 8543 3496 8549 3548
rect 8729 3496 8735 3548
rect 8543 3483 8550 3496
rect 8728 3483 8735 3496
rect 8543 3431 8549 3483
rect 8729 3431 8735 3483
rect 8543 3418 8550 3431
rect 8728 3418 8735 3431
rect 8543 3366 8549 3418
rect 8729 3366 8735 3418
rect 8543 3353 8550 3366
rect 8728 3353 8735 3366
rect 8543 3301 8549 3353
rect 8729 3301 8735 3353
rect 8543 3288 8550 3301
rect 8728 3288 8735 3301
rect 8543 3236 8549 3288
rect 8729 3236 8735 3288
rect 8543 3223 8550 3236
rect 8728 3223 8735 3236
rect 8543 3171 8549 3223
rect 8729 3171 8735 3223
rect 8543 3158 8550 3171
rect 8728 3158 8735 3171
rect 8543 3106 8549 3158
rect 8729 3106 8735 3158
rect 8543 3093 8550 3106
rect 8728 3093 8735 3106
rect 8543 3041 8549 3093
rect 8601 3041 8613 3092
rect 8665 3041 8677 3092
rect 8729 3041 8735 3093
rect 8543 3040 8735 3041
rect 8543 3028 8550 3040
rect 8728 3028 8735 3040
rect 8543 2976 8549 3028
rect 8729 2976 8735 3028
rect 8543 2963 8550 2976
rect 8728 2963 8735 2976
rect 8543 2911 8549 2963
rect 8729 2911 8735 2963
rect 8543 2898 8550 2911
rect 8728 2898 8735 2911
rect 8543 2846 8549 2898
rect 8729 2846 8735 2898
rect 8543 2833 8550 2846
rect 8728 2833 8735 2846
rect 8543 2781 8549 2833
rect 8729 2781 8735 2833
rect 8543 2768 8550 2781
rect 8728 2768 8735 2781
rect 8543 2716 8549 2768
rect 8729 2716 8735 2768
rect 8543 2703 8550 2716
rect 8728 2703 8735 2716
rect 8543 2651 8549 2703
rect 8729 2651 8735 2703
rect 8543 2638 8550 2651
rect 8728 2638 8735 2651
rect 8543 2586 8549 2638
rect 8729 2586 8735 2638
rect 8543 2574 8550 2586
rect 8728 2574 8735 2586
rect 8543 2573 8735 2574
rect 8543 2521 8549 2573
rect 8601 2521 8613 2573
rect 8665 2521 8677 2573
rect 8729 2521 8735 2573
rect 8543 2508 8550 2521
rect 8584 2508 8622 2521
rect 8656 2508 8694 2521
rect 8728 2508 8735 2521
rect 8543 2456 8549 2508
rect 8601 2456 8613 2508
rect 8665 2456 8677 2508
rect 8729 2456 8735 2508
rect 8543 2449 8622 2456
rect 8656 2449 8735 2456
rect 8543 2443 8550 2449
rect 8728 2443 8735 2449
rect 8543 2391 8549 2443
rect 8729 2391 8735 2443
rect 8543 2378 8550 2391
rect 8728 2378 8735 2391
rect 8543 2326 8549 2378
rect 8729 2326 8735 2378
rect 8543 2313 8550 2326
rect 8728 2313 8735 2326
rect 8543 2261 8549 2313
rect 8729 2261 8735 2313
rect 8543 2248 8550 2261
rect 8728 2248 8735 2261
rect 8543 2196 8549 2248
rect 8729 2196 8735 2248
rect 8543 2183 8550 2196
rect 8728 2183 8735 2196
rect 8543 2131 8549 2183
rect 8729 2131 8735 2183
rect 8543 2118 8550 2131
rect 8728 2118 8735 2131
rect 8543 2066 8549 2118
rect 8729 2066 8735 2118
rect 8543 2053 8550 2066
rect 8728 2053 8735 2066
rect 8543 2001 8549 2053
rect 8729 2001 8735 2053
rect 8543 1987 8550 2001
rect 8728 1987 8735 2001
rect 8543 1935 8549 1987
rect 8729 1935 8735 1987
rect 8543 1921 8550 1935
rect 8728 1921 8735 1935
rect 8543 1869 8549 1921
rect 8729 1869 8735 1921
rect 8543 1855 8550 1869
rect 8728 1855 8735 1869
rect 8543 1803 8549 1855
rect 8729 1803 8735 1855
rect 8543 1789 8550 1803
rect 8728 1789 8735 1803
rect 8543 1737 8549 1789
rect 8729 1737 8735 1789
rect 8543 1723 8550 1737
rect 8728 1723 8735 1737
rect 8543 1671 8549 1723
rect 8729 1671 8735 1723
rect 8543 1657 8550 1671
rect 8728 1657 8735 1671
rect 8543 1605 8549 1657
rect 8729 1605 8735 1657
rect 8543 1591 8550 1605
rect 8728 1591 8735 1605
rect 8543 1539 8549 1591
rect 8729 1539 8735 1591
rect 8543 1525 8550 1539
rect 8728 1525 8735 1539
rect 8543 1473 8549 1525
rect 8601 1473 8613 1491
rect 8665 1473 8677 1491
rect 8729 1473 8735 1525
rect 8543 1467 8735 1473
rect 9039 4068 9231 4074
rect 9039 4016 9045 4068
rect 9097 4016 9109 4068
rect 9161 4016 9173 4068
rect 9225 4016 9231 4068
rect 9039 4003 9231 4016
rect 9039 3951 9045 4003
rect 9097 3951 9109 4003
rect 9161 3951 9173 4003
rect 9225 3951 9231 4003
rect 9039 3938 9231 3951
rect 9039 3886 9045 3938
rect 9097 3886 9109 3938
rect 9161 3886 9173 3938
rect 9225 3886 9231 3938
rect 9039 3880 9046 3886
rect 9080 3880 9118 3886
rect 9152 3880 9190 3886
rect 9224 3880 9231 3886
rect 9039 3873 9231 3880
rect 9039 3821 9045 3873
rect 9097 3821 9109 3873
rect 9161 3821 9173 3873
rect 9225 3821 9231 3873
rect 9039 3808 9046 3821
rect 9080 3808 9118 3821
rect 9152 3808 9190 3821
rect 9224 3808 9231 3821
rect 9039 3756 9045 3808
rect 9097 3756 9109 3808
rect 9161 3756 9173 3808
rect 9225 3756 9231 3808
rect 9039 3743 9046 3756
rect 9080 3743 9118 3756
rect 9152 3743 9190 3756
rect 9224 3743 9231 3756
rect 9039 3691 9045 3743
rect 9097 3691 9109 3743
rect 9161 3691 9173 3743
rect 9225 3691 9231 3743
rect 9039 3678 9046 3691
rect 9080 3678 9118 3691
rect 9152 3678 9190 3691
rect 9224 3678 9231 3691
rect 9039 3626 9045 3678
rect 9097 3626 9109 3678
rect 9161 3626 9173 3678
rect 9225 3626 9231 3678
rect 9039 3618 9231 3626
rect 9039 3613 9046 3618
rect 9080 3613 9118 3618
rect 9152 3613 9190 3618
rect 9224 3613 9231 3618
rect 9039 3561 9045 3613
rect 9097 3561 9109 3613
rect 9161 3561 9173 3613
rect 9225 3561 9231 3613
rect 9039 3548 9231 3561
rect 9039 3496 9045 3548
rect 9097 3496 9109 3548
rect 9161 3496 9173 3548
rect 9225 3496 9231 3548
rect 9039 3483 9231 3496
rect 9039 3431 9045 3483
rect 9097 3431 9109 3483
rect 9161 3431 9173 3483
rect 9225 3431 9231 3483
rect 9039 3418 9231 3431
rect 9039 3366 9045 3418
rect 9097 3366 9109 3418
rect 9161 3366 9173 3418
rect 9225 3366 9231 3418
rect 9039 3362 9046 3366
rect 9080 3362 9118 3366
rect 9152 3362 9190 3366
rect 9224 3362 9231 3366
rect 9039 3353 9231 3362
rect 9039 3301 9045 3353
rect 9097 3301 9109 3353
rect 9161 3301 9173 3353
rect 9225 3301 9231 3353
rect 9039 3288 9046 3301
rect 9080 3288 9118 3301
rect 9152 3288 9190 3301
rect 9224 3288 9231 3301
rect 9039 3236 9045 3288
rect 9097 3236 9109 3288
rect 9161 3236 9173 3288
rect 9225 3236 9231 3288
rect 9039 3223 9046 3236
rect 9080 3223 9118 3236
rect 9152 3223 9190 3236
rect 9224 3223 9231 3236
rect 9039 3171 9045 3223
rect 9097 3171 9109 3223
rect 9161 3171 9173 3223
rect 9225 3171 9231 3223
rect 9039 3158 9046 3171
rect 9080 3158 9118 3171
rect 9152 3158 9190 3171
rect 9224 3158 9231 3171
rect 9039 3106 9045 3158
rect 9097 3106 9109 3158
rect 9161 3106 9173 3158
rect 9225 3106 9231 3158
rect 9039 3100 9231 3106
rect 9039 3093 9046 3100
rect 9080 3093 9118 3100
rect 9152 3093 9190 3100
rect 9224 3093 9231 3100
rect 9039 3041 9045 3093
rect 9097 3041 9109 3093
rect 9161 3041 9173 3093
rect 9225 3041 9231 3093
rect 9039 3028 9231 3041
rect 9039 2976 9045 3028
rect 9097 2976 9109 3028
rect 9161 2976 9173 3028
rect 9225 2976 9231 3028
rect 9039 2963 9231 2976
rect 9039 2911 9045 2963
rect 9097 2911 9109 2963
rect 9161 2911 9173 2963
rect 9225 2911 9231 2963
rect 9039 2898 9231 2911
rect 9039 2846 9045 2898
rect 9097 2846 9109 2898
rect 9161 2846 9173 2898
rect 9225 2846 9231 2898
rect 9039 2844 9046 2846
rect 9080 2844 9118 2846
rect 9152 2844 9190 2846
rect 9224 2844 9231 2846
rect 9039 2833 9231 2844
rect 9039 2781 9045 2833
rect 9097 2781 9109 2833
rect 9161 2781 9173 2833
rect 9225 2781 9231 2833
rect 9039 2770 9046 2781
rect 9080 2770 9118 2781
rect 9152 2770 9190 2781
rect 9224 2770 9231 2781
rect 9039 2768 9231 2770
rect 9039 2716 9045 2768
rect 9097 2716 9109 2768
rect 9161 2716 9173 2768
rect 9225 2716 9231 2768
rect 9039 2703 9046 2716
rect 9080 2703 9118 2716
rect 9152 2703 9190 2716
rect 9224 2703 9231 2716
rect 9039 2651 9045 2703
rect 9097 2651 9109 2703
rect 9161 2651 9173 2703
rect 9225 2651 9231 2703
rect 9039 2638 9046 2651
rect 9080 2638 9118 2651
rect 9152 2638 9190 2651
rect 9224 2638 9231 2651
rect 9039 2586 9045 2638
rect 9097 2586 9109 2638
rect 9161 2586 9173 2638
rect 9225 2586 9231 2638
rect 9039 2582 9231 2586
rect 9039 2573 9046 2582
rect 9080 2573 9118 2582
rect 9152 2573 9190 2582
rect 9224 2573 9231 2582
rect 9039 2521 9045 2573
rect 9097 2521 9109 2573
rect 9161 2521 9173 2573
rect 9225 2521 9231 2573
rect 9039 2508 9231 2521
rect 9039 2456 9045 2508
rect 9097 2456 9109 2508
rect 9161 2456 9173 2508
rect 9225 2456 9231 2508
rect 9039 2443 9231 2456
rect 9039 2391 9045 2443
rect 9097 2391 9109 2443
rect 9161 2391 9173 2443
rect 9225 2391 9231 2443
rect 9039 2378 9231 2391
rect 9039 2326 9045 2378
rect 9097 2326 9109 2378
rect 9161 2326 9173 2378
rect 9225 2326 9231 2378
rect 9039 2313 9231 2326
rect 9039 2261 9045 2313
rect 9097 2261 9109 2313
rect 9161 2261 9173 2313
rect 9225 2261 9231 2313
rect 9039 2252 9046 2261
rect 9080 2252 9118 2261
rect 9152 2252 9190 2261
rect 9224 2252 9231 2261
rect 9039 2248 9231 2252
rect 9039 2196 9045 2248
rect 9097 2196 9109 2248
rect 9161 2196 9173 2248
rect 9225 2196 9231 2248
rect 9039 2183 9046 2196
rect 9080 2183 9118 2196
rect 9152 2183 9190 2196
rect 9224 2183 9231 2196
rect 9039 2131 9045 2183
rect 9097 2131 9109 2183
rect 9161 2131 9173 2183
rect 9225 2131 9231 2183
rect 9039 2118 9046 2131
rect 9080 2118 9118 2131
rect 9152 2118 9190 2131
rect 9224 2118 9231 2131
rect 9039 2066 9045 2118
rect 9097 2066 9109 2118
rect 9161 2066 9173 2118
rect 9225 2066 9231 2118
rect 9039 2064 9231 2066
rect 9039 2053 9046 2064
rect 9080 2053 9118 2064
rect 9152 2053 9190 2064
rect 9224 2053 9231 2064
rect 9039 2001 9045 2053
rect 9097 2001 9109 2053
rect 9161 2001 9173 2053
rect 9225 2001 9231 2053
rect 9039 1990 9231 2001
rect 9039 1987 9046 1990
rect 9080 1987 9118 1990
rect 9152 1987 9190 1990
rect 9224 1987 9231 1990
rect 9039 1935 9045 1987
rect 9097 1935 9109 1987
rect 9161 1935 9173 1987
rect 9225 1935 9231 1987
rect 9039 1921 9231 1935
rect 9039 1869 9045 1921
rect 9097 1869 9109 1921
rect 9161 1869 9173 1921
rect 9225 1869 9231 1921
rect 9039 1855 9231 1869
rect 9039 1803 9045 1855
rect 9097 1803 9109 1855
rect 9161 1803 9173 1855
rect 9225 1803 9231 1855
rect 9039 1789 9231 1803
rect 9039 1737 9045 1789
rect 9097 1737 9109 1789
rect 9161 1737 9173 1789
rect 9225 1737 9231 1789
rect 9039 1734 9046 1737
rect 9080 1734 9118 1737
rect 9152 1734 9190 1737
rect 9224 1734 9231 1737
rect 9039 1723 9231 1734
rect 9039 1671 9045 1723
rect 9097 1671 9109 1723
rect 9161 1671 9173 1723
rect 9225 1671 9231 1723
rect 9039 1660 9046 1671
rect 9080 1660 9118 1671
rect 9152 1660 9190 1671
rect 9224 1660 9231 1671
rect 9039 1657 9231 1660
rect 9039 1605 9045 1657
rect 9097 1605 9109 1657
rect 9161 1605 9173 1657
rect 9225 1605 9231 1657
rect 9039 1591 9046 1605
rect 9080 1591 9118 1605
rect 9152 1591 9190 1605
rect 9224 1591 9231 1605
rect 9039 1539 9045 1591
rect 9097 1539 9109 1591
rect 9161 1539 9173 1591
rect 9225 1539 9231 1591
rect 9039 1525 9046 1539
rect 9080 1525 9118 1539
rect 9152 1525 9190 1539
rect 9224 1525 9231 1539
rect 9039 1473 9045 1525
rect 9097 1473 9109 1525
rect 9161 1473 9173 1525
rect 9225 1473 9231 1525
rect 9039 1467 9231 1473
rect 9535 4068 9727 4074
rect 9535 4016 9541 4068
rect 9593 4050 9605 4068
rect 9657 4050 9669 4068
rect 9721 4016 9727 4068
rect 9535 4003 9542 4016
rect 9720 4003 9727 4016
rect 9535 3951 9541 4003
rect 9721 3951 9727 4003
rect 9535 3938 9542 3951
rect 9720 3938 9727 3951
rect 9535 3886 9541 3938
rect 9721 3886 9727 3938
rect 9535 3873 9542 3886
rect 9720 3873 9727 3886
rect 9535 3821 9541 3873
rect 9721 3821 9727 3873
rect 9535 3808 9542 3821
rect 9720 3808 9727 3821
rect 9535 3756 9541 3808
rect 9721 3756 9727 3808
rect 9535 3743 9542 3756
rect 9720 3743 9727 3756
rect 9535 3691 9541 3743
rect 9721 3691 9727 3743
rect 9535 3678 9542 3691
rect 9720 3678 9727 3691
rect 9535 3626 9541 3678
rect 9721 3626 9727 3678
rect 9535 3613 9542 3626
rect 9720 3613 9727 3626
rect 9535 3561 9541 3613
rect 9721 3561 9727 3613
rect 9535 3548 9542 3561
rect 9720 3548 9727 3561
rect 9535 3496 9541 3548
rect 9721 3496 9727 3548
rect 9535 3483 9542 3496
rect 9720 3483 9727 3496
rect 9535 3431 9541 3483
rect 9721 3431 9727 3483
rect 9535 3418 9542 3431
rect 9720 3418 9727 3431
rect 9535 3366 9541 3418
rect 9721 3366 9727 3418
rect 9535 3353 9542 3366
rect 9720 3353 9727 3366
rect 9535 3301 9541 3353
rect 9721 3301 9727 3353
rect 9535 3288 9542 3301
rect 9720 3288 9727 3301
rect 9535 3236 9541 3288
rect 9721 3236 9727 3288
rect 9535 3223 9542 3236
rect 9720 3223 9727 3236
rect 9535 3171 9541 3223
rect 9721 3171 9727 3223
rect 9535 3158 9542 3171
rect 9720 3158 9727 3171
rect 9535 3106 9541 3158
rect 9721 3106 9727 3158
rect 9535 3093 9542 3106
rect 9720 3093 9727 3106
rect 9535 3041 9541 3093
rect 9593 3041 9605 3092
rect 9657 3041 9669 3092
rect 9721 3041 9727 3093
rect 9535 3040 9727 3041
rect 9535 3028 9542 3040
rect 9720 3028 9727 3040
rect 9535 2976 9541 3028
rect 9721 2976 9727 3028
rect 9535 2963 9542 2976
rect 9720 2963 9727 2976
rect 9535 2911 9541 2963
rect 9721 2911 9727 2963
rect 9535 2898 9542 2911
rect 9720 2898 9727 2911
rect 9535 2846 9541 2898
rect 9721 2846 9727 2898
rect 9535 2833 9542 2846
rect 9720 2833 9727 2846
rect 9535 2781 9541 2833
rect 9721 2781 9727 2833
rect 9535 2768 9542 2781
rect 9720 2768 9727 2781
rect 9535 2716 9541 2768
rect 9721 2716 9727 2768
rect 9535 2703 9542 2716
rect 9720 2703 9727 2716
rect 9535 2651 9541 2703
rect 9721 2651 9727 2703
rect 9535 2638 9542 2651
rect 9720 2638 9727 2651
rect 9535 2586 9541 2638
rect 9721 2586 9727 2638
rect 9535 2574 9542 2586
rect 9720 2574 9727 2586
rect 9535 2573 9727 2574
rect 9535 2521 9541 2573
rect 9593 2521 9605 2573
rect 9657 2521 9669 2573
rect 9721 2521 9727 2573
rect 9535 2508 9542 2521
rect 9576 2508 9614 2521
rect 9648 2508 9686 2521
rect 9720 2508 9727 2521
rect 9535 2456 9541 2508
rect 9593 2456 9605 2508
rect 9657 2456 9669 2508
rect 9721 2456 9727 2508
rect 9535 2449 9614 2456
rect 9648 2449 9727 2456
rect 9535 2443 9542 2449
rect 9720 2443 9727 2449
rect 9535 2391 9541 2443
rect 9721 2391 9727 2443
rect 9535 2378 9542 2391
rect 9720 2378 9727 2391
rect 9535 2326 9541 2378
rect 9721 2326 9727 2378
rect 9535 2313 9542 2326
rect 9720 2313 9727 2326
rect 9535 2261 9541 2313
rect 9721 2261 9727 2313
rect 9535 2248 9542 2261
rect 9720 2248 9727 2261
rect 9535 2196 9541 2248
rect 9721 2196 9727 2248
rect 9535 2183 9542 2196
rect 9720 2183 9727 2196
rect 9535 2131 9541 2183
rect 9721 2131 9727 2183
rect 9535 2118 9542 2131
rect 9720 2118 9727 2131
rect 9535 2066 9541 2118
rect 9721 2066 9727 2118
rect 9535 2053 9542 2066
rect 9720 2053 9727 2066
rect 9535 2001 9541 2053
rect 9721 2001 9727 2053
rect 9535 1987 9542 2001
rect 9720 1987 9727 2001
rect 9535 1935 9541 1987
rect 9721 1935 9727 1987
rect 9535 1921 9542 1935
rect 9720 1921 9727 1935
rect 9535 1869 9541 1921
rect 9721 1869 9727 1921
rect 9535 1855 9542 1869
rect 9720 1855 9727 1869
rect 9535 1803 9541 1855
rect 9721 1803 9727 1855
rect 9535 1789 9542 1803
rect 9720 1789 9727 1803
rect 9535 1737 9541 1789
rect 9721 1737 9727 1789
rect 9535 1723 9542 1737
rect 9720 1723 9727 1737
rect 9535 1671 9541 1723
rect 9721 1671 9727 1723
rect 9535 1657 9542 1671
rect 9720 1657 9727 1671
rect 9535 1605 9541 1657
rect 9721 1605 9727 1657
rect 9535 1591 9542 1605
rect 9720 1591 9727 1605
rect 9535 1539 9541 1591
rect 9721 1539 9727 1591
rect 9535 1525 9542 1539
rect 9720 1525 9727 1539
rect 9535 1473 9541 1525
rect 9593 1473 9605 1491
rect 9657 1473 9669 1491
rect 9721 1473 9727 1525
rect 9535 1467 9727 1473
rect 10031 4068 10223 4074
rect 10031 4016 10037 4068
rect 10089 4016 10101 4068
rect 10153 4016 10165 4068
rect 10217 4016 10223 4068
rect 10031 4003 10223 4016
rect 10031 3951 10037 4003
rect 10089 3951 10101 4003
rect 10153 3951 10165 4003
rect 10217 3951 10223 4003
rect 10031 3938 10223 3951
rect 10031 3886 10037 3938
rect 10089 3886 10101 3938
rect 10153 3886 10165 3938
rect 10217 3886 10223 3938
rect 10031 3880 10038 3886
rect 10072 3880 10110 3886
rect 10144 3880 10182 3886
rect 10216 3880 10223 3886
rect 10031 3873 10223 3880
rect 10031 3821 10037 3873
rect 10089 3821 10101 3873
rect 10153 3821 10165 3873
rect 10217 3821 10223 3873
rect 10031 3808 10038 3821
rect 10072 3808 10110 3821
rect 10144 3808 10182 3821
rect 10216 3808 10223 3821
rect 10031 3756 10037 3808
rect 10089 3756 10101 3808
rect 10153 3756 10165 3808
rect 10217 3756 10223 3808
rect 10031 3743 10038 3756
rect 10072 3743 10110 3756
rect 10144 3743 10182 3756
rect 10216 3743 10223 3756
rect 10031 3691 10037 3743
rect 10089 3691 10101 3743
rect 10153 3691 10165 3743
rect 10217 3691 10223 3743
rect 10031 3678 10038 3691
rect 10072 3678 10110 3691
rect 10144 3678 10182 3691
rect 10216 3678 10223 3691
rect 10031 3626 10037 3678
rect 10089 3626 10101 3678
rect 10153 3626 10165 3678
rect 10217 3626 10223 3678
rect 10031 3618 10223 3626
rect 10031 3613 10038 3618
rect 10072 3613 10110 3618
rect 10144 3613 10182 3618
rect 10216 3613 10223 3618
rect 10031 3561 10037 3613
rect 10089 3561 10101 3613
rect 10153 3561 10165 3613
rect 10217 3561 10223 3613
rect 10031 3548 10223 3561
rect 10031 3496 10037 3548
rect 10089 3496 10101 3548
rect 10153 3496 10165 3548
rect 10217 3496 10223 3548
rect 10031 3483 10223 3496
rect 10031 3431 10037 3483
rect 10089 3431 10101 3483
rect 10153 3431 10165 3483
rect 10217 3431 10223 3483
rect 10031 3418 10223 3431
rect 10031 3366 10037 3418
rect 10089 3366 10101 3418
rect 10153 3366 10165 3418
rect 10217 3366 10223 3418
rect 10031 3362 10038 3366
rect 10072 3362 10110 3366
rect 10144 3362 10182 3366
rect 10216 3362 10223 3366
rect 10031 3353 10223 3362
rect 10031 3301 10037 3353
rect 10089 3301 10101 3353
rect 10153 3301 10165 3353
rect 10217 3301 10223 3353
rect 10031 3288 10038 3301
rect 10072 3288 10110 3301
rect 10144 3288 10182 3301
rect 10216 3288 10223 3301
rect 10031 3236 10037 3288
rect 10089 3236 10101 3288
rect 10153 3236 10165 3288
rect 10217 3236 10223 3288
rect 10031 3223 10038 3236
rect 10072 3223 10110 3236
rect 10144 3223 10182 3236
rect 10216 3223 10223 3236
rect 10031 3171 10037 3223
rect 10089 3171 10101 3223
rect 10153 3171 10165 3223
rect 10217 3171 10223 3223
rect 10031 3158 10038 3171
rect 10072 3158 10110 3171
rect 10144 3158 10182 3171
rect 10216 3158 10223 3171
rect 10031 3106 10037 3158
rect 10089 3106 10101 3158
rect 10153 3106 10165 3158
rect 10217 3106 10223 3158
rect 10031 3100 10223 3106
rect 10031 3093 10038 3100
rect 10072 3093 10110 3100
rect 10144 3093 10182 3100
rect 10216 3093 10223 3100
rect 10031 3041 10037 3093
rect 10089 3041 10101 3093
rect 10153 3041 10165 3093
rect 10217 3041 10223 3093
rect 10031 3028 10223 3041
rect 10031 2976 10037 3028
rect 10089 2976 10101 3028
rect 10153 2976 10165 3028
rect 10217 2976 10223 3028
rect 10031 2963 10223 2976
rect 10031 2911 10037 2963
rect 10089 2911 10101 2963
rect 10153 2911 10165 2963
rect 10217 2911 10223 2963
rect 10031 2898 10223 2911
rect 10031 2846 10037 2898
rect 10089 2846 10101 2898
rect 10153 2846 10165 2898
rect 10217 2846 10223 2898
rect 10031 2844 10038 2846
rect 10072 2844 10110 2846
rect 10144 2844 10182 2846
rect 10216 2844 10223 2846
rect 10031 2833 10223 2844
rect 10031 2781 10037 2833
rect 10089 2781 10101 2833
rect 10153 2781 10165 2833
rect 10217 2781 10223 2833
rect 10031 2770 10038 2781
rect 10072 2770 10110 2781
rect 10144 2770 10182 2781
rect 10216 2770 10223 2781
rect 10031 2768 10223 2770
rect 10031 2716 10037 2768
rect 10089 2716 10101 2768
rect 10153 2716 10165 2768
rect 10217 2716 10223 2768
rect 10031 2703 10038 2716
rect 10072 2703 10110 2716
rect 10144 2703 10182 2716
rect 10216 2703 10223 2716
rect 10031 2651 10037 2703
rect 10089 2651 10101 2703
rect 10153 2651 10165 2703
rect 10217 2651 10223 2703
rect 10031 2638 10038 2651
rect 10072 2638 10110 2651
rect 10144 2638 10182 2651
rect 10216 2638 10223 2651
rect 10031 2586 10037 2638
rect 10089 2586 10101 2638
rect 10153 2586 10165 2638
rect 10217 2586 10223 2638
rect 10031 2582 10223 2586
rect 10031 2573 10038 2582
rect 10072 2573 10110 2582
rect 10144 2573 10182 2582
rect 10216 2573 10223 2582
rect 10031 2521 10037 2573
rect 10089 2521 10101 2573
rect 10153 2521 10165 2573
rect 10217 2521 10223 2573
rect 10031 2508 10223 2521
rect 10031 2456 10037 2508
rect 10089 2456 10101 2508
rect 10153 2456 10165 2508
rect 10217 2456 10223 2508
rect 10031 2443 10223 2456
rect 10031 2391 10037 2443
rect 10089 2391 10101 2443
rect 10153 2391 10165 2443
rect 10217 2391 10223 2443
rect 10031 2378 10223 2391
rect 10031 2326 10037 2378
rect 10089 2326 10101 2378
rect 10153 2326 10165 2378
rect 10217 2326 10223 2378
rect 10031 2313 10223 2326
rect 10031 2261 10037 2313
rect 10089 2261 10101 2313
rect 10153 2261 10165 2313
rect 10217 2261 10223 2313
rect 10031 2252 10038 2261
rect 10072 2252 10110 2261
rect 10144 2252 10182 2261
rect 10216 2252 10223 2261
rect 10031 2248 10223 2252
rect 10031 2196 10037 2248
rect 10089 2196 10101 2248
rect 10153 2196 10165 2248
rect 10217 2196 10223 2248
rect 10031 2183 10038 2196
rect 10072 2183 10110 2196
rect 10144 2183 10182 2196
rect 10216 2183 10223 2196
rect 10031 2131 10037 2183
rect 10089 2131 10101 2183
rect 10153 2131 10165 2183
rect 10217 2131 10223 2183
rect 10031 2118 10038 2131
rect 10072 2118 10110 2131
rect 10144 2118 10182 2131
rect 10216 2118 10223 2131
rect 10031 2066 10037 2118
rect 10089 2066 10101 2118
rect 10153 2066 10165 2118
rect 10217 2066 10223 2118
rect 10031 2064 10223 2066
rect 10031 2053 10038 2064
rect 10072 2053 10110 2064
rect 10144 2053 10182 2064
rect 10216 2053 10223 2064
rect 10031 2001 10037 2053
rect 10089 2001 10101 2053
rect 10153 2001 10165 2053
rect 10217 2001 10223 2053
rect 10031 1990 10223 2001
rect 10031 1987 10038 1990
rect 10072 1987 10110 1990
rect 10144 1987 10182 1990
rect 10216 1987 10223 1990
rect 10031 1935 10037 1987
rect 10089 1935 10101 1987
rect 10153 1935 10165 1987
rect 10217 1935 10223 1987
rect 10031 1921 10223 1935
rect 10031 1869 10037 1921
rect 10089 1869 10101 1921
rect 10153 1869 10165 1921
rect 10217 1869 10223 1921
rect 10031 1855 10223 1869
rect 10031 1803 10037 1855
rect 10089 1803 10101 1855
rect 10153 1803 10165 1855
rect 10217 1803 10223 1855
rect 10031 1789 10223 1803
rect 10031 1737 10037 1789
rect 10089 1737 10101 1789
rect 10153 1737 10165 1789
rect 10217 1737 10223 1789
rect 10031 1734 10038 1737
rect 10072 1734 10110 1737
rect 10144 1734 10182 1737
rect 10216 1734 10223 1737
rect 10031 1723 10223 1734
rect 10031 1671 10037 1723
rect 10089 1671 10101 1723
rect 10153 1671 10165 1723
rect 10217 1671 10223 1723
rect 10031 1660 10038 1671
rect 10072 1660 10110 1671
rect 10144 1660 10182 1671
rect 10216 1660 10223 1671
rect 10031 1657 10223 1660
rect 10031 1605 10037 1657
rect 10089 1605 10101 1657
rect 10153 1605 10165 1657
rect 10217 1605 10223 1657
rect 10031 1591 10038 1605
rect 10072 1591 10110 1605
rect 10144 1591 10182 1605
rect 10216 1591 10223 1605
rect 10031 1539 10037 1591
rect 10089 1539 10101 1591
rect 10153 1539 10165 1591
rect 10217 1539 10223 1591
rect 10031 1525 10038 1539
rect 10072 1525 10110 1539
rect 10144 1525 10182 1539
rect 10216 1525 10223 1539
rect 10031 1473 10037 1525
rect 10089 1473 10101 1525
rect 10153 1473 10165 1525
rect 10217 1473 10223 1525
rect 10031 1467 10223 1473
rect 10527 4068 10719 4074
rect 10527 4016 10533 4068
rect 10585 4050 10597 4068
rect 10649 4050 10661 4068
rect 10713 4016 10719 4068
rect 10527 4003 10534 4016
rect 10712 4003 10719 4016
rect 10527 3951 10533 4003
rect 10713 3951 10719 4003
rect 10527 3938 10534 3951
rect 10712 3938 10719 3951
rect 10527 3886 10533 3938
rect 10713 3886 10719 3938
rect 10527 3873 10534 3886
rect 10712 3873 10719 3886
rect 10527 3821 10533 3873
rect 10713 3821 10719 3873
rect 10527 3808 10534 3821
rect 10712 3808 10719 3821
rect 10527 3756 10533 3808
rect 10713 3756 10719 3808
rect 10527 3743 10534 3756
rect 10712 3743 10719 3756
rect 10527 3691 10533 3743
rect 10713 3691 10719 3743
rect 10527 3678 10534 3691
rect 10712 3678 10719 3691
rect 10527 3626 10533 3678
rect 10713 3626 10719 3678
rect 10527 3613 10534 3626
rect 10712 3613 10719 3626
rect 10527 3561 10533 3613
rect 10713 3561 10719 3613
rect 10527 3548 10534 3561
rect 10712 3548 10719 3561
rect 10527 3496 10533 3548
rect 10713 3496 10719 3548
rect 10527 3483 10534 3496
rect 10712 3483 10719 3496
rect 10527 3431 10533 3483
rect 10713 3431 10719 3483
rect 10527 3418 10534 3431
rect 10712 3418 10719 3431
rect 10527 3366 10533 3418
rect 10713 3366 10719 3418
rect 10527 3353 10534 3366
rect 10712 3353 10719 3366
rect 10527 3301 10533 3353
rect 10713 3301 10719 3353
rect 10527 3288 10534 3301
rect 10712 3288 10719 3301
rect 10527 3236 10533 3288
rect 10713 3236 10719 3288
rect 10527 3223 10534 3236
rect 10712 3223 10719 3236
rect 10527 3171 10533 3223
rect 10713 3171 10719 3223
rect 10527 3158 10534 3171
rect 10712 3158 10719 3171
rect 10527 3106 10533 3158
rect 10713 3106 10719 3158
rect 10527 3093 10534 3106
rect 10712 3093 10719 3106
rect 10527 3041 10533 3093
rect 10585 3041 10597 3092
rect 10649 3041 10661 3092
rect 10713 3041 10719 3093
rect 10527 3037 10719 3041
rect 10527 3028 10534 3037
rect 10568 3028 10606 3037
rect 10640 3028 10678 3037
rect 10712 3028 10719 3037
rect 10527 2976 10533 3028
rect 10585 2976 10597 3028
rect 10649 2976 10661 3028
rect 10713 2976 10719 3028
rect 10527 2963 10719 2976
rect 10527 2911 10533 2963
rect 10585 2911 10597 2963
rect 10649 2911 10661 2963
rect 10713 2911 10719 2963
rect 10527 2898 10719 2911
rect 10527 2846 10533 2898
rect 10585 2846 10597 2898
rect 10649 2846 10661 2898
rect 10713 2846 10719 2898
rect 10527 2837 10534 2846
rect 10568 2837 10606 2846
rect 10640 2837 10678 2846
rect 10712 2837 10719 2846
rect 10527 2833 10719 2837
rect 10527 2781 10533 2833
rect 10585 2781 10597 2833
rect 10649 2781 10661 2833
rect 10713 2781 10719 2833
rect 10527 2768 10534 2781
rect 10568 2768 10606 2781
rect 10640 2768 10678 2781
rect 10712 2768 10719 2781
rect 10527 2716 10533 2768
rect 10585 2716 10597 2768
rect 10649 2716 10661 2768
rect 10713 2716 10719 2768
rect 10527 2703 10719 2716
rect 10527 2651 10533 2703
rect 10585 2651 10597 2703
rect 10649 2651 10661 2703
rect 10713 2651 10719 2703
rect 10527 2638 10719 2651
rect 10527 2586 10533 2638
rect 10585 2586 10597 2638
rect 10649 2586 10661 2638
rect 10713 2586 10719 2638
rect 10527 2585 10534 2586
rect 10568 2585 10606 2586
rect 10640 2585 10678 2586
rect 10712 2585 10719 2586
rect 10527 2573 10719 2585
rect 10527 2521 10533 2573
rect 10585 2521 10597 2573
rect 10649 2521 10661 2573
rect 10713 2521 10719 2573
rect 10527 2508 10534 2521
rect 10568 2508 10606 2521
rect 10640 2508 10678 2521
rect 10712 2508 10719 2521
rect 10527 2456 10533 2508
rect 10585 2456 10597 2508
rect 10649 2456 10661 2508
rect 10713 2456 10719 2508
rect 10527 2449 10606 2456
rect 10640 2449 10719 2456
rect 10527 2443 10534 2449
rect 10712 2443 10719 2449
rect 10527 2391 10533 2443
rect 10713 2391 10719 2443
rect 10527 2378 10534 2391
rect 10712 2378 10719 2391
rect 10527 2326 10533 2378
rect 10713 2326 10719 2378
rect 10527 2313 10534 2326
rect 10712 2313 10719 2326
rect 10527 2261 10533 2313
rect 10713 2261 10719 2313
rect 10527 2248 10534 2261
rect 10712 2248 10719 2261
rect 10527 2196 10533 2248
rect 10713 2196 10719 2248
rect 10527 2183 10534 2196
rect 10712 2183 10719 2196
rect 10527 2131 10533 2183
rect 10713 2131 10719 2183
rect 10527 2118 10534 2131
rect 10712 2118 10719 2131
rect 10527 2066 10533 2118
rect 10713 2066 10719 2118
rect 10527 2053 10534 2066
rect 10712 2053 10719 2066
rect 10527 2001 10533 2053
rect 10713 2001 10719 2053
rect 10527 1987 10534 2001
rect 10712 1987 10719 2001
rect 10527 1935 10533 1987
rect 10713 1935 10719 1987
rect 10527 1921 10534 1935
rect 10712 1921 10719 1935
rect 10527 1869 10533 1921
rect 10713 1869 10719 1921
rect 10527 1855 10534 1869
rect 10712 1855 10719 1869
rect 10527 1803 10533 1855
rect 10713 1803 10719 1855
rect 10527 1789 10534 1803
rect 10712 1789 10719 1803
rect 10527 1737 10533 1789
rect 10713 1737 10719 1789
rect 10527 1723 10534 1737
rect 10712 1723 10719 1737
rect 10527 1671 10533 1723
rect 10713 1671 10719 1723
rect 10527 1657 10534 1671
rect 10712 1657 10719 1671
rect 10527 1605 10533 1657
rect 10713 1605 10719 1657
rect 10527 1591 10534 1605
rect 10712 1591 10719 1605
rect 10527 1539 10533 1591
rect 10713 1539 10719 1591
rect 10527 1525 10534 1539
rect 10712 1525 10719 1539
rect 10527 1473 10533 1525
rect 10585 1473 10597 1491
rect 10649 1473 10661 1491
rect 10713 1473 10719 1525
rect 10527 1467 10719 1473
rect 11023 4068 11215 4074
rect 11023 4016 11029 4068
rect 11081 4016 11093 4068
rect 11145 4016 11157 4068
rect 11209 4016 11215 4068
rect 11023 4003 11215 4016
rect 11023 3951 11029 4003
rect 11081 3951 11093 4003
rect 11145 3951 11157 4003
rect 11209 3951 11215 4003
rect 11023 3938 11215 3951
rect 11023 3886 11029 3938
rect 11081 3886 11093 3938
rect 11145 3886 11157 3938
rect 11209 3886 11215 3938
rect 11023 3880 11030 3886
rect 11064 3880 11102 3886
rect 11136 3880 11174 3886
rect 11208 3880 11215 3886
rect 11023 3873 11215 3880
rect 11023 3821 11029 3873
rect 11081 3821 11093 3873
rect 11145 3821 11157 3873
rect 11209 3821 11215 3873
rect 11023 3808 11030 3821
rect 11064 3808 11102 3821
rect 11136 3808 11174 3821
rect 11208 3808 11215 3821
rect 11023 3756 11029 3808
rect 11081 3756 11093 3808
rect 11145 3756 11157 3808
rect 11209 3756 11215 3808
rect 11023 3743 11030 3756
rect 11064 3743 11102 3756
rect 11136 3743 11174 3756
rect 11208 3743 11215 3756
rect 11023 3691 11029 3743
rect 11081 3691 11093 3743
rect 11145 3691 11157 3743
rect 11209 3691 11215 3743
rect 11023 3678 11030 3691
rect 11064 3678 11102 3691
rect 11136 3678 11174 3691
rect 11208 3678 11215 3691
rect 11023 3626 11029 3678
rect 11081 3626 11093 3678
rect 11145 3626 11157 3678
rect 11209 3626 11215 3678
rect 11023 3618 11215 3626
rect 11023 3613 11030 3618
rect 11064 3613 11102 3618
rect 11136 3613 11174 3618
rect 11208 3613 11215 3618
rect 11023 3561 11029 3613
rect 11081 3561 11093 3613
rect 11145 3561 11157 3613
rect 11209 3561 11215 3613
rect 11023 3548 11215 3561
rect 11023 3496 11029 3548
rect 11081 3496 11093 3548
rect 11145 3496 11157 3548
rect 11209 3496 11215 3548
rect 11023 3483 11215 3496
rect 11023 3431 11029 3483
rect 11081 3431 11093 3483
rect 11145 3431 11157 3483
rect 11209 3431 11215 3483
rect 11023 3418 11215 3431
rect 11023 3366 11029 3418
rect 11081 3366 11093 3418
rect 11145 3366 11157 3418
rect 11209 3366 11215 3418
rect 11023 3362 11030 3366
rect 11064 3362 11102 3366
rect 11136 3362 11174 3366
rect 11208 3362 11215 3366
rect 11023 3353 11215 3362
rect 11023 3301 11029 3353
rect 11081 3301 11093 3353
rect 11145 3301 11157 3353
rect 11209 3301 11215 3353
rect 11023 3288 11030 3301
rect 11064 3288 11102 3301
rect 11136 3288 11174 3301
rect 11208 3288 11215 3301
rect 11023 3236 11029 3288
rect 11081 3236 11093 3288
rect 11145 3236 11157 3288
rect 11209 3236 11215 3288
rect 11023 3223 11030 3236
rect 11064 3223 11102 3236
rect 11136 3223 11174 3236
rect 11208 3223 11215 3236
rect 11023 3171 11029 3223
rect 11081 3171 11093 3223
rect 11145 3171 11157 3223
rect 11209 3171 11215 3223
rect 11023 3158 11030 3171
rect 11064 3158 11102 3171
rect 11136 3158 11174 3171
rect 11208 3158 11215 3171
rect 11023 3106 11029 3158
rect 11081 3106 11093 3158
rect 11145 3106 11157 3158
rect 11209 3106 11215 3158
rect 11023 3100 11215 3106
rect 11023 3093 11030 3100
rect 11064 3093 11102 3100
rect 11136 3093 11174 3100
rect 11208 3093 11215 3100
rect 11023 3041 11029 3093
rect 11081 3041 11093 3093
rect 11145 3041 11157 3093
rect 11209 3041 11215 3093
rect 11023 3028 11215 3041
rect 11023 2976 11029 3028
rect 11081 2976 11093 3028
rect 11145 2976 11157 3028
rect 11209 2976 11215 3028
rect 11023 2963 11215 2976
rect 11023 2911 11029 2963
rect 11081 2911 11093 2963
rect 11145 2911 11157 2963
rect 11209 2911 11215 2963
rect 11023 2898 11215 2911
rect 11023 2846 11029 2898
rect 11081 2846 11093 2898
rect 11145 2846 11157 2898
rect 11209 2846 11215 2898
rect 11023 2844 11030 2846
rect 11064 2844 11102 2846
rect 11136 2844 11174 2846
rect 11208 2844 11215 2846
rect 11023 2833 11215 2844
rect 11023 2781 11029 2833
rect 11081 2781 11093 2833
rect 11145 2781 11157 2833
rect 11209 2781 11215 2833
rect 11023 2770 11030 2781
rect 11064 2770 11102 2781
rect 11136 2770 11174 2781
rect 11208 2770 11215 2781
rect 11023 2768 11215 2770
rect 11023 2716 11029 2768
rect 11081 2716 11093 2768
rect 11145 2716 11157 2768
rect 11209 2716 11215 2768
rect 11023 2703 11030 2716
rect 11064 2703 11102 2716
rect 11136 2703 11174 2716
rect 11208 2703 11215 2716
rect 11023 2651 11029 2703
rect 11081 2651 11093 2703
rect 11145 2651 11157 2703
rect 11209 2651 11215 2703
rect 11023 2638 11030 2651
rect 11064 2638 11102 2651
rect 11136 2638 11174 2651
rect 11208 2638 11215 2651
rect 11023 2586 11029 2638
rect 11081 2586 11093 2638
rect 11145 2586 11157 2638
rect 11209 2586 11215 2638
rect 11023 2582 11215 2586
rect 11023 2573 11030 2582
rect 11064 2573 11102 2582
rect 11136 2573 11174 2582
rect 11208 2573 11215 2582
rect 11023 2521 11029 2573
rect 11081 2521 11093 2573
rect 11145 2521 11157 2573
rect 11209 2521 11215 2573
rect 11023 2508 11215 2521
rect 11023 2456 11029 2508
rect 11081 2456 11093 2508
rect 11145 2456 11157 2508
rect 11209 2456 11215 2508
rect 11023 2443 11215 2456
rect 11023 2391 11029 2443
rect 11081 2391 11093 2443
rect 11145 2391 11157 2443
rect 11209 2391 11215 2443
rect 11023 2378 11215 2391
rect 11023 2326 11029 2378
rect 11081 2326 11093 2378
rect 11145 2326 11157 2378
rect 11209 2326 11215 2378
rect 11023 2313 11215 2326
rect 11023 2261 11029 2313
rect 11081 2261 11093 2313
rect 11145 2261 11157 2313
rect 11209 2261 11215 2313
rect 11023 2252 11030 2261
rect 11064 2252 11102 2261
rect 11136 2252 11174 2261
rect 11208 2252 11215 2261
rect 11023 2248 11215 2252
rect 11023 2196 11029 2248
rect 11081 2196 11093 2248
rect 11145 2196 11157 2248
rect 11209 2196 11215 2248
rect 11023 2183 11030 2196
rect 11064 2183 11102 2196
rect 11136 2183 11174 2196
rect 11208 2183 11215 2196
rect 11023 2131 11029 2183
rect 11081 2131 11093 2183
rect 11145 2131 11157 2183
rect 11209 2131 11215 2183
rect 11023 2118 11030 2131
rect 11064 2118 11102 2131
rect 11136 2118 11174 2131
rect 11208 2118 11215 2131
rect 11023 2066 11029 2118
rect 11081 2066 11093 2118
rect 11145 2066 11157 2118
rect 11209 2066 11215 2118
rect 11023 2064 11215 2066
rect 11023 2053 11030 2064
rect 11064 2053 11102 2064
rect 11136 2053 11174 2064
rect 11208 2053 11215 2064
rect 11023 2001 11029 2053
rect 11081 2001 11093 2053
rect 11145 2001 11157 2053
rect 11209 2001 11215 2053
rect 11023 1990 11215 2001
rect 11023 1987 11030 1990
rect 11064 1987 11102 1990
rect 11136 1987 11174 1990
rect 11208 1987 11215 1990
rect 11023 1935 11029 1987
rect 11081 1935 11093 1987
rect 11145 1935 11157 1987
rect 11209 1935 11215 1987
rect 11023 1921 11215 1935
rect 11023 1869 11029 1921
rect 11081 1869 11093 1921
rect 11145 1869 11157 1921
rect 11209 1869 11215 1921
rect 11023 1855 11215 1869
rect 11023 1803 11029 1855
rect 11081 1803 11093 1855
rect 11145 1803 11157 1855
rect 11209 1803 11215 1855
rect 11023 1789 11215 1803
rect 11023 1737 11029 1789
rect 11081 1737 11093 1789
rect 11145 1737 11157 1789
rect 11209 1737 11215 1789
rect 11023 1734 11030 1737
rect 11064 1734 11102 1737
rect 11136 1734 11174 1737
rect 11208 1734 11215 1737
rect 11023 1723 11215 1734
rect 11023 1671 11029 1723
rect 11081 1671 11093 1723
rect 11145 1671 11157 1723
rect 11209 1671 11215 1723
rect 11023 1660 11030 1671
rect 11064 1660 11102 1671
rect 11136 1660 11174 1671
rect 11208 1660 11215 1671
rect 11023 1657 11215 1660
rect 11023 1605 11029 1657
rect 11081 1605 11093 1657
rect 11145 1605 11157 1657
rect 11209 1605 11215 1657
rect 11023 1591 11030 1605
rect 11064 1591 11102 1605
rect 11136 1591 11174 1605
rect 11208 1591 11215 1605
rect 11023 1539 11029 1591
rect 11081 1539 11093 1591
rect 11145 1539 11157 1591
rect 11209 1539 11215 1591
rect 11023 1525 11030 1539
rect 11064 1525 11102 1539
rect 11136 1525 11174 1539
rect 11208 1525 11215 1539
rect 11023 1473 11029 1525
rect 11081 1473 11093 1525
rect 11145 1473 11157 1525
rect 11209 1473 11215 1525
rect 11023 1467 11215 1473
rect 11519 4068 11711 4074
rect 11519 4016 11525 4068
rect 11577 4050 11589 4068
rect 11641 4050 11653 4068
rect 11705 4016 11711 4068
rect 11519 4003 11526 4016
rect 11704 4003 11711 4016
rect 11519 3951 11525 4003
rect 11705 3951 11711 4003
rect 11519 3938 11526 3951
rect 11704 3938 11711 3951
rect 11519 3886 11525 3938
rect 11705 3886 11711 3938
rect 11519 3873 11526 3886
rect 11704 3873 11711 3886
rect 11519 3821 11525 3873
rect 11705 3821 11711 3873
rect 11519 3808 11526 3821
rect 11704 3808 11711 3821
rect 11519 3756 11525 3808
rect 11705 3756 11711 3808
rect 11519 3743 11526 3756
rect 11704 3743 11711 3756
rect 11519 3691 11525 3743
rect 11705 3691 11711 3743
rect 11519 3678 11526 3691
rect 11704 3678 11711 3691
rect 11519 3626 11525 3678
rect 11705 3626 11711 3678
rect 11519 3613 11526 3626
rect 11704 3613 11711 3626
rect 11519 3561 11525 3613
rect 11705 3561 11711 3613
rect 11519 3548 11526 3561
rect 11704 3548 11711 3561
rect 11519 3496 11525 3548
rect 11705 3496 11711 3548
rect 11519 3483 11526 3496
rect 11704 3483 11711 3496
rect 11519 3431 11525 3483
rect 11705 3431 11711 3483
rect 11519 3418 11526 3431
rect 11704 3418 11711 3431
rect 11519 3366 11525 3418
rect 11705 3366 11711 3418
rect 11519 3353 11526 3366
rect 11704 3353 11711 3366
rect 11519 3301 11525 3353
rect 11705 3301 11711 3353
rect 11519 3288 11526 3301
rect 11704 3288 11711 3301
rect 11519 3236 11525 3288
rect 11705 3236 11711 3288
rect 11519 3223 11526 3236
rect 11704 3223 11711 3236
rect 11519 3171 11525 3223
rect 11705 3171 11711 3223
rect 11519 3158 11526 3171
rect 11704 3158 11711 3171
rect 11519 3106 11525 3158
rect 11705 3106 11711 3158
rect 11519 3093 11526 3106
rect 11704 3093 11711 3106
rect 11519 3041 11525 3093
rect 11577 3041 11589 3092
rect 11641 3041 11653 3092
rect 11705 3041 11711 3093
rect 11519 3037 11711 3041
rect 11519 3028 11526 3037
rect 11560 3028 11598 3037
rect 11632 3028 11670 3037
rect 11704 3028 11711 3037
rect 11519 2976 11525 3028
rect 11577 2976 11589 3028
rect 11641 2976 11653 3028
rect 11705 2976 11711 3028
rect 11519 2963 11711 2976
rect 11519 2911 11525 2963
rect 11577 2911 11589 2963
rect 11641 2911 11653 2963
rect 11705 2911 11711 2963
rect 11519 2898 11711 2911
rect 11519 2846 11525 2898
rect 11577 2846 11589 2898
rect 11641 2846 11653 2898
rect 11705 2846 11711 2898
rect 11519 2837 11526 2846
rect 11560 2837 11598 2846
rect 11632 2837 11670 2846
rect 11704 2837 11711 2846
rect 11519 2833 11711 2837
rect 11519 2781 11525 2833
rect 11577 2781 11589 2833
rect 11641 2781 11653 2833
rect 11705 2781 11711 2833
rect 11519 2768 11526 2781
rect 11560 2768 11598 2781
rect 11632 2768 11670 2781
rect 11704 2768 11711 2781
rect 11519 2716 11525 2768
rect 11577 2716 11589 2768
rect 11641 2716 11653 2768
rect 11705 2716 11711 2768
rect 11519 2703 11711 2716
rect 11519 2651 11525 2703
rect 11577 2651 11589 2703
rect 11641 2651 11653 2703
rect 11705 2651 11711 2703
rect 11519 2638 11711 2651
rect 11519 2586 11525 2638
rect 11577 2586 11589 2638
rect 11641 2586 11653 2638
rect 11705 2586 11711 2638
rect 11519 2585 11526 2586
rect 11560 2585 11598 2586
rect 11632 2585 11670 2586
rect 11704 2585 11711 2586
rect 11519 2573 11711 2585
rect 11519 2521 11525 2573
rect 11577 2521 11589 2573
rect 11641 2521 11653 2573
rect 11705 2521 11711 2573
rect 11519 2508 11526 2521
rect 11560 2508 11598 2521
rect 11632 2508 11670 2521
rect 11704 2508 11711 2521
rect 11519 2456 11525 2508
rect 11577 2456 11589 2508
rect 11641 2456 11653 2508
rect 11705 2456 11711 2508
rect 11519 2449 11598 2456
rect 11632 2449 11711 2456
rect 11519 2443 11526 2449
rect 11704 2443 11711 2449
rect 11519 2391 11525 2443
rect 11705 2391 11711 2443
rect 11519 2378 11526 2391
rect 11704 2378 11711 2391
rect 11519 2326 11525 2378
rect 11705 2326 11711 2378
rect 11519 2313 11526 2326
rect 11704 2313 11711 2326
rect 11519 2261 11525 2313
rect 11705 2261 11711 2313
rect 11519 2248 11526 2261
rect 11704 2248 11711 2261
rect 11519 2196 11525 2248
rect 11705 2196 11711 2248
rect 11519 2183 11526 2196
rect 11704 2183 11711 2196
rect 11519 2131 11525 2183
rect 11705 2131 11711 2183
rect 11519 2118 11526 2131
rect 11704 2118 11711 2131
rect 11519 2066 11525 2118
rect 11705 2066 11711 2118
rect 11519 2053 11526 2066
rect 11704 2053 11711 2066
rect 11519 2001 11525 2053
rect 11705 2001 11711 2053
rect 11519 1987 11526 2001
rect 11704 1987 11711 2001
rect 11519 1935 11525 1987
rect 11705 1935 11711 1987
rect 11519 1921 11526 1935
rect 11704 1921 11711 1935
rect 11519 1869 11525 1921
rect 11705 1869 11711 1921
rect 11519 1855 11526 1869
rect 11704 1855 11711 1869
rect 11519 1803 11525 1855
rect 11705 1803 11711 1855
rect 11519 1789 11526 1803
rect 11704 1789 11711 1803
rect 11519 1737 11525 1789
rect 11705 1737 11711 1789
rect 11519 1723 11526 1737
rect 11704 1723 11711 1737
rect 11519 1671 11525 1723
rect 11705 1671 11711 1723
rect 11519 1657 11526 1671
rect 11704 1657 11711 1671
rect 11519 1605 11525 1657
rect 11705 1605 11711 1657
rect 11519 1591 11526 1605
rect 11704 1591 11711 1605
rect 11519 1539 11525 1591
rect 11705 1539 11711 1591
rect 11519 1525 11526 1539
rect 11704 1525 11711 1539
rect 11519 1473 11525 1525
rect 11577 1473 11589 1491
rect 11641 1473 11653 1491
rect 11705 1473 11711 1525
rect 11519 1467 11711 1473
rect 12015 4068 12207 4074
rect 12015 4016 12021 4068
rect 12073 4016 12085 4068
rect 12137 4016 12149 4068
rect 12201 4016 12207 4068
rect 12015 4003 12207 4016
rect 12015 3951 12021 4003
rect 12073 3951 12085 4003
rect 12137 3951 12149 4003
rect 12201 3951 12207 4003
rect 12015 3938 12207 3951
rect 12015 3886 12021 3938
rect 12073 3886 12085 3938
rect 12137 3886 12149 3938
rect 12201 3886 12207 3938
rect 12015 3880 12022 3886
rect 12056 3880 12094 3886
rect 12128 3880 12166 3886
rect 12200 3880 12207 3886
rect 12015 3873 12207 3880
rect 12015 3821 12021 3873
rect 12073 3821 12085 3873
rect 12137 3821 12149 3873
rect 12201 3821 12207 3873
rect 12015 3808 12022 3821
rect 12056 3808 12094 3821
rect 12128 3808 12166 3821
rect 12200 3808 12207 3821
rect 12015 3756 12021 3808
rect 12073 3756 12085 3808
rect 12137 3756 12149 3808
rect 12201 3756 12207 3808
rect 12015 3743 12022 3756
rect 12056 3743 12094 3756
rect 12128 3743 12166 3756
rect 12200 3743 12207 3756
rect 12015 3691 12021 3743
rect 12073 3691 12085 3743
rect 12137 3691 12149 3743
rect 12201 3691 12207 3743
rect 12015 3678 12022 3691
rect 12056 3678 12094 3691
rect 12128 3678 12166 3691
rect 12200 3678 12207 3691
rect 12015 3626 12021 3678
rect 12073 3626 12085 3678
rect 12137 3626 12149 3678
rect 12201 3626 12207 3678
rect 12015 3618 12207 3626
rect 12015 3613 12022 3618
rect 12056 3613 12094 3618
rect 12128 3613 12166 3618
rect 12200 3613 12207 3618
rect 12015 3561 12021 3613
rect 12073 3561 12085 3613
rect 12137 3561 12149 3613
rect 12201 3561 12207 3613
rect 12015 3548 12207 3561
rect 12015 3496 12021 3548
rect 12073 3496 12085 3548
rect 12137 3496 12149 3548
rect 12201 3496 12207 3548
rect 12015 3483 12207 3496
rect 12015 3431 12021 3483
rect 12073 3431 12085 3483
rect 12137 3431 12149 3483
rect 12201 3431 12207 3483
rect 12015 3418 12207 3431
rect 12015 3366 12021 3418
rect 12073 3366 12085 3418
rect 12137 3366 12149 3418
rect 12201 3366 12207 3418
rect 12015 3362 12022 3366
rect 12056 3362 12094 3366
rect 12128 3362 12166 3366
rect 12200 3362 12207 3366
rect 12015 3353 12207 3362
rect 12015 3301 12021 3353
rect 12073 3301 12085 3353
rect 12137 3301 12149 3353
rect 12201 3301 12207 3353
rect 12015 3288 12022 3301
rect 12056 3288 12094 3301
rect 12128 3288 12166 3301
rect 12200 3288 12207 3301
rect 12015 3236 12021 3288
rect 12073 3236 12085 3288
rect 12137 3236 12149 3288
rect 12201 3236 12207 3288
rect 12015 3223 12022 3236
rect 12056 3223 12094 3236
rect 12128 3223 12166 3236
rect 12200 3223 12207 3236
rect 12015 3171 12021 3223
rect 12073 3171 12085 3223
rect 12137 3171 12149 3223
rect 12201 3171 12207 3223
rect 12015 3158 12022 3171
rect 12056 3158 12094 3171
rect 12128 3158 12166 3171
rect 12200 3158 12207 3171
rect 12015 3106 12021 3158
rect 12073 3106 12085 3158
rect 12137 3106 12149 3158
rect 12201 3106 12207 3158
rect 12015 3100 12207 3106
rect 12015 3093 12022 3100
rect 12056 3093 12094 3100
rect 12128 3093 12166 3100
rect 12200 3093 12207 3100
rect 12015 3041 12021 3093
rect 12073 3041 12085 3093
rect 12137 3041 12149 3093
rect 12201 3041 12207 3093
rect 12015 3028 12207 3041
rect 12015 2976 12021 3028
rect 12073 2976 12085 3028
rect 12137 2976 12149 3028
rect 12201 2976 12207 3028
rect 12015 2963 12207 2976
rect 12015 2911 12021 2963
rect 12073 2911 12085 2963
rect 12137 2911 12149 2963
rect 12201 2911 12207 2963
rect 12015 2898 12207 2911
rect 12015 2846 12021 2898
rect 12073 2846 12085 2898
rect 12137 2846 12149 2898
rect 12201 2846 12207 2898
rect 12015 2844 12022 2846
rect 12056 2844 12094 2846
rect 12128 2844 12166 2846
rect 12200 2844 12207 2846
rect 12015 2833 12207 2844
rect 12015 2781 12021 2833
rect 12073 2781 12085 2833
rect 12137 2781 12149 2833
rect 12201 2781 12207 2833
rect 12015 2770 12022 2781
rect 12056 2770 12094 2781
rect 12128 2770 12166 2781
rect 12200 2770 12207 2781
rect 12015 2768 12207 2770
rect 12015 2716 12021 2768
rect 12073 2716 12085 2768
rect 12137 2716 12149 2768
rect 12201 2716 12207 2768
rect 12015 2703 12022 2716
rect 12056 2703 12094 2716
rect 12128 2703 12166 2716
rect 12200 2703 12207 2716
rect 12015 2651 12021 2703
rect 12073 2651 12085 2703
rect 12137 2651 12149 2703
rect 12201 2651 12207 2703
rect 12015 2638 12022 2651
rect 12056 2638 12094 2651
rect 12128 2638 12166 2651
rect 12200 2638 12207 2651
rect 12015 2586 12021 2638
rect 12073 2586 12085 2638
rect 12137 2586 12149 2638
rect 12201 2586 12207 2638
rect 12015 2582 12207 2586
rect 12015 2573 12022 2582
rect 12056 2573 12094 2582
rect 12128 2573 12166 2582
rect 12200 2573 12207 2582
rect 12015 2521 12021 2573
rect 12073 2521 12085 2573
rect 12137 2521 12149 2573
rect 12201 2521 12207 2573
rect 12015 2508 12207 2521
rect 12015 2456 12021 2508
rect 12073 2456 12085 2508
rect 12137 2456 12149 2508
rect 12201 2456 12207 2508
rect 12015 2443 12207 2456
rect 12015 2391 12021 2443
rect 12073 2391 12085 2443
rect 12137 2391 12149 2443
rect 12201 2391 12207 2443
rect 12015 2378 12207 2391
rect 12015 2326 12021 2378
rect 12073 2326 12085 2378
rect 12137 2326 12149 2378
rect 12201 2326 12207 2378
rect 12015 2313 12207 2326
rect 12015 2261 12021 2313
rect 12073 2261 12085 2313
rect 12137 2261 12149 2313
rect 12201 2261 12207 2313
rect 12015 2252 12022 2261
rect 12056 2252 12094 2261
rect 12128 2252 12166 2261
rect 12200 2252 12207 2261
rect 12015 2248 12207 2252
rect 12015 2196 12021 2248
rect 12073 2196 12085 2248
rect 12137 2196 12149 2248
rect 12201 2196 12207 2248
rect 12015 2183 12022 2196
rect 12056 2183 12094 2196
rect 12128 2183 12166 2196
rect 12200 2183 12207 2196
rect 12015 2131 12021 2183
rect 12073 2131 12085 2183
rect 12137 2131 12149 2183
rect 12201 2131 12207 2183
rect 12015 2118 12022 2131
rect 12056 2118 12094 2131
rect 12128 2118 12166 2131
rect 12200 2118 12207 2131
rect 12015 2066 12021 2118
rect 12073 2066 12085 2118
rect 12137 2066 12149 2118
rect 12201 2066 12207 2118
rect 12015 2064 12207 2066
rect 12015 2053 12022 2064
rect 12056 2053 12094 2064
rect 12128 2053 12166 2064
rect 12200 2053 12207 2064
rect 12015 2001 12021 2053
rect 12073 2001 12085 2053
rect 12137 2001 12149 2053
rect 12201 2001 12207 2053
rect 12015 1990 12207 2001
rect 12015 1987 12022 1990
rect 12056 1987 12094 1990
rect 12128 1987 12166 1990
rect 12200 1987 12207 1990
rect 12015 1935 12021 1987
rect 12073 1935 12085 1987
rect 12137 1935 12149 1987
rect 12201 1935 12207 1987
rect 12015 1921 12207 1935
rect 12015 1869 12021 1921
rect 12073 1869 12085 1921
rect 12137 1869 12149 1921
rect 12201 1869 12207 1921
rect 12015 1855 12207 1869
rect 12015 1803 12021 1855
rect 12073 1803 12085 1855
rect 12137 1803 12149 1855
rect 12201 1803 12207 1855
rect 12015 1789 12207 1803
rect 12015 1737 12021 1789
rect 12073 1737 12085 1789
rect 12137 1737 12149 1789
rect 12201 1737 12207 1789
rect 12015 1734 12022 1737
rect 12056 1734 12094 1737
rect 12128 1734 12166 1737
rect 12200 1734 12207 1737
rect 12015 1723 12207 1734
rect 12015 1671 12021 1723
rect 12073 1671 12085 1723
rect 12137 1671 12149 1723
rect 12201 1671 12207 1723
rect 12015 1660 12022 1671
rect 12056 1660 12094 1671
rect 12128 1660 12166 1671
rect 12200 1660 12207 1671
rect 12015 1657 12207 1660
rect 12015 1605 12021 1657
rect 12073 1605 12085 1657
rect 12137 1605 12149 1657
rect 12201 1605 12207 1657
rect 12015 1591 12022 1605
rect 12056 1591 12094 1605
rect 12128 1591 12166 1605
rect 12200 1591 12207 1605
rect 12015 1539 12021 1591
rect 12073 1539 12085 1591
rect 12137 1539 12149 1591
rect 12201 1539 12207 1591
rect 12015 1525 12022 1539
rect 12056 1525 12094 1539
rect 12128 1525 12166 1539
rect 12200 1525 12207 1539
rect 12015 1473 12021 1525
rect 12073 1473 12085 1525
rect 12137 1473 12149 1525
rect 12201 1473 12207 1525
rect 12015 1467 12207 1473
rect 12511 4068 12703 4074
rect 12511 4016 12517 4068
rect 12569 4050 12581 4068
rect 12633 4050 12645 4068
rect 12697 4016 12703 4068
rect 12511 4003 12518 4016
rect 12696 4003 12703 4016
rect 12511 3951 12517 4003
rect 12697 3951 12703 4003
rect 12511 3938 12518 3951
rect 12696 3938 12703 3951
rect 12511 3886 12517 3938
rect 12697 3886 12703 3938
rect 12511 3873 12518 3886
rect 12696 3873 12703 3886
rect 12511 3821 12517 3873
rect 12697 3821 12703 3873
rect 12511 3808 12518 3821
rect 12696 3808 12703 3821
rect 12511 3756 12517 3808
rect 12697 3756 12703 3808
rect 12511 3743 12518 3756
rect 12696 3743 12703 3756
rect 12511 3691 12517 3743
rect 12697 3691 12703 3743
rect 12511 3678 12518 3691
rect 12696 3678 12703 3691
rect 12511 3626 12517 3678
rect 12697 3626 12703 3678
rect 12511 3613 12518 3626
rect 12696 3613 12703 3626
rect 12511 3561 12517 3613
rect 12697 3561 12703 3613
rect 12511 3548 12518 3561
rect 12696 3548 12703 3561
rect 12511 3496 12517 3548
rect 12697 3496 12703 3548
rect 12511 3483 12518 3496
rect 12696 3483 12703 3496
rect 12511 3431 12517 3483
rect 12697 3431 12703 3483
rect 12511 3418 12518 3431
rect 12696 3418 12703 3431
rect 12511 3366 12517 3418
rect 12697 3366 12703 3418
rect 12511 3353 12518 3366
rect 12696 3353 12703 3366
rect 12511 3301 12517 3353
rect 12697 3301 12703 3353
rect 12511 3288 12518 3301
rect 12696 3288 12703 3301
rect 12511 3236 12517 3288
rect 12697 3236 12703 3288
rect 12511 3223 12518 3236
rect 12696 3223 12703 3236
rect 12511 3171 12517 3223
rect 12697 3171 12703 3223
rect 12511 3158 12518 3171
rect 12696 3158 12703 3171
rect 12511 3106 12517 3158
rect 12697 3106 12703 3158
rect 12511 3093 12518 3106
rect 12696 3093 12703 3106
rect 12511 3041 12517 3093
rect 12569 3041 12581 3092
rect 12633 3041 12645 3092
rect 12697 3041 12703 3093
rect 12511 3038 12703 3041
rect 12511 3028 12518 3038
rect 12552 3028 12590 3038
rect 12624 3028 12662 3038
rect 12696 3028 12703 3038
rect 12511 2976 12517 3028
rect 12569 2976 12581 3028
rect 12633 2976 12645 3028
rect 12697 2976 12703 3028
rect 12511 2963 12703 2976
rect 12511 2911 12517 2963
rect 12569 2911 12581 2963
rect 12633 2911 12645 2963
rect 12697 2911 12703 2963
rect 12511 2898 12703 2911
rect 12511 2846 12517 2898
rect 12569 2846 12581 2898
rect 12633 2846 12645 2898
rect 12697 2846 12703 2898
rect 12511 2837 12518 2846
rect 12552 2837 12590 2846
rect 12624 2837 12662 2846
rect 12696 2837 12703 2846
rect 12511 2833 12703 2837
rect 12511 2781 12517 2833
rect 12569 2781 12581 2833
rect 12633 2781 12645 2833
rect 12697 2781 12703 2833
rect 12511 2768 12518 2781
rect 12552 2768 12590 2781
rect 12624 2768 12662 2781
rect 12696 2768 12703 2781
rect 12511 2716 12517 2768
rect 12569 2716 12581 2768
rect 12633 2716 12645 2768
rect 12697 2716 12703 2768
rect 12511 2703 12703 2716
rect 12511 2651 12517 2703
rect 12569 2651 12581 2703
rect 12633 2651 12645 2703
rect 12697 2651 12703 2703
rect 12511 2638 12703 2651
rect 12511 2586 12517 2638
rect 12569 2586 12581 2638
rect 12633 2586 12645 2638
rect 12697 2586 12703 2638
rect 12511 2585 12518 2586
rect 12552 2585 12590 2586
rect 12624 2585 12662 2586
rect 12696 2585 12703 2586
rect 12511 2573 12703 2585
rect 12511 2521 12517 2573
rect 12569 2521 12581 2573
rect 12633 2521 12645 2573
rect 12697 2521 12703 2573
rect 12511 2508 12518 2521
rect 12552 2508 12590 2521
rect 12624 2508 12662 2521
rect 12696 2508 12703 2521
rect 12511 2456 12517 2508
rect 12569 2456 12581 2508
rect 12633 2456 12645 2508
rect 12697 2456 12703 2508
rect 12511 2449 12590 2456
rect 12624 2449 12703 2456
rect 12511 2443 12518 2449
rect 12696 2443 12703 2449
rect 12511 2391 12517 2443
rect 12697 2391 12703 2443
rect 12511 2378 12518 2391
rect 12696 2378 12703 2391
rect 12511 2326 12517 2378
rect 12697 2326 12703 2378
rect 12511 2313 12518 2326
rect 12696 2313 12703 2326
rect 12511 2261 12517 2313
rect 12697 2261 12703 2313
rect 12511 2248 12518 2261
rect 12696 2248 12703 2261
rect 12511 2196 12517 2248
rect 12697 2196 12703 2248
rect 12511 2183 12518 2196
rect 12696 2183 12703 2196
rect 12511 2131 12517 2183
rect 12697 2131 12703 2183
rect 12511 2118 12518 2131
rect 12696 2118 12703 2131
rect 12511 2066 12517 2118
rect 12697 2066 12703 2118
rect 12511 2053 12518 2066
rect 12696 2053 12703 2066
rect 12511 2001 12517 2053
rect 12697 2001 12703 2053
rect 12511 1987 12518 2001
rect 12696 1987 12703 2001
rect 12511 1935 12517 1987
rect 12697 1935 12703 1987
rect 12511 1921 12518 1935
rect 12696 1921 12703 1935
rect 12511 1869 12517 1921
rect 12697 1869 12703 1921
rect 12511 1855 12518 1869
rect 12696 1855 12703 1869
rect 12511 1803 12517 1855
rect 12697 1803 12703 1855
rect 12511 1789 12518 1803
rect 12696 1789 12703 1803
rect 12511 1737 12517 1789
rect 12697 1737 12703 1789
rect 12511 1723 12518 1737
rect 12696 1723 12703 1737
rect 12511 1671 12517 1723
rect 12697 1671 12703 1723
rect 12511 1657 12518 1671
rect 12696 1657 12703 1671
rect 12511 1605 12517 1657
rect 12697 1605 12703 1657
rect 12511 1591 12518 1605
rect 12696 1591 12703 1605
rect 12511 1539 12517 1591
rect 12697 1539 12703 1591
rect 12511 1525 12518 1539
rect 12696 1525 12703 1539
rect 12511 1473 12517 1525
rect 12569 1473 12581 1491
rect 12633 1473 12645 1491
rect 12697 1473 12703 1525
rect 12511 1467 12703 1473
rect 13007 4068 13199 4074
rect 13007 4016 13013 4068
rect 13065 4016 13077 4068
rect 13129 4016 13141 4068
rect 13193 4016 13199 4068
rect 13007 4003 13199 4016
rect 13007 3951 13013 4003
rect 13065 3951 13077 4003
rect 13129 3951 13141 4003
rect 13193 3951 13199 4003
rect 13007 3938 13199 3951
rect 13007 3886 13013 3938
rect 13065 3886 13077 3938
rect 13129 3886 13141 3938
rect 13193 3886 13199 3938
rect 13007 3880 13014 3886
rect 13048 3880 13086 3886
rect 13120 3880 13158 3886
rect 13192 3880 13199 3886
rect 13007 3873 13199 3880
rect 13007 3821 13013 3873
rect 13065 3821 13077 3873
rect 13129 3821 13141 3873
rect 13193 3821 13199 3873
rect 13007 3808 13014 3821
rect 13048 3808 13086 3821
rect 13120 3808 13158 3821
rect 13192 3808 13199 3821
rect 13007 3756 13013 3808
rect 13065 3756 13077 3808
rect 13129 3756 13141 3808
rect 13193 3756 13199 3808
rect 13007 3743 13014 3756
rect 13048 3743 13086 3756
rect 13120 3743 13158 3756
rect 13192 3743 13199 3756
rect 13007 3691 13013 3743
rect 13065 3691 13077 3743
rect 13129 3691 13141 3743
rect 13193 3691 13199 3743
rect 13007 3678 13014 3691
rect 13048 3678 13086 3691
rect 13120 3678 13158 3691
rect 13192 3678 13199 3691
rect 13007 3626 13013 3678
rect 13065 3626 13077 3678
rect 13129 3626 13141 3678
rect 13193 3626 13199 3678
rect 13007 3618 13199 3626
rect 13007 3613 13014 3618
rect 13048 3613 13086 3618
rect 13120 3613 13158 3618
rect 13192 3613 13199 3618
rect 13007 3561 13013 3613
rect 13065 3561 13077 3613
rect 13129 3561 13141 3613
rect 13193 3561 13199 3613
rect 13007 3548 13199 3561
rect 13007 3496 13013 3548
rect 13065 3496 13077 3548
rect 13129 3496 13141 3548
rect 13193 3496 13199 3548
rect 13007 3483 13199 3496
rect 13007 3431 13013 3483
rect 13065 3431 13077 3483
rect 13129 3431 13141 3483
rect 13193 3431 13199 3483
rect 13007 3418 13199 3431
rect 13007 3366 13013 3418
rect 13065 3366 13077 3418
rect 13129 3366 13141 3418
rect 13193 3366 13199 3418
rect 13007 3362 13014 3366
rect 13048 3362 13086 3366
rect 13120 3362 13158 3366
rect 13192 3362 13199 3366
rect 13007 3353 13199 3362
rect 13007 3301 13013 3353
rect 13065 3301 13077 3353
rect 13129 3301 13141 3353
rect 13193 3301 13199 3353
rect 13007 3288 13014 3301
rect 13048 3288 13086 3301
rect 13120 3288 13158 3301
rect 13192 3288 13199 3301
rect 13007 3236 13013 3288
rect 13065 3236 13077 3288
rect 13129 3236 13141 3288
rect 13193 3236 13199 3288
rect 13007 3223 13014 3236
rect 13048 3223 13086 3236
rect 13120 3223 13158 3236
rect 13192 3223 13199 3236
rect 13007 3171 13013 3223
rect 13065 3171 13077 3223
rect 13129 3171 13141 3223
rect 13193 3171 13199 3223
rect 13007 3158 13014 3171
rect 13048 3158 13086 3171
rect 13120 3158 13158 3171
rect 13192 3158 13199 3171
rect 13007 3106 13013 3158
rect 13065 3106 13077 3158
rect 13129 3106 13141 3158
rect 13193 3106 13199 3158
rect 13007 3100 13199 3106
rect 13007 3093 13014 3100
rect 13048 3093 13086 3100
rect 13120 3093 13158 3100
rect 13192 3093 13199 3100
rect 13007 3041 13013 3093
rect 13065 3041 13077 3093
rect 13129 3041 13141 3093
rect 13193 3041 13199 3093
rect 13007 3028 13199 3041
rect 13007 2976 13013 3028
rect 13065 2976 13077 3028
rect 13129 2976 13141 3028
rect 13193 2976 13199 3028
rect 13007 2963 13199 2976
rect 13007 2911 13013 2963
rect 13065 2911 13077 2963
rect 13129 2911 13141 2963
rect 13193 2911 13199 2963
rect 13007 2898 13199 2911
rect 13007 2846 13013 2898
rect 13065 2846 13077 2898
rect 13129 2846 13141 2898
rect 13193 2846 13199 2898
rect 13007 2844 13014 2846
rect 13048 2844 13086 2846
rect 13120 2844 13158 2846
rect 13192 2844 13199 2846
rect 13007 2833 13199 2844
rect 13007 2781 13013 2833
rect 13065 2781 13077 2833
rect 13129 2781 13141 2833
rect 13193 2781 13199 2833
rect 13007 2770 13014 2781
rect 13048 2770 13086 2781
rect 13120 2770 13158 2781
rect 13192 2770 13199 2781
rect 13007 2768 13199 2770
rect 13007 2716 13013 2768
rect 13065 2716 13077 2768
rect 13129 2716 13141 2768
rect 13193 2716 13199 2768
rect 13007 2703 13014 2716
rect 13048 2703 13086 2716
rect 13120 2703 13158 2716
rect 13192 2703 13199 2716
rect 13007 2651 13013 2703
rect 13065 2651 13077 2703
rect 13129 2651 13141 2703
rect 13193 2651 13199 2703
rect 13007 2638 13014 2651
rect 13048 2638 13086 2651
rect 13120 2638 13158 2651
rect 13192 2638 13199 2651
rect 13007 2586 13013 2638
rect 13065 2586 13077 2638
rect 13129 2586 13141 2638
rect 13193 2586 13199 2638
rect 13007 2582 13199 2586
rect 13007 2573 13014 2582
rect 13048 2573 13086 2582
rect 13120 2573 13158 2582
rect 13192 2573 13199 2582
rect 13007 2521 13013 2573
rect 13065 2521 13077 2573
rect 13129 2521 13141 2573
rect 13193 2521 13199 2573
rect 13007 2508 13199 2521
rect 13007 2456 13013 2508
rect 13065 2456 13077 2508
rect 13129 2456 13141 2508
rect 13193 2456 13199 2508
rect 13007 2443 13199 2456
rect 13007 2391 13013 2443
rect 13065 2391 13077 2443
rect 13129 2391 13141 2443
rect 13193 2391 13199 2443
rect 13007 2378 13199 2391
rect 13007 2326 13013 2378
rect 13065 2326 13077 2378
rect 13129 2326 13141 2378
rect 13193 2326 13199 2378
rect 13007 2313 13199 2326
rect 13007 2261 13013 2313
rect 13065 2261 13077 2313
rect 13129 2261 13141 2313
rect 13193 2261 13199 2313
rect 13007 2252 13014 2261
rect 13048 2252 13086 2261
rect 13120 2252 13158 2261
rect 13192 2252 13199 2261
rect 13007 2248 13199 2252
rect 13007 2196 13013 2248
rect 13065 2196 13077 2248
rect 13129 2196 13141 2248
rect 13193 2196 13199 2248
rect 13007 2183 13014 2196
rect 13048 2183 13086 2196
rect 13120 2183 13158 2196
rect 13192 2183 13199 2196
rect 13007 2131 13013 2183
rect 13065 2131 13077 2183
rect 13129 2131 13141 2183
rect 13193 2131 13199 2183
rect 13007 2118 13014 2131
rect 13048 2118 13086 2131
rect 13120 2118 13158 2131
rect 13192 2118 13199 2131
rect 13007 2066 13013 2118
rect 13065 2066 13077 2118
rect 13129 2066 13141 2118
rect 13193 2066 13199 2118
rect 13007 2064 13199 2066
rect 13007 2053 13014 2064
rect 13048 2053 13086 2064
rect 13120 2053 13158 2064
rect 13192 2053 13199 2064
rect 13007 2001 13013 2053
rect 13065 2001 13077 2053
rect 13129 2001 13141 2053
rect 13193 2001 13199 2053
rect 13007 1990 13199 2001
rect 13007 1987 13014 1990
rect 13048 1987 13086 1990
rect 13120 1987 13158 1990
rect 13192 1987 13199 1990
rect 13007 1935 13013 1987
rect 13065 1935 13077 1987
rect 13129 1935 13141 1987
rect 13193 1935 13199 1987
rect 13007 1921 13199 1935
rect 13007 1869 13013 1921
rect 13065 1869 13077 1921
rect 13129 1869 13141 1921
rect 13193 1869 13199 1921
rect 13007 1855 13199 1869
rect 13007 1803 13013 1855
rect 13065 1803 13077 1855
rect 13129 1803 13141 1855
rect 13193 1803 13199 1855
rect 13007 1789 13199 1803
rect 13007 1737 13013 1789
rect 13065 1737 13077 1789
rect 13129 1737 13141 1789
rect 13193 1737 13199 1789
rect 13007 1734 13014 1737
rect 13048 1734 13086 1737
rect 13120 1734 13158 1737
rect 13192 1734 13199 1737
rect 13007 1723 13199 1734
rect 13007 1671 13013 1723
rect 13065 1671 13077 1723
rect 13129 1671 13141 1723
rect 13193 1671 13199 1723
rect 13007 1660 13014 1671
rect 13048 1660 13086 1671
rect 13120 1660 13158 1671
rect 13192 1660 13199 1671
rect 13007 1657 13199 1660
rect 13007 1605 13013 1657
rect 13065 1605 13077 1657
rect 13129 1605 13141 1657
rect 13193 1605 13199 1657
rect 13007 1591 13014 1605
rect 13048 1591 13086 1605
rect 13120 1591 13158 1605
rect 13192 1591 13199 1605
rect 13007 1539 13013 1591
rect 13065 1539 13077 1591
rect 13129 1539 13141 1591
rect 13193 1539 13199 1591
rect 13007 1525 13014 1539
rect 13048 1525 13086 1539
rect 13120 1525 13158 1539
rect 13192 1525 13199 1539
rect 13007 1473 13013 1525
rect 13065 1473 13077 1525
rect 13129 1473 13141 1525
rect 13193 1473 13199 1525
rect 13007 1467 13199 1473
rect 13503 4068 13695 4074
rect 13503 4016 13509 4068
rect 13561 4050 13573 4068
rect 13625 4050 13637 4068
rect 13689 4016 13695 4068
rect 13503 4003 13510 4016
rect 13688 4003 13695 4016
rect 13503 3951 13509 4003
rect 13689 3951 13695 4003
rect 13503 3938 13510 3951
rect 13688 3938 13695 3951
rect 13503 3886 13509 3938
rect 13689 3886 13695 3938
rect 13503 3873 13510 3886
rect 13688 3873 13695 3886
rect 13503 3821 13509 3873
rect 13689 3821 13695 3873
rect 13503 3808 13510 3821
rect 13688 3808 13695 3821
rect 13503 3756 13509 3808
rect 13689 3756 13695 3808
rect 13503 3743 13510 3756
rect 13688 3743 13695 3756
rect 13503 3691 13509 3743
rect 13689 3691 13695 3743
rect 13503 3678 13510 3691
rect 13688 3678 13695 3691
rect 13503 3626 13509 3678
rect 13689 3626 13695 3678
rect 13503 3613 13510 3626
rect 13688 3613 13695 3626
rect 13503 3561 13509 3613
rect 13689 3561 13695 3613
rect 13503 3548 13510 3561
rect 13688 3548 13695 3561
rect 13503 3496 13509 3548
rect 13689 3496 13695 3548
rect 13503 3483 13510 3496
rect 13688 3483 13695 3496
rect 13503 3431 13509 3483
rect 13689 3431 13695 3483
rect 13503 3418 13510 3431
rect 13688 3418 13695 3431
rect 13503 3366 13509 3418
rect 13689 3366 13695 3418
rect 13503 3353 13510 3366
rect 13688 3353 13695 3366
rect 13503 3301 13509 3353
rect 13689 3301 13695 3353
rect 13503 3288 13510 3301
rect 13688 3288 13695 3301
rect 13503 3236 13509 3288
rect 13689 3236 13695 3288
rect 13503 3223 13510 3236
rect 13688 3223 13695 3236
rect 13503 3171 13509 3223
rect 13689 3171 13695 3223
rect 13503 3158 13510 3171
rect 13688 3158 13695 3171
rect 13503 3106 13509 3158
rect 13689 3106 13695 3158
rect 13503 3093 13510 3106
rect 13688 3093 13695 3106
rect 13503 3041 13509 3093
rect 13561 3041 13573 3092
rect 13625 3041 13637 3092
rect 13689 3041 13695 3093
rect 13503 3040 13695 3041
rect 13503 3028 13510 3040
rect 13688 3028 13695 3040
rect 13503 2976 13509 3028
rect 13689 2976 13695 3028
rect 13503 2963 13510 2976
rect 13688 2963 13695 2976
rect 13503 2911 13509 2963
rect 13689 2911 13695 2963
rect 13503 2898 13510 2911
rect 13688 2898 13695 2911
rect 13503 2846 13509 2898
rect 13689 2846 13695 2898
rect 13503 2833 13510 2846
rect 13688 2833 13695 2846
rect 13503 2781 13509 2833
rect 13689 2781 13695 2833
rect 13503 2768 13510 2781
rect 13688 2768 13695 2781
rect 13503 2716 13509 2768
rect 13689 2716 13695 2768
rect 13503 2703 13510 2716
rect 13688 2703 13695 2716
rect 13503 2651 13509 2703
rect 13689 2651 13695 2703
rect 13503 2638 13510 2651
rect 13688 2638 13695 2651
rect 13503 2586 13509 2638
rect 13689 2586 13695 2638
rect 13503 2574 13510 2586
rect 13688 2574 13695 2586
rect 13503 2573 13695 2574
rect 13503 2521 13509 2573
rect 13561 2521 13573 2573
rect 13625 2521 13637 2573
rect 13689 2521 13695 2573
rect 13503 2508 13510 2521
rect 13544 2508 13582 2521
rect 13616 2508 13654 2521
rect 13688 2508 13695 2521
rect 13503 2456 13509 2508
rect 13561 2456 13573 2508
rect 13625 2456 13637 2508
rect 13689 2456 13695 2508
rect 13503 2449 13582 2456
rect 13616 2449 13695 2456
rect 13503 2443 13510 2449
rect 13688 2443 13695 2449
rect 13503 2391 13509 2443
rect 13689 2391 13695 2443
rect 13503 2378 13510 2391
rect 13688 2378 13695 2391
rect 13503 2326 13509 2378
rect 13689 2326 13695 2378
rect 13503 2313 13510 2326
rect 13688 2313 13695 2326
rect 13503 2261 13509 2313
rect 13689 2261 13695 2313
rect 13503 2248 13510 2261
rect 13688 2248 13695 2261
rect 13503 2196 13509 2248
rect 13689 2196 13695 2248
rect 13503 2183 13510 2196
rect 13688 2183 13695 2196
rect 13503 2131 13509 2183
rect 13689 2131 13695 2183
rect 13503 2118 13510 2131
rect 13688 2118 13695 2131
rect 13503 2066 13509 2118
rect 13689 2066 13695 2118
rect 13503 2053 13510 2066
rect 13688 2053 13695 2066
rect 13503 2001 13509 2053
rect 13689 2001 13695 2053
rect 13503 1987 13510 2001
rect 13688 1987 13695 2001
rect 13503 1935 13509 1987
rect 13689 1935 13695 1987
rect 13503 1921 13510 1935
rect 13688 1921 13695 1935
rect 13503 1869 13509 1921
rect 13689 1869 13695 1921
rect 13503 1855 13510 1869
rect 13688 1855 13695 1869
rect 13503 1803 13509 1855
rect 13689 1803 13695 1855
rect 13503 1789 13510 1803
rect 13688 1789 13695 1803
rect 13503 1737 13509 1789
rect 13689 1737 13695 1789
rect 13503 1723 13510 1737
rect 13688 1723 13695 1737
rect 13503 1671 13509 1723
rect 13689 1671 13695 1723
rect 13503 1657 13510 1671
rect 13688 1657 13695 1671
rect 13503 1605 13509 1657
rect 13689 1605 13695 1657
rect 13503 1591 13510 1605
rect 13688 1591 13695 1605
rect 13503 1539 13509 1591
rect 13689 1539 13695 1591
rect 13503 1525 13510 1539
rect 13688 1525 13695 1539
rect 13503 1473 13509 1525
rect 13561 1473 13573 1491
rect 13625 1473 13637 1491
rect 13689 1473 13695 1525
rect 13503 1467 13695 1473
rect 14000 4068 14226 4074
rect 14000 4062 14037 4068
rect 14089 4062 14105 4068
rect 14000 2732 14006 4062
rect 14157 4016 14173 4068
rect 14225 4016 14226 4068
rect 14112 4003 14226 4016
rect 14157 3951 14173 4003
rect 14225 3951 14226 4003
rect 14112 3938 14226 3951
rect 14157 3886 14173 3938
rect 14225 3886 14226 3938
rect 14112 3873 14226 3886
rect 14157 3821 14173 3873
rect 14225 3821 14226 3873
rect 14112 3808 14226 3821
rect 14157 3756 14173 3808
rect 14225 3756 14226 3808
rect 14112 3743 14226 3756
rect 14157 3691 14173 3743
rect 14225 3691 14226 3743
rect 14112 3678 14226 3691
rect 14157 3626 14173 3678
rect 14225 3626 14226 3678
rect 14112 3613 14226 3626
rect 14157 3561 14173 3613
rect 14225 3561 14226 3613
rect 14112 3548 14226 3561
rect 14157 3496 14173 3548
rect 14225 3496 14226 3548
rect 14112 3483 14226 3496
rect 14157 3431 14173 3483
rect 14225 3431 14226 3483
rect 14112 3418 14226 3431
rect 14157 3366 14173 3418
rect 14225 3366 14226 3418
rect 14112 3353 14226 3366
rect 14157 3301 14173 3353
rect 14225 3301 14226 3353
rect 14112 3288 14226 3301
rect 14157 3236 14173 3288
rect 14225 3236 14226 3288
rect 14112 3223 14226 3236
rect 14157 3171 14173 3223
rect 14225 3171 14226 3223
rect 14112 3158 14226 3171
rect 14157 3106 14173 3158
rect 14225 3106 14226 3158
rect 14112 3093 14226 3106
rect 14157 3041 14173 3093
rect 14225 3041 14226 3093
rect 14112 3028 14226 3041
rect 14157 2976 14173 3028
rect 14225 2976 14226 3028
rect 14112 2963 14226 2976
rect 14157 2911 14173 2963
rect 14225 2911 14226 2963
rect 14112 2898 14226 2911
rect 14157 2846 14173 2898
rect 14225 2846 14226 2898
rect 14112 2833 14226 2846
rect 14157 2781 14173 2833
rect 14225 2781 14226 2833
rect 14112 2768 14226 2781
rect 14000 2716 14037 2732
rect 14089 2716 14105 2732
rect 14157 2716 14173 2768
rect 14225 2716 14226 2768
rect 14000 2703 14226 2716
rect 14000 2693 14037 2703
rect 14089 2693 14105 2703
rect 14000 2659 14006 2693
rect 14000 2651 14037 2659
rect 14089 2651 14105 2659
rect 14157 2651 14173 2703
rect 14225 2651 14226 2703
rect 14000 2638 14226 2651
rect 14000 2620 14037 2638
rect 14089 2620 14105 2638
rect 14000 2586 14006 2620
rect 14157 2586 14173 2638
rect 14225 2586 14226 2638
rect 14000 2573 14226 2586
rect 14000 2547 14037 2573
rect 14089 2547 14105 2573
rect 14000 2513 14006 2547
rect 14157 2521 14173 2573
rect 14225 2521 14226 2573
rect 14040 2513 14078 2521
rect 14112 2513 14226 2521
rect 14000 2508 14226 2513
rect 14000 2474 14037 2508
rect 14089 2474 14105 2508
rect 14000 2440 14006 2474
rect 14157 2456 14173 2508
rect 14225 2456 14226 2508
rect 14040 2443 14078 2456
rect 14112 2443 14226 2456
rect 14000 2401 14037 2440
rect 14089 2401 14105 2440
rect 14000 2367 14006 2401
rect 14157 2391 14173 2443
rect 14225 2391 14226 2443
rect 14040 2378 14078 2391
rect 14112 2378 14226 2391
rect 14000 2328 14037 2367
rect 14089 2328 14105 2367
rect 14000 2294 14006 2328
rect 14157 2326 14173 2378
rect 14225 2326 14226 2378
rect 14040 2313 14078 2326
rect 14112 2313 14226 2326
rect 14000 2261 14037 2294
rect 14089 2261 14105 2294
rect 14157 2261 14173 2313
rect 14225 2261 14226 2313
rect 14000 2255 14226 2261
rect 14000 2221 14006 2255
rect 14040 2248 14078 2255
rect 14112 2248 14226 2255
rect 14000 2196 14037 2221
rect 14089 2196 14105 2221
rect 14157 2196 14173 2248
rect 14225 2196 14226 2248
rect 14000 2183 14226 2196
rect 14000 2182 14037 2183
rect 14089 2182 14105 2183
rect 14000 2148 14006 2182
rect 14000 2131 14037 2148
rect 14089 2131 14105 2148
rect 14157 2131 14173 2183
rect 14225 2131 14226 2183
rect 14000 2118 14226 2131
rect 14000 2109 14037 2118
rect 14089 2109 14105 2118
rect 14000 2075 14006 2109
rect 14000 2066 14037 2075
rect 14089 2066 14105 2075
rect 14157 2066 14173 2118
rect 14225 2066 14226 2118
rect 14000 2053 14226 2066
rect 14000 2036 14037 2053
rect 14089 2036 14105 2053
rect 14000 2002 14006 2036
rect 14000 2001 14037 2002
rect 14089 2001 14105 2002
rect 14157 2001 14173 2053
rect 14225 2001 14226 2053
rect 14000 1987 14226 2001
rect 14000 1963 14037 1987
rect 14089 1963 14105 1987
rect 14000 1929 14006 1963
rect 14157 1935 14173 1987
rect 14225 1935 14226 1987
rect 14040 1929 14078 1935
rect 14112 1929 14226 1935
rect 14000 1921 14226 1929
rect 14000 1890 14037 1921
rect 14089 1890 14105 1921
rect 14000 1856 14006 1890
rect 14157 1869 14173 1921
rect 14225 1869 14226 1921
rect 14040 1856 14078 1869
rect 14112 1856 14226 1869
rect 14000 1855 14226 1856
rect 14000 1817 14037 1855
rect 14089 1817 14105 1855
rect 14000 1783 14006 1817
rect 14157 1803 14173 1855
rect 14225 1803 14226 1855
rect 14040 1789 14078 1803
rect 14112 1789 14226 1803
rect 14000 1744 14037 1783
rect 14089 1744 14105 1783
rect 14000 1710 14006 1744
rect 14157 1737 14173 1789
rect 14225 1737 14226 1789
rect 14040 1723 14078 1737
rect 14112 1723 14226 1737
rect 14000 1671 14037 1710
rect 14089 1671 14105 1710
rect 14157 1671 14173 1723
rect 14225 1671 14226 1723
rect 14000 1637 14006 1671
rect 14040 1657 14078 1671
rect 14112 1657 14226 1671
rect 14000 1605 14037 1637
rect 14089 1605 14105 1637
rect 14157 1605 14173 1657
rect 14225 1605 14226 1657
rect 14000 1598 14226 1605
rect 14000 1564 14006 1598
rect 14040 1591 14078 1598
rect 14112 1591 14226 1598
rect 14000 1539 14037 1564
rect 14089 1539 14105 1564
rect 14157 1539 14173 1591
rect 14225 1539 14226 1591
rect 14000 1525 14226 1539
rect 14000 1491 14006 1525
rect 14000 1473 14037 1491
rect 14089 1473 14105 1491
rect 14157 1473 14173 1525
rect 14225 1473 14226 1525
rect 14000 1467 14226 1473
rect 14400 4068 14510 4083
rect 14544 4068 14582 4086
rect 14616 4068 14628 4086
rect 14452 4044 14488 4068
rect 14544 4052 14576 4068
rect 14465 4016 14488 4044
rect 14540 4016 14576 4052
rect 14400 4010 14431 4016
rect 14465 4013 14628 4016
rect 14465 4010 14510 4013
rect 14400 4003 14510 4010
rect 14544 4003 14582 4013
rect 14616 4003 14628 4013
rect 14452 3971 14488 4003
rect 14544 3979 14576 4003
rect 14465 3951 14488 3971
rect 14540 3951 14576 3979
rect 14400 3938 14431 3951
rect 14465 3940 14628 3951
rect 14465 3938 14510 3940
rect 14544 3938 14582 3940
rect 14616 3938 14628 3940
rect 14465 3937 14488 3938
rect 14452 3898 14488 3937
rect 14544 3906 14576 3938
rect 14465 3886 14488 3898
rect 14540 3886 14576 3906
rect 14400 3873 14431 3886
rect 14465 3873 14628 3886
rect 14465 3864 14488 3873
rect 14540 3867 14576 3873
rect 14452 3825 14488 3864
rect 14544 3833 14576 3867
rect 14465 3821 14488 3825
rect 14540 3821 14576 3833
rect 14400 3808 14431 3821
rect 14465 3808 14628 3821
rect 14465 3791 14488 3808
rect 14540 3794 14576 3808
rect 14452 3756 14488 3791
rect 14544 3760 14576 3794
rect 14540 3756 14576 3760
rect 14400 3752 14628 3756
rect 14400 3743 14431 3752
rect 14465 3743 14628 3752
rect 14465 3718 14488 3743
rect 14540 3721 14576 3743
rect 14452 3691 14488 3718
rect 14544 3691 14576 3721
rect 14400 3687 14510 3691
rect 14544 3687 14582 3691
rect 14616 3687 14628 3691
rect 14400 3679 14628 3687
rect 14400 3678 14431 3679
rect 14465 3678 14628 3679
rect 14465 3645 14488 3678
rect 14540 3648 14576 3678
rect 14452 3626 14488 3645
rect 14544 3626 14576 3648
rect 14400 3614 14510 3626
rect 14544 3614 14582 3626
rect 14616 3614 14628 3626
rect 14400 3613 14628 3614
rect 14452 3606 14488 3613
rect 14465 3572 14488 3606
rect 14540 3575 14576 3613
rect 14452 3561 14488 3572
rect 14544 3561 14576 3575
rect 14400 3548 14510 3561
rect 14544 3548 14582 3561
rect 14616 3548 14628 3561
rect 14452 3533 14488 3548
rect 14544 3541 14576 3548
rect 14465 3499 14488 3533
rect 14540 3502 14576 3541
rect 14452 3496 14488 3499
rect 14544 3496 14576 3502
rect 14400 3483 14510 3496
rect 14544 3483 14582 3496
rect 14616 3483 14628 3496
rect 14452 3460 14488 3483
rect 14544 3468 14576 3483
rect 14465 3431 14488 3460
rect 14540 3431 14576 3468
rect 14400 3426 14431 3431
rect 14465 3429 14628 3431
rect 14465 3426 14510 3429
rect 14400 3418 14510 3426
rect 14544 3418 14582 3429
rect 14616 3418 14628 3429
rect 14452 3387 14488 3418
rect 14544 3395 14576 3418
rect 14465 3366 14488 3387
rect 14540 3366 14576 3395
rect 14400 3353 14431 3366
rect 14465 3356 14628 3366
rect 14465 3353 14510 3356
rect 14544 3353 14582 3356
rect 14616 3353 14628 3356
rect 14452 3314 14488 3353
rect 14544 3322 14576 3353
rect 14465 3301 14488 3314
rect 14540 3301 14576 3322
rect 14400 3288 14431 3301
rect 14465 3288 14628 3301
rect 14465 3280 14488 3288
rect 14540 3283 14576 3288
rect 14452 3241 14488 3280
rect 14544 3249 14576 3283
rect 14465 3236 14488 3241
rect 14540 3236 14576 3249
rect 14400 3223 14431 3236
rect 14465 3223 14628 3236
rect 14465 3207 14488 3223
rect 14540 3210 14576 3223
rect 14452 3171 14488 3207
rect 14544 3176 14576 3210
rect 14540 3171 14576 3176
rect 14400 3168 14628 3171
rect 14400 3158 14431 3168
rect 14465 3158 14628 3168
rect 14465 3134 14488 3158
rect 14540 3137 14576 3158
rect 14452 3106 14488 3134
rect 14544 3106 14576 3137
rect 14400 3103 14510 3106
rect 14544 3103 14582 3106
rect 14616 3103 14628 3106
rect 14400 3095 14628 3103
rect 14400 3093 14431 3095
rect 14465 3093 14628 3095
rect 14465 3061 14488 3093
rect 14540 3064 14576 3093
rect 14452 3041 14488 3061
rect 14544 3041 14576 3064
rect 14400 3030 14510 3041
rect 14544 3030 14582 3041
rect 14616 3030 14628 3041
rect 14400 3028 14628 3030
rect 14452 3022 14488 3028
rect 14465 2988 14488 3022
rect 14540 2991 14576 3028
rect 14452 2976 14488 2988
rect 14544 2976 14576 2991
rect 14400 2963 14510 2976
rect 14544 2963 14582 2976
rect 14616 2963 14628 2976
rect 14452 2949 14488 2963
rect 14544 2957 14576 2963
rect 14465 2915 14488 2949
rect 14540 2918 14576 2957
rect 14452 2911 14488 2915
rect 14544 2911 14576 2918
rect 14400 2898 14510 2911
rect 14544 2898 14582 2911
rect 14616 2898 14628 2911
rect 14452 2876 14488 2898
rect 14544 2884 14576 2898
rect 14465 2846 14488 2876
rect 14540 2846 14576 2884
rect 14400 2842 14431 2846
rect 14465 2845 14628 2846
rect 14465 2842 14510 2845
rect 14400 2833 14510 2842
rect 14544 2833 14582 2845
rect 14616 2833 14628 2845
rect 14452 2803 14488 2833
rect 14544 2811 14576 2833
rect 14465 2781 14488 2803
rect 14540 2781 14576 2811
rect 14400 2769 14431 2781
rect 14465 2772 14628 2781
rect 14465 2769 14510 2772
rect 14400 2768 14510 2769
rect 14544 2768 14582 2772
rect 14616 2768 14628 2772
rect 14452 2730 14488 2768
rect 14544 2738 14576 2768
rect 14465 2716 14488 2730
rect 14540 2716 14576 2738
rect 14400 2703 14431 2716
rect 14465 2703 14628 2716
rect 14465 2696 14488 2703
rect 14540 2699 14576 2703
rect 14452 2657 14488 2696
rect 14544 2665 14576 2699
rect 14465 2651 14488 2657
rect 14540 2651 14576 2665
rect 14400 2638 14431 2651
rect 14465 2638 14628 2651
rect 14465 2623 14488 2638
rect 14540 2626 14576 2638
rect 14452 2586 14488 2623
rect 14544 2592 14576 2626
rect 14540 2586 14576 2592
rect 14400 2584 14628 2586
rect 14400 2573 14431 2584
rect 14465 2573 14628 2584
rect 14465 2550 14488 2573
rect 14540 2553 14576 2573
rect 14452 2521 14488 2550
rect 14544 2521 14576 2553
rect 14400 2519 14510 2521
rect 14544 2519 14582 2521
rect 14616 2519 14628 2521
rect 14400 2511 14628 2519
rect 14400 2508 14431 2511
rect 14465 2508 14628 2511
rect 14465 2477 14488 2508
rect 14540 2480 14576 2508
rect 14452 2456 14488 2477
rect 14544 2456 14576 2480
rect 14400 2446 14510 2456
rect 14544 2446 14582 2456
rect 14616 2446 14628 2456
rect 14400 2443 14628 2446
rect 14452 2438 14488 2443
rect 14465 2404 14488 2438
rect 14540 2407 14576 2443
rect 14452 2391 14488 2404
rect 14544 2391 14576 2407
rect 14400 2378 14510 2391
rect 14544 2378 14582 2391
rect 14616 2378 14628 2391
rect 14452 2365 14488 2378
rect 14544 2373 14576 2378
rect 14465 2331 14488 2365
rect 14540 2334 14576 2373
rect 14452 2326 14488 2331
rect 14544 2326 14576 2334
rect 14400 2313 14510 2326
rect 14544 2313 14582 2326
rect 14616 2313 14628 2326
rect 14452 2292 14488 2313
rect 14544 2300 14576 2313
rect 14465 2261 14488 2292
rect 14540 2261 14576 2300
rect 14400 2258 14431 2261
rect 14465 2260 14628 2261
rect 14465 2258 14510 2260
rect 14400 2248 14510 2258
rect 14544 2248 14582 2260
rect 14616 2248 14628 2260
rect 14452 2219 14488 2248
rect 14544 2226 14576 2248
rect 14465 2196 14488 2219
rect 14540 2196 14576 2226
rect 14400 2185 14431 2196
rect 14465 2186 14628 2196
rect 14465 2185 14510 2186
rect 14400 2183 14510 2185
rect 14544 2183 14582 2186
rect 14616 2183 14628 2186
rect 14452 2146 14488 2183
rect 14544 2152 14576 2183
rect 14465 2131 14488 2146
rect 14540 2131 14576 2152
rect 14400 2118 14431 2131
rect 14465 2118 14628 2131
rect 14465 2112 14488 2118
rect 14540 2112 14576 2118
rect 14452 2073 14488 2112
rect 14544 2078 14576 2112
rect 14465 2066 14488 2073
rect 14540 2066 14576 2078
rect 14400 2053 14431 2066
rect 14465 2053 14628 2066
rect 14465 2039 14488 2053
rect 14452 2001 14488 2039
rect 14540 2038 14576 2053
rect 14544 2004 14576 2038
rect 14540 2001 14576 2004
rect 14400 2000 14628 2001
rect 14400 1987 14431 2000
rect 14465 1987 14628 2000
rect 14465 1966 14488 1987
rect 14452 1935 14488 1966
rect 14540 1964 14576 1987
rect 14544 1935 14576 1964
rect 14400 1930 14510 1935
rect 14544 1930 14582 1935
rect 14616 1930 14628 1935
rect 14400 1927 14628 1930
rect 14400 1921 14431 1927
rect 14465 1921 14628 1927
rect 14465 1893 14488 1921
rect 14452 1869 14488 1893
rect 14540 1890 14576 1921
rect 14544 1869 14576 1890
rect 14400 1856 14510 1869
rect 14544 1856 14582 1869
rect 14616 1856 14628 1869
rect 14400 1855 14628 1856
rect 14452 1854 14488 1855
rect 14465 1820 14488 1854
rect 14452 1803 14488 1820
rect 14540 1816 14576 1855
rect 14544 1803 14576 1816
rect 14400 1789 14510 1803
rect 14544 1789 14582 1803
rect 14616 1789 14628 1803
rect 14452 1781 14488 1789
rect 14544 1782 14576 1789
rect 14465 1747 14488 1781
rect 14452 1737 14488 1747
rect 14540 1742 14576 1782
rect 14544 1737 14576 1742
rect 14400 1723 14510 1737
rect 14544 1723 14582 1737
rect 14616 1723 14628 1737
rect 14452 1708 14488 1723
rect 14544 1708 14576 1723
rect 14465 1674 14488 1708
rect 14452 1671 14488 1674
rect 14540 1671 14576 1708
rect 14400 1668 14628 1671
rect 14400 1657 14510 1668
rect 14544 1657 14582 1668
rect 14616 1657 14628 1668
rect 14452 1635 14488 1657
rect 14465 1605 14488 1635
rect 14544 1634 14576 1657
rect 14540 1605 14576 1634
rect 14400 1601 14431 1605
rect 14465 1601 14628 1605
rect 14400 1594 14628 1601
rect 14400 1591 14510 1594
rect 14544 1591 14582 1594
rect 14616 1591 14628 1594
rect 14452 1562 14488 1591
rect 14465 1539 14488 1562
rect 14544 1560 14576 1591
rect 14540 1539 14576 1560
rect 14400 1528 14431 1539
rect 14465 1528 14628 1539
rect 14400 1525 14628 1528
rect 14452 1489 14488 1525
rect 14540 1520 14576 1525
rect 14465 1473 14488 1489
rect 14544 1486 14576 1520
rect 14540 1473 14576 1486
rect 575 1419 803 1455
rect 575 1385 587 1419
rect 621 1385 659 1419
rect 693 1416 803 1419
rect 693 1385 733 1416
rect 575 1382 733 1385
rect 767 1382 803 1416
rect 575 1342 803 1382
rect 575 1330 733 1342
rect 575 1296 587 1330
rect 621 1296 659 1330
rect 693 1308 733 1330
rect 767 1308 803 1342
rect 14400 1455 14431 1473
rect 14465 1455 14628 1473
rect 14400 1446 14628 1455
rect 14400 1416 14510 1446
rect 14400 1382 14431 1416
rect 14465 1412 14510 1416
rect 14544 1412 14582 1446
rect 14616 1412 14628 1446
rect 14465 1382 14628 1412
rect 14400 1372 14628 1382
rect 14400 1342 14510 1372
tri 803 1308 832 1337 sw
tri 14390 1308 14400 1318 se
rect 14400 1308 14431 1342
rect 14465 1338 14510 1342
rect 14544 1338 14582 1372
rect 14616 1338 14628 1372
rect 14465 1308 14628 1338
rect 693 1298 832 1308
tri 832 1298 842 1308 sw
tri 14380 1298 14390 1308 se
rect 14390 1298 14628 1308
rect 693 1296 842 1298
rect 575 1268 842 1296
tri 842 1268 872 1298 sw
tri 14350 1268 14380 1298 se
rect 14380 1268 14510 1298
rect 575 1241 733 1268
rect 575 1207 587 1241
rect 621 1207 659 1241
rect 693 1234 733 1241
rect 767 1234 872 1268
tri 872 1234 906 1268 sw
tri 14316 1234 14350 1268 se
rect 14350 1234 14431 1268
rect 14465 1264 14510 1268
rect 14544 1264 14582 1298
rect 14616 1264 14628 1298
rect 14465 1234 14628 1264
rect 693 1224 906 1234
tri 906 1224 916 1234 sw
tri 14306 1224 14316 1234 se
rect 14316 1224 14628 1234
rect 693 1207 916 1224
rect 575 1194 916 1207
tri 916 1194 946 1224 sw
tri 14276 1194 14306 1224 se
rect 14306 1194 14510 1224
rect 575 1160 733 1194
rect 767 1160 946 1194
tri 946 1160 980 1194 sw
tri 14242 1160 14276 1194 se
rect 14276 1160 14431 1194
rect 14465 1190 14510 1194
rect 14544 1190 14582 1224
rect 14616 1190 14628 1224
rect 14465 1160 14628 1190
rect 575 1141 980 1160
tri 980 1141 999 1160 sw
tri 14230 1148 14242 1160 se
rect 14242 1148 14628 1160
tri 14223 1141 14230 1148 se
rect 14230 1141 14628 1148
rect 575 1128 999 1141
tri 999 1128 1012 1141 sw
tri 14210 1128 14223 1141 se
rect 14223 1128 14628 1141
rect 575 1116 14628 1128
rect 575 1114 767 1116
tri 575 1082 607 1114 ne
rect 607 1082 767 1114
rect 801 1082 840 1116
rect 874 1082 913 1116
rect 947 1082 986 1116
rect 1020 1082 1059 1116
rect 1093 1082 1132 1116
rect 1166 1082 1205 1116
rect 1239 1082 1278 1116
rect 1312 1082 1351 1116
rect 1385 1082 1424 1116
rect 1458 1082 1497 1116
rect 1531 1082 1570 1116
rect 1604 1082 1643 1116
rect 1677 1082 1716 1116
rect 1750 1082 1789 1116
rect 1823 1082 1862 1116
rect 1896 1082 1935 1116
rect 1969 1082 2008 1116
rect 2042 1082 2081 1116
rect 2115 1082 2154 1116
rect 2188 1082 2227 1116
rect 2261 1082 2300 1116
rect 2334 1082 2373 1116
rect 2407 1082 2446 1116
rect 2480 1082 2519 1116
rect 2553 1082 2592 1116
rect 2626 1082 2665 1116
rect 2699 1082 2738 1116
rect 267 1054 409 1055
rect 59 1016 409 1054
tri 607 1044 645 1082 ne
rect 645 1044 2738 1082
rect 59 982 233 1016
rect 267 982 369 1016
rect 403 982 409 1016
tri 645 1010 679 1044 ne
rect 679 1010 767 1044
rect 801 1010 840 1044
rect 874 1010 913 1044
rect 947 1010 986 1044
rect 1020 1010 1059 1044
rect 1093 1010 1132 1044
rect 1166 1010 1205 1044
rect 1239 1010 1278 1044
rect 1312 1010 1351 1044
rect 1385 1010 1424 1044
rect 1458 1010 1497 1044
rect 1531 1010 1570 1044
rect 1604 1010 1643 1044
rect 1677 1010 1716 1044
rect 1750 1010 1789 1044
rect 1823 1010 1862 1044
rect 1896 1010 1935 1044
rect 1969 1010 2008 1044
rect 2042 1010 2081 1044
rect 2115 1010 2154 1044
rect 2188 1010 2227 1044
rect 2261 1010 2300 1044
rect 2334 1010 2373 1044
rect 2407 1010 2446 1044
rect 2480 1010 2519 1044
rect 2553 1010 2592 1044
rect 2626 1010 2665 1044
rect 2699 1010 2738 1044
rect 14436 1114 14628 1116
rect 14436 1111 14625 1114
tri 14625 1111 14628 1114 nw
rect 14818 4819 15117 4849
rect 14818 4785 14833 4819
rect 14867 4811 15117 4819
rect 14867 4785 14969 4811
rect 14818 4777 14969 4785
rect 15003 4777 15117 4811
rect 14818 4747 15117 4777
rect 14818 4713 14833 4747
rect 14867 4739 15117 4747
rect 14867 4713 14969 4739
rect 14818 4705 14969 4713
rect 15003 4705 15117 4739
rect 14818 4675 15117 4705
rect 14818 4641 14833 4675
rect 14867 4667 15117 4675
rect 14867 4641 14969 4667
rect 14818 4633 14969 4641
rect 15003 4633 15117 4667
rect 14818 4603 15117 4633
rect 14818 4569 14833 4603
rect 14867 4595 15117 4603
rect 14867 4569 14969 4595
rect 14818 4561 14969 4569
rect 15003 4561 15117 4595
rect 14818 4531 15117 4561
rect 14818 4497 14833 4531
rect 14867 4523 15117 4531
rect 14867 4497 14969 4523
rect 14818 4489 14969 4497
rect 15003 4489 15117 4523
rect 14818 4459 15117 4489
rect 14818 4425 14833 4459
rect 14867 4451 15117 4459
rect 14867 4425 14969 4451
rect 14818 4417 14969 4425
rect 15003 4417 15117 4451
rect 14818 4387 15117 4417
rect 14818 4353 14833 4387
rect 14867 4379 15117 4387
rect 14867 4353 14969 4379
rect 14818 4345 14969 4353
rect 15003 4345 15117 4379
rect 14818 4314 15117 4345
rect 14818 4280 14833 4314
rect 14867 4307 15117 4314
rect 14867 4280 14969 4307
rect 14818 4273 14969 4280
rect 15003 4273 15117 4307
rect 14818 4241 15117 4273
rect 14818 4207 14833 4241
rect 14867 4235 15117 4241
rect 14867 4207 14969 4235
rect 14818 4201 14969 4207
rect 15003 4201 15117 4235
rect 14818 4168 15117 4201
rect 14818 4134 14833 4168
rect 14867 4163 15117 4168
rect 14867 4134 14969 4163
rect 14818 4129 14969 4134
rect 15003 4129 15117 4163
rect 14818 4095 15117 4129
rect 14818 4061 14833 4095
rect 14867 4091 15117 4095
rect 14867 4061 14969 4091
rect 14818 4057 14969 4061
rect 15003 4057 15117 4091
rect 14818 4022 15117 4057
rect 14818 3988 14833 4022
rect 14867 4019 15117 4022
rect 14867 3988 14969 4019
rect 14818 3985 14969 3988
rect 15003 3985 15117 4019
rect 14818 3949 15117 3985
rect 14818 3915 14833 3949
rect 14867 3947 15117 3949
rect 14867 3915 14969 3947
rect 14818 3913 14969 3915
rect 15003 3913 15117 3947
rect 14818 3876 15117 3913
rect 14818 3842 14833 3876
rect 14867 3875 15117 3876
rect 14867 3842 14969 3875
rect 14818 3841 14969 3842
rect 15003 3841 15117 3875
rect 14818 3803 15117 3841
rect 14818 3769 14833 3803
rect 14867 3769 14969 3803
rect 15003 3769 15117 3803
rect 14818 3731 15117 3769
rect 14818 3730 14969 3731
rect 14818 3696 14833 3730
rect 14867 3697 14969 3730
rect 15003 3697 15117 3731
rect 14867 3696 15117 3697
rect 14818 3659 15117 3696
rect 14818 3657 14969 3659
rect 14818 3623 14833 3657
rect 14867 3625 14969 3657
rect 15003 3625 15117 3659
rect 14867 3623 15117 3625
rect 14818 3587 15117 3623
rect 14818 3584 14969 3587
rect 14818 3550 14833 3584
rect 14867 3553 14969 3584
rect 15003 3553 15117 3587
rect 14867 3550 15117 3553
rect 14818 3515 15117 3550
rect 14818 3511 14969 3515
rect 14818 3477 14833 3511
rect 14867 3481 14969 3511
rect 15003 3481 15117 3515
rect 14867 3477 15117 3481
rect 14818 3443 15117 3477
rect 14818 3438 14969 3443
rect 14818 3404 14833 3438
rect 14867 3409 14969 3438
rect 15003 3409 15117 3443
rect 14867 3404 15117 3409
rect 14818 3371 15117 3404
rect 14818 3365 14969 3371
rect 14818 3331 14833 3365
rect 14867 3337 14969 3365
rect 15003 3337 15117 3371
rect 14867 3331 15117 3337
rect 14818 3299 15117 3331
rect 14818 3292 14969 3299
rect 14818 3258 14833 3292
rect 14867 3265 14969 3292
rect 15003 3265 15117 3299
rect 14867 3258 15117 3265
rect 14818 3227 15117 3258
rect 14818 3219 14969 3227
rect 14818 3185 14833 3219
rect 14867 3193 14969 3219
rect 15003 3193 15117 3227
rect 14867 3185 15117 3193
rect 14818 3155 15117 3185
rect 14818 3146 14969 3155
rect 14818 3112 14833 3146
rect 14867 3121 14969 3146
rect 15003 3121 15117 3155
rect 14867 3112 15117 3121
rect 14818 3082 15117 3112
rect 14818 3073 14969 3082
rect 14818 3039 14833 3073
rect 14867 3048 14969 3073
rect 15003 3048 15117 3082
rect 14867 3039 15117 3048
rect 14818 3009 15117 3039
rect 14818 3000 14969 3009
rect 14818 2966 14833 3000
rect 14867 2975 14969 3000
rect 15003 2975 15117 3009
rect 14867 2966 15117 2975
rect 14818 2936 15117 2966
rect 14818 2927 14969 2936
rect 14818 2893 14833 2927
rect 14867 2902 14969 2927
rect 15003 2902 15117 2936
rect 14867 2893 15117 2902
rect 14818 2863 15117 2893
rect 14818 2854 14969 2863
rect 14818 2820 14833 2854
rect 14867 2829 14969 2854
rect 15003 2829 15117 2863
rect 14867 2820 15117 2829
rect 14818 2790 15117 2820
rect 14818 2781 14969 2790
rect 14818 2747 14833 2781
rect 14867 2756 14969 2781
rect 15003 2756 15117 2790
rect 14867 2747 15117 2756
rect 14818 2717 15117 2747
rect 14818 2708 14969 2717
rect 14818 2674 14833 2708
rect 14867 2683 14969 2708
rect 15003 2683 15117 2717
rect 14867 2674 15117 2683
rect 14818 2644 15117 2674
rect 14818 2635 14969 2644
rect 14818 2601 14833 2635
rect 14867 2610 14969 2635
rect 15003 2610 15117 2644
rect 14867 2601 15117 2610
rect 14818 2571 15117 2601
rect 14818 2562 14969 2571
rect 14818 2528 14833 2562
rect 14867 2537 14969 2562
rect 15003 2537 15117 2571
rect 14867 2528 15117 2537
rect 14818 2498 15117 2528
rect 14818 2489 14969 2498
rect 14818 2455 14833 2489
rect 14867 2464 14969 2489
rect 15003 2464 15117 2498
rect 14867 2455 15117 2464
rect 14818 2425 15117 2455
rect 14818 2416 14969 2425
rect 14818 2382 14833 2416
rect 14867 2391 14969 2416
rect 15003 2391 15117 2425
rect 14867 2382 15117 2391
rect 14818 2352 15117 2382
rect 14818 2343 14969 2352
rect 14818 2309 14833 2343
rect 14867 2318 14969 2343
rect 15003 2318 15117 2352
rect 14867 2309 15117 2318
rect 14818 2279 15117 2309
rect 14818 2270 14969 2279
rect 14818 2236 14833 2270
rect 14867 2245 14969 2270
rect 15003 2245 15117 2279
rect 14867 2236 15117 2245
rect 14818 2206 15117 2236
rect 14818 2197 14969 2206
rect 14818 2163 14833 2197
rect 14867 2172 14969 2197
rect 15003 2172 15117 2206
rect 14867 2163 15117 2172
rect 14818 2133 15117 2163
rect 14818 2124 14969 2133
rect 14818 2090 14833 2124
rect 14867 2099 14969 2124
rect 15003 2099 15117 2133
rect 14867 2090 15117 2099
rect 14818 2060 15117 2090
rect 14818 2051 14969 2060
rect 14818 2017 14833 2051
rect 14867 2026 14969 2051
rect 15003 2026 15117 2060
rect 14867 2017 15117 2026
rect 14818 1987 15117 2017
rect 14818 1978 14969 1987
rect 14818 1944 14833 1978
rect 14867 1953 14969 1978
rect 15003 1953 15117 1987
rect 14867 1944 15117 1953
rect 14818 1914 15117 1944
rect 14818 1905 14969 1914
rect 14818 1871 14833 1905
rect 14867 1880 14969 1905
rect 15003 1880 15117 1914
rect 14867 1871 15117 1880
rect 14818 1841 15117 1871
rect 14818 1832 14969 1841
rect 14818 1798 14833 1832
rect 14867 1807 14969 1832
rect 15003 1807 15117 1841
rect 14867 1798 15117 1807
rect 14818 1768 15117 1798
rect 14818 1759 14969 1768
rect 14818 1725 14833 1759
rect 14867 1734 14969 1759
rect 15003 1734 15117 1768
rect 14867 1725 15117 1734
rect 14818 1695 15117 1725
rect 14818 1686 14969 1695
rect 14818 1652 14833 1686
rect 14867 1661 14969 1686
rect 15003 1661 15117 1695
rect 14867 1652 15117 1661
rect 14818 1622 15117 1652
rect 14818 1613 14969 1622
rect 14818 1579 14833 1613
rect 14867 1588 14969 1613
rect 15003 1588 15117 1622
rect 14867 1579 15117 1588
rect 14818 1549 15117 1579
rect 14818 1540 14969 1549
rect 14818 1506 14833 1540
rect 14867 1515 14969 1540
rect 15003 1515 15117 1549
rect 14867 1506 15117 1515
rect 14818 1476 15117 1506
rect 14818 1467 14969 1476
rect 14818 1433 14833 1467
rect 14867 1442 14969 1467
rect 15003 1442 15117 1476
rect 14867 1433 15117 1442
rect 14818 1403 15117 1433
rect 14818 1394 14969 1403
rect 14818 1360 14833 1394
rect 14867 1369 14969 1394
rect 15003 1369 15117 1403
rect 14867 1360 15117 1369
rect 14818 1330 15117 1360
rect 14818 1321 14969 1330
rect 14818 1287 14833 1321
rect 14867 1296 14969 1321
rect 15003 1296 15117 1330
rect 14867 1287 15117 1296
rect 14818 1257 15117 1287
rect 14818 1248 14969 1257
rect 14818 1214 14833 1248
rect 14867 1223 14969 1248
rect 15003 1223 15117 1257
rect 14867 1214 15117 1223
rect 14818 1184 15117 1214
rect 14818 1175 14969 1184
rect 14818 1141 14833 1175
rect 14867 1150 14969 1175
rect 15003 1150 15117 1184
rect 14867 1141 15117 1150
rect 14818 1111 15117 1141
rect 14436 1102 14616 1111
tri 14616 1102 14625 1111 nw
rect 14818 1102 14969 1111
rect 14436 1068 14582 1102
tri 14582 1068 14616 1102 nw
rect 14818 1068 14833 1102
rect 14867 1077 14969 1102
rect 15003 1077 15117 1111
rect 14867 1068 15117 1077
rect 14436 1038 14552 1068
tri 14552 1038 14582 1068 nw
rect 14818 1038 15117 1068
rect 14436 1029 14543 1038
tri 14543 1029 14552 1038 nw
rect 14818 1029 14969 1038
rect 14436 1010 14512 1029
tri 679 998 691 1010 ne
rect 691 998 14512 1010
tri 14512 998 14543 1029 nw
rect 59 944 409 982
rect 59 910 233 944
rect 267 910 369 944
rect 403 910 409 944
rect 59 872 409 910
rect 59 838 233 872
rect 267 838 369 872
rect 403 849 409 872
rect 14818 995 14833 1029
rect 14867 1004 14969 1029
rect 15003 1004 15117 1038
rect 14867 995 15117 1004
rect 14818 965 15117 995
rect 14818 956 14969 965
rect 14818 922 14833 956
rect 14867 931 14969 956
rect 15003 931 15117 965
rect 14867 922 15117 931
rect 14818 892 15117 922
rect 14818 883 14969 892
tri 409 849 420 860 sw
rect 14818 849 14833 883
rect 14867 858 14969 883
rect 15003 858 15117 892
rect 14867 849 15117 858
rect 403 838 420 849
tri 420 838 431 849 sw
rect 59 819 431 838
tri 431 819 450 838 sw
tri 14799 819 14818 838 se
rect 14818 819 15117 849
rect 59 810 450 819
tri 450 810 459 819 sw
tri 14790 810 14799 819 se
rect 14799 810 14969 819
rect 59 776 459 810
tri 459 776 493 810 sw
tri 14756 776 14790 810 se
rect 14790 776 14833 810
rect 14867 785 14969 810
rect 15003 785 15117 819
rect 14867 776 15117 785
rect 59 762 493 776
rect 59 728 212 762
rect 246 749 493 762
rect 246 728 348 749
rect 59 715 348 728
rect 382 746 493 749
tri 493 746 523 776 sw
tri 14726 746 14756 776 se
rect 14756 746 15117 776
rect 382 737 523 746
tri 523 737 532 746 sw
tri 14717 737 14726 746 se
rect 14726 737 14969 746
rect 382 715 532 737
rect 59 703 532 715
tri 532 703 566 737 sw
tri 14683 703 14717 737 se
rect 14717 703 14833 737
rect 14867 712 14969 737
rect 15003 712 15117 746
rect 14867 703 15117 712
rect 59 684 566 703
rect 59 650 212 684
rect 246 676 566 684
tri 566 676 593 703 sw
tri 14656 676 14683 703 se
rect 14683 676 15117 703
rect 246 673 15117 676
rect 246 664 14969 673
rect 246 650 348 664
rect 59 630 348 650
rect 382 630 421 664
rect 455 630 494 664
rect 528 630 567 664
rect 601 630 640 664
rect 674 630 713 664
rect 747 630 786 664
rect 820 630 859 664
rect 893 630 932 664
rect 966 630 1005 664
rect 1039 630 1078 664
rect 1112 630 1151 664
rect 1185 630 1224 664
rect 1258 630 1297 664
rect 1331 630 1369 664
rect 1403 630 1441 664
rect 1475 630 1513 664
rect 1547 630 1585 664
rect 1619 630 1657 664
rect 1691 630 1729 664
rect 1763 630 1801 664
rect 1835 630 1873 664
rect 1907 630 1945 664
rect 1979 630 2017 664
rect 2051 630 2089 664
rect 2123 630 2161 664
rect 2195 630 2233 664
rect 2267 630 2305 664
rect 2339 630 2377 664
rect 2411 630 2449 664
rect 2483 630 2521 664
rect 2555 630 2593 664
rect 2627 630 2665 664
rect 2699 630 2737 664
rect 2771 630 2809 664
rect 2843 630 2881 664
rect 2915 630 2953 664
rect 2987 630 3025 664
rect 3059 630 3097 664
rect 3131 630 3169 664
rect 3203 630 3241 664
rect 3275 630 3313 664
rect 3347 630 3385 664
rect 3419 630 3457 664
rect 3491 630 3529 664
rect 3563 630 3601 664
rect 3635 630 3673 664
rect 3707 630 3745 664
rect 3779 630 3817 664
rect 3851 630 3889 664
rect 3923 630 3961 664
rect 3995 630 4033 664
rect 4067 630 4105 664
rect 4139 630 4177 664
rect 4211 630 4249 664
rect 4283 630 4321 664
rect 4355 630 4393 664
rect 4427 630 4465 664
rect 4499 630 4537 664
rect 4571 630 4609 664
rect 4643 630 4681 664
rect 4715 630 4753 664
rect 4787 630 4825 664
rect 4859 630 4897 664
rect 4931 630 4969 664
rect 5003 630 5041 664
rect 5075 630 5113 664
rect 5147 630 5185 664
rect 5219 630 5257 664
rect 5291 630 5329 664
rect 5363 630 5401 664
rect 5435 630 5473 664
rect 5507 630 5545 664
rect 5579 630 5617 664
rect 5651 630 5689 664
rect 5723 630 5761 664
rect 5795 630 5833 664
rect 5867 630 5905 664
rect 5939 630 5977 664
rect 6011 630 6049 664
rect 6083 630 6121 664
rect 6155 630 6193 664
rect 6227 630 6265 664
rect 6299 630 6337 664
rect 6371 630 6409 664
rect 6443 630 6481 664
rect 6515 630 6553 664
rect 6587 630 6625 664
rect 6659 630 6697 664
rect 6731 630 6769 664
rect 6803 630 6841 664
rect 6875 630 6913 664
rect 6947 630 6985 664
rect 7019 630 7057 664
rect 7091 630 7129 664
rect 7163 630 7201 664
rect 7235 630 7273 664
rect 7307 630 7345 664
rect 7379 630 7417 664
rect 7451 630 7489 664
rect 7523 630 7561 664
rect 7595 630 7633 664
rect 7667 630 7705 664
rect 7739 630 7777 664
rect 7811 630 7849 664
rect 7883 630 7921 664
rect 7955 630 7993 664
rect 8027 630 8065 664
rect 8099 630 8137 664
rect 8171 630 8209 664
rect 8243 630 8281 664
rect 8315 630 8353 664
rect 8387 630 8425 664
rect 8459 630 8497 664
rect 8531 630 8569 664
rect 8603 630 8641 664
rect 8675 630 8713 664
rect 8747 630 8785 664
rect 8819 630 8857 664
rect 8891 630 8929 664
rect 8963 630 9001 664
rect 9035 630 9073 664
rect 9107 630 9145 664
rect 9179 630 9217 664
rect 9251 630 9289 664
rect 9323 630 9361 664
rect 9395 630 9433 664
rect 9467 630 9505 664
rect 9539 630 9577 664
rect 9611 630 9649 664
rect 9683 630 9721 664
rect 9755 630 9793 664
rect 9827 630 9865 664
rect 9899 630 9937 664
rect 9971 630 10009 664
rect 10043 630 10081 664
rect 10115 630 10153 664
rect 10187 630 10225 664
rect 10259 630 10297 664
rect 10331 630 10369 664
rect 10403 630 10441 664
rect 10475 630 10513 664
rect 10547 630 10585 664
rect 10619 630 10657 664
rect 10691 630 10729 664
rect 10763 630 10801 664
rect 10835 630 10873 664
rect 10907 630 10945 664
rect 10979 630 11017 664
rect 11051 630 11089 664
rect 11123 630 11161 664
rect 11195 630 11233 664
rect 11267 630 11305 664
rect 11339 630 11377 664
rect 11411 630 11449 664
rect 11483 630 11521 664
rect 11555 630 11593 664
rect 11627 630 11665 664
rect 11699 630 11737 664
rect 11771 630 11809 664
rect 11843 630 11881 664
rect 11915 630 11953 664
rect 11987 630 12025 664
rect 12059 630 12097 664
rect 12131 630 12169 664
rect 12203 630 12241 664
rect 12275 630 12313 664
rect 12347 630 12385 664
rect 12419 630 12457 664
rect 12491 630 12529 664
rect 12563 630 12601 664
rect 12635 630 12673 664
rect 12707 630 12745 664
rect 12779 630 12817 664
rect 12851 630 12889 664
rect 12923 630 12961 664
rect 12995 630 13033 664
rect 13067 630 13105 664
rect 13139 630 13177 664
rect 13211 630 13249 664
rect 13283 630 13321 664
rect 13355 630 13393 664
rect 13427 630 13465 664
rect 13499 630 13537 664
rect 13571 630 13609 664
rect 13643 630 13681 664
rect 13715 630 13753 664
rect 13787 630 13825 664
rect 13859 630 13897 664
rect 13931 630 13969 664
rect 14003 630 14041 664
rect 14075 630 14113 664
rect 14147 630 14185 664
rect 14219 630 14257 664
rect 14291 630 14329 664
rect 14363 630 14401 664
rect 14435 630 14473 664
rect 14507 630 14545 664
rect 14579 630 14617 664
rect 14651 630 14689 664
rect 14723 630 14761 664
rect 14795 630 14833 664
rect 14867 639 14969 664
rect 15003 639 15117 673
rect 14867 630 15117 639
rect 59 606 15117 630
rect 59 572 212 606
rect 246 600 15117 606
rect 246 572 14969 600
rect 59 566 14969 572
rect 15003 566 15117 600
rect 59 528 15117 566
rect 59 494 284 528
rect 318 494 357 528
rect 391 494 430 528
rect 464 494 503 528
rect 537 494 576 528
rect 610 494 649 528
rect 683 494 722 528
rect 756 494 795 528
rect 829 494 868 528
rect 902 494 941 528
rect 975 494 1014 528
rect 1048 494 1087 528
rect 1121 494 1160 528
rect 1194 494 1233 528
rect 1267 494 1306 528
rect 1340 494 1379 528
rect 1413 494 1452 528
rect 1486 494 1525 528
rect 1559 494 1598 528
rect 1632 494 1671 528
rect 1705 494 1744 528
rect 1778 494 1817 528
rect 1851 494 1890 528
rect 1924 494 1963 528
rect 1997 494 2036 528
rect 2070 494 2109 528
rect 2143 494 2182 528
rect 2216 494 2255 528
rect 2289 494 2328 528
rect 2362 494 2401 528
rect 2435 494 2474 528
rect 2508 494 2547 528
rect 2581 494 2620 528
rect 2654 494 2693 528
rect 2727 494 2766 528
rect 2800 494 2839 528
rect 2873 494 2912 528
rect 2946 494 2985 528
rect 3019 494 3058 528
rect 3092 494 3131 528
rect 3165 494 3204 528
rect 3238 494 3277 528
rect 3311 494 3350 528
rect 3384 494 3423 528
rect 3457 494 3496 528
rect 3530 494 3569 528
rect 3603 494 3642 528
rect 3676 494 3715 528
rect 3749 494 3788 528
rect 3822 494 3861 528
rect 3895 494 3934 528
rect 3968 494 4007 528
rect 4041 494 4080 528
rect 4114 494 4153 528
rect 4187 494 4226 528
rect 4260 494 4299 528
rect 4333 494 4372 528
rect 4406 494 4445 528
rect 4479 494 4518 528
rect 4552 494 4591 528
rect 4625 494 4664 528
rect 4698 494 4737 528
rect 4771 494 4810 528
rect 4844 494 4883 528
rect 4917 494 4956 528
rect 4990 494 5029 528
rect 5063 494 5102 528
rect 5136 494 5175 528
rect 5209 494 5248 528
rect 5282 494 5321 528
rect 5355 494 5393 528
rect 5427 494 5465 528
rect 5499 494 5537 528
rect 5571 494 5609 528
rect 5643 494 5681 528
rect 5715 494 5753 528
rect 5787 494 5825 528
rect 5859 494 5897 528
rect 5931 494 5969 528
rect 6003 494 6041 528
rect 6075 494 6113 528
rect 6147 494 6185 528
rect 6219 494 6257 528
rect 6291 494 6329 528
rect 6363 494 6401 528
rect 6435 494 6473 528
rect 6507 494 6545 528
rect 6579 494 6617 528
rect 6651 494 6689 528
rect 6723 494 6761 528
rect 6795 494 6833 528
rect 6867 494 6905 528
rect 6939 494 6977 528
rect 7011 494 7049 528
rect 7083 494 7121 528
rect 7155 494 7193 528
rect 7227 494 7265 528
rect 7299 494 7337 528
rect 7371 494 7409 528
rect 7443 494 7481 528
rect 7515 494 7553 528
rect 7587 494 7625 528
rect 7659 494 7697 528
rect 7731 494 7769 528
rect 7803 494 7841 528
rect 7875 494 7913 528
rect 7947 494 7985 528
rect 8019 494 8057 528
rect 8091 494 8129 528
rect 8163 494 8201 528
rect 8235 494 8273 528
rect 8307 494 8345 528
rect 8379 494 8417 528
rect 8451 494 8489 528
rect 8523 494 8561 528
rect 8595 494 8633 528
rect 8667 494 8705 528
rect 8739 494 8777 528
rect 8811 494 8849 528
rect 8883 494 8921 528
rect 8955 494 8993 528
rect 9027 494 9065 528
rect 9099 494 9137 528
rect 9171 494 9209 528
rect 9243 494 9281 528
rect 9315 494 9353 528
rect 9387 494 9425 528
rect 9459 494 9497 528
rect 9531 494 9569 528
rect 9603 494 9641 528
rect 9675 494 9713 528
rect 9747 494 9785 528
rect 9819 494 9857 528
rect 9891 494 9929 528
rect 9963 494 10001 528
rect 10035 494 10073 528
rect 10107 494 10145 528
rect 10179 494 10217 528
rect 10251 494 10289 528
rect 10323 494 10361 528
rect 10395 494 10433 528
rect 10467 494 10505 528
rect 10539 494 10577 528
rect 10611 494 10649 528
rect 10683 494 10721 528
rect 10755 494 10793 528
rect 10827 494 10865 528
rect 10899 494 10937 528
rect 10971 494 11009 528
rect 11043 494 11081 528
rect 11115 494 11153 528
rect 11187 494 11225 528
rect 11259 494 11297 528
rect 11331 494 11369 528
rect 11403 494 11441 528
rect 11475 494 11513 528
rect 11547 494 11585 528
rect 11619 494 11657 528
rect 11691 494 11729 528
rect 11763 494 11801 528
rect 11835 494 11873 528
rect 11907 494 11945 528
rect 11979 494 12017 528
rect 12051 494 12089 528
rect 12123 494 12161 528
rect 12195 494 12233 528
rect 12267 494 12305 528
rect 12339 494 12377 528
rect 12411 494 12449 528
rect 12483 494 12521 528
rect 12555 494 12593 528
rect 12627 494 12665 528
rect 12699 494 12737 528
rect 12771 494 12809 528
rect 12843 494 12881 528
rect 12915 494 12953 528
rect 12987 494 13025 528
rect 13059 494 13097 528
rect 13131 494 13169 528
rect 13203 494 13241 528
rect 13275 494 13313 528
rect 13347 494 13385 528
rect 13419 494 13457 528
rect 13491 494 13529 528
rect 13563 494 13601 528
rect 13635 494 13673 528
rect 13707 494 13745 528
rect 13779 494 13817 528
rect 13851 494 13889 528
rect 13923 494 13961 528
rect 13995 494 14033 528
rect 14067 494 14105 528
rect 14139 494 14177 528
rect 14211 494 14249 528
rect 14283 494 14321 528
rect 14355 494 14393 528
rect 14427 494 14465 528
rect 14499 494 14537 528
rect 14571 494 14609 528
rect 14643 494 14681 528
rect 14715 494 14753 528
rect 14787 494 14825 528
rect 14859 494 14897 528
rect 14931 494 15117 528
rect 59 473 15117 494
<< via1 >>
rect 575 4050 587 4068
rect 587 4050 621 4068
rect 621 4050 627 4068
rect 663 4050 693 4068
rect 693 4050 715 4068
rect 575 4016 627 4050
rect 663 4016 715 4050
rect 751 4044 803 4068
rect 751 4016 767 4044
rect 767 4016 803 4044
rect 575 3977 587 4003
rect 587 3977 621 4003
rect 621 3977 627 4003
rect 663 3977 693 4003
rect 693 3977 715 4003
rect 575 3951 627 3977
rect 663 3951 715 3977
rect 751 3971 803 4003
rect 751 3951 767 3971
rect 767 3951 803 3971
rect 575 3904 587 3938
rect 587 3904 621 3938
rect 621 3904 627 3938
rect 663 3904 693 3938
rect 693 3904 715 3938
rect 751 3937 767 3938
rect 767 3937 803 3938
rect 575 3886 627 3904
rect 663 3886 715 3904
rect 751 3898 803 3937
rect 751 3886 767 3898
rect 767 3886 803 3898
rect 575 3865 627 3873
rect 663 3865 715 3873
rect 575 3831 587 3865
rect 587 3831 621 3865
rect 621 3831 627 3865
rect 663 3831 693 3865
rect 693 3831 715 3865
rect 751 3864 767 3873
rect 767 3864 803 3873
rect 575 3821 627 3831
rect 663 3821 715 3831
rect 751 3825 803 3864
rect 751 3821 767 3825
rect 767 3821 803 3825
rect 575 3792 627 3808
rect 663 3792 715 3808
rect 575 3758 587 3792
rect 587 3758 621 3792
rect 621 3758 627 3792
rect 663 3758 693 3792
rect 693 3758 715 3792
rect 751 3791 767 3808
rect 767 3791 803 3808
rect 575 3756 627 3758
rect 663 3756 715 3758
rect 751 3756 803 3791
rect 575 3719 627 3743
rect 663 3719 715 3743
rect 575 3691 587 3719
rect 587 3691 621 3719
rect 621 3691 627 3719
rect 663 3691 693 3719
rect 693 3691 715 3719
rect 751 3718 767 3743
rect 767 3718 803 3743
rect 751 3691 803 3718
rect 575 3646 627 3678
rect 663 3646 715 3678
rect 575 3626 587 3646
rect 587 3626 621 3646
rect 621 3626 627 3646
rect 663 3626 693 3646
rect 693 3626 715 3646
rect 751 3645 767 3678
rect 767 3645 803 3678
rect 751 3626 803 3645
rect 575 3612 587 3613
rect 587 3612 621 3613
rect 621 3612 627 3613
rect 663 3612 693 3613
rect 693 3612 715 3613
rect 575 3573 627 3612
rect 663 3573 715 3612
rect 751 3606 803 3613
rect 575 3561 587 3573
rect 587 3561 621 3573
rect 621 3561 627 3573
rect 663 3561 693 3573
rect 693 3561 715 3573
rect 751 3572 767 3606
rect 767 3572 803 3606
rect 751 3561 803 3572
rect 575 3539 587 3548
rect 587 3539 621 3548
rect 621 3539 627 3548
rect 663 3539 693 3548
rect 693 3539 715 3548
rect 575 3500 627 3539
rect 663 3500 715 3539
rect 751 3533 803 3548
rect 575 3496 587 3500
rect 587 3496 621 3500
rect 621 3496 627 3500
rect 663 3496 693 3500
rect 693 3496 715 3500
rect 751 3499 767 3533
rect 767 3499 803 3533
rect 751 3496 803 3499
rect 575 3466 587 3483
rect 587 3466 621 3483
rect 621 3466 627 3483
rect 663 3466 693 3483
rect 693 3466 715 3483
rect 575 3431 627 3466
rect 663 3431 715 3466
rect 751 3460 803 3483
rect 751 3431 767 3460
rect 767 3431 803 3460
rect 575 3393 587 3418
rect 587 3393 621 3418
rect 621 3393 627 3418
rect 663 3393 693 3418
rect 693 3393 715 3418
rect 575 3366 627 3393
rect 663 3366 715 3393
rect 751 3387 803 3418
rect 751 3366 767 3387
rect 767 3366 803 3387
rect 575 3320 587 3353
rect 587 3320 621 3353
rect 621 3320 627 3353
rect 663 3320 693 3353
rect 693 3320 715 3353
rect 575 3301 627 3320
rect 663 3301 715 3320
rect 751 3314 803 3353
rect 751 3301 767 3314
rect 767 3301 803 3314
rect 575 3281 627 3288
rect 663 3281 715 3288
rect 575 3247 587 3281
rect 587 3247 621 3281
rect 621 3247 627 3281
rect 663 3247 693 3281
rect 693 3247 715 3281
rect 751 3280 767 3288
rect 767 3280 803 3288
rect 575 3236 627 3247
rect 663 3236 715 3247
rect 751 3241 803 3280
rect 751 3236 767 3241
rect 767 3236 803 3241
rect 575 3208 627 3223
rect 663 3208 715 3223
rect 575 3174 587 3208
rect 587 3174 621 3208
rect 621 3174 627 3208
rect 663 3174 693 3208
rect 693 3174 715 3208
rect 751 3207 767 3223
rect 767 3207 803 3223
rect 575 3171 627 3174
rect 663 3171 715 3174
rect 751 3171 803 3207
rect 575 3135 627 3158
rect 663 3135 715 3158
rect 575 3106 587 3135
rect 587 3106 621 3135
rect 621 3106 627 3135
rect 663 3106 693 3135
rect 693 3106 715 3135
rect 751 3134 767 3158
rect 767 3134 803 3158
rect 751 3106 803 3134
rect 575 3062 627 3093
rect 663 3062 715 3093
rect 575 3041 587 3062
rect 587 3041 621 3062
rect 621 3041 627 3062
rect 663 3041 693 3062
rect 693 3041 715 3062
rect 751 3061 767 3093
rect 767 3061 803 3093
rect 751 3041 803 3061
rect 575 2989 627 3028
rect 663 2989 715 3028
rect 751 3022 803 3028
rect 575 2976 587 2989
rect 587 2976 621 2989
rect 621 2976 627 2989
rect 663 2976 693 2989
rect 693 2976 715 2989
rect 751 2988 767 3022
rect 767 2988 803 3022
rect 751 2976 803 2988
rect 575 2955 587 2963
rect 587 2955 621 2963
rect 621 2955 627 2963
rect 663 2955 693 2963
rect 693 2955 715 2963
rect 575 2916 627 2955
rect 663 2916 715 2955
rect 751 2949 803 2963
rect 575 2911 587 2916
rect 587 2911 621 2916
rect 621 2911 627 2916
rect 663 2911 693 2916
rect 693 2911 715 2916
rect 751 2915 767 2949
rect 767 2915 803 2949
rect 751 2911 803 2915
rect 575 2882 587 2898
rect 587 2882 621 2898
rect 621 2882 627 2898
rect 663 2882 693 2898
rect 693 2882 715 2898
rect 575 2846 627 2882
rect 663 2846 715 2882
rect 751 2876 803 2898
rect 751 2846 767 2876
rect 767 2846 803 2876
rect 575 2809 587 2833
rect 587 2809 621 2833
rect 621 2809 627 2833
rect 663 2809 693 2833
rect 693 2809 715 2833
rect 575 2781 627 2809
rect 663 2781 715 2809
rect 751 2803 803 2833
rect 751 2781 767 2803
rect 767 2781 803 2803
rect 575 2736 587 2768
rect 587 2736 621 2768
rect 621 2736 627 2768
rect 663 2736 693 2768
rect 693 2736 715 2768
rect 575 2716 627 2736
rect 663 2716 715 2736
rect 751 2730 803 2768
rect 751 2716 767 2730
rect 767 2716 803 2730
rect 575 2697 627 2703
rect 663 2697 715 2703
rect 575 2663 587 2697
rect 587 2663 621 2697
rect 621 2663 627 2697
rect 663 2663 693 2697
rect 693 2663 715 2697
rect 751 2696 767 2703
rect 767 2696 803 2703
rect 575 2651 627 2663
rect 663 2651 715 2663
rect 751 2657 803 2696
rect 751 2651 767 2657
rect 767 2651 803 2657
rect 575 2624 627 2638
rect 663 2624 715 2638
rect 575 2590 587 2624
rect 587 2590 621 2624
rect 621 2590 627 2624
rect 663 2590 693 2624
rect 693 2590 715 2624
rect 751 2623 767 2638
rect 767 2623 803 2638
rect 575 2586 627 2590
rect 663 2586 715 2590
rect 751 2586 803 2623
rect 575 2551 627 2573
rect 663 2551 715 2573
rect 575 2521 587 2551
rect 587 2521 621 2551
rect 621 2521 627 2551
rect 663 2521 693 2551
rect 693 2521 715 2551
rect 751 2550 767 2573
rect 767 2550 803 2573
rect 751 2521 803 2550
rect 575 2478 627 2508
rect 663 2478 715 2508
rect 575 2456 587 2478
rect 587 2456 621 2478
rect 621 2456 627 2478
rect 663 2456 693 2478
rect 693 2456 715 2478
rect 751 2477 767 2508
rect 767 2477 803 2508
rect 751 2456 803 2477
rect 575 2405 627 2443
rect 663 2405 715 2443
rect 751 2438 803 2443
rect 575 2391 587 2405
rect 587 2391 621 2405
rect 621 2391 627 2405
rect 663 2391 693 2405
rect 693 2391 715 2405
rect 751 2404 767 2438
rect 767 2404 803 2438
rect 751 2391 803 2404
rect 575 2371 587 2378
rect 587 2371 621 2378
rect 621 2371 627 2378
rect 663 2371 693 2378
rect 693 2371 715 2378
rect 575 2332 627 2371
rect 663 2332 715 2371
rect 751 2365 803 2378
rect 575 2326 587 2332
rect 587 2326 621 2332
rect 621 2326 627 2332
rect 663 2326 693 2332
rect 693 2326 715 2332
rect 751 2331 767 2365
rect 767 2331 803 2365
rect 751 2326 803 2331
rect 575 2298 587 2313
rect 587 2298 621 2313
rect 621 2298 627 2313
rect 663 2298 693 2313
rect 693 2298 715 2313
rect 575 2261 627 2298
rect 663 2261 715 2298
rect 751 2292 803 2313
rect 751 2261 767 2292
rect 767 2261 803 2292
rect 575 2225 587 2248
rect 587 2225 621 2248
rect 621 2225 627 2248
rect 663 2225 693 2248
rect 693 2225 715 2248
rect 575 2196 627 2225
rect 663 2196 715 2225
rect 751 2219 803 2248
rect 751 2196 767 2219
rect 767 2196 803 2219
rect 575 2152 587 2183
rect 587 2152 621 2183
rect 621 2152 627 2183
rect 663 2152 693 2183
rect 693 2152 715 2183
rect 575 2131 627 2152
rect 663 2131 715 2152
rect 751 2146 803 2183
rect 751 2131 767 2146
rect 767 2131 803 2146
rect 575 2113 627 2118
rect 663 2113 715 2118
rect 575 2079 587 2113
rect 587 2079 621 2113
rect 621 2079 627 2113
rect 663 2079 693 2113
rect 693 2079 715 2113
rect 751 2112 767 2118
rect 767 2112 803 2118
rect 575 2066 627 2079
rect 663 2066 715 2079
rect 751 2073 803 2112
rect 751 2066 767 2073
rect 767 2066 803 2073
rect 575 2040 627 2053
rect 663 2040 715 2053
rect 575 2006 587 2040
rect 587 2006 621 2040
rect 621 2006 627 2040
rect 663 2006 693 2040
rect 693 2006 715 2040
rect 751 2039 767 2053
rect 767 2039 803 2053
rect 575 2001 627 2006
rect 663 2001 715 2006
rect 751 2001 803 2039
rect 575 1967 627 1987
rect 663 1967 715 1987
rect 575 1935 587 1967
rect 587 1935 621 1967
rect 621 1935 627 1967
rect 663 1935 693 1967
rect 693 1935 715 1967
rect 751 1966 767 1987
rect 767 1966 803 1987
rect 751 1935 803 1966
rect 575 1894 627 1921
rect 663 1894 715 1921
rect 575 1869 587 1894
rect 587 1869 621 1894
rect 621 1869 627 1894
rect 663 1869 693 1894
rect 693 1869 715 1894
rect 751 1893 767 1921
rect 767 1893 803 1921
rect 751 1869 803 1893
rect 575 1821 627 1855
rect 663 1821 715 1855
rect 751 1854 803 1855
rect 575 1803 587 1821
rect 587 1803 621 1821
rect 621 1803 627 1821
rect 663 1803 693 1821
rect 693 1803 715 1821
rect 751 1820 767 1854
rect 767 1820 803 1854
rect 751 1803 803 1820
rect 575 1787 587 1789
rect 587 1787 621 1789
rect 621 1787 627 1789
rect 663 1787 693 1789
rect 693 1787 715 1789
rect 575 1748 627 1787
rect 663 1748 715 1787
rect 751 1781 803 1789
rect 575 1737 587 1748
rect 587 1737 621 1748
rect 621 1737 627 1748
rect 663 1737 693 1748
rect 693 1737 715 1748
rect 751 1747 767 1781
rect 767 1747 803 1781
rect 751 1737 803 1747
rect 575 1714 587 1723
rect 587 1714 621 1723
rect 621 1714 627 1723
rect 663 1714 693 1723
rect 693 1714 715 1723
rect 575 1675 627 1714
rect 663 1675 715 1714
rect 751 1708 803 1723
rect 575 1671 587 1675
rect 587 1671 621 1675
rect 621 1671 627 1675
rect 663 1671 693 1675
rect 693 1671 715 1675
rect 751 1674 767 1708
rect 767 1674 803 1708
rect 751 1671 803 1674
rect 575 1641 587 1657
rect 587 1641 621 1657
rect 621 1641 627 1657
rect 663 1641 693 1657
rect 693 1641 715 1657
rect 575 1605 627 1641
rect 663 1605 715 1641
rect 751 1635 803 1657
rect 751 1605 767 1635
rect 767 1605 803 1635
rect 575 1568 587 1591
rect 587 1568 621 1591
rect 621 1568 627 1591
rect 663 1568 693 1591
rect 693 1568 715 1591
rect 575 1539 627 1568
rect 663 1539 715 1568
rect 751 1562 803 1591
rect 751 1539 767 1562
rect 767 1539 803 1562
rect 575 1495 587 1525
rect 587 1495 621 1525
rect 621 1495 627 1525
rect 663 1495 693 1525
rect 693 1495 715 1525
rect 575 1473 627 1495
rect 663 1473 715 1495
rect 751 1489 803 1525
rect 751 1473 767 1489
rect 767 1473 803 1489
rect 1109 4062 1161 4068
rect 1109 4028 1110 4062
rect 1110 4028 1144 4062
rect 1144 4028 1161 4062
rect 1109 4016 1161 4028
rect 1173 4062 1225 4068
rect 1173 4028 1182 4062
rect 1182 4028 1216 4062
rect 1216 4028 1225 4062
rect 1173 4016 1225 4028
rect 1237 4062 1289 4068
rect 1237 4028 1254 4062
rect 1254 4028 1288 4062
rect 1288 4028 1289 4062
rect 1237 4016 1289 4028
rect 1109 3988 1161 4003
rect 1109 3954 1110 3988
rect 1110 3954 1144 3988
rect 1144 3954 1161 3988
rect 1109 3951 1161 3954
rect 1173 3988 1225 4003
rect 1173 3954 1182 3988
rect 1182 3954 1216 3988
rect 1216 3954 1225 3988
rect 1173 3951 1225 3954
rect 1237 3988 1289 4003
rect 1237 3954 1254 3988
rect 1254 3954 1288 3988
rect 1288 3954 1289 3988
rect 1237 3951 1289 3954
rect 1109 3914 1161 3938
rect 1109 3886 1110 3914
rect 1110 3886 1144 3914
rect 1144 3886 1161 3914
rect 1173 3914 1225 3938
rect 1173 3886 1182 3914
rect 1182 3886 1216 3914
rect 1216 3886 1225 3914
rect 1237 3914 1289 3938
rect 1237 3886 1254 3914
rect 1254 3886 1288 3914
rect 1288 3886 1289 3914
rect 1109 3840 1161 3873
rect 1109 3821 1110 3840
rect 1110 3821 1144 3840
rect 1144 3821 1161 3840
rect 1173 3840 1225 3873
rect 1173 3821 1182 3840
rect 1182 3821 1216 3840
rect 1216 3821 1225 3840
rect 1237 3840 1289 3873
rect 1237 3821 1254 3840
rect 1254 3821 1288 3840
rect 1288 3821 1289 3840
rect 1109 3806 1110 3808
rect 1110 3806 1144 3808
rect 1144 3806 1161 3808
rect 1109 3766 1161 3806
rect 1109 3756 1110 3766
rect 1110 3756 1144 3766
rect 1144 3756 1161 3766
rect 1173 3806 1182 3808
rect 1182 3806 1216 3808
rect 1216 3806 1225 3808
rect 1173 3766 1225 3806
rect 1173 3756 1182 3766
rect 1182 3756 1216 3766
rect 1216 3756 1225 3766
rect 1237 3806 1254 3808
rect 1254 3806 1288 3808
rect 1288 3806 1289 3808
rect 1237 3766 1289 3806
rect 1237 3756 1254 3766
rect 1254 3756 1288 3766
rect 1288 3756 1289 3766
rect 1109 3732 1110 3743
rect 1110 3732 1144 3743
rect 1144 3732 1161 3743
rect 1109 3692 1161 3732
rect 1109 3691 1110 3692
rect 1110 3691 1144 3692
rect 1144 3691 1161 3692
rect 1173 3732 1182 3743
rect 1182 3732 1216 3743
rect 1216 3732 1225 3743
rect 1173 3692 1225 3732
rect 1173 3691 1182 3692
rect 1182 3691 1216 3692
rect 1216 3691 1225 3692
rect 1237 3732 1254 3743
rect 1254 3732 1288 3743
rect 1288 3732 1289 3743
rect 1237 3692 1289 3732
rect 1237 3691 1254 3692
rect 1254 3691 1288 3692
rect 1288 3691 1289 3692
rect 1109 3658 1110 3678
rect 1110 3658 1144 3678
rect 1144 3658 1161 3678
rect 1109 3626 1161 3658
rect 1173 3658 1182 3678
rect 1182 3658 1216 3678
rect 1216 3658 1225 3678
rect 1173 3626 1225 3658
rect 1237 3658 1254 3678
rect 1254 3658 1288 3678
rect 1288 3658 1289 3678
rect 1237 3626 1289 3658
rect 1109 3584 1110 3613
rect 1110 3584 1144 3613
rect 1144 3584 1161 3613
rect 1109 3561 1161 3584
rect 1173 3584 1182 3613
rect 1182 3584 1216 3613
rect 1216 3584 1225 3613
rect 1173 3561 1225 3584
rect 1237 3584 1254 3613
rect 1254 3584 1288 3613
rect 1288 3584 1289 3613
rect 1237 3561 1289 3584
rect 1109 3544 1161 3548
rect 1109 3510 1110 3544
rect 1110 3510 1144 3544
rect 1144 3510 1161 3544
rect 1109 3496 1161 3510
rect 1173 3544 1225 3548
rect 1173 3510 1182 3544
rect 1182 3510 1216 3544
rect 1216 3510 1225 3544
rect 1173 3496 1225 3510
rect 1237 3544 1289 3548
rect 1237 3510 1254 3544
rect 1254 3510 1288 3544
rect 1288 3510 1289 3544
rect 1237 3496 1289 3510
rect 1109 3470 1161 3483
rect 1109 3436 1110 3470
rect 1110 3436 1144 3470
rect 1144 3436 1161 3470
rect 1109 3431 1161 3436
rect 1173 3470 1225 3483
rect 1173 3436 1182 3470
rect 1182 3436 1216 3470
rect 1216 3436 1225 3470
rect 1173 3431 1225 3436
rect 1237 3470 1289 3483
rect 1237 3436 1254 3470
rect 1254 3436 1288 3470
rect 1288 3436 1289 3470
rect 1237 3431 1289 3436
rect 1109 3396 1161 3418
rect 1109 3366 1110 3396
rect 1110 3366 1144 3396
rect 1144 3366 1161 3396
rect 1173 3396 1225 3418
rect 1173 3366 1182 3396
rect 1182 3366 1216 3396
rect 1216 3366 1225 3396
rect 1237 3396 1289 3418
rect 1237 3366 1254 3396
rect 1254 3366 1288 3396
rect 1288 3366 1289 3396
rect 1109 3322 1161 3353
rect 1109 3301 1110 3322
rect 1110 3301 1144 3322
rect 1144 3301 1161 3322
rect 1173 3322 1225 3353
rect 1173 3301 1182 3322
rect 1182 3301 1216 3322
rect 1216 3301 1225 3322
rect 1237 3322 1289 3353
rect 1237 3301 1254 3322
rect 1254 3301 1288 3322
rect 1288 3301 1289 3322
rect 1109 3248 1161 3288
rect 1109 3236 1110 3248
rect 1110 3236 1144 3248
rect 1144 3236 1161 3248
rect 1173 3248 1225 3288
rect 1173 3236 1182 3248
rect 1182 3236 1216 3248
rect 1216 3236 1225 3248
rect 1237 3248 1289 3288
rect 1237 3236 1254 3248
rect 1254 3236 1288 3248
rect 1288 3236 1289 3248
rect 1109 3214 1110 3223
rect 1110 3214 1144 3223
rect 1144 3214 1161 3223
rect 1109 3174 1161 3214
rect 1109 3171 1110 3174
rect 1110 3171 1144 3174
rect 1144 3171 1161 3174
rect 1173 3214 1182 3223
rect 1182 3214 1216 3223
rect 1216 3214 1225 3223
rect 1173 3174 1225 3214
rect 1173 3171 1182 3174
rect 1182 3171 1216 3174
rect 1216 3171 1225 3174
rect 1237 3214 1254 3223
rect 1254 3214 1288 3223
rect 1288 3214 1289 3223
rect 1237 3174 1289 3214
rect 1237 3171 1254 3174
rect 1254 3171 1288 3174
rect 1288 3171 1289 3174
rect 1109 3140 1110 3158
rect 1110 3140 1144 3158
rect 1144 3140 1161 3158
rect 1109 3106 1161 3140
rect 1173 3140 1182 3158
rect 1182 3140 1216 3158
rect 1216 3140 1225 3158
rect 1173 3106 1225 3140
rect 1237 3140 1254 3158
rect 1254 3140 1288 3158
rect 1288 3140 1289 3158
rect 1237 3106 1289 3140
rect 1109 3066 1110 3093
rect 1110 3066 1144 3093
rect 1144 3066 1161 3093
rect 1109 3041 1161 3066
rect 1173 3066 1182 3093
rect 1182 3066 1216 3093
rect 1216 3066 1225 3093
rect 1173 3041 1225 3066
rect 1237 3066 1254 3093
rect 1254 3066 1288 3093
rect 1288 3066 1289 3093
rect 1237 3041 1289 3066
rect 1109 3026 1161 3028
rect 1109 2992 1110 3026
rect 1110 2992 1144 3026
rect 1144 2992 1161 3026
rect 1109 2976 1161 2992
rect 1173 3026 1225 3028
rect 1173 2992 1182 3026
rect 1182 2992 1216 3026
rect 1216 2992 1225 3026
rect 1173 2976 1225 2992
rect 1237 3026 1289 3028
rect 1237 2992 1254 3026
rect 1254 2992 1288 3026
rect 1288 2992 1289 3026
rect 1237 2976 1289 2992
rect 1109 2952 1161 2963
rect 1109 2918 1110 2952
rect 1110 2918 1144 2952
rect 1144 2918 1161 2952
rect 1109 2911 1161 2918
rect 1173 2952 1225 2963
rect 1173 2918 1182 2952
rect 1182 2918 1216 2952
rect 1216 2918 1225 2952
rect 1173 2911 1225 2918
rect 1237 2952 1289 2963
rect 1237 2918 1254 2952
rect 1254 2918 1288 2952
rect 1288 2918 1289 2952
rect 1237 2911 1289 2918
rect 1109 2878 1161 2898
rect 1109 2846 1110 2878
rect 1110 2846 1144 2878
rect 1144 2846 1161 2878
rect 1173 2878 1225 2898
rect 1173 2846 1182 2878
rect 1182 2846 1216 2878
rect 1216 2846 1225 2878
rect 1237 2878 1289 2898
rect 1237 2846 1254 2878
rect 1254 2846 1288 2878
rect 1288 2846 1289 2878
rect 1109 2804 1161 2833
rect 1109 2781 1110 2804
rect 1110 2781 1144 2804
rect 1144 2781 1161 2804
rect 1173 2804 1225 2833
rect 1173 2781 1182 2804
rect 1182 2781 1216 2804
rect 1216 2781 1225 2804
rect 1237 2804 1289 2833
rect 1237 2781 1254 2804
rect 1254 2781 1288 2804
rect 1288 2781 1289 2804
rect 1109 2730 1161 2768
rect 1109 2716 1110 2730
rect 1110 2716 1144 2730
rect 1144 2716 1161 2730
rect 1173 2730 1225 2768
rect 1173 2716 1182 2730
rect 1182 2716 1216 2730
rect 1216 2716 1225 2730
rect 1237 2730 1289 2768
rect 1237 2716 1254 2730
rect 1254 2716 1288 2730
rect 1288 2716 1289 2730
rect 1109 2696 1110 2703
rect 1110 2696 1144 2703
rect 1144 2696 1161 2703
rect 1109 2656 1161 2696
rect 1109 2651 1110 2656
rect 1110 2651 1144 2656
rect 1144 2651 1161 2656
rect 1173 2696 1182 2703
rect 1182 2696 1216 2703
rect 1216 2696 1225 2703
rect 1173 2656 1225 2696
rect 1173 2651 1182 2656
rect 1182 2651 1216 2656
rect 1216 2651 1225 2656
rect 1237 2696 1254 2703
rect 1254 2696 1288 2703
rect 1288 2696 1289 2703
rect 1237 2656 1289 2696
rect 1237 2651 1254 2656
rect 1254 2651 1288 2656
rect 1288 2651 1289 2656
rect 1109 2622 1110 2638
rect 1110 2622 1144 2638
rect 1144 2622 1161 2638
rect 1109 2586 1161 2622
rect 1173 2622 1182 2638
rect 1182 2622 1216 2638
rect 1216 2622 1225 2638
rect 1173 2586 1225 2622
rect 1237 2622 1254 2638
rect 1254 2622 1288 2638
rect 1288 2622 1289 2638
rect 1237 2586 1289 2622
rect 1109 2548 1110 2573
rect 1110 2548 1144 2573
rect 1144 2548 1161 2573
rect 1109 2521 1161 2548
rect 1173 2548 1182 2573
rect 1182 2548 1216 2573
rect 1216 2548 1225 2573
rect 1173 2521 1225 2548
rect 1237 2548 1254 2573
rect 1254 2548 1288 2573
rect 1288 2548 1289 2573
rect 1237 2521 1289 2548
rect 1109 2474 1110 2508
rect 1110 2474 1144 2508
rect 1144 2474 1161 2508
rect 1109 2456 1161 2474
rect 1173 2474 1182 2508
rect 1182 2474 1216 2508
rect 1216 2474 1225 2508
rect 1173 2456 1225 2474
rect 1237 2474 1254 2508
rect 1254 2474 1288 2508
rect 1288 2474 1289 2508
rect 1237 2456 1289 2474
rect 1109 2434 1161 2443
rect 1109 2400 1110 2434
rect 1110 2400 1144 2434
rect 1144 2400 1161 2434
rect 1109 2391 1161 2400
rect 1173 2434 1225 2443
rect 1173 2400 1182 2434
rect 1182 2400 1216 2434
rect 1216 2400 1225 2434
rect 1173 2391 1225 2400
rect 1237 2434 1289 2443
rect 1237 2400 1254 2434
rect 1254 2400 1288 2434
rect 1288 2400 1289 2434
rect 1237 2391 1289 2400
rect 1109 2360 1161 2378
rect 1109 2326 1110 2360
rect 1110 2326 1144 2360
rect 1144 2326 1161 2360
rect 1173 2360 1225 2378
rect 1173 2326 1182 2360
rect 1182 2326 1216 2360
rect 1216 2326 1225 2360
rect 1237 2360 1289 2378
rect 1237 2326 1254 2360
rect 1254 2326 1288 2360
rect 1288 2326 1289 2360
rect 1109 2286 1161 2313
rect 1109 2261 1110 2286
rect 1110 2261 1144 2286
rect 1144 2261 1161 2286
rect 1173 2286 1225 2313
rect 1173 2261 1182 2286
rect 1182 2261 1216 2286
rect 1216 2261 1225 2286
rect 1237 2286 1289 2313
rect 1237 2261 1254 2286
rect 1254 2261 1288 2286
rect 1288 2261 1289 2286
rect 1109 2212 1161 2248
rect 1109 2196 1110 2212
rect 1110 2196 1144 2212
rect 1144 2196 1161 2212
rect 1173 2212 1225 2248
rect 1173 2196 1182 2212
rect 1182 2196 1216 2212
rect 1216 2196 1225 2212
rect 1237 2212 1289 2248
rect 1237 2196 1254 2212
rect 1254 2196 1288 2212
rect 1288 2196 1289 2212
rect 1109 2178 1110 2183
rect 1110 2178 1144 2183
rect 1144 2178 1161 2183
rect 1109 2138 1161 2178
rect 1109 2131 1110 2138
rect 1110 2131 1144 2138
rect 1144 2131 1161 2138
rect 1173 2178 1182 2183
rect 1182 2178 1216 2183
rect 1216 2178 1225 2183
rect 1173 2138 1225 2178
rect 1173 2131 1182 2138
rect 1182 2131 1216 2138
rect 1216 2131 1225 2138
rect 1237 2178 1254 2183
rect 1254 2178 1288 2183
rect 1288 2178 1289 2183
rect 1237 2138 1289 2178
rect 1237 2131 1254 2138
rect 1254 2131 1288 2138
rect 1288 2131 1289 2138
rect 1109 2104 1110 2118
rect 1110 2104 1144 2118
rect 1144 2104 1161 2118
rect 1109 2066 1161 2104
rect 1173 2104 1182 2118
rect 1182 2104 1216 2118
rect 1216 2104 1225 2118
rect 1173 2066 1225 2104
rect 1237 2104 1254 2118
rect 1254 2104 1288 2118
rect 1288 2104 1289 2118
rect 1237 2066 1289 2104
rect 1109 2030 1110 2053
rect 1110 2030 1144 2053
rect 1144 2030 1161 2053
rect 1109 2001 1161 2030
rect 1173 2030 1182 2053
rect 1182 2030 1216 2053
rect 1216 2030 1225 2053
rect 1173 2001 1225 2030
rect 1237 2030 1254 2053
rect 1254 2030 1288 2053
rect 1288 2030 1289 2053
rect 1237 2001 1289 2030
rect 1109 1956 1110 1987
rect 1110 1956 1144 1987
rect 1144 1956 1161 1987
rect 1109 1935 1161 1956
rect 1173 1956 1182 1987
rect 1182 1956 1216 1987
rect 1216 1956 1225 1987
rect 1173 1935 1225 1956
rect 1237 1956 1254 1987
rect 1254 1956 1288 1987
rect 1288 1956 1289 1987
rect 1237 1935 1289 1956
rect 1109 1916 1161 1921
rect 1109 1882 1110 1916
rect 1110 1882 1144 1916
rect 1144 1882 1161 1916
rect 1109 1869 1161 1882
rect 1173 1916 1225 1921
rect 1173 1882 1182 1916
rect 1182 1882 1216 1916
rect 1216 1882 1225 1916
rect 1173 1869 1225 1882
rect 1237 1916 1289 1921
rect 1237 1882 1254 1916
rect 1254 1882 1288 1916
rect 1288 1882 1289 1916
rect 1237 1869 1289 1882
rect 1109 1842 1161 1855
rect 1109 1808 1110 1842
rect 1110 1808 1144 1842
rect 1144 1808 1161 1842
rect 1109 1803 1161 1808
rect 1173 1842 1225 1855
rect 1173 1808 1182 1842
rect 1182 1808 1216 1842
rect 1216 1808 1225 1842
rect 1173 1803 1225 1808
rect 1237 1842 1289 1855
rect 1237 1808 1254 1842
rect 1254 1808 1288 1842
rect 1288 1808 1289 1842
rect 1237 1803 1289 1808
rect 1109 1768 1161 1789
rect 1109 1737 1110 1768
rect 1110 1737 1144 1768
rect 1144 1737 1161 1768
rect 1173 1768 1225 1789
rect 1173 1737 1182 1768
rect 1182 1737 1216 1768
rect 1216 1737 1225 1768
rect 1237 1768 1289 1789
rect 1237 1737 1254 1768
rect 1254 1737 1288 1768
rect 1288 1737 1289 1768
rect 1109 1694 1161 1723
rect 1109 1671 1110 1694
rect 1110 1671 1144 1694
rect 1144 1671 1161 1694
rect 1173 1694 1225 1723
rect 1173 1671 1182 1694
rect 1182 1671 1216 1694
rect 1216 1671 1225 1694
rect 1237 1694 1289 1723
rect 1237 1671 1254 1694
rect 1254 1671 1288 1694
rect 1288 1671 1289 1694
rect 1109 1620 1161 1657
rect 1109 1605 1110 1620
rect 1110 1605 1144 1620
rect 1144 1605 1161 1620
rect 1173 1620 1225 1657
rect 1173 1605 1182 1620
rect 1182 1605 1216 1620
rect 1216 1605 1225 1620
rect 1237 1620 1289 1657
rect 1237 1605 1254 1620
rect 1254 1605 1288 1620
rect 1288 1605 1289 1620
rect 1109 1586 1110 1591
rect 1110 1586 1144 1591
rect 1144 1586 1161 1591
rect 1109 1545 1161 1586
rect 1109 1539 1110 1545
rect 1110 1539 1144 1545
rect 1144 1539 1161 1545
rect 1173 1586 1182 1591
rect 1182 1586 1216 1591
rect 1216 1586 1225 1591
rect 1173 1545 1225 1586
rect 1173 1539 1182 1545
rect 1182 1539 1216 1545
rect 1216 1539 1225 1545
rect 1237 1586 1254 1591
rect 1254 1586 1288 1591
rect 1288 1586 1289 1591
rect 1237 1545 1289 1586
rect 1237 1539 1254 1545
rect 1254 1539 1288 1545
rect 1288 1539 1289 1545
rect 1109 1511 1110 1525
rect 1110 1511 1144 1525
rect 1144 1511 1161 1525
rect 1109 1473 1161 1511
rect 1173 1511 1182 1525
rect 1182 1511 1216 1525
rect 1216 1511 1225 1525
rect 1173 1473 1225 1511
rect 1237 1511 1254 1525
rect 1254 1511 1288 1525
rect 1288 1511 1289 1525
rect 1237 1473 1289 1511
rect 1605 4050 1657 4068
rect 1669 4062 1721 4068
rect 1669 4050 1678 4062
rect 1678 4050 1712 4062
rect 1712 4050 1721 4062
rect 1733 4050 1785 4068
rect 1605 4016 1606 4050
rect 1606 4016 1657 4050
rect 1669 4016 1721 4050
rect 1733 4016 1784 4050
rect 1784 4016 1785 4050
rect 1605 3951 1606 4003
rect 1606 3951 1657 4003
rect 1669 3951 1721 4003
rect 1733 3951 1784 4003
rect 1784 3951 1785 4003
rect 1605 3886 1606 3938
rect 1606 3886 1657 3938
rect 1669 3886 1721 3938
rect 1733 3886 1784 3938
rect 1784 3886 1785 3938
rect 1605 3821 1606 3873
rect 1606 3821 1657 3873
rect 1669 3821 1721 3873
rect 1733 3821 1784 3873
rect 1784 3821 1785 3873
rect 1605 3756 1606 3808
rect 1606 3756 1657 3808
rect 1669 3756 1721 3808
rect 1733 3756 1784 3808
rect 1784 3756 1785 3808
rect 1605 3691 1606 3743
rect 1606 3691 1657 3743
rect 1669 3691 1721 3743
rect 1733 3691 1784 3743
rect 1784 3691 1785 3743
rect 1605 3626 1606 3678
rect 1606 3626 1657 3678
rect 1669 3626 1721 3678
rect 1733 3626 1784 3678
rect 1784 3626 1785 3678
rect 1605 3561 1606 3613
rect 1606 3561 1657 3613
rect 1669 3561 1721 3613
rect 1733 3561 1784 3613
rect 1784 3561 1785 3613
rect 1605 3496 1606 3548
rect 1606 3496 1657 3548
rect 1669 3496 1721 3548
rect 1733 3496 1784 3548
rect 1784 3496 1785 3548
rect 1605 3431 1606 3483
rect 1606 3431 1657 3483
rect 1669 3431 1721 3483
rect 1733 3431 1784 3483
rect 1784 3431 1785 3483
rect 1605 3366 1606 3418
rect 1606 3366 1657 3418
rect 1669 3366 1721 3418
rect 1733 3366 1784 3418
rect 1784 3366 1785 3418
rect 1605 3301 1606 3353
rect 1606 3301 1657 3353
rect 1669 3301 1721 3353
rect 1733 3301 1784 3353
rect 1784 3301 1785 3353
rect 1605 3236 1606 3288
rect 1606 3236 1657 3288
rect 1669 3236 1721 3288
rect 1733 3236 1784 3288
rect 1784 3236 1785 3288
rect 1605 3171 1606 3223
rect 1606 3171 1657 3223
rect 1669 3171 1721 3223
rect 1733 3171 1784 3223
rect 1784 3171 1785 3223
rect 1605 3106 1606 3158
rect 1606 3106 1657 3158
rect 1669 3106 1721 3158
rect 1733 3106 1784 3158
rect 1784 3106 1785 3158
rect 1605 3080 1606 3093
rect 1606 3092 1657 3093
rect 1669 3092 1721 3093
rect 1733 3092 1784 3093
rect 1606 3080 1640 3092
rect 1640 3080 1657 3092
rect 1605 3041 1657 3080
rect 1669 3041 1721 3092
rect 1733 3080 1750 3092
rect 1750 3080 1784 3092
rect 1784 3080 1785 3093
rect 1733 3041 1785 3080
rect 1605 2976 1606 3028
rect 1606 2976 1657 3028
rect 1669 2976 1721 3028
rect 1733 2976 1784 3028
rect 1784 2976 1785 3028
rect 1605 2911 1606 2963
rect 1606 2911 1657 2963
rect 1669 2911 1721 2963
rect 1733 2911 1784 2963
rect 1784 2911 1785 2963
rect 1605 2846 1606 2898
rect 1606 2846 1657 2898
rect 1669 2846 1721 2898
rect 1733 2846 1784 2898
rect 1784 2846 1785 2898
rect 1605 2781 1606 2833
rect 1606 2781 1657 2833
rect 1669 2781 1721 2833
rect 1733 2781 1784 2833
rect 1784 2781 1785 2833
rect 1605 2716 1606 2768
rect 1606 2716 1657 2768
rect 1669 2716 1721 2768
rect 1733 2716 1784 2768
rect 1784 2716 1785 2768
rect 1605 2651 1606 2703
rect 1606 2651 1657 2703
rect 1669 2651 1721 2703
rect 1733 2651 1784 2703
rect 1784 2651 1785 2703
rect 1605 2586 1606 2638
rect 1606 2586 1657 2638
rect 1669 2586 1721 2638
rect 1733 2586 1784 2638
rect 1784 2586 1785 2638
rect 1605 2535 1657 2573
rect 1605 2521 1606 2535
rect 1606 2521 1640 2535
rect 1640 2521 1657 2535
rect 1669 2535 1721 2573
rect 1669 2521 1678 2535
rect 1678 2521 1712 2535
rect 1712 2521 1721 2535
rect 1733 2535 1785 2573
rect 1733 2521 1750 2535
rect 1750 2521 1784 2535
rect 1784 2521 1785 2535
rect 1605 2501 1606 2508
rect 1606 2501 1640 2508
rect 1640 2501 1657 2508
rect 1605 2456 1657 2501
rect 1669 2501 1678 2508
rect 1678 2501 1712 2508
rect 1712 2501 1721 2508
rect 1669 2461 1721 2501
rect 1669 2456 1678 2461
rect 1678 2456 1712 2461
rect 1712 2456 1721 2461
rect 1733 2501 1750 2508
rect 1750 2501 1784 2508
rect 1784 2501 1785 2508
rect 1733 2456 1785 2501
rect 1605 2391 1606 2443
rect 1606 2391 1657 2443
rect 1669 2391 1721 2443
rect 1733 2391 1784 2443
rect 1784 2391 1785 2443
rect 1605 2326 1606 2378
rect 1606 2326 1657 2378
rect 1669 2326 1721 2378
rect 1733 2326 1784 2378
rect 1784 2326 1785 2378
rect 1605 2261 1606 2313
rect 1606 2261 1657 2313
rect 1669 2261 1721 2313
rect 1733 2261 1784 2313
rect 1784 2261 1785 2313
rect 1605 2196 1606 2248
rect 1606 2196 1657 2248
rect 1669 2196 1721 2248
rect 1733 2196 1784 2248
rect 1784 2196 1785 2248
rect 1605 2131 1606 2183
rect 1606 2131 1657 2183
rect 1669 2131 1721 2183
rect 1733 2131 1784 2183
rect 1784 2131 1785 2183
rect 1605 2066 1606 2118
rect 1606 2066 1657 2118
rect 1669 2066 1721 2118
rect 1733 2066 1784 2118
rect 1784 2066 1785 2118
rect 1605 2001 1606 2053
rect 1606 2001 1657 2053
rect 1669 2001 1721 2053
rect 1733 2001 1784 2053
rect 1784 2001 1785 2053
rect 1605 1935 1606 1987
rect 1606 1935 1657 1987
rect 1669 1935 1721 1987
rect 1733 1935 1784 1987
rect 1784 1935 1785 1987
rect 1605 1869 1606 1921
rect 1606 1869 1657 1921
rect 1669 1869 1721 1921
rect 1733 1869 1784 1921
rect 1784 1869 1785 1921
rect 1605 1803 1606 1855
rect 1606 1803 1657 1855
rect 1669 1803 1721 1855
rect 1733 1803 1784 1855
rect 1784 1803 1785 1855
rect 1605 1737 1606 1789
rect 1606 1737 1657 1789
rect 1669 1737 1721 1789
rect 1733 1737 1784 1789
rect 1784 1737 1785 1789
rect 1605 1671 1606 1723
rect 1606 1671 1657 1723
rect 1669 1671 1721 1723
rect 1733 1671 1784 1723
rect 1784 1671 1785 1723
rect 1605 1605 1606 1657
rect 1606 1605 1657 1657
rect 1669 1605 1721 1657
rect 1733 1605 1784 1657
rect 1784 1605 1785 1657
rect 1605 1539 1606 1591
rect 1606 1539 1657 1591
rect 1669 1539 1721 1591
rect 1733 1539 1784 1591
rect 1784 1539 1785 1591
rect 1605 1479 1606 1525
rect 1606 1491 1657 1525
rect 1669 1491 1721 1525
rect 1733 1491 1784 1525
rect 1606 1479 1640 1491
rect 1640 1479 1657 1491
rect 1605 1473 1657 1479
rect 1669 1473 1721 1491
rect 1733 1479 1750 1491
rect 1750 1479 1784 1491
rect 1784 1479 1785 1525
rect 1733 1473 1785 1479
rect 2101 4062 2153 4068
rect 2101 4028 2102 4062
rect 2102 4028 2136 4062
rect 2136 4028 2153 4062
rect 2101 4016 2153 4028
rect 2165 4062 2217 4068
rect 2165 4028 2174 4062
rect 2174 4028 2208 4062
rect 2208 4028 2217 4062
rect 2165 4016 2217 4028
rect 2229 4062 2281 4068
rect 2229 4028 2246 4062
rect 2246 4028 2280 4062
rect 2280 4028 2281 4062
rect 2229 4016 2281 4028
rect 2101 3988 2153 4003
rect 2101 3954 2102 3988
rect 2102 3954 2136 3988
rect 2136 3954 2153 3988
rect 2101 3951 2153 3954
rect 2165 3988 2217 4003
rect 2165 3954 2174 3988
rect 2174 3954 2208 3988
rect 2208 3954 2217 3988
rect 2165 3951 2217 3954
rect 2229 3988 2281 4003
rect 2229 3954 2246 3988
rect 2246 3954 2280 3988
rect 2280 3954 2281 3988
rect 2229 3951 2281 3954
rect 2101 3914 2153 3938
rect 2101 3886 2102 3914
rect 2102 3886 2136 3914
rect 2136 3886 2153 3914
rect 2165 3914 2217 3938
rect 2165 3886 2174 3914
rect 2174 3886 2208 3914
rect 2208 3886 2217 3914
rect 2229 3914 2281 3938
rect 2229 3886 2246 3914
rect 2246 3886 2280 3914
rect 2280 3886 2281 3914
rect 2101 3840 2153 3873
rect 2101 3821 2102 3840
rect 2102 3821 2136 3840
rect 2136 3821 2153 3840
rect 2165 3840 2217 3873
rect 2165 3821 2174 3840
rect 2174 3821 2208 3840
rect 2208 3821 2217 3840
rect 2229 3840 2281 3873
rect 2229 3821 2246 3840
rect 2246 3821 2280 3840
rect 2280 3821 2281 3840
rect 2101 3806 2102 3808
rect 2102 3806 2136 3808
rect 2136 3806 2153 3808
rect 2101 3766 2153 3806
rect 2101 3756 2102 3766
rect 2102 3756 2136 3766
rect 2136 3756 2153 3766
rect 2165 3806 2174 3808
rect 2174 3806 2208 3808
rect 2208 3806 2217 3808
rect 2165 3766 2217 3806
rect 2165 3756 2174 3766
rect 2174 3756 2208 3766
rect 2208 3756 2217 3766
rect 2229 3806 2246 3808
rect 2246 3806 2280 3808
rect 2280 3806 2281 3808
rect 2229 3766 2281 3806
rect 2229 3756 2246 3766
rect 2246 3756 2280 3766
rect 2280 3756 2281 3766
rect 2101 3732 2102 3743
rect 2102 3732 2136 3743
rect 2136 3732 2153 3743
rect 2101 3692 2153 3732
rect 2101 3691 2102 3692
rect 2102 3691 2136 3692
rect 2136 3691 2153 3692
rect 2165 3732 2174 3743
rect 2174 3732 2208 3743
rect 2208 3732 2217 3743
rect 2165 3692 2217 3732
rect 2165 3691 2174 3692
rect 2174 3691 2208 3692
rect 2208 3691 2217 3692
rect 2229 3732 2246 3743
rect 2246 3732 2280 3743
rect 2280 3732 2281 3743
rect 2229 3692 2281 3732
rect 2229 3691 2246 3692
rect 2246 3691 2280 3692
rect 2280 3691 2281 3692
rect 2101 3658 2102 3678
rect 2102 3658 2136 3678
rect 2136 3658 2153 3678
rect 2101 3626 2153 3658
rect 2165 3658 2174 3678
rect 2174 3658 2208 3678
rect 2208 3658 2217 3678
rect 2165 3626 2217 3658
rect 2229 3658 2246 3678
rect 2246 3658 2280 3678
rect 2280 3658 2281 3678
rect 2229 3626 2281 3658
rect 2101 3584 2102 3613
rect 2102 3584 2136 3613
rect 2136 3584 2153 3613
rect 2101 3561 2153 3584
rect 2165 3584 2174 3613
rect 2174 3584 2208 3613
rect 2208 3584 2217 3613
rect 2165 3561 2217 3584
rect 2229 3584 2246 3613
rect 2246 3584 2280 3613
rect 2280 3584 2281 3613
rect 2229 3561 2281 3584
rect 2101 3544 2153 3548
rect 2101 3510 2102 3544
rect 2102 3510 2136 3544
rect 2136 3510 2153 3544
rect 2101 3496 2153 3510
rect 2165 3544 2217 3548
rect 2165 3510 2174 3544
rect 2174 3510 2208 3544
rect 2208 3510 2217 3544
rect 2165 3496 2217 3510
rect 2229 3544 2281 3548
rect 2229 3510 2246 3544
rect 2246 3510 2280 3544
rect 2280 3510 2281 3544
rect 2229 3496 2281 3510
rect 2101 3470 2153 3483
rect 2101 3436 2102 3470
rect 2102 3436 2136 3470
rect 2136 3436 2153 3470
rect 2101 3431 2153 3436
rect 2165 3470 2217 3483
rect 2165 3436 2174 3470
rect 2174 3436 2208 3470
rect 2208 3436 2217 3470
rect 2165 3431 2217 3436
rect 2229 3470 2281 3483
rect 2229 3436 2246 3470
rect 2246 3436 2280 3470
rect 2280 3436 2281 3470
rect 2229 3431 2281 3436
rect 2101 3396 2153 3418
rect 2101 3366 2102 3396
rect 2102 3366 2136 3396
rect 2136 3366 2153 3396
rect 2165 3396 2217 3418
rect 2165 3366 2174 3396
rect 2174 3366 2208 3396
rect 2208 3366 2217 3396
rect 2229 3396 2281 3418
rect 2229 3366 2246 3396
rect 2246 3366 2280 3396
rect 2280 3366 2281 3396
rect 2101 3322 2153 3353
rect 2101 3301 2102 3322
rect 2102 3301 2136 3322
rect 2136 3301 2153 3322
rect 2165 3322 2217 3353
rect 2165 3301 2174 3322
rect 2174 3301 2208 3322
rect 2208 3301 2217 3322
rect 2229 3322 2281 3353
rect 2229 3301 2246 3322
rect 2246 3301 2280 3322
rect 2280 3301 2281 3322
rect 2101 3248 2153 3288
rect 2101 3236 2102 3248
rect 2102 3236 2136 3248
rect 2136 3236 2153 3248
rect 2165 3248 2217 3288
rect 2165 3236 2174 3248
rect 2174 3236 2208 3248
rect 2208 3236 2217 3248
rect 2229 3248 2281 3288
rect 2229 3236 2246 3248
rect 2246 3236 2280 3248
rect 2280 3236 2281 3248
rect 2101 3214 2102 3223
rect 2102 3214 2136 3223
rect 2136 3214 2153 3223
rect 2101 3174 2153 3214
rect 2101 3171 2102 3174
rect 2102 3171 2136 3174
rect 2136 3171 2153 3174
rect 2165 3214 2174 3223
rect 2174 3214 2208 3223
rect 2208 3214 2217 3223
rect 2165 3174 2217 3214
rect 2165 3171 2174 3174
rect 2174 3171 2208 3174
rect 2208 3171 2217 3174
rect 2229 3214 2246 3223
rect 2246 3214 2280 3223
rect 2280 3214 2281 3223
rect 2229 3174 2281 3214
rect 2229 3171 2246 3174
rect 2246 3171 2280 3174
rect 2280 3171 2281 3174
rect 2101 3140 2102 3158
rect 2102 3140 2136 3158
rect 2136 3140 2153 3158
rect 2101 3106 2153 3140
rect 2165 3140 2174 3158
rect 2174 3140 2208 3158
rect 2208 3140 2217 3158
rect 2165 3106 2217 3140
rect 2229 3140 2246 3158
rect 2246 3140 2280 3158
rect 2280 3140 2281 3158
rect 2229 3106 2281 3140
rect 2101 3066 2102 3093
rect 2102 3066 2136 3093
rect 2136 3066 2153 3093
rect 2101 3041 2153 3066
rect 2165 3066 2174 3093
rect 2174 3066 2208 3093
rect 2208 3066 2217 3093
rect 2165 3041 2217 3066
rect 2229 3066 2246 3093
rect 2246 3066 2280 3093
rect 2280 3066 2281 3093
rect 2229 3041 2281 3066
rect 2101 3026 2153 3028
rect 2101 2992 2102 3026
rect 2102 2992 2136 3026
rect 2136 2992 2153 3026
rect 2101 2976 2153 2992
rect 2165 3026 2217 3028
rect 2165 2992 2174 3026
rect 2174 2992 2208 3026
rect 2208 2992 2217 3026
rect 2165 2976 2217 2992
rect 2229 3026 2281 3028
rect 2229 2992 2246 3026
rect 2246 2992 2280 3026
rect 2280 2992 2281 3026
rect 2229 2976 2281 2992
rect 2101 2952 2153 2963
rect 2101 2918 2102 2952
rect 2102 2918 2136 2952
rect 2136 2918 2153 2952
rect 2101 2911 2153 2918
rect 2165 2952 2217 2963
rect 2165 2918 2174 2952
rect 2174 2918 2208 2952
rect 2208 2918 2217 2952
rect 2165 2911 2217 2918
rect 2229 2952 2281 2963
rect 2229 2918 2246 2952
rect 2246 2918 2280 2952
rect 2280 2918 2281 2952
rect 2229 2911 2281 2918
rect 2101 2878 2153 2898
rect 2101 2846 2102 2878
rect 2102 2846 2136 2878
rect 2136 2846 2153 2878
rect 2165 2878 2217 2898
rect 2165 2846 2174 2878
rect 2174 2846 2208 2878
rect 2208 2846 2217 2878
rect 2229 2878 2281 2898
rect 2229 2846 2246 2878
rect 2246 2846 2280 2878
rect 2280 2846 2281 2878
rect 2101 2804 2153 2833
rect 2101 2781 2102 2804
rect 2102 2781 2136 2804
rect 2136 2781 2153 2804
rect 2165 2804 2217 2833
rect 2165 2781 2174 2804
rect 2174 2781 2208 2804
rect 2208 2781 2217 2804
rect 2229 2804 2281 2833
rect 2229 2781 2246 2804
rect 2246 2781 2280 2804
rect 2280 2781 2281 2804
rect 2101 2730 2153 2768
rect 2101 2716 2102 2730
rect 2102 2716 2136 2730
rect 2136 2716 2153 2730
rect 2165 2730 2217 2768
rect 2165 2716 2174 2730
rect 2174 2716 2208 2730
rect 2208 2716 2217 2730
rect 2229 2730 2281 2768
rect 2229 2716 2246 2730
rect 2246 2716 2280 2730
rect 2280 2716 2281 2730
rect 2101 2696 2102 2703
rect 2102 2696 2136 2703
rect 2136 2696 2153 2703
rect 2101 2656 2153 2696
rect 2101 2651 2102 2656
rect 2102 2651 2136 2656
rect 2136 2651 2153 2656
rect 2165 2696 2174 2703
rect 2174 2696 2208 2703
rect 2208 2696 2217 2703
rect 2165 2656 2217 2696
rect 2165 2651 2174 2656
rect 2174 2651 2208 2656
rect 2208 2651 2217 2656
rect 2229 2696 2246 2703
rect 2246 2696 2280 2703
rect 2280 2696 2281 2703
rect 2229 2656 2281 2696
rect 2229 2651 2246 2656
rect 2246 2651 2280 2656
rect 2280 2651 2281 2656
rect 2101 2622 2102 2638
rect 2102 2622 2136 2638
rect 2136 2622 2153 2638
rect 2101 2586 2153 2622
rect 2165 2622 2174 2638
rect 2174 2622 2208 2638
rect 2208 2622 2217 2638
rect 2165 2586 2217 2622
rect 2229 2622 2246 2638
rect 2246 2622 2280 2638
rect 2280 2622 2281 2638
rect 2229 2586 2281 2622
rect 2101 2548 2102 2573
rect 2102 2548 2136 2573
rect 2136 2548 2153 2573
rect 2101 2521 2153 2548
rect 2165 2548 2174 2573
rect 2174 2548 2208 2573
rect 2208 2548 2217 2573
rect 2165 2521 2217 2548
rect 2229 2548 2246 2573
rect 2246 2548 2280 2573
rect 2280 2548 2281 2573
rect 2229 2521 2281 2548
rect 2101 2474 2102 2508
rect 2102 2474 2136 2508
rect 2136 2474 2153 2508
rect 2101 2456 2153 2474
rect 2165 2474 2174 2508
rect 2174 2474 2208 2508
rect 2208 2474 2217 2508
rect 2165 2456 2217 2474
rect 2229 2474 2246 2508
rect 2246 2474 2280 2508
rect 2280 2474 2281 2508
rect 2229 2456 2281 2474
rect 2101 2434 2153 2443
rect 2101 2400 2102 2434
rect 2102 2400 2136 2434
rect 2136 2400 2153 2434
rect 2101 2391 2153 2400
rect 2165 2434 2217 2443
rect 2165 2400 2174 2434
rect 2174 2400 2208 2434
rect 2208 2400 2217 2434
rect 2165 2391 2217 2400
rect 2229 2434 2281 2443
rect 2229 2400 2246 2434
rect 2246 2400 2280 2434
rect 2280 2400 2281 2434
rect 2229 2391 2281 2400
rect 2101 2360 2153 2378
rect 2101 2326 2102 2360
rect 2102 2326 2136 2360
rect 2136 2326 2153 2360
rect 2165 2360 2217 2378
rect 2165 2326 2174 2360
rect 2174 2326 2208 2360
rect 2208 2326 2217 2360
rect 2229 2360 2281 2378
rect 2229 2326 2246 2360
rect 2246 2326 2280 2360
rect 2280 2326 2281 2360
rect 2101 2286 2153 2313
rect 2101 2261 2102 2286
rect 2102 2261 2136 2286
rect 2136 2261 2153 2286
rect 2165 2286 2217 2313
rect 2165 2261 2174 2286
rect 2174 2261 2208 2286
rect 2208 2261 2217 2286
rect 2229 2286 2281 2313
rect 2229 2261 2246 2286
rect 2246 2261 2280 2286
rect 2280 2261 2281 2286
rect 2101 2212 2153 2248
rect 2101 2196 2102 2212
rect 2102 2196 2136 2212
rect 2136 2196 2153 2212
rect 2165 2212 2217 2248
rect 2165 2196 2174 2212
rect 2174 2196 2208 2212
rect 2208 2196 2217 2212
rect 2229 2212 2281 2248
rect 2229 2196 2246 2212
rect 2246 2196 2280 2212
rect 2280 2196 2281 2212
rect 2101 2178 2102 2183
rect 2102 2178 2136 2183
rect 2136 2178 2153 2183
rect 2101 2138 2153 2178
rect 2101 2131 2102 2138
rect 2102 2131 2136 2138
rect 2136 2131 2153 2138
rect 2165 2178 2174 2183
rect 2174 2178 2208 2183
rect 2208 2178 2217 2183
rect 2165 2138 2217 2178
rect 2165 2131 2174 2138
rect 2174 2131 2208 2138
rect 2208 2131 2217 2138
rect 2229 2178 2246 2183
rect 2246 2178 2280 2183
rect 2280 2178 2281 2183
rect 2229 2138 2281 2178
rect 2229 2131 2246 2138
rect 2246 2131 2280 2138
rect 2280 2131 2281 2138
rect 2101 2104 2102 2118
rect 2102 2104 2136 2118
rect 2136 2104 2153 2118
rect 2101 2066 2153 2104
rect 2165 2104 2174 2118
rect 2174 2104 2208 2118
rect 2208 2104 2217 2118
rect 2165 2066 2217 2104
rect 2229 2104 2246 2118
rect 2246 2104 2280 2118
rect 2280 2104 2281 2118
rect 2229 2066 2281 2104
rect 2101 2030 2102 2053
rect 2102 2030 2136 2053
rect 2136 2030 2153 2053
rect 2101 2001 2153 2030
rect 2165 2030 2174 2053
rect 2174 2030 2208 2053
rect 2208 2030 2217 2053
rect 2165 2001 2217 2030
rect 2229 2030 2246 2053
rect 2246 2030 2280 2053
rect 2280 2030 2281 2053
rect 2229 2001 2281 2030
rect 2101 1956 2102 1987
rect 2102 1956 2136 1987
rect 2136 1956 2153 1987
rect 2101 1935 2153 1956
rect 2165 1956 2174 1987
rect 2174 1956 2208 1987
rect 2208 1956 2217 1987
rect 2165 1935 2217 1956
rect 2229 1956 2246 1987
rect 2246 1956 2280 1987
rect 2280 1956 2281 1987
rect 2229 1935 2281 1956
rect 2101 1916 2153 1921
rect 2101 1882 2102 1916
rect 2102 1882 2136 1916
rect 2136 1882 2153 1916
rect 2101 1869 2153 1882
rect 2165 1916 2217 1921
rect 2165 1882 2174 1916
rect 2174 1882 2208 1916
rect 2208 1882 2217 1916
rect 2165 1869 2217 1882
rect 2229 1916 2281 1921
rect 2229 1882 2246 1916
rect 2246 1882 2280 1916
rect 2280 1882 2281 1916
rect 2229 1869 2281 1882
rect 2101 1842 2153 1855
rect 2101 1808 2102 1842
rect 2102 1808 2136 1842
rect 2136 1808 2153 1842
rect 2101 1803 2153 1808
rect 2165 1842 2217 1855
rect 2165 1808 2174 1842
rect 2174 1808 2208 1842
rect 2208 1808 2217 1842
rect 2165 1803 2217 1808
rect 2229 1842 2281 1855
rect 2229 1808 2246 1842
rect 2246 1808 2280 1842
rect 2280 1808 2281 1842
rect 2229 1803 2281 1808
rect 2101 1768 2153 1789
rect 2101 1737 2102 1768
rect 2102 1737 2136 1768
rect 2136 1737 2153 1768
rect 2165 1768 2217 1789
rect 2165 1737 2174 1768
rect 2174 1737 2208 1768
rect 2208 1737 2217 1768
rect 2229 1768 2281 1789
rect 2229 1737 2246 1768
rect 2246 1737 2280 1768
rect 2280 1737 2281 1768
rect 2101 1694 2153 1723
rect 2101 1671 2102 1694
rect 2102 1671 2136 1694
rect 2136 1671 2153 1694
rect 2165 1694 2217 1723
rect 2165 1671 2174 1694
rect 2174 1671 2208 1694
rect 2208 1671 2217 1694
rect 2229 1694 2281 1723
rect 2229 1671 2246 1694
rect 2246 1671 2280 1694
rect 2280 1671 2281 1694
rect 2101 1620 2153 1657
rect 2101 1605 2102 1620
rect 2102 1605 2136 1620
rect 2136 1605 2153 1620
rect 2165 1620 2217 1657
rect 2165 1605 2174 1620
rect 2174 1605 2208 1620
rect 2208 1605 2217 1620
rect 2229 1620 2281 1657
rect 2229 1605 2246 1620
rect 2246 1605 2280 1620
rect 2280 1605 2281 1620
rect 2101 1586 2102 1591
rect 2102 1586 2136 1591
rect 2136 1586 2153 1591
rect 2101 1545 2153 1586
rect 2101 1539 2102 1545
rect 2102 1539 2136 1545
rect 2136 1539 2153 1545
rect 2165 1586 2174 1591
rect 2174 1586 2208 1591
rect 2208 1586 2217 1591
rect 2165 1545 2217 1586
rect 2165 1539 2174 1545
rect 2174 1539 2208 1545
rect 2208 1539 2217 1545
rect 2229 1586 2246 1591
rect 2246 1586 2280 1591
rect 2280 1586 2281 1591
rect 2229 1545 2281 1586
rect 2229 1539 2246 1545
rect 2246 1539 2280 1545
rect 2280 1539 2281 1545
rect 2101 1511 2102 1525
rect 2102 1511 2136 1525
rect 2136 1511 2153 1525
rect 2101 1473 2153 1511
rect 2165 1511 2174 1525
rect 2174 1511 2208 1525
rect 2208 1511 2217 1525
rect 2165 1473 2217 1511
rect 2229 1511 2246 1525
rect 2246 1511 2280 1525
rect 2280 1511 2281 1525
rect 2229 1473 2281 1511
rect 2597 4050 2649 4068
rect 2661 4062 2713 4068
rect 2661 4050 2670 4062
rect 2670 4050 2704 4062
rect 2704 4050 2713 4062
rect 2725 4050 2777 4068
rect 2597 4016 2598 4050
rect 2598 4016 2649 4050
rect 2661 4016 2713 4050
rect 2725 4016 2776 4050
rect 2776 4016 2777 4050
rect 2597 3951 2598 4003
rect 2598 3951 2649 4003
rect 2661 3951 2713 4003
rect 2725 3951 2776 4003
rect 2776 3951 2777 4003
rect 2597 3886 2598 3938
rect 2598 3886 2649 3938
rect 2661 3886 2713 3938
rect 2725 3886 2776 3938
rect 2776 3886 2777 3938
rect 2597 3821 2598 3873
rect 2598 3821 2649 3873
rect 2661 3821 2713 3873
rect 2725 3821 2776 3873
rect 2776 3821 2777 3873
rect 2597 3756 2598 3808
rect 2598 3756 2649 3808
rect 2661 3756 2713 3808
rect 2725 3756 2776 3808
rect 2776 3756 2777 3808
rect 2597 3691 2598 3743
rect 2598 3691 2649 3743
rect 2661 3691 2713 3743
rect 2725 3691 2776 3743
rect 2776 3691 2777 3743
rect 2597 3626 2598 3678
rect 2598 3626 2649 3678
rect 2661 3626 2713 3678
rect 2725 3626 2776 3678
rect 2776 3626 2777 3678
rect 2597 3561 2598 3613
rect 2598 3561 2649 3613
rect 2661 3561 2713 3613
rect 2725 3561 2776 3613
rect 2776 3561 2777 3613
rect 2597 3496 2598 3548
rect 2598 3496 2649 3548
rect 2661 3496 2713 3548
rect 2725 3496 2776 3548
rect 2776 3496 2777 3548
rect 2597 3431 2598 3483
rect 2598 3431 2649 3483
rect 2661 3431 2713 3483
rect 2725 3431 2776 3483
rect 2776 3431 2777 3483
rect 2597 3366 2598 3418
rect 2598 3366 2649 3418
rect 2661 3366 2713 3418
rect 2725 3366 2776 3418
rect 2776 3366 2777 3418
rect 2597 3301 2598 3353
rect 2598 3301 2649 3353
rect 2661 3301 2713 3353
rect 2725 3301 2776 3353
rect 2776 3301 2777 3353
rect 2597 3236 2598 3288
rect 2598 3236 2649 3288
rect 2661 3236 2713 3288
rect 2725 3236 2776 3288
rect 2776 3236 2777 3288
rect 2597 3171 2598 3223
rect 2598 3171 2649 3223
rect 2661 3171 2713 3223
rect 2725 3171 2776 3223
rect 2776 3171 2777 3223
rect 2597 3106 2598 3158
rect 2598 3106 2649 3158
rect 2661 3106 2713 3158
rect 2725 3106 2776 3158
rect 2776 3106 2777 3158
rect 2597 3080 2598 3093
rect 2598 3092 2649 3093
rect 2661 3092 2713 3093
rect 2725 3092 2776 3093
rect 2598 3080 2632 3092
rect 2632 3080 2649 3092
rect 2597 3041 2649 3080
rect 2661 3041 2713 3092
rect 2725 3080 2742 3092
rect 2742 3080 2776 3092
rect 2776 3080 2777 3093
rect 2725 3041 2777 3080
rect 2597 2976 2598 3028
rect 2598 2976 2649 3028
rect 2661 2976 2713 3028
rect 2725 2976 2776 3028
rect 2776 2976 2777 3028
rect 2597 2911 2598 2963
rect 2598 2911 2649 2963
rect 2661 2911 2713 2963
rect 2725 2911 2776 2963
rect 2776 2911 2777 2963
rect 2597 2846 2598 2898
rect 2598 2846 2649 2898
rect 2661 2846 2713 2898
rect 2725 2846 2776 2898
rect 2776 2846 2777 2898
rect 2597 2781 2598 2833
rect 2598 2781 2649 2833
rect 2661 2781 2713 2833
rect 2725 2781 2776 2833
rect 2776 2781 2777 2833
rect 2597 2716 2598 2768
rect 2598 2716 2649 2768
rect 2661 2716 2713 2768
rect 2725 2716 2776 2768
rect 2776 2716 2777 2768
rect 2597 2651 2598 2703
rect 2598 2651 2649 2703
rect 2661 2651 2713 2703
rect 2725 2651 2776 2703
rect 2776 2651 2777 2703
rect 2597 2586 2598 2638
rect 2598 2586 2649 2638
rect 2661 2586 2713 2638
rect 2725 2586 2776 2638
rect 2776 2586 2777 2638
rect 2597 2535 2649 2573
rect 2597 2521 2598 2535
rect 2598 2521 2632 2535
rect 2632 2521 2649 2535
rect 2661 2535 2713 2573
rect 2661 2521 2670 2535
rect 2670 2521 2704 2535
rect 2704 2521 2713 2535
rect 2725 2535 2777 2573
rect 2725 2521 2742 2535
rect 2742 2521 2776 2535
rect 2776 2521 2777 2535
rect 2597 2501 2598 2508
rect 2598 2501 2632 2508
rect 2632 2501 2649 2508
rect 2597 2456 2649 2501
rect 2661 2501 2670 2508
rect 2670 2501 2704 2508
rect 2704 2501 2713 2508
rect 2661 2461 2713 2501
rect 2661 2456 2670 2461
rect 2670 2456 2704 2461
rect 2704 2456 2713 2461
rect 2725 2501 2742 2508
rect 2742 2501 2776 2508
rect 2776 2501 2777 2508
rect 2725 2456 2777 2501
rect 2597 2391 2598 2443
rect 2598 2391 2649 2443
rect 2661 2391 2713 2443
rect 2725 2391 2776 2443
rect 2776 2391 2777 2443
rect 2597 2326 2598 2378
rect 2598 2326 2649 2378
rect 2661 2326 2713 2378
rect 2725 2326 2776 2378
rect 2776 2326 2777 2378
rect 2597 2261 2598 2313
rect 2598 2261 2649 2313
rect 2661 2261 2713 2313
rect 2725 2261 2776 2313
rect 2776 2261 2777 2313
rect 2597 2196 2598 2248
rect 2598 2196 2649 2248
rect 2661 2196 2713 2248
rect 2725 2196 2776 2248
rect 2776 2196 2777 2248
rect 2597 2131 2598 2183
rect 2598 2131 2649 2183
rect 2661 2131 2713 2183
rect 2725 2131 2776 2183
rect 2776 2131 2777 2183
rect 2597 2066 2598 2118
rect 2598 2066 2649 2118
rect 2661 2066 2713 2118
rect 2725 2066 2776 2118
rect 2776 2066 2777 2118
rect 2597 2001 2598 2053
rect 2598 2001 2649 2053
rect 2661 2001 2713 2053
rect 2725 2001 2776 2053
rect 2776 2001 2777 2053
rect 2597 1935 2598 1987
rect 2598 1935 2649 1987
rect 2661 1935 2713 1987
rect 2725 1935 2776 1987
rect 2776 1935 2777 1987
rect 2597 1869 2598 1921
rect 2598 1869 2649 1921
rect 2661 1869 2713 1921
rect 2725 1869 2776 1921
rect 2776 1869 2777 1921
rect 2597 1803 2598 1855
rect 2598 1803 2649 1855
rect 2661 1803 2713 1855
rect 2725 1803 2776 1855
rect 2776 1803 2777 1855
rect 2597 1737 2598 1789
rect 2598 1737 2649 1789
rect 2661 1737 2713 1789
rect 2725 1737 2776 1789
rect 2776 1737 2777 1789
rect 2597 1671 2598 1723
rect 2598 1671 2649 1723
rect 2661 1671 2713 1723
rect 2725 1671 2776 1723
rect 2776 1671 2777 1723
rect 2597 1605 2598 1657
rect 2598 1605 2649 1657
rect 2661 1605 2713 1657
rect 2725 1605 2776 1657
rect 2776 1605 2777 1657
rect 2597 1539 2598 1591
rect 2598 1539 2649 1591
rect 2661 1539 2713 1591
rect 2725 1539 2776 1591
rect 2776 1539 2777 1591
rect 2597 1479 2598 1525
rect 2598 1491 2649 1525
rect 2661 1491 2713 1525
rect 2725 1491 2776 1525
rect 2598 1479 2632 1491
rect 2632 1479 2649 1491
rect 2597 1473 2649 1479
rect 2661 1473 2713 1491
rect 2725 1479 2742 1491
rect 2742 1479 2776 1491
rect 2776 1479 2777 1525
rect 2725 1473 2777 1479
rect 3093 4062 3145 4068
rect 3093 4028 3094 4062
rect 3094 4028 3128 4062
rect 3128 4028 3145 4062
rect 3093 4016 3145 4028
rect 3157 4062 3209 4068
rect 3157 4028 3166 4062
rect 3166 4028 3200 4062
rect 3200 4028 3209 4062
rect 3157 4016 3209 4028
rect 3221 4062 3273 4068
rect 3221 4028 3238 4062
rect 3238 4028 3272 4062
rect 3272 4028 3273 4062
rect 3221 4016 3273 4028
rect 3093 3988 3145 4003
rect 3093 3954 3094 3988
rect 3094 3954 3128 3988
rect 3128 3954 3145 3988
rect 3093 3951 3145 3954
rect 3157 3988 3209 4003
rect 3157 3954 3166 3988
rect 3166 3954 3200 3988
rect 3200 3954 3209 3988
rect 3157 3951 3209 3954
rect 3221 3988 3273 4003
rect 3221 3954 3238 3988
rect 3238 3954 3272 3988
rect 3272 3954 3273 3988
rect 3221 3951 3273 3954
rect 3093 3914 3145 3938
rect 3093 3886 3094 3914
rect 3094 3886 3128 3914
rect 3128 3886 3145 3914
rect 3157 3914 3209 3938
rect 3157 3886 3166 3914
rect 3166 3886 3200 3914
rect 3200 3886 3209 3914
rect 3221 3914 3273 3938
rect 3221 3886 3238 3914
rect 3238 3886 3272 3914
rect 3272 3886 3273 3914
rect 3093 3840 3145 3873
rect 3093 3821 3094 3840
rect 3094 3821 3128 3840
rect 3128 3821 3145 3840
rect 3157 3840 3209 3873
rect 3157 3821 3166 3840
rect 3166 3821 3200 3840
rect 3200 3821 3209 3840
rect 3221 3840 3273 3873
rect 3221 3821 3238 3840
rect 3238 3821 3272 3840
rect 3272 3821 3273 3840
rect 3093 3806 3094 3808
rect 3094 3806 3128 3808
rect 3128 3806 3145 3808
rect 3093 3766 3145 3806
rect 3093 3756 3094 3766
rect 3094 3756 3128 3766
rect 3128 3756 3145 3766
rect 3157 3806 3166 3808
rect 3166 3806 3200 3808
rect 3200 3806 3209 3808
rect 3157 3766 3209 3806
rect 3157 3756 3166 3766
rect 3166 3756 3200 3766
rect 3200 3756 3209 3766
rect 3221 3806 3238 3808
rect 3238 3806 3272 3808
rect 3272 3806 3273 3808
rect 3221 3766 3273 3806
rect 3221 3756 3238 3766
rect 3238 3756 3272 3766
rect 3272 3756 3273 3766
rect 3093 3732 3094 3743
rect 3094 3732 3128 3743
rect 3128 3732 3145 3743
rect 3093 3692 3145 3732
rect 3093 3691 3094 3692
rect 3094 3691 3128 3692
rect 3128 3691 3145 3692
rect 3157 3732 3166 3743
rect 3166 3732 3200 3743
rect 3200 3732 3209 3743
rect 3157 3692 3209 3732
rect 3157 3691 3166 3692
rect 3166 3691 3200 3692
rect 3200 3691 3209 3692
rect 3221 3732 3238 3743
rect 3238 3732 3272 3743
rect 3272 3732 3273 3743
rect 3221 3692 3273 3732
rect 3221 3691 3238 3692
rect 3238 3691 3272 3692
rect 3272 3691 3273 3692
rect 3093 3658 3094 3678
rect 3094 3658 3128 3678
rect 3128 3658 3145 3678
rect 3093 3626 3145 3658
rect 3157 3658 3166 3678
rect 3166 3658 3200 3678
rect 3200 3658 3209 3678
rect 3157 3626 3209 3658
rect 3221 3658 3238 3678
rect 3238 3658 3272 3678
rect 3272 3658 3273 3678
rect 3221 3626 3273 3658
rect 3093 3584 3094 3613
rect 3094 3584 3128 3613
rect 3128 3584 3145 3613
rect 3093 3561 3145 3584
rect 3157 3584 3166 3613
rect 3166 3584 3200 3613
rect 3200 3584 3209 3613
rect 3157 3561 3209 3584
rect 3221 3584 3238 3613
rect 3238 3584 3272 3613
rect 3272 3584 3273 3613
rect 3221 3561 3273 3584
rect 3093 3544 3145 3548
rect 3093 3510 3094 3544
rect 3094 3510 3128 3544
rect 3128 3510 3145 3544
rect 3093 3496 3145 3510
rect 3157 3544 3209 3548
rect 3157 3510 3166 3544
rect 3166 3510 3200 3544
rect 3200 3510 3209 3544
rect 3157 3496 3209 3510
rect 3221 3544 3273 3548
rect 3221 3510 3238 3544
rect 3238 3510 3272 3544
rect 3272 3510 3273 3544
rect 3221 3496 3273 3510
rect 3093 3470 3145 3483
rect 3093 3436 3094 3470
rect 3094 3436 3128 3470
rect 3128 3436 3145 3470
rect 3093 3431 3145 3436
rect 3157 3470 3209 3483
rect 3157 3436 3166 3470
rect 3166 3436 3200 3470
rect 3200 3436 3209 3470
rect 3157 3431 3209 3436
rect 3221 3470 3273 3483
rect 3221 3436 3238 3470
rect 3238 3436 3272 3470
rect 3272 3436 3273 3470
rect 3221 3431 3273 3436
rect 3093 3396 3145 3418
rect 3093 3366 3094 3396
rect 3094 3366 3128 3396
rect 3128 3366 3145 3396
rect 3157 3396 3209 3418
rect 3157 3366 3166 3396
rect 3166 3366 3200 3396
rect 3200 3366 3209 3396
rect 3221 3396 3273 3418
rect 3221 3366 3238 3396
rect 3238 3366 3272 3396
rect 3272 3366 3273 3396
rect 3093 3322 3145 3353
rect 3093 3301 3094 3322
rect 3094 3301 3128 3322
rect 3128 3301 3145 3322
rect 3157 3322 3209 3353
rect 3157 3301 3166 3322
rect 3166 3301 3200 3322
rect 3200 3301 3209 3322
rect 3221 3322 3273 3353
rect 3221 3301 3238 3322
rect 3238 3301 3272 3322
rect 3272 3301 3273 3322
rect 3093 3248 3145 3288
rect 3093 3236 3094 3248
rect 3094 3236 3128 3248
rect 3128 3236 3145 3248
rect 3157 3248 3209 3288
rect 3157 3236 3166 3248
rect 3166 3236 3200 3248
rect 3200 3236 3209 3248
rect 3221 3248 3273 3288
rect 3221 3236 3238 3248
rect 3238 3236 3272 3248
rect 3272 3236 3273 3248
rect 3093 3214 3094 3223
rect 3094 3214 3128 3223
rect 3128 3214 3145 3223
rect 3093 3174 3145 3214
rect 3093 3171 3094 3174
rect 3094 3171 3128 3174
rect 3128 3171 3145 3174
rect 3157 3214 3166 3223
rect 3166 3214 3200 3223
rect 3200 3214 3209 3223
rect 3157 3174 3209 3214
rect 3157 3171 3166 3174
rect 3166 3171 3200 3174
rect 3200 3171 3209 3174
rect 3221 3214 3238 3223
rect 3238 3214 3272 3223
rect 3272 3214 3273 3223
rect 3221 3174 3273 3214
rect 3221 3171 3238 3174
rect 3238 3171 3272 3174
rect 3272 3171 3273 3174
rect 3093 3140 3094 3158
rect 3094 3140 3128 3158
rect 3128 3140 3145 3158
rect 3093 3106 3145 3140
rect 3157 3140 3166 3158
rect 3166 3140 3200 3158
rect 3200 3140 3209 3158
rect 3157 3106 3209 3140
rect 3221 3140 3238 3158
rect 3238 3140 3272 3158
rect 3272 3140 3273 3158
rect 3221 3106 3273 3140
rect 3093 3066 3094 3093
rect 3094 3066 3128 3093
rect 3128 3066 3145 3093
rect 3093 3041 3145 3066
rect 3157 3066 3166 3093
rect 3166 3066 3200 3093
rect 3200 3066 3209 3093
rect 3157 3041 3209 3066
rect 3221 3066 3238 3093
rect 3238 3066 3272 3093
rect 3272 3066 3273 3093
rect 3221 3041 3273 3066
rect 3093 3026 3145 3028
rect 3093 2992 3094 3026
rect 3094 2992 3128 3026
rect 3128 2992 3145 3026
rect 3093 2976 3145 2992
rect 3157 3026 3209 3028
rect 3157 2992 3166 3026
rect 3166 2992 3200 3026
rect 3200 2992 3209 3026
rect 3157 2976 3209 2992
rect 3221 3026 3273 3028
rect 3221 2992 3238 3026
rect 3238 2992 3272 3026
rect 3272 2992 3273 3026
rect 3221 2976 3273 2992
rect 3093 2952 3145 2963
rect 3093 2918 3094 2952
rect 3094 2918 3128 2952
rect 3128 2918 3145 2952
rect 3093 2911 3145 2918
rect 3157 2952 3209 2963
rect 3157 2918 3166 2952
rect 3166 2918 3200 2952
rect 3200 2918 3209 2952
rect 3157 2911 3209 2918
rect 3221 2952 3273 2963
rect 3221 2918 3238 2952
rect 3238 2918 3272 2952
rect 3272 2918 3273 2952
rect 3221 2911 3273 2918
rect 3093 2878 3145 2898
rect 3093 2846 3094 2878
rect 3094 2846 3128 2878
rect 3128 2846 3145 2878
rect 3157 2878 3209 2898
rect 3157 2846 3166 2878
rect 3166 2846 3200 2878
rect 3200 2846 3209 2878
rect 3221 2878 3273 2898
rect 3221 2846 3238 2878
rect 3238 2846 3272 2878
rect 3272 2846 3273 2878
rect 3093 2804 3145 2833
rect 3093 2781 3094 2804
rect 3094 2781 3128 2804
rect 3128 2781 3145 2804
rect 3157 2804 3209 2833
rect 3157 2781 3166 2804
rect 3166 2781 3200 2804
rect 3200 2781 3209 2804
rect 3221 2804 3273 2833
rect 3221 2781 3238 2804
rect 3238 2781 3272 2804
rect 3272 2781 3273 2804
rect 3093 2730 3145 2768
rect 3093 2716 3094 2730
rect 3094 2716 3128 2730
rect 3128 2716 3145 2730
rect 3157 2730 3209 2768
rect 3157 2716 3166 2730
rect 3166 2716 3200 2730
rect 3200 2716 3209 2730
rect 3221 2730 3273 2768
rect 3221 2716 3238 2730
rect 3238 2716 3272 2730
rect 3272 2716 3273 2730
rect 3093 2696 3094 2703
rect 3094 2696 3128 2703
rect 3128 2696 3145 2703
rect 3093 2656 3145 2696
rect 3093 2651 3094 2656
rect 3094 2651 3128 2656
rect 3128 2651 3145 2656
rect 3157 2696 3166 2703
rect 3166 2696 3200 2703
rect 3200 2696 3209 2703
rect 3157 2656 3209 2696
rect 3157 2651 3166 2656
rect 3166 2651 3200 2656
rect 3200 2651 3209 2656
rect 3221 2696 3238 2703
rect 3238 2696 3272 2703
rect 3272 2696 3273 2703
rect 3221 2656 3273 2696
rect 3221 2651 3238 2656
rect 3238 2651 3272 2656
rect 3272 2651 3273 2656
rect 3093 2622 3094 2638
rect 3094 2622 3128 2638
rect 3128 2622 3145 2638
rect 3093 2586 3145 2622
rect 3157 2622 3166 2638
rect 3166 2622 3200 2638
rect 3200 2622 3209 2638
rect 3157 2586 3209 2622
rect 3221 2622 3238 2638
rect 3238 2622 3272 2638
rect 3272 2622 3273 2638
rect 3221 2586 3273 2622
rect 3093 2548 3094 2573
rect 3094 2548 3128 2573
rect 3128 2548 3145 2573
rect 3093 2521 3145 2548
rect 3157 2548 3166 2573
rect 3166 2548 3200 2573
rect 3200 2548 3209 2573
rect 3157 2521 3209 2548
rect 3221 2548 3238 2573
rect 3238 2548 3272 2573
rect 3272 2548 3273 2573
rect 3221 2521 3273 2548
rect 3093 2474 3094 2508
rect 3094 2474 3128 2508
rect 3128 2474 3145 2508
rect 3093 2456 3145 2474
rect 3157 2474 3166 2508
rect 3166 2474 3200 2508
rect 3200 2474 3209 2508
rect 3157 2456 3209 2474
rect 3221 2474 3238 2508
rect 3238 2474 3272 2508
rect 3272 2474 3273 2508
rect 3221 2456 3273 2474
rect 3093 2434 3145 2443
rect 3093 2400 3094 2434
rect 3094 2400 3128 2434
rect 3128 2400 3145 2434
rect 3093 2391 3145 2400
rect 3157 2434 3209 2443
rect 3157 2400 3166 2434
rect 3166 2400 3200 2434
rect 3200 2400 3209 2434
rect 3157 2391 3209 2400
rect 3221 2434 3273 2443
rect 3221 2400 3238 2434
rect 3238 2400 3272 2434
rect 3272 2400 3273 2434
rect 3221 2391 3273 2400
rect 3093 2360 3145 2378
rect 3093 2326 3094 2360
rect 3094 2326 3128 2360
rect 3128 2326 3145 2360
rect 3157 2360 3209 2378
rect 3157 2326 3166 2360
rect 3166 2326 3200 2360
rect 3200 2326 3209 2360
rect 3221 2360 3273 2378
rect 3221 2326 3238 2360
rect 3238 2326 3272 2360
rect 3272 2326 3273 2360
rect 3093 2286 3145 2313
rect 3093 2261 3094 2286
rect 3094 2261 3128 2286
rect 3128 2261 3145 2286
rect 3157 2286 3209 2313
rect 3157 2261 3166 2286
rect 3166 2261 3200 2286
rect 3200 2261 3209 2286
rect 3221 2286 3273 2313
rect 3221 2261 3238 2286
rect 3238 2261 3272 2286
rect 3272 2261 3273 2286
rect 3093 2212 3145 2248
rect 3093 2196 3094 2212
rect 3094 2196 3128 2212
rect 3128 2196 3145 2212
rect 3157 2212 3209 2248
rect 3157 2196 3166 2212
rect 3166 2196 3200 2212
rect 3200 2196 3209 2212
rect 3221 2212 3273 2248
rect 3221 2196 3238 2212
rect 3238 2196 3272 2212
rect 3272 2196 3273 2212
rect 3093 2178 3094 2183
rect 3094 2178 3128 2183
rect 3128 2178 3145 2183
rect 3093 2138 3145 2178
rect 3093 2131 3094 2138
rect 3094 2131 3128 2138
rect 3128 2131 3145 2138
rect 3157 2178 3166 2183
rect 3166 2178 3200 2183
rect 3200 2178 3209 2183
rect 3157 2138 3209 2178
rect 3157 2131 3166 2138
rect 3166 2131 3200 2138
rect 3200 2131 3209 2138
rect 3221 2178 3238 2183
rect 3238 2178 3272 2183
rect 3272 2178 3273 2183
rect 3221 2138 3273 2178
rect 3221 2131 3238 2138
rect 3238 2131 3272 2138
rect 3272 2131 3273 2138
rect 3093 2104 3094 2118
rect 3094 2104 3128 2118
rect 3128 2104 3145 2118
rect 3093 2066 3145 2104
rect 3157 2104 3166 2118
rect 3166 2104 3200 2118
rect 3200 2104 3209 2118
rect 3157 2066 3209 2104
rect 3221 2104 3238 2118
rect 3238 2104 3272 2118
rect 3272 2104 3273 2118
rect 3221 2066 3273 2104
rect 3093 2030 3094 2053
rect 3094 2030 3128 2053
rect 3128 2030 3145 2053
rect 3093 2001 3145 2030
rect 3157 2030 3166 2053
rect 3166 2030 3200 2053
rect 3200 2030 3209 2053
rect 3157 2001 3209 2030
rect 3221 2030 3238 2053
rect 3238 2030 3272 2053
rect 3272 2030 3273 2053
rect 3221 2001 3273 2030
rect 3093 1956 3094 1987
rect 3094 1956 3128 1987
rect 3128 1956 3145 1987
rect 3093 1935 3145 1956
rect 3157 1956 3166 1987
rect 3166 1956 3200 1987
rect 3200 1956 3209 1987
rect 3157 1935 3209 1956
rect 3221 1956 3238 1987
rect 3238 1956 3272 1987
rect 3272 1956 3273 1987
rect 3221 1935 3273 1956
rect 3093 1916 3145 1921
rect 3093 1882 3094 1916
rect 3094 1882 3128 1916
rect 3128 1882 3145 1916
rect 3093 1869 3145 1882
rect 3157 1916 3209 1921
rect 3157 1882 3166 1916
rect 3166 1882 3200 1916
rect 3200 1882 3209 1916
rect 3157 1869 3209 1882
rect 3221 1916 3273 1921
rect 3221 1882 3238 1916
rect 3238 1882 3272 1916
rect 3272 1882 3273 1916
rect 3221 1869 3273 1882
rect 3093 1842 3145 1855
rect 3093 1808 3094 1842
rect 3094 1808 3128 1842
rect 3128 1808 3145 1842
rect 3093 1803 3145 1808
rect 3157 1842 3209 1855
rect 3157 1808 3166 1842
rect 3166 1808 3200 1842
rect 3200 1808 3209 1842
rect 3157 1803 3209 1808
rect 3221 1842 3273 1855
rect 3221 1808 3238 1842
rect 3238 1808 3272 1842
rect 3272 1808 3273 1842
rect 3221 1803 3273 1808
rect 3093 1768 3145 1789
rect 3093 1737 3094 1768
rect 3094 1737 3128 1768
rect 3128 1737 3145 1768
rect 3157 1768 3209 1789
rect 3157 1737 3166 1768
rect 3166 1737 3200 1768
rect 3200 1737 3209 1768
rect 3221 1768 3273 1789
rect 3221 1737 3238 1768
rect 3238 1737 3272 1768
rect 3272 1737 3273 1768
rect 3093 1694 3145 1723
rect 3093 1671 3094 1694
rect 3094 1671 3128 1694
rect 3128 1671 3145 1694
rect 3157 1694 3209 1723
rect 3157 1671 3166 1694
rect 3166 1671 3200 1694
rect 3200 1671 3209 1694
rect 3221 1694 3273 1723
rect 3221 1671 3238 1694
rect 3238 1671 3272 1694
rect 3272 1671 3273 1694
rect 3093 1620 3145 1657
rect 3093 1605 3094 1620
rect 3094 1605 3128 1620
rect 3128 1605 3145 1620
rect 3157 1620 3209 1657
rect 3157 1605 3166 1620
rect 3166 1605 3200 1620
rect 3200 1605 3209 1620
rect 3221 1620 3273 1657
rect 3221 1605 3238 1620
rect 3238 1605 3272 1620
rect 3272 1605 3273 1620
rect 3093 1586 3094 1591
rect 3094 1586 3128 1591
rect 3128 1586 3145 1591
rect 3093 1545 3145 1586
rect 3093 1539 3094 1545
rect 3094 1539 3128 1545
rect 3128 1539 3145 1545
rect 3157 1586 3166 1591
rect 3166 1586 3200 1591
rect 3200 1586 3209 1591
rect 3157 1545 3209 1586
rect 3157 1539 3166 1545
rect 3166 1539 3200 1545
rect 3200 1539 3209 1545
rect 3221 1586 3238 1591
rect 3238 1586 3272 1591
rect 3272 1586 3273 1591
rect 3221 1545 3273 1586
rect 3221 1539 3238 1545
rect 3238 1539 3272 1545
rect 3272 1539 3273 1545
rect 3093 1511 3094 1525
rect 3094 1511 3128 1525
rect 3128 1511 3145 1525
rect 3093 1473 3145 1511
rect 3157 1511 3166 1525
rect 3166 1511 3200 1525
rect 3200 1511 3209 1525
rect 3157 1473 3209 1511
rect 3221 1511 3238 1525
rect 3238 1511 3272 1525
rect 3272 1511 3273 1525
rect 3221 1473 3273 1511
rect 3589 4050 3641 4068
rect 3653 4062 3705 4068
rect 3653 4050 3662 4062
rect 3662 4050 3696 4062
rect 3696 4050 3705 4062
rect 3717 4050 3769 4068
rect 3589 4016 3590 4050
rect 3590 4016 3641 4050
rect 3653 4016 3705 4050
rect 3717 4016 3768 4050
rect 3768 4016 3769 4050
rect 3589 3951 3590 4003
rect 3590 3951 3641 4003
rect 3653 3951 3705 4003
rect 3717 3951 3768 4003
rect 3768 3951 3769 4003
rect 3589 3886 3590 3938
rect 3590 3886 3641 3938
rect 3653 3886 3705 3938
rect 3717 3886 3768 3938
rect 3768 3886 3769 3938
rect 3589 3821 3590 3873
rect 3590 3821 3641 3873
rect 3653 3821 3705 3873
rect 3717 3821 3768 3873
rect 3768 3821 3769 3873
rect 3589 3756 3590 3808
rect 3590 3756 3641 3808
rect 3653 3756 3705 3808
rect 3717 3756 3768 3808
rect 3768 3756 3769 3808
rect 3589 3691 3590 3743
rect 3590 3691 3641 3743
rect 3653 3691 3705 3743
rect 3717 3691 3768 3743
rect 3768 3691 3769 3743
rect 3589 3626 3590 3678
rect 3590 3626 3641 3678
rect 3653 3626 3705 3678
rect 3717 3626 3768 3678
rect 3768 3626 3769 3678
rect 3589 3561 3590 3613
rect 3590 3561 3641 3613
rect 3653 3561 3705 3613
rect 3717 3561 3768 3613
rect 3768 3561 3769 3613
rect 3589 3496 3590 3548
rect 3590 3496 3641 3548
rect 3653 3496 3705 3548
rect 3717 3496 3768 3548
rect 3768 3496 3769 3548
rect 3589 3431 3590 3483
rect 3590 3431 3641 3483
rect 3653 3431 3705 3483
rect 3717 3431 3768 3483
rect 3768 3431 3769 3483
rect 3589 3366 3590 3418
rect 3590 3366 3641 3418
rect 3653 3366 3705 3418
rect 3717 3366 3768 3418
rect 3768 3366 3769 3418
rect 3589 3301 3590 3353
rect 3590 3301 3641 3353
rect 3653 3301 3705 3353
rect 3717 3301 3768 3353
rect 3768 3301 3769 3353
rect 3589 3236 3590 3288
rect 3590 3236 3641 3288
rect 3653 3236 3705 3288
rect 3717 3236 3768 3288
rect 3768 3236 3769 3288
rect 3589 3171 3590 3223
rect 3590 3171 3641 3223
rect 3653 3171 3705 3223
rect 3717 3171 3768 3223
rect 3768 3171 3769 3223
rect 3589 3106 3590 3158
rect 3590 3106 3641 3158
rect 3653 3106 3705 3158
rect 3717 3106 3768 3158
rect 3768 3106 3769 3158
rect 3589 3080 3590 3093
rect 3590 3092 3641 3093
rect 3653 3092 3705 3093
rect 3717 3092 3768 3093
rect 3590 3080 3624 3092
rect 3624 3080 3641 3092
rect 3589 3041 3641 3080
rect 3653 3041 3705 3092
rect 3717 3080 3734 3092
rect 3734 3080 3768 3092
rect 3768 3080 3769 3093
rect 3717 3041 3769 3080
rect 3589 2976 3590 3028
rect 3590 2976 3641 3028
rect 3653 2976 3705 3028
rect 3717 2976 3768 3028
rect 3768 2976 3769 3028
rect 3589 2911 3590 2963
rect 3590 2911 3641 2963
rect 3653 2911 3705 2963
rect 3717 2911 3768 2963
rect 3768 2911 3769 2963
rect 3589 2846 3590 2898
rect 3590 2846 3641 2898
rect 3653 2846 3705 2898
rect 3717 2846 3768 2898
rect 3768 2846 3769 2898
rect 3589 2781 3590 2833
rect 3590 2781 3641 2833
rect 3653 2781 3705 2833
rect 3717 2781 3768 2833
rect 3768 2781 3769 2833
rect 3589 2716 3590 2768
rect 3590 2716 3641 2768
rect 3653 2716 3705 2768
rect 3717 2716 3768 2768
rect 3768 2716 3769 2768
rect 3589 2651 3590 2703
rect 3590 2651 3641 2703
rect 3653 2651 3705 2703
rect 3717 2651 3768 2703
rect 3768 2651 3769 2703
rect 3589 2586 3590 2638
rect 3590 2586 3641 2638
rect 3653 2586 3705 2638
rect 3717 2586 3768 2638
rect 3768 2586 3769 2638
rect 3589 2535 3641 2573
rect 3589 2521 3590 2535
rect 3590 2521 3624 2535
rect 3624 2521 3641 2535
rect 3653 2535 3705 2573
rect 3653 2521 3662 2535
rect 3662 2521 3696 2535
rect 3696 2521 3705 2535
rect 3717 2535 3769 2573
rect 3717 2521 3734 2535
rect 3734 2521 3768 2535
rect 3768 2521 3769 2535
rect 3589 2501 3590 2508
rect 3590 2501 3624 2508
rect 3624 2501 3641 2508
rect 3589 2456 3641 2501
rect 3653 2501 3662 2508
rect 3662 2501 3696 2508
rect 3696 2501 3705 2508
rect 3653 2461 3705 2501
rect 3653 2456 3662 2461
rect 3662 2456 3696 2461
rect 3696 2456 3705 2461
rect 3717 2501 3734 2508
rect 3734 2501 3768 2508
rect 3768 2501 3769 2508
rect 3717 2456 3769 2501
rect 3589 2391 3590 2443
rect 3590 2391 3641 2443
rect 3653 2391 3705 2443
rect 3717 2391 3768 2443
rect 3768 2391 3769 2443
rect 3589 2326 3590 2378
rect 3590 2326 3641 2378
rect 3653 2326 3705 2378
rect 3717 2326 3768 2378
rect 3768 2326 3769 2378
rect 3589 2261 3590 2313
rect 3590 2261 3641 2313
rect 3653 2261 3705 2313
rect 3717 2261 3768 2313
rect 3768 2261 3769 2313
rect 3589 2196 3590 2248
rect 3590 2196 3641 2248
rect 3653 2196 3705 2248
rect 3717 2196 3768 2248
rect 3768 2196 3769 2248
rect 3589 2131 3590 2183
rect 3590 2131 3641 2183
rect 3653 2131 3705 2183
rect 3717 2131 3768 2183
rect 3768 2131 3769 2183
rect 3589 2066 3590 2118
rect 3590 2066 3641 2118
rect 3653 2066 3705 2118
rect 3717 2066 3768 2118
rect 3768 2066 3769 2118
rect 3589 2001 3590 2053
rect 3590 2001 3641 2053
rect 3653 2001 3705 2053
rect 3717 2001 3768 2053
rect 3768 2001 3769 2053
rect 3589 1935 3590 1987
rect 3590 1935 3641 1987
rect 3653 1935 3705 1987
rect 3717 1935 3768 1987
rect 3768 1935 3769 1987
rect 3589 1869 3590 1921
rect 3590 1869 3641 1921
rect 3653 1869 3705 1921
rect 3717 1869 3768 1921
rect 3768 1869 3769 1921
rect 3589 1803 3590 1855
rect 3590 1803 3641 1855
rect 3653 1803 3705 1855
rect 3717 1803 3768 1855
rect 3768 1803 3769 1855
rect 3589 1737 3590 1789
rect 3590 1737 3641 1789
rect 3653 1737 3705 1789
rect 3717 1737 3768 1789
rect 3768 1737 3769 1789
rect 3589 1671 3590 1723
rect 3590 1671 3641 1723
rect 3653 1671 3705 1723
rect 3717 1671 3768 1723
rect 3768 1671 3769 1723
rect 3589 1605 3590 1657
rect 3590 1605 3641 1657
rect 3653 1605 3705 1657
rect 3717 1605 3768 1657
rect 3768 1605 3769 1657
rect 3589 1539 3590 1591
rect 3590 1539 3641 1591
rect 3653 1539 3705 1591
rect 3717 1539 3768 1591
rect 3768 1539 3769 1591
rect 3589 1479 3590 1525
rect 3590 1491 3641 1525
rect 3653 1491 3705 1525
rect 3717 1491 3768 1525
rect 3590 1479 3624 1491
rect 3624 1479 3641 1491
rect 3589 1473 3641 1479
rect 3653 1473 3705 1491
rect 3717 1479 3734 1491
rect 3734 1479 3768 1491
rect 3768 1479 3769 1525
rect 3717 1473 3769 1479
rect 4085 4062 4137 4068
rect 4085 4028 4086 4062
rect 4086 4028 4120 4062
rect 4120 4028 4137 4062
rect 4085 4016 4137 4028
rect 4149 4062 4201 4068
rect 4149 4028 4158 4062
rect 4158 4028 4192 4062
rect 4192 4028 4201 4062
rect 4149 4016 4201 4028
rect 4213 4062 4265 4068
rect 4213 4028 4230 4062
rect 4230 4028 4264 4062
rect 4264 4028 4265 4062
rect 4213 4016 4265 4028
rect 4085 3988 4137 4003
rect 4085 3954 4086 3988
rect 4086 3954 4120 3988
rect 4120 3954 4137 3988
rect 4085 3951 4137 3954
rect 4149 3988 4201 4003
rect 4149 3954 4158 3988
rect 4158 3954 4192 3988
rect 4192 3954 4201 3988
rect 4149 3951 4201 3954
rect 4213 3988 4265 4003
rect 4213 3954 4230 3988
rect 4230 3954 4264 3988
rect 4264 3954 4265 3988
rect 4213 3951 4265 3954
rect 4085 3914 4137 3938
rect 4085 3886 4086 3914
rect 4086 3886 4120 3914
rect 4120 3886 4137 3914
rect 4149 3914 4201 3938
rect 4149 3886 4158 3914
rect 4158 3886 4192 3914
rect 4192 3886 4201 3914
rect 4213 3914 4265 3938
rect 4213 3886 4230 3914
rect 4230 3886 4264 3914
rect 4264 3886 4265 3914
rect 4085 3840 4137 3873
rect 4085 3821 4086 3840
rect 4086 3821 4120 3840
rect 4120 3821 4137 3840
rect 4149 3840 4201 3873
rect 4149 3821 4158 3840
rect 4158 3821 4192 3840
rect 4192 3821 4201 3840
rect 4213 3840 4265 3873
rect 4213 3821 4230 3840
rect 4230 3821 4264 3840
rect 4264 3821 4265 3840
rect 4085 3806 4086 3808
rect 4086 3806 4120 3808
rect 4120 3806 4137 3808
rect 4085 3766 4137 3806
rect 4085 3756 4086 3766
rect 4086 3756 4120 3766
rect 4120 3756 4137 3766
rect 4149 3806 4158 3808
rect 4158 3806 4192 3808
rect 4192 3806 4201 3808
rect 4149 3766 4201 3806
rect 4149 3756 4158 3766
rect 4158 3756 4192 3766
rect 4192 3756 4201 3766
rect 4213 3806 4230 3808
rect 4230 3806 4264 3808
rect 4264 3806 4265 3808
rect 4213 3766 4265 3806
rect 4213 3756 4230 3766
rect 4230 3756 4264 3766
rect 4264 3756 4265 3766
rect 4085 3732 4086 3743
rect 4086 3732 4120 3743
rect 4120 3732 4137 3743
rect 4085 3692 4137 3732
rect 4085 3691 4086 3692
rect 4086 3691 4120 3692
rect 4120 3691 4137 3692
rect 4149 3732 4158 3743
rect 4158 3732 4192 3743
rect 4192 3732 4201 3743
rect 4149 3692 4201 3732
rect 4149 3691 4158 3692
rect 4158 3691 4192 3692
rect 4192 3691 4201 3692
rect 4213 3732 4230 3743
rect 4230 3732 4264 3743
rect 4264 3732 4265 3743
rect 4213 3692 4265 3732
rect 4213 3691 4230 3692
rect 4230 3691 4264 3692
rect 4264 3691 4265 3692
rect 4085 3658 4086 3678
rect 4086 3658 4120 3678
rect 4120 3658 4137 3678
rect 4085 3626 4137 3658
rect 4149 3658 4158 3678
rect 4158 3658 4192 3678
rect 4192 3658 4201 3678
rect 4149 3626 4201 3658
rect 4213 3658 4230 3678
rect 4230 3658 4264 3678
rect 4264 3658 4265 3678
rect 4213 3626 4265 3658
rect 4085 3584 4086 3613
rect 4086 3584 4120 3613
rect 4120 3584 4137 3613
rect 4085 3561 4137 3584
rect 4149 3584 4158 3613
rect 4158 3584 4192 3613
rect 4192 3584 4201 3613
rect 4149 3561 4201 3584
rect 4213 3584 4230 3613
rect 4230 3584 4264 3613
rect 4264 3584 4265 3613
rect 4213 3561 4265 3584
rect 4085 3544 4137 3548
rect 4085 3510 4086 3544
rect 4086 3510 4120 3544
rect 4120 3510 4137 3544
rect 4085 3496 4137 3510
rect 4149 3544 4201 3548
rect 4149 3510 4158 3544
rect 4158 3510 4192 3544
rect 4192 3510 4201 3544
rect 4149 3496 4201 3510
rect 4213 3544 4265 3548
rect 4213 3510 4230 3544
rect 4230 3510 4264 3544
rect 4264 3510 4265 3544
rect 4213 3496 4265 3510
rect 4085 3470 4137 3483
rect 4085 3436 4086 3470
rect 4086 3436 4120 3470
rect 4120 3436 4137 3470
rect 4085 3431 4137 3436
rect 4149 3470 4201 3483
rect 4149 3436 4158 3470
rect 4158 3436 4192 3470
rect 4192 3436 4201 3470
rect 4149 3431 4201 3436
rect 4213 3470 4265 3483
rect 4213 3436 4230 3470
rect 4230 3436 4264 3470
rect 4264 3436 4265 3470
rect 4213 3431 4265 3436
rect 4085 3396 4137 3418
rect 4085 3366 4086 3396
rect 4086 3366 4120 3396
rect 4120 3366 4137 3396
rect 4149 3396 4201 3418
rect 4149 3366 4158 3396
rect 4158 3366 4192 3396
rect 4192 3366 4201 3396
rect 4213 3396 4265 3418
rect 4213 3366 4230 3396
rect 4230 3366 4264 3396
rect 4264 3366 4265 3396
rect 4085 3322 4137 3353
rect 4085 3301 4086 3322
rect 4086 3301 4120 3322
rect 4120 3301 4137 3322
rect 4149 3322 4201 3353
rect 4149 3301 4158 3322
rect 4158 3301 4192 3322
rect 4192 3301 4201 3322
rect 4213 3322 4265 3353
rect 4213 3301 4230 3322
rect 4230 3301 4264 3322
rect 4264 3301 4265 3322
rect 4085 3248 4137 3288
rect 4085 3236 4086 3248
rect 4086 3236 4120 3248
rect 4120 3236 4137 3248
rect 4149 3248 4201 3288
rect 4149 3236 4158 3248
rect 4158 3236 4192 3248
rect 4192 3236 4201 3248
rect 4213 3248 4265 3288
rect 4213 3236 4230 3248
rect 4230 3236 4264 3248
rect 4264 3236 4265 3248
rect 4085 3214 4086 3223
rect 4086 3214 4120 3223
rect 4120 3214 4137 3223
rect 4085 3174 4137 3214
rect 4085 3171 4086 3174
rect 4086 3171 4120 3174
rect 4120 3171 4137 3174
rect 4149 3214 4158 3223
rect 4158 3214 4192 3223
rect 4192 3214 4201 3223
rect 4149 3174 4201 3214
rect 4149 3171 4158 3174
rect 4158 3171 4192 3174
rect 4192 3171 4201 3174
rect 4213 3214 4230 3223
rect 4230 3214 4264 3223
rect 4264 3214 4265 3223
rect 4213 3174 4265 3214
rect 4213 3171 4230 3174
rect 4230 3171 4264 3174
rect 4264 3171 4265 3174
rect 4085 3140 4086 3158
rect 4086 3140 4120 3158
rect 4120 3140 4137 3158
rect 4085 3106 4137 3140
rect 4149 3140 4158 3158
rect 4158 3140 4192 3158
rect 4192 3140 4201 3158
rect 4149 3106 4201 3140
rect 4213 3140 4230 3158
rect 4230 3140 4264 3158
rect 4264 3140 4265 3158
rect 4213 3106 4265 3140
rect 4085 3066 4086 3093
rect 4086 3066 4120 3093
rect 4120 3066 4137 3093
rect 4085 3041 4137 3066
rect 4149 3066 4158 3093
rect 4158 3066 4192 3093
rect 4192 3066 4201 3093
rect 4149 3041 4201 3066
rect 4213 3066 4230 3093
rect 4230 3066 4264 3093
rect 4264 3066 4265 3093
rect 4213 3041 4265 3066
rect 4085 3026 4137 3028
rect 4085 2992 4086 3026
rect 4086 2992 4120 3026
rect 4120 2992 4137 3026
rect 4085 2976 4137 2992
rect 4149 3026 4201 3028
rect 4149 2992 4158 3026
rect 4158 2992 4192 3026
rect 4192 2992 4201 3026
rect 4149 2976 4201 2992
rect 4213 3026 4265 3028
rect 4213 2992 4230 3026
rect 4230 2992 4264 3026
rect 4264 2992 4265 3026
rect 4213 2976 4265 2992
rect 4085 2952 4137 2963
rect 4085 2918 4086 2952
rect 4086 2918 4120 2952
rect 4120 2918 4137 2952
rect 4085 2911 4137 2918
rect 4149 2952 4201 2963
rect 4149 2918 4158 2952
rect 4158 2918 4192 2952
rect 4192 2918 4201 2952
rect 4149 2911 4201 2918
rect 4213 2952 4265 2963
rect 4213 2918 4230 2952
rect 4230 2918 4264 2952
rect 4264 2918 4265 2952
rect 4213 2911 4265 2918
rect 4085 2878 4137 2898
rect 4085 2846 4086 2878
rect 4086 2846 4120 2878
rect 4120 2846 4137 2878
rect 4149 2878 4201 2898
rect 4149 2846 4158 2878
rect 4158 2846 4192 2878
rect 4192 2846 4201 2878
rect 4213 2878 4265 2898
rect 4213 2846 4230 2878
rect 4230 2846 4264 2878
rect 4264 2846 4265 2878
rect 4085 2804 4137 2833
rect 4085 2781 4086 2804
rect 4086 2781 4120 2804
rect 4120 2781 4137 2804
rect 4149 2804 4201 2833
rect 4149 2781 4158 2804
rect 4158 2781 4192 2804
rect 4192 2781 4201 2804
rect 4213 2804 4265 2833
rect 4213 2781 4230 2804
rect 4230 2781 4264 2804
rect 4264 2781 4265 2804
rect 4085 2730 4137 2768
rect 4085 2716 4086 2730
rect 4086 2716 4120 2730
rect 4120 2716 4137 2730
rect 4149 2730 4201 2768
rect 4149 2716 4158 2730
rect 4158 2716 4192 2730
rect 4192 2716 4201 2730
rect 4213 2730 4265 2768
rect 4213 2716 4230 2730
rect 4230 2716 4264 2730
rect 4264 2716 4265 2730
rect 4085 2696 4086 2703
rect 4086 2696 4120 2703
rect 4120 2696 4137 2703
rect 4085 2656 4137 2696
rect 4085 2651 4086 2656
rect 4086 2651 4120 2656
rect 4120 2651 4137 2656
rect 4149 2696 4158 2703
rect 4158 2696 4192 2703
rect 4192 2696 4201 2703
rect 4149 2656 4201 2696
rect 4149 2651 4158 2656
rect 4158 2651 4192 2656
rect 4192 2651 4201 2656
rect 4213 2696 4230 2703
rect 4230 2696 4264 2703
rect 4264 2696 4265 2703
rect 4213 2656 4265 2696
rect 4213 2651 4230 2656
rect 4230 2651 4264 2656
rect 4264 2651 4265 2656
rect 4085 2622 4086 2638
rect 4086 2622 4120 2638
rect 4120 2622 4137 2638
rect 4085 2586 4137 2622
rect 4149 2622 4158 2638
rect 4158 2622 4192 2638
rect 4192 2622 4201 2638
rect 4149 2586 4201 2622
rect 4213 2622 4230 2638
rect 4230 2622 4264 2638
rect 4264 2622 4265 2638
rect 4213 2586 4265 2622
rect 4085 2548 4086 2573
rect 4086 2548 4120 2573
rect 4120 2548 4137 2573
rect 4085 2521 4137 2548
rect 4149 2548 4158 2573
rect 4158 2548 4192 2573
rect 4192 2548 4201 2573
rect 4149 2521 4201 2548
rect 4213 2548 4230 2573
rect 4230 2548 4264 2573
rect 4264 2548 4265 2573
rect 4213 2521 4265 2548
rect 4085 2474 4086 2508
rect 4086 2474 4120 2508
rect 4120 2474 4137 2508
rect 4085 2456 4137 2474
rect 4149 2474 4158 2508
rect 4158 2474 4192 2508
rect 4192 2474 4201 2508
rect 4149 2456 4201 2474
rect 4213 2474 4230 2508
rect 4230 2474 4264 2508
rect 4264 2474 4265 2508
rect 4213 2456 4265 2474
rect 4085 2434 4137 2443
rect 4085 2400 4086 2434
rect 4086 2400 4120 2434
rect 4120 2400 4137 2434
rect 4085 2391 4137 2400
rect 4149 2434 4201 2443
rect 4149 2400 4158 2434
rect 4158 2400 4192 2434
rect 4192 2400 4201 2434
rect 4149 2391 4201 2400
rect 4213 2434 4265 2443
rect 4213 2400 4230 2434
rect 4230 2400 4264 2434
rect 4264 2400 4265 2434
rect 4213 2391 4265 2400
rect 4085 2360 4137 2378
rect 4085 2326 4086 2360
rect 4086 2326 4120 2360
rect 4120 2326 4137 2360
rect 4149 2360 4201 2378
rect 4149 2326 4158 2360
rect 4158 2326 4192 2360
rect 4192 2326 4201 2360
rect 4213 2360 4265 2378
rect 4213 2326 4230 2360
rect 4230 2326 4264 2360
rect 4264 2326 4265 2360
rect 4085 2286 4137 2313
rect 4085 2261 4086 2286
rect 4086 2261 4120 2286
rect 4120 2261 4137 2286
rect 4149 2286 4201 2313
rect 4149 2261 4158 2286
rect 4158 2261 4192 2286
rect 4192 2261 4201 2286
rect 4213 2286 4265 2313
rect 4213 2261 4230 2286
rect 4230 2261 4264 2286
rect 4264 2261 4265 2286
rect 4085 2212 4137 2248
rect 4085 2196 4086 2212
rect 4086 2196 4120 2212
rect 4120 2196 4137 2212
rect 4149 2212 4201 2248
rect 4149 2196 4158 2212
rect 4158 2196 4192 2212
rect 4192 2196 4201 2212
rect 4213 2212 4265 2248
rect 4213 2196 4230 2212
rect 4230 2196 4264 2212
rect 4264 2196 4265 2212
rect 4085 2178 4086 2183
rect 4086 2178 4120 2183
rect 4120 2178 4137 2183
rect 4085 2138 4137 2178
rect 4085 2131 4086 2138
rect 4086 2131 4120 2138
rect 4120 2131 4137 2138
rect 4149 2178 4158 2183
rect 4158 2178 4192 2183
rect 4192 2178 4201 2183
rect 4149 2138 4201 2178
rect 4149 2131 4158 2138
rect 4158 2131 4192 2138
rect 4192 2131 4201 2138
rect 4213 2178 4230 2183
rect 4230 2178 4264 2183
rect 4264 2178 4265 2183
rect 4213 2138 4265 2178
rect 4213 2131 4230 2138
rect 4230 2131 4264 2138
rect 4264 2131 4265 2138
rect 4085 2104 4086 2118
rect 4086 2104 4120 2118
rect 4120 2104 4137 2118
rect 4085 2066 4137 2104
rect 4149 2104 4158 2118
rect 4158 2104 4192 2118
rect 4192 2104 4201 2118
rect 4149 2066 4201 2104
rect 4213 2104 4230 2118
rect 4230 2104 4264 2118
rect 4264 2104 4265 2118
rect 4213 2066 4265 2104
rect 4085 2030 4086 2053
rect 4086 2030 4120 2053
rect 4120 2030 4137 2053
rect 4085 2001 4137 2030
rect 4149 2030 4158 2053
rect 4158 2030 4192 2053
rect 4192 2030 4201 2053
rect 4149 2001 4201 2030
rect 4213 2030 4230 2053
rect 4230 2030 4264 2053
rect 4264 2030 4265 2053
rect 4213 2001 4265 2030
rect 4085 1956 4086 1987
rect 4086 1956 4120 1987
rect 4120 1956 4137 1987
rect 4085 1935 4137 1956
rect 4149 1956 4158 1987
rect 4158 1956 4192 1987
rect 4192 1956 4201 1987
rect 4149 1935 4201 1956
rect 4213 1956 4230 1987
rect 4230 1956 4264 1987
rect 4264 1956 4265 1987
rect 4213 1935 4265 1956
rect 4085 1916 4137 1921
rect 4085 1882 4086 1916
rect 4086 1882 4120 1916
rect 4120 1882 4137 1916
rect 4085 1869 4137 1882
rect 4149 1916 4201 1921
rect 4149 1882 4158 1916
rect 4158 1882 4192 1916
rect 4192 1882 4201 1916
rect 4149 1869 4201 1882
rect 4213 1916 4265 1921
rect 4213 1882 4230 1916
rect 4230 1882 4264 1916
rect 4264 1882 4265 1916
rect 4213 1869 4265 1882
rect 4085 1842 4137 1855
rect 4085 1808 4086 1842
rect 4086 1808 4120 1842
rect 4120 1808 4137 1842
rect 4085 1803 4137 1808
rect 4149 1842 4201 1855
rect 4149 1808 4158 1842
rect 4158 1808 4192 1842
rect 4192 1808 4201 1842
rect 4149 1803 4201 1808
rect 4213 1842 4265 1855
rect 4213 1808 4230 1842
rect 4230 1808 4264 1842
rect 4264 1808 4265 1842
rect 4213 1803 4265 1808
rect 4085 1768 4137 1789
rect 4085 1737 4086 1768
rect 4086 1737 4120 1768
rect 4120 1737 4137 1768
rect 4149 1768 4201 1789
rect 4149 1737 4158 1768
rect 4158 1737 4192 1768
rect 4192 1737 4201 1768
rect 4213 1768 4265 1789
rect 4213 1737 4230 1768
rect 4230 1737 4264 1768
rect 4264 1737 4265 1768
rect 4085 1694 4137 1723
rect 4085 1671 4086 1694
rect 4086 1671 4120 1694
rect 4120 1671 4137 1694
rect 4149 1694 4201 1723
rect 4149 1671 4158 1694
rect 4158 1671 4192 1694
rect 4192 1671 4201 1694
rect 4213 1694 4265 1723
rect 4213 1671 4230 1694
rect 4230 1671 4264 1694
rect 4264 1671 4265 1694
rect 4085 1620 4137 1657
rect 4085 1605 4086 1620
rect 4086 1605 4120 1620
rect 4120 1605 4137 1620
rect 4149 1620 4201 1657
rect 4149 1605 4158 1620
rect 4158 1605 4192 1620
rect 4192 1605 4201 1620
rect 4213 1620 4265 1657
rect 4213 1605 4230 1620
rect 4230 1605 4264 1620
rect 4264 1605 4265 1620
rect 4085 1586 4086 1591
rect 4086 1586 4120 1591
rect 4120 1586 4137 1591
rect 4085 1545 4137 1586
rect 4085 1539 4086 1545
rect 4086 1539 4120 1545
rect 4120 1539 4137 1545
rect 4149 1586 4158 1591
rect 4158 1586 4192 1591
rect 4192 1586 4201 1591
rect 4149 1545 4201 1586
rect 4149 1539 4158 1545
rect 4158 1539 4192 1545
rect 4192 1539 4201 1545
rect 4213 1586 4230 1591
rect 4230 1586 4264 1591
rect 4264 1586 4265 1591
rect 4213 1545 4265 1586
rect 4213 1539 4230 1545
rect 4230 1539 4264 1545
rect 4264 1539 4265 1545
rect 4085 1511 4086 1525
rect 4086 1511 4120 1525
rect 4120 1511 4137 1525
rect 4085 1473 4137 1511
rect 4149 1511 4158 1525
rect 4158 1511 4192 1525
rect 4192 1511 4201 1525
rect 4149 1473 4201 1511
rect 4213 1511 4230 1525
rect 4230 1511 4264 1525
rect 4264 1511 4265 1525
rect 4213 1473 4265 1511
rect 4581 4050 4633 4068
rect 4645 4062 4697 4068
rect 4645 4050 4654 4062
rect 4654 4050 4688 4062
rect 4688 4050 4697 4062
rect 4709 4050 4761 4068
rect 4581 4016 4582 4050
rect 4582 4016 4633 4050
rect 4645 4016 4697 4050
rect 4709 4016 4760 4050
rect 4760 4016 4761 4050
rect 4581 3951 4582 4003
rect 4582 3951 4633 4003
rect 4645 3951 4697 4003
rect 4709 3951 4760 4003
rect 4760 3951 4761 4003
rect 4581 3886 4582 3938
rect 4582 3886 4633 3938
rect 4645 3886 4697 3938
rect 4709 3886 4760 3938
rect 4760 3886 4761 3938
rect 4581 3821 4582 3873
rect 4582 3821 4633 3873
rect 4645 3821 4697 3873
rect 4709 3821 4760 3873
rect 4760 3821 4761 3873
rect 4581 3756 4582 3808
rect 4582 3756 4633 3808
rect 4645 3756 4697 3808
rect 4709 3756 4760 3808
rect 4760 3756 4761 3808
rect 4581 3691 4582 3743
rect 4582 3691 4633 3743
rect 4645 3691 4697 3743
rect 4709 3691 4760 3743
rect 4760 3691 4761 3743
rect 4581 3626 4582 3678
rect 4582 3626 4633 3678
rect 4645 3626 4697 3678
rect 4709 3626 4760 3678
rect 4760 3626 4761 3678
rect 4581 3561 4582 3613
rect 4582 3561 4633 3613
rect 4645 3561 4697 3613
rect 4709 3561 4760 3613
rect 4760 3561 4761 3613
rect 4581 3496 4582 3548
rect 4582 3496 4633 3548
rect 4645 3496 4697 3548
rect 4709 3496 4760 3548
rect 4760 3496 4761 3548
rect 4581 3431 4582 3483
rect 4582 3431 4633 3483
rect 4645 3431 4697 3483
rect 4709 3431 4760 3483
rect 4760 3431 4761 3483
rect 4581 3366 4582 3418
rect 4582 3366 4633 3418
rect 4645 3366 4697 3418
rect 4709 3366 4760 3418
rect 4760 3366 4761 3418
rect 4581 3301 4582 3353
rect 4582 3301 4633 3353
rect 4645 3301 4697 3353
rect 4709 3301 4760 3353
rect 4760 3301 4761 3353
rect 4581 3236 4582 3288
rect 4582 3236 4633 3288
rect 4645 3236 4697 3288
rect 4709 3236 4760 3288
rect 4760 3236 4761 3288
rect 4581 3171 4582 3223
rect 4582 3171 4633 3223
rect 4645 3171 4697 3223
rect 4709 3171 4760 3223
rect 4760 3171 4761 3223
rect 4581 3106 4582 3158
rect 4582 3106 4633 3158
rect 4645 3106 4697 3158
rect 4709 3106 4760 3158
rect 4760 3106 4761 3158
rect 4581 3080 4582 3093
rect 4582 3092 4633 3093
rect 4645 3092 4697 3093
rect 4709 3092 4760 3093
rect 4582 3080 4616 3092
rect 4616 3080 4633 3092
rect 4581 3041 4633 3080
rect 4645 3041 4697 3092
rect 4709 3080 4726 3092
rect 4726 3080 4760 3092
rect 4760 3080 4761 3093
rect 4709 3041 4761 3080
rect 4581 2976 4582 3028
rect 4582 2976 4633 3028
rect 4645 2976 4697 3028
rect 4709 2976 4760 3028
rect 4760 2976 4761 3028
rect 4581 2911 4582 2963
rect 4582 2911 4633 2963
rect 4645 2911 4697 2963
rect 4709 2911 4760 2963
rect 4760 2911 4761 2963
rect 4581 2846 4582 2898
rect 4582 2846 4633 2898
rect 4645 2846 4697 2898
rect 4709 2846 4760 2898
rect 4760 2846 4761 2898
rect 4581 2781 4582 2833
rect 4582 2781 4633 2833
rect 4645 2781 4697 2833
rect 4709 2781 4760 2833
rect 4760 2781 4761 2833
rect 4581 2716 4582 2768
rect 4582 2716 4633 2768
rect 4645 2716 4697 2768
rect 4709 2716 4760 2768
rect 4760 2716 4761 2768
rect 4581 2651 4582 2703
rect 4582 2651 4633 2703
rect 4645 2651 4697 2703
rect 4709 2651 4760 2703
rect 4760 2651 4761 2703
rect 4581 2586 4582 2638
rect 4582 2586 4633 2638
rect 4645 2586 4697 2638
rect 4709 2586 4760 2638
rect 4760 2586 4761 2638
rect 4581 2535 4633 2573
rect 4581 2521 4582 2535
rect 4582 2521 4616 2535
rect 4616 2521 4633 2535
rect 4645 2535 4697 2573
rect 4645 2521 4654 2535
rect 4654 2521 4688 2535
rect 4688 2521 4697 2535
rect 4709 2535 4761 2573
rect 4709 2521 4726 2535
rect 4726 2521 4760 2535
rect 4760 2521 4761 2535
rect 4581 2501 4582 2508
rect 4582 2501 4616 2508
rect 4616 2501 4633 2508
rect 4581 2456 4633 2501
rect 4645 2501 4654 2508
rect 4654 2501 4688 2508
rect 4688 2501 4697 2508
rect 4645 2461 4697 2501
rect 4645 2456 4654 2461
rect 4654 2456 4688 2461
rect 4688 2456 4697 2461
rect 4709 2501 4726 2508
rect 4726 2501 4760 2508
rect 4760 2501 4761 2508
rect 4709 2456 4761 2501
rect 4581 2391 4582 2443
rect 4582 2391 4633 2443
rect 4645 2391 4697 2443
rect 4709 2391 4760 2443
rect 4760 2391 4761 2443
rect 4581 2326 4582 2378
rect 4582 2326 4633 2378
rect 4645 2326 4697 2378
rect 4709 2326 4760 2378
rect 4760 2326 4761 2378
rect 4581 2261 4582 2313
rect 4582 2261 4633 2313
rect 4645 2261 4697 2313
rect 4709 2261 4760 2313
rect 4760 2261 4761 2313
rect 4581 2196 4582 2248
rect 4582 2196 4633 2248
rect 4645 2196 4697 2248
rect 4709 2196 4760 2248
rect 4760 2196 4761 2248
rect 4581 2131 4582 2183
rect 4582 2131 4633 2183
rect 4645 2131 4697 2183
rect 4709 2131 4760 2183
rect 4760 2131 4761 2183
rect 4581 2066 4582 2118
rect 4582 2066 4633 2118
rect 4645 2066 4697 2118
rect 4709 2066 4760 2118
rect 4760 2066 4761 2118
rect 4581 2001 4582 2053
rect 4582 2001 4633 2053
rect 4645 2001 4697 2053
rect 4709 2001 4760 2053
rect 4760 2001 4761 2053
rect 4581 1935 4582 1987
rect 4582 1935 4633 1987
rect 4645 1935 4697 1987
rect 4709 1935 4760 1987
rect 4760 1935 4761 1987
rect 4581 1869 4582 1921
rect 4582 1869 4633 1921
rect 4645 1869 4697 1921
rect 4709 1869 4760 1921
rect 4760 1869 4761 1921
rect 4581 1803 4582 1855
rect 4582 1803 4633 1855
rect 4645 1803 4697 1855
rect 4709 1803 4760 1855
rect 4760 1803 4761 1855
rect 4581 1737 4582 1789
rect 4582 1737 4633 1789
rect 4645 1737 4697 1789
rect 4709 1737 4760 1789
rect 4760 1737 4761 1789
rect 4581 1671 4582 1723
rect 4582 1671 4633 1723
rect 4645 1671 4697 1723
rect 4709 1671 4760 1723
rect 4760 1671 4761 1723
rect 4581 1605 4582 1657
rect 4582 1605 4633 1657
rect 4645 1605 4697 1657
rect 4709 1605 4760 1657
rect 4760 1605 4761 1657
rect 4581 1539 4582 1591
rect 4582 1539 4633 1591
rect 4645 1539 4697 1591
rect 4709 1539 4760 1591
rect 4760 1539 4761 1591
rect 4581 1479 4582 1525
rect 4582 1491 4633 1525
rect 4645 1491 4697 1525
rect 4709 1491 4760 1525
rect 4582 1479 4616 1491
rect 4616 1479 4633 1491
rect 4581 1473 4633 1479
rect 4645 1473 4697 1491
rect 4709 1479 4726 1491
rect 4726 1479 4760 1491
rect 4760 1479 4761 1525
rect 4709 1473 4761 1479
rect 5077 4062 5129 4068
rect 5077 4028 5078 4062
rect 5078 4028 5112 4062
rect 5112 4028 5129 4062
rect 5077 4016 5129 4028
rect 5141 4062 5193 4068
rect 5141 4028 5150 4062
rect 5150 4028 5184 4062
rect 5184 4028 5193 4062
rect 5141 4016 5193 4028
rect 5205 4062 5257 4068
rect 5205 4028 5222 4062
rect 5222 4028 5256 4062
rect 5256 4028 5257 4062
rect 5205 4016 5257 4028
rect 5077 3988 5129 4003
rect 5077 3954 5078 3988
rect 5078 3954 5112 3988
rect 5112 3954 5129 3988
rect 5077 3951 5129 3954
rect 5141 3988 5193 4003
rect 5141 3954 5150 3988
rect 5150 3954 5184 3988
rect 5184 3954 5193 3988
rect 5141 3951 5193 3954
rect 5205 3988 5257 4003
rect 5205 3954 5222 3988
rect 5222 3954 5256 3988
rect 5256 3954 5257 3988
rect 5205 3951 5257 3954
rect 5077 3914 5129 3938
rect 5077 3886 5078 3914
rect 5078 3886 5112 3914
rect 5112 3886 5129 3914
rect 5141 3914 5193 3938
rect 5141 3886 5150 3914
rect 5150 3886 5184 3914
rect 5184 3886 5193 3914
rect 5205 3914 5257 3938
rect 5205 3886 5222 3914
rect 5222 3886 5256 3914
rect 5256 3886 5257 3914
rect 5077 3840 5129 3873
rect 5077 3821 5078 3840
rect 5078 3821 5112 3840
rect 5112 3821 5129 3840
rect 5141 3840 5193 3873
rect 5141 3821 5150 3840
rect 5150 3821 5184 3840
rect 5184 3821 5193 3840
rect 5205 3840 5257 3873
rect 5205 3821 5222 3840
rect 5222 3821 5256 3840
rect 5256 3821 5257 3840
rect 5077 3806 5078 3808
rect 5078 3806 5112 3808
rect 5112 3806 5129 3808
rect 5077 3766 5129 3806
rect 5077 3756 5078 3766
rect 5078 3756 5112 3766
rect 5112 3756 5129 3766
rect 5141 3806 5150 3808
rect 5150 3806 5184 3808
rect 5184 3806 5193 3808
rect 5141 3766 5193 3806
rect 5141 3756 5150 3766
rect 5150 3756 5184 3766
rect 5184 3756 5193 3766
rect 5205 3806 5222 3808
rect 5222 3806 5256 3808
rect 5256 3806 5257 3808
rect 5205 3766 5257 3806
rect 5205 3756 5222 3766
rect 5222 3756 5256 3766
rect 5256 3756 5257 3766
rect 5077 3732 5078 3743
rect 5078 3732 5112 3743
rect 5112 3732 5129 3743
rect 5077 3692 5129 3732
rect 5077 3691 5078 3692
rect 5078 3691 5112 3692
rect 5112 3691 5129 3692
rect 5141 3732 5150 3743
rect 5150 3732 5184 3743
rect 5184 3732 5193 3743
rect 5141 3692 5193 3732
rect 5141 3691 5150 3692
rect 5150 3691 5184 3692
rect 5184 3691 5193 3692
rect 5205 3732 5222 3743
rect 5222 3732 5256 3743
rect 5256 3732 5257 3743
rect 5205 3692 5257 3732
rect 5205 3691 5222 3692
rect 5222 3691 5256 3692
rect 5256 3691 5257 3692
rect 5077 3658 5078 3678
rect 5078 3658 5112 3678
rect 5112 3658 5129 3678
rect 5077 3626 5129 3658
rect 5141 3658 5150 3678
rect 5150 3658 5184 3678
rect 5184 3658 5193 3678
rect 5141 3626 5193 3658
rect 5205 3658 5222 3678
rect 5222 3658 5256 3678
rect 5256 3658 5257 3678
rect 5205 3626 5257 3658
rect 5077 3584 5078 3613
rect 5078 3584 5112 3613
rect 5112 3584 5129 3613
rect 5077 3561 5129 3584
rect 5141 3584 5150 3613
rect 5150 3584 5184 3613
rect 5184 3584 5193 3613
rect 5141 3561 5193 3584
rect 5205 3584 5222 3613
rect 5222 3584 5256 3613
rect 5256 3584 5257 3613
rect 5205 3561 5257 3584
rect 5077 3544 5129 3548
rect 5077 3510 5078 3544
rect 5078 3510 5112 3544
rect 5112 3510 5129 3544
rect 5077 3496 5129 3510
rect 5141 3544 5193 3548
rect 5141 3510 5150 3544
rect 5150 3510 5184 3544
rect 5184 3510 5193 3544
rect 5141 3496 5193 3510
rect 5205 3544 5257 3548
rect 5205 3510 5222 3544
rect 5222 3510 5256 3544
rect 5256 3510 5257 3544
rect 5205 3496 5257 3510
rect 5077 3470 5129 3483
rect 5077 3436 5078 3470
rect 5078 3436 5112 3470
rect 5112 3436 5129 3470
rect 5077 3431 5129 3436
rect 5141 3470 5193 3483
rect 5141 3436 5150 3470
rect 5150 3436 5184 3470
rect 5184 3436 5193 3470
rect 5141 3431 5193 3436
rect 5205 3470 5257 3483
rect 5205 3436 5222 3470
rect 5222 3436 5256 3470
rect 5256 3436 5257 3470
rect 5205 3431 5257 3436
rect 5077 3396 5129 3418
rect 5077 3366 5078 3396
rect 5078 3366 5112 3396
rect 5112 3366 5129 3396
rect 5141 3396 5193 3418
rect 5141 3366 5150 3396
rect 5150 3366 5184 3396
rect 5184 3366 5193 3396
rect 5205 3396 5257 3418
rect 5205 3366 5222 3396
rect 5222 3366 5256 3396
rect 5256 3366 5257 3396
rect 5077 3322 5129 3353
rect 5077 3301 5078 3322
rect 5078 3301 5112 3322
rect 5112 3301 5129 3322
rect 5141 3322 5193 3353
rect 5141 3301 5150 3322
rect 5150 3301 5184 3322
rect 5184 3301 5193 3322
rect 5205 3322 5257 3353
rect 5205 3301 5222 3322
rect 5222 3301 5256 3322
rect 5256 3301 5257 3322
rect 5077 3248 5129 3288
rect 5077 3236 5078 3248
rect 5078 3236 5112 3248
rect 5112 3236 5129 3248
rect 5141 3248 5193 3288
rect 5141 3236 5150 3248
rect 5150 3236 5184 3248
rect 5184 3236 5193 3248
rect 5205 3248 5257 3288
rect 5205 3236 5222 3248
rect 5222 3236 5256 3248
rect 5256 3236 5257 3248
rect 5077 3214 5078 3223
rect 5078 3214 5112 3223
rect 5112 3214 5129 3223
rect 5077 3174 5129 3214
rect 5077 3171 5078 3174
rect 5078 3171 5112 3174
rect 5112 3171 5129 3174
rect 5141 3214 5150 3223
rect 5150 3214 5184 3223
rect 5184 3214 5193 3223
rect 5141 3174 5193 3214
rect 5141 3171 5150 3174
rect 5150 3171 5184 3174
rect 5184 3171 5193 3174
rect 5205 3214 5222 3223
rect 5222 3214 5256 3223
rect 5256 3214 5257 3223
rect 5205 3174 5257 3214
rect 5205 3171 5222 3174
rect 5222 3171 5256 3174
rect 5256 3171 5257 3174
rect 5077 3140 5078 3158
rect 5078 3140 5112 3158
rect 5112 3140 5129 3158
rect 5077 3106 5129 3140
rect 5141 3140 5150 3158
rect 5150 3140 5184 3158
rect 5184 3140 5193 3158
rect 5141 3106 5193 3140
rect 5205 3140 5222 3158
rect 5222 3140 5256 3158
rect 5256 3140 5257 3158
rect 5205 3106 5257 3140
rect 5077 3066 5078 3093
rect 5078 3066 5112 3093
rect 5112 3066 5129 3093
rect 5077 3041 5129 3066
rect 5141 3066 5150 3093
rect 5150 3066 5184 3093
rect 5184 3066 5193 3093
rect 5141 3041 5193 3066
rect 5205 3066 5222 3093
rect 5222 3066 5256 3093
rect 5256 3066 5257 3093
rect 5205 3041 5257 3066
rect 5077 3026 5129 3028
rect 5077 2992 5078 3026
rect 5078 2992 5112 3026
rect 5112 2992 5129 3026
rect 5077 2976 5129 2992
rect 5141 3026 5193 3028
rect 5141 2992 5150 3026
rect 5150 2992 5184 3026
rect 5184 2992 5193 3026
rect 5141 2976 5193 2992
rect 5205 3026 5257 3028
rect 5205 2992 5222 3026
rect 5222 2992 5256 3026
rect 5256 2992 5257 3026
rect 5205 2976 5257 2992
rect 5077 2952 5129 2963
rect 5077 2918 5078 2952
rect 5078 2918 5112 2952
rect 5112 2918 5129 2952
rect 5077 2911 5129 2918
rect 5141 2952 5193 2963
rect 5141 2918 5150 2952
rect 5150 2918 5184 2952
rect 5184 2918 5193 2952
rect 5141 2911 5193 2918
rect 5205 2952 5257 2963
rect 5205 2918 5222 2952
rect 5222 2918 5256 2952
rect 5256 2918 5257 2952
rect 5205 2911 5257 2918
rect 5077 2878 5129 2898
rect 5077 2846 5078 2878
rect 5078 2846 5112 2878
rect 5112 2846 5129 2878
rect 5141 2878 5193 2898
rect 5141 2846 5150 2878
rect 5150 2846 5184 2878
rect 5184 2846 5193 2878
rect 5205 2878 5257 2898
rect 5205 2846 5222 2878
rect 5222 2846 5256 2878
rect 5256 2846 5257 2878
rect 5077 2804 5129 2833
rect 5077 2781 5078 2804
rect 5078 2781 5112 2804
rect 5112 2781 5129 2804
rect 5141 2804 5193 2833
rect 5141 2781 5150 2804
rect 5150 2781 5184 2804
rect 5184 2781 5193 2804
rect 5205 2804 5257 2833
rect 5205 2781 5222 2804
rect 5222 2781 5256 2804
rect 5256 2781 5257 2804
rect 5077 2730 5129 2768
rect 5077 2716 5078 2730
rect 5078 2716 5112 2730
rect 5112 2716 5129 2730
rect 5141 2730 5193 2768
rect 5141 2716 5150 2730
rect 5150 2716 5184 2730
rect 5184 2716 5193 2730
rect 5205 2730 5257 2768
rect 5205 2716 5222 2730
rect 5222 2716 5256 2730
rect 5256 2716 5257 2730
rect 5077 2696 5078 2703
rect 5078 2696 5112 2703
rect 5112 2696 5129 2703
rect 5077 2656 5129 2696
rect 5077 2651 5078 2656
rect 5078 2651 5112 2656
rect 5112 2651 5129 2656
rect 5141 2696 5150 2703
rect 5150 2696 5184 2703
rect 5184 2696 5193 2703
rect 5141 2656 5193 2696
rect 5141 2651 5150 2656
rect 5150 2651 5184 2656
rect 5184 2651 5193 2656
rect 5205 2696 5222 2703
rect 5222 2696 5256 2703
rect 5256 2696 5257 2703
rect 5205 2656 5257 2696
rect 5205 2651 5222 2656
rect 5222 2651 5256 2656
rect 5256 2651 5257 2656
rect 5077 2622 5078 2638
rect 5078 2622 5112 2638
rect 5112 2622 5129 2638
rect 5077 2586 5129 2622
rect 5141 2622 5150 2638
rect 5150 2622 5184 2638
rect 5184 2622 5193 2638
rect 5141 2586 5193 2622
rect 5205 2622 5222 2638
rect 5222 2622 5256 2638
rect 5256 2622 5257 2638
rect 5205 2586 5257 2622
rect 5077 2548 5078 2573
rect 5078 2548 5112 2573
rect 5112 2548 5129 2573
rect 5077 2521 5129 2548
rect 5141 2548 5150 2573
rect 5150 2548 5184 2573
rect 5184 2548 5193 2573
rect 5141 2521 5193 2548
rect 5205 2548 5222 2573
rect 5222 2548 5256 2573
rect 5256 2548 5257 2573
rect 5205 2521 5257 2548
rect 5077 2474 5078 2508
rect 5078 2474 5112 2508
rect 5112 2474 5129 2508
rect 5077 2456 5129 2474
rect 5141 2474 5150 2508
rect 5150 2474 5184 2508
rect 5184 2474 5193 2508
rect 5141 2456 5193 2474
rect 5205 2474 5222 2508
rect 5222 2474 5256 2508
rect 5256 2474 5257 2508
rect 5205 2456 5257 2474
rect 5077 2434 5129 2443
rect 5077 2400 5078 2434
rect 5078 2400 5112 2434
rect 5112 2400 5129 2434
rect 5077 2391 5129 2400
rect 5141 2434 5193 2443
rect 5141 2400 5150 2434
rect 5150 2400 5184 2434
rect 5184 2400 5193 2434
rect 5141 2391 5193 2400
rect 5205 2434 5257 2443
rect 5205 2400 5222 2434
rect 5222 2400 5256 2434
rect 5256 2400 5257 2434
rect 5205 2391 5257 2400
rect 5077 2360 5129 2378
rect 5077 2326 5078 2360
rect 5078 2326 5112 2360
rect 5112 2326 5129 2360
rect 5141 2360 5193 2378
rect 5141 2326 5150 2360
rect 5150 2326 5184 2360
rect 5184 2326 5193 2360
rect 5205 2360 5257 2378
rect 5205 2326 5222 2360
rect 5222 2326 5256 2360
rect 5256 2326 5257 2360
rect 5077 2286 5129 2313
rect 5077 2261 5078 2286
rect 5078 2261 5112 2286
rect 5112 2261 5129 2286
rect 5141 2286 5193 2313
rect 5141 2261 5150 2286
rect 5150 2261 5184 2286
rect 5184 2261 5193 2286
rect 5205 2286 5257 2313
rect 5205 2261 5222 2286
rect 5222 2261 5256 2286
rect 5256 2261 5257 2286
rect 5077 2212 5129 2248
rect 5077 2196 5078 2212
rect 5078 2196 5112 2212
rect 5112 2196 5129 2212
rect 5141 2212 5193 2248
rect 5141 2196 5150 2212
rect 5150 2196 5184 2212
rect 5184 2196 5193 2212
rect 5205 2212 5257 2248
rect 5205 2196 5222 2212
rect 5222 2196 5256 2212
rect 5256 2196 5257 2212
rect 5077 2178 5078 2183
rect 5078 2178 5112 2183
rect 5112 2178 5129 2183
rect 5077 2138 5129 2178
rect 5077 2131 5078 2138
rect 5078 2131 5112 2138
rect 5112 2131 5129 2138
rect 5141 2178 5150 2183
rect 5150 2178 5184 2183
rect 5184 2178 5193 2183
rect 5141 2138 5193 2178
rect 5141 2131 5150 2138
rect 5150 2131 5184 2138
rect 5184 2131 5193 2138
rect 5205 2178 5222 2183
rect 5222 2178 5256 2183
rect 5256 2178 5257 2183
rect 5205 2138 5257 2178
rect 5205 2131 5222 2138
rect 5222 2131 5256 2138
rect 5256 2131 5257 2138
rect 5077 2104 5078 2118
rect 5078 2104 5112 2118
rect 5112 2104 5129 2118
rect 5077 2066 5129 2104
rect 5141 2104 5150 2118
rect 5150 2104 5184 2118
rect 5184 2104 5193 2118
rect 5141 2066 5193 2104
rect 5205 2104 5222 2118
rect 5222 2104 5256 2118
rect 5256 2104 5257 2118
rect 5205 2066 5257 2104
rect 5077 2030 5078 2053
rect 5078 2030 5112 2053
rect 5112 2030 5129 2053
rect 5077 2001 5129 2030
rect 5141 2030 5150 2053
rect 5150 2030 5184 2053
rect 5184 2030 5193 2053
rect 5141 2001 5193 2030
rect 5205 2030 5222 2053
rect 5222 2030 5256 2053
rect 5256 2030 5257 2053
rect 5205 2001 5257 2030
rect 5077 1956 5078 1987
rect 5078 1956 5112 1987
rect 5112 1956 5129 1987
rect 5077 1935 5129 1956
rect 5141 1956 5150 1987
rect 5150 1956 5184 1987
rect 5184 1956 5193 1987
rect 5141 1935 5193 1956
rect 5205 1956 5222 1987
rect 5222 1956 5256 1987
rect 5256 1956 5257 1987
rect 5205 1935 5257 1956
rect 5077 1916 5129 1921
rect 5077 1882 5078 1916
rect 5078 1882 5112 1916
rect 5112 1882 5129 1916
rect 5077 1869 5129 1882
rect 5141 1916 5193 1921
rect 5141 1882 5150 1916
rect 5150 1882 5184 1916
rect 5184 1882 5193 1916
rect 5141 1869 5193 1882
rect 5205 1916 5257 1921
rect 5205 1882 5222 1916
rect 5222 1882 5256 1916
rect 5256 1882 5257 1916
rect 5205 1869 5257 1882
rect 5077 1842 5129 1855
rect 5077 1808 5078 1842
rect 5078 1808 5112 1842
rect 5112 1808 5129 1842
rect 5077 1803 5129 1808
rect 5141 1842 5193 1855
rect 5141 1808 5150 1842
rect 5150 1808 5184 1842
rect 5184 1808 5193 1842
rect 5141 1803 5193 1808
rect 5205 1842 5257 1855
rect 5205 1808 5222 1842
rect 5222 1808 5256 1842
rect 5256 1808 5257 1842
rect 5205 1803 5257 1808
rect 5077 1768 5129 1789
rect 5077 1737 5078 1768
rect 5078 1737 5112 1768
rect 5112 1737 5129 1768
rect 5141 1768 5193 1789
rect 5141 1737 5150 1768
rect 5150 1737 5184 1768
rect 5184 1737 5193 1768
rect 5205 1768 5257 1789
rect 5205 1737 5222 1768
rect 5222 1737 5256 1768
rect 5256 1737 5257 1768
rect 5077 1694 5129 1723
rect 5077 1671 5078 1694
rect 5078 1671 5112 1694
rect 5112 1671 5129 1694
rect 5141 1694 5193 1723
rect 5141 1671 5150 1694
rect 5150 1671 5184 1694
rect 5184 1671 5193 1694
rect 5205 1694 5257 1723
rect 5205 1671 5222 1694
rect 5222 1671 5256 1694
rect 5256 1671 5257 1694
rect 5077 1620 5129 1657
rect 5077 1605 5078 1620
rect 5078 1605 5112 1620
rect 5112 1605 5129 1620
rect 5141 1620 5193 1657
rect 5141 1605 5150 1620
rect 5150 1605 5184 1620
rect 5184 1605 5193 1620
rect 5205 1620 5257 1657
rect 5205 1605 5222 1620
rect 5222 1605 5256 1620
rect 5256 1605 5257 1620
rect 5077 1586 5078 1591
rect 5078 1586 5112 1591
rect 5112 1586 5129 1591
rect 5077 1545 5129 1586
rect 5077 1539 5078 1545
rect 5078 1539 5112 1545
rect 5112 1539 5129 1545
rect 5141 1586 5150 1591
rect 5150 1586 5184 1591
rect 5184 1586 5193 1591
rect 5141 1545 5193 1586
rect 5141 1539 5150 1545
rect 5150 1539 5184 1545
rect 5184 1539 5193 1545
rect 5205 1586 5222 1591
rect 5222 1586 5256 1591
rect 5256 1586 5257 1591
rect 5205 1545 5257 1586
rect 5205 1539 5222 1545
rect 5222 1539 5256 1545
rect 5256 1539 5257 1545
rect 5077 1511 5078 1525
rect 5078 1511 5112 1525
rect 5112 1511 5129 1525
rect 5077 1473 5129 1511
rect 5141 1511 5150 1525
rect 5150 1511 5184 1525
rect 5184 1511 5193 1525
rect 5141 1473 5193 1511
rect 5205 1511 5222 1525
rect 5222 1511 5256 1525
rect 5256 1511 5257 1525
rect 5205 1473 5257 1511
rect 5573 4050 5625 4068
rect 5637 4062 5689 4068
rect 5637 4050 5646 4062
rect 5646 4050 5680 4062
rect 5680 4050 5689 4062
rect 5701 4050 5753 4068
rect 5573 4016 5574 4050
rect 5574 4016 5625 4050
rect 5637 4016 5689 4050
rect 5701 4016 5752 4050
rect 5752 4016 5753 4050
rect 5573 3951 5574 4003
rect 5574 3951 5625 4003
rect 5637 3951 5689 4003
rect 5701 3951 5752 4003
rect 5752 3951 5753 4003
rect 5573 3886 5574 3938
rect 5574 3886 5625 3938
rect 5637 3886 5689 3938
rect 5701 3886 5752 3938
rect 5752 3886 5753 3938
rect 5573 3821 5574 3873
rect 5574 3821 5625 3873
rect 5637 3821 5689 3873
rect 5701 3821 5752 3873
rect 5752 3821 5753 3873
rect 5573 3756 5574 3808
rect 5574 3756 5625 3808
rect 5637 3756 5689 3808
rect 5701 3756 5752 3808
rect 5752 3756 5753 3808
rect 5573 3691 5574 3743
rect 5574 3691 5625 3743
rect 5637 3691 5689 3743
rect 5701 3691 5752 3743
rect 5752 3691 5753 3743
rect 5573 3626 5574 3678
rect 5574 3626 5625 3678
rect 5637 3626 5689 3678
rect 5701 3626 5752 3678
rect 5752 3626 5753 3678
rect 5573 3561 5574 3613
rect 5574 3561 5625 3613
rect 5637 3561 5689 3613
rect 5701 3561 5752 3613
rect 5752 3561 5753 3613
rect 5573 3496 5574 3548
rect 5574 3496 5625 3548
rect 5637 3496 5689 3548
rect 5701 3496 5752 3548
rect 5752 3496 5753 3548
rect 5573 3431 5574 3483
rect 5574 3431 5625 3483
rect 5637 3431 5689 3483
rect 5701 3431 5752 3483
rect 5752 3431 5753 3483
rect 5573 3366 5574 3418
rect 5574 3366 5625 3418
rect 5637 3366 5689 3418
rect 5701 3366 5752 3418
rect 5752 3366 5753 3418
rect 5573 3301 5574 3353
rect 5574 3301 5625 3353
rect 5637 3301 5689 3353
rect 5701 3301 5752 3353
rect 5752 3301 5753 3353
rect 5573 3236 5574 3288
rect 5574 3236 5625 3288
rect 5637 3236 5689 3288
rect 5701 3236 5752 3288
rect 5752 3236 5753 3288
rect 5573 3171 5574 3223
rect 5574 3171 5625 3223
rect 5637 3171 5689 3223
rect 5701 3171 5752 3223
rect 5752 3171 5753 3223
rect 5573 3106 5574 3158
rect 5574 3106 5625 3158
rect 5637 3106 5689 3158
rect 5701 3106 5752 3158
rect 5752 3106 5753 3158
rect 5573 3080 5574 3093
rect 5574 3092 5625 3093
rect 5637 3092 5689 3093
rect 5701 3092 5752 3093
rect 5574 3080 5608 3092
rect 5608 3080 5625 3092
rect 5573 3041 5625 3080
rect 5637 3041 5689 3092
rect 5701 3080 5718 3092
rect 5718 3080 5752 3092
rect 5752 3080 5753 3093
rect 5701 3041 5753 3080
rect 5573 2976 5574 3028
rect 5574 2976 5625 3028
rect 5637 2976 5689 3028
rect 5701 2976 5752 3028
rect 5752 2976 5753 3028
rect 5573 2911 5574 2963
rect 5574 2911 5625 2963
rect 5637 2911 5689 2963
rect 5701 2911 5752 2963
rect 5752 2911 5753 2963
rect 5573 2846 5574 2898
rect 5574 2846 5625 2898
rect 5637 2846 5689 2898
rect 5701 2846 5752 2898
rect 5752 2846 5753 2898
rect 5573 2781 5574 2833
rect 5574 2781 5625 2833
rect 5637 2781 5689 2833
rect 5701 2781 5752 2833
rect 5752 2781 5753 2833
rect 5573 2716 5574 2768
rect 5574 2716 5625 2768
rect 5637 2716 5689 2768
rect 5701 2716 5752 2768
rect 5752 2716 5753 2768
rect 5573 2651 5574 2703
rect 5574 2651 5625 2703
rect 5637 2651 5689 2703
rect 5701 2651 5752 2703
rect 5752 2651 5753 2703
rect 5573 2586 5574 2638
rect 5574 2586 5625 2638
rect 5637 2586 5689 2638
rect 5701 2586 5752 2638
rect 5752 2586 5753 2638
rect 5573 2535 5625 2573
rect 5573 2521 5574 2535
rect 5574 2521 5608 2535
rect 5608 2521 5625 2535
rect 5637 2535 5689 2573
rect 5637 2521 5646 2535
rect 5646 2521 5680 2535
rect 5680 2521 5689 2535
rect 5701 2535 5753 2573
rect 5701 2521 5718 2535
rect 5718 2521 5752 2535
rect 5752 2521 5753 2535
rect 5573 2501 5574 2508
rect 5574 2501 5608 2508
rect 5608 2501 5625 2508
rect 5573 2456 5625 2501
rect 5637 2501 5646 2508
rect 5646 2501 5680 2508
rect 5680 2501 5689 2508
rect 5637 2461 5689 2501
rect 5637 2456 5646 2461
rect 5646 2456 5680 2461
rect 5680 2456 5689 2461
rect 5701 2501 5718 2508
rect 5718 2501 5752 2508
rect 5752 2501 5753 2508
rect 5701 2456 5753 2501
rect 5573 2391 5574 2443
rect 5574 2391 5625 2443
rect 5637 2391 5689 2443
rect 5701 2391 5752 2443
rect 5752 2391 5753 2443
rect 5573 2326 5574 2378
rect 5574 2326 5625 2378
rect 5637 2326 5689 2378
rect 5701 2326 5752 2378
rect 5752 2326 5753 2378
rect 5573 2261 5574 2313
rect 5574 2261 5625 2313
rect 5637 2261 5689 2313
rect 5701 2261 5752 2313
rect 5752 2261 5753 2313
rect 5573 2196 5574 2248
rect 5574 2196 5625 2248
rect 5637 2196 5689 2248
rect 5701 2196 5752 2248
rect 5752 2196 5753 2248
rect 5573 2131 5574 2183
rect 5574 2131 5625 2183
rect 5637 2131 5689 2183
rect 5701 2131 5752 2183
rect 5752 2131 5753 2183
rect 5573 2066 5574 2118
rect 5574 2066 5625 2118
rect 5637 2066 5689 2118
rect 5701 2066 5752 2118
rect 5752 2066 5753 2118
rect 5573 2001 5574 2053
rect 5574 2001 5625 2053
rect 5637 2001 5689 2053
rect 5701 2001 5752 2053
rect 5752 2001 5753 2053
rect 5573 1935 5574 1987
rect 5574 1935 5625 1987
rect 5637 1935 5689 1987
rect 5701 1935 5752 1987
rect 5752 1935 5753 1987
rect 5573 1869 5574 1921
rect 5574 1869 5625 1921
rect 5637 1869 5689 1921
rect 5701 1869 5752 1921
rect 5752 1869 5753 1921
rect 5573 1803 5574 1855
rect 5574 1803 5625 1855
rect 5637 1803 5689 1855
rect 5701 1803 5752 1855
rect 5752 1803 5753 1855
rect 5573 1737 5574 1789
rect 5574 1737 5625 1789
rect 5637 1737 5689 1789
rect 5701 1737 5752 1789
rect 5752 1737 5753 1789
rect 5573 1671 5574 1723
rect 5574 1671 5625 1723
rect 5637 1671 5689 1723
rect 5701 1671 5752 1723
rect 5752 1671 5753 1723
rect 5573 1605 5574 1657
rect 5574 1605 5625 1657
rect 5637 1605 5689 1657
rect 5701 1605 5752 1657
rect 5752 1605 5753 1657
rect 5573 1539 5574 1591
rect 5574 1539 5625 1591
rect 5637 1539 5689 1591
rect 5701 1539 5752 1591
rect 5752 1539 5753 1591
rect 5573 1479 5574 1525
rect 5574 1491 5625 1525
rect 5637 1491 5689 1525
rect 5701 1491 5752 1525
rect 5574 1479 5608 1491
rect 5608 1479 5625 1491
rect 5573 1473 5625 1479
rect 5637 1473 5689 1491
rect 5701 1479 5718 1491
rect 5718 1479 5752 1491
rect 5752 1479 5753 1525
rect 5701 1473 5753 1479
rect 6069 4062 6121 4068
rect 6069 4028 6070 4062
rect 6070 4028 6104 4062
rect 6104 4028 6121 4062
rect 6069 4016 6121 4028
rect 6133 4062 6185 4068
rect 6133 4028 6142 4062
rect 6142 4028 6176 4062
rect 6176 4028 6185 4062
rect 6133 4016 6185 4028
rect 6197 4062 6249 4068
rect 6197 4028 6214 4062
rect 6214 4028 6248 4062
rect 6248 4028 6249 4062
rect 6197 4016 6249 4028
rect 6069 3988 6121 4003
rect 6069 3954 6070 3988
rect 6070 3954 6104 3988
rect 6104 3954 6121 3988
rect 6069 3951 6121 3954
rect 6133 3988 6185 4003
rect 6133 3954 6142 3988
rect 6142 3954 6176 3988
rect 6176 3954 6185 3988
rect 6133 3951 6185 3954
rect 6197 3988 6249 4003
rect 6197 3954 6214 3988
rect 6214 3954 6248 3988
rect 6248 3954 6249 3988
rect 6197 3951 6249 3954
rect 6069 3914 6121 3938
rect 6069 3886 6070 3914
rect 6070 3886 6104 3914
rect 6104 3886 6121 3914
rect 6133 3914 6185 3938
rect 6133 3886 6142 3914
rect 6142 3886 6176 3914
rect 6176 3886 6185 3914
rect 6197 3914 6249 3938
rect 6197 3886 6214 3914
rect 6214 3886 6248 3914
rect 6248 3886 6249 3914
rect 6069 3840 6121 3873
rect 6069 3821 6070 3840
rect 6070 3821 6104 3840
rect 6104 3821 6121 3840
rect 6133 3840 6185 3873
rect 6133 3821 6142 3840
rect 6142 3821 6176 3840
rect 6176 3821 6185 3840
rect 6197 3840 6249 3873
rect 6197 3821 6214 3840
rect 6214 3821 6248 3840
rect 6248 3821 6249 3840
rect 6069 3806 6070 3808
rect 6070 3806 6104 3808
rect 6104 3806 6121 3808
rect 6069 3766 6121 3806
rect 6069 3756 6070 3766
rect 6070 3756 6104 3766
rect 6104 3756 6121 3766
rect 6133 3806 6142 3808
rect 6142 3806 6176 3808
rect 6176 3806 6185 3808
rect 6133 3766 6185 3806
rect 6133 3756 6142 3766
rect 6142 3756 6176 3766
rect 6176 3756 6185 3766
rect 6197 3806 6214 3808
rect 6214 3806 6248 3808
rect 6248 3806 6249 3808
rect 6197 3766 6249 3806
rect 6197 3756 6214 3766
rect 6214 3756 6248 3766
rect 6248 3756 6249 3766
rect 6069 3732 6070 3743
rect 6070 3732 6104 3743
rect 6104 3732 6121 3743
rect 6069 3692 6121 3732
rect 6069 3691 6070 3692
rect 6070 3691 6104 3692
rect 6104 3691 6121 3692
rect 6133 3732 6142 3743
rect 6142 3732 6176 3743
rect 6176 3732 6185 3743
rect 6133 3692 6185 3732
rect 6133 3691 6142 3692
rect 6142 3691 6176 3692
rect 6176 3691 6185 3692
rect 6197 3732 6214 3743
rect 6214 3732 6248 3743
rect 6248 3732 6249 3743
rect 6197 3692 6249 3732
rect 6197 3691 6214 3692
rect 6214 3691 6248 3692
rect 6248 3691 6249 3692
rect 6069 3658 6070 3678
rect 6070 3658 6104 3678
rect 6104 3658 6121 3678
rect 6069 3626 6121 3658
rect 6133 3658 6142 3678
rect 6142 3658 6176 3678
rect 6176 3658 6185 3678
rect 6133 3626 6185 3658
rect 6197 3658 6214 3678
rect 6214 3658 6248 3678
rect 6248 3658 6249 3678
rect 6197 3626 6249 3658
rect 6069 3584 6070 3613
rect 6070 3584 6104 3613
rect 6104 3584 6121 3613
rect 6069 3561 6121 3584
rect 6133 3584 6142 3613
rect 6142 3584 6176 3613
rect 6176 3584 6185 3613
rect 6133 3561 6185 3584
rect 6197 3584 6214 3613
rect 6214 3584 6248 3613
rect 6248 3584 6249 3613
rect 6197 3561 6249 3584
rect 6069 3544 6121 3548
rect 6069 3510 6070 3544
rect 6070 3510 6104 3544
rect 6104 3510 6121 3544
rect 6069 3496 6121 3510
rect 6133 3544 6185 3548
rect 6133 3510 6142 3544
rect 6142 3510 6176 3544
rect 6176 3510 6185 3544
rect 6133 3496 6185 3510
rect 6197 3544 6249 3548
rect 6197 3510 6214 3544
rect 6214 3510 6248 3544
rect 6248 3510 6249 3544
rect 6197 3496 6249 3510
rect 6069 3470 6121 3483
rect 6069 3436 6070 3470
rect 6070 3436 6104 3470
rect 6104 3436 6121 3470
rect 6069 3431 6121 3436
rect 6133 3470 6185 3483
rect 6133 3436 6142 3470
rect 6142 3436 6176 3470
rect 6176 3436 6185 3470
rect 6133 3431 6185 3436
rect 6197 3470 6249 3483
rect 6197 3436 6214 3470
rect 6214 3436 6248 3470
rect 6248 3436 6249 3470
rect 6197 3431 6249 3436
rect 6069 3396 6121 3418
rect 6069 3366 6070 3396
rect 6070 3366 6104 3396
rect 6104 3366 6121 3396
rect 6133 3396 6185 3418
rect 6133 3366 6142 3396
rect 6142 3366 6176 3396
rect 6176 3366 6185 3396
rect 6197 3396 6249 3418
rect 6197 3366 6214 3396
rect 6214 3366 6248 3396
rect 6248 3366 6249 3396
rect 6069 3322 6121 3353
rect 6069 3301 6070 3322
rect 6070 3301 6104 3322
rect 6104 3301 6121 3322
rect 6133 3322 6185 3353
rect 6133 3301 6142 3322
rect 6142 3301 6176 3322
rect 6176 3301 6185 3322
rect 6197 3322 6249 3353
rect 6197 3301 6214 3322
rect 6214 3301 6248 3322
rect 6248 3301 6249 3322
rect 6069 3248 6121 3288
rect 6069 3236 6070 3248
rect 6070 3236 6104 3248
rect 6104 3236 6121 3248
rect 6133 3248 6185 3288
rect 6133 3236 6142 3248
rect 6142 3236 6176 3248
rect 6176 3236 6185 3248
rect 6197 3248 6249 3288
rect 6197 3236 6214 3248
rect 6214 3236 6248 3248
rect 6248 3236 6249 3248
rect 6069 3214 6070 3223
rect 6070 3214 6104 3223
rect 6104 3214 6121 3223
rect 6069 3174 6121 3214
rect 6069 3171 6070 3174
rect 6070 3171 6104 3174
rect 6104 3171 6121 3174
rect 6133 3214 6142 3223
rect 6142 3214 6176 3223
rect 6176 3214 6185 3223
rect 6133 3174 6185 3214
rect 6133 3171 6142 3174
rect 6142 3171 6176 3174
rect 6176 3171 6185 3174
rect 6197 3214 6214 3223
rect 6214 3214 6248 3223
rect 6248 3214 6249 3223
rect 6197 3174 6249 3214
rect 6197 3171 6214 3174
rect 6214 3171 6248 3174
rect 6248 3171 6249 3174
rect 6069 3140 6070 3158
rect 6070 3140 6104 3158
rect 6104 3140 6121 3158
rect 6069 3106 6121 3140
rect 6133 3140 6142 3158
rect 6142 3140 6176 3158
rect 6176 3140 6185 3158
rect 6133 3106 6185 3140
rect 6197 3140 6214 3158
rect 6214 3140 6248 3158
rect 6248 3140 6249 3158
rect 6197 3106 6249 3140
rect 6069 3066 6070 3093
rect 6070 3066 6104 3093
rect 6104 3066 6121 3093
rect 6069 3041 6121 3066
rect 6133 3066 6142 3093
rect 6142 3066 6176 3093
rect 6176 3066 6185 3093
rect 6133 3041 6185 3066
rect 6197 3066 6214 3093
rect 6214 3066 6248 3093
rect 6248 3066 6249 3093
rect 6197 3041 6249 3066
rect 6069 3026 6121 3028
rect 6069 2992 6070 3026
rect 6070 2992 6104 3026
rect 6104 2992 6121 3026
rect 6069 2976 6121 2992
rect 6133 3026 6185 3028
rect 6133 2992 6142 3026
rect 6142 2992 6176 3026
rect 6176 2992 6185 3026
rect 6133 2976 6185 2992
rect 6197 3026 6249 3028
rect 6197 2992 6214 3026
rect 6214 2992 6248 3026
rect 6248 2992 6249 3026
rect 6197 2976 6249 2992
rect 6069 2952 6121 2963
rect 6069 2918 6070 2952
rect 6070 2918 6104 2952
rect 6104 2918 6121 2952
rect 6069 2911 6121 2918
rect 6133 2952 6185 2963
rect 6133 2918 6142 2952
rect 6142 2918 6176 2952
rect 6176 2918 6185 2952
rect 6133 2911 6185 2918
rect 6197 2952 6249 2963
rect 6197 2918 6214 2952
rect 6214 2918 6248 2952
rect 6248 2918 6249 2952
rect 6197 2911 6249 2918
rect 6069 2878 6121 2898
rect 6069 2846 6070 2878
rect 6070 2846 6104 2878
rect 6104 2846 6121 2878
rect 6133 2878 6185 2898
rect 6133 2846 6142 2878
rect 6142 2846 6176 2878
rect 6176 2846 6185 2878
rect 6197 2878 6249 2898
rect 6197 2846 6214 2878
rect 6214 2846 6248 2878
rect 6248 2846 6249 2878
rect 6069 2804 6121 2833
rect 6069 2781 6070 2804
rect 6070 2781 6104 2804
rect 6104 2781 6121 2804
rect 6133 2804 6185 2833
rect 6133 2781 6142 2804
rect 6142 2781 6176 2804
rect 6176 2781 6185 2804
rect 6197 2804 6249 2833
rect 6197 2781 6214 2804
rect 6214 2781 6248 2804
rect 6248 2781 6249 2804
rect 6069 2730 6121 2768
rect 6069 2716 6070 2730
rect 6070 2716 6104 2730
rect 6104 2716 6121 2730
rect 6133 2730 6185 2768
rect 6133 2716 6142 2730
rect 6142 2716 6176 2730
rect 6176 2716 6185 2730
rect 6197 2730 6249 2768
rect 6197 2716 6214 2730
rect 6214 2716 6248 2730
rect 6248 2716 6249 2730
rect 6069 2696 6070 2703
rect 6070 2696 6104 2703
rect 6104 2696 6121 2703
rect 6069 2656 6121 2696
rect 6069 2651 6070 2656
rect 6070 2651 6104 2656
rect 6104 2651 6121 2656
rect 6133 2696 6142 2703
rect 6142 2696 6176 2703
rect 6176 2696 6185 2703
rect 6133 2656 6185 2696
rect 6133 2651 6142 2656
rect 6142 2651 6176 2656
rect 6176 2651 6185 2656
rect 6197 2696 6214 2703
rect 6214 2696 6248 2703
rect 6248 2696 6249 2703
rect 6197 2656 6249 2696
rect 6197 2651 6214 2656
rect 6214 2651 6248 2656
rect 6248 2651 6249 2656
rect 6069 2622 6070 2638
rect 6070 2622 6104 2638
rect 6104 2622 6121 2638
rect 6069 2586 6121 2622
rect 6133 2622 6142 2638
rect 6142 2622 6176 2638
rect 6176 2622 6185 2638
rect 6133 2586 6185 2622
rect 6197 2622 6214 2638
rect 6214 2622 6248 2638
rect 6248 2622 6249 2638
rect 6197 2586 6249 2622
rect 6069 2548 6070 2573
rect 6070 2548 6104 2573
rect 6104 2548 6121 2573
rect 6069 2521 6121 2548
rect 6133 2548 6142 2573
rect 6142 2548 6176 2573
rect 6176 2548 6185 2573
rect 6133 2521 6185 2548
rect 6197 2548 6214 2573
rect 6214 2548 6248 2573
rect 6248 2548 6249 2573
rect 6197 2521 6249 2548
rect 6069 2474 6070 2508
rect 6070 2474 6104 2508
rect 6104 2474 6121 2508
rect 6069 2456 6121 2474
rect 6133 2474 6142 2508
rect 6142 2474 6176 2508
rect 6176 2474 6185 2508
rect 6133 2456 6185 2474
rect 6197 2474 6214 2508
rect 6214 2474 6248 2508
rect 6248 2474 6249 2508
rect 6197 2456 6249 2474
rect 6069 2434 6121 2443
rect 6069 2400 6070 2434
rect 6070 2400 6104 2434
rect 6104 2400 6121 2434
rect 6069 2391 6121 2400
rect 6133 2434 6185 2443
rect 6133 2400 6142 2434
rect 6142 2400 6176 2434
rect 6176 2400 6185 2434
rect 6133 2391 6185 2400
rect 6197 2434 6249 2443
rect 6197 2400 6214 2434
rect 6214 2400 6248 2434
rect 6248 2400 6249 2434
rect 6197 2391 6249 2400
rect 6069 2360 6121 2378
rect 6069 2326 6070 2360
rect 6070 2326 6104 2360
rect 6104 2326 6121 2360
rect 6133 2360 6185 2378
rect 6133 2326 6142 2360
rect 6142 2326 6176 2360
rect 6176 2326 6185 2360
rect 6197 2360 6249 2378
rect 6197 2326 6214 2360
rect 6214 2326 6248 2360
rect 6248 2326 6249 2360
rect 6069 2286 6121 2313
rect 6069 2261 6070 2286
rect 6070 2261 6104 2286
rect 6104 2261 6121 2286
rect 6133 2286 6185 2313
rect 6133 2261 6142 2286
rect 6142 2261 6176 2286
rect 6176 2261 6185 2286
rect 6197 2286 6249 2313
rect 6197 2261 6214 2286
rect 6214 2261 6248 2286
rect 6248 2261 6249 2286
rect 6069 2212 6121 2248
rect 6069 2196 6070 2212
rect 6070 2196 6104 2212
rect 6104 2196 6121 2212
rect 6133 2212 6185 2248
rect 6133 2196 6142 2212
rect 6142 2196 6176 2212
rect 6176 2196 6185 2212
rect 6197 2212 6249 2248
rect 6197 2196 6214 2212
rect 6214 2196 6248 2212
rect 6248 2196 6249 2212
rect 6069 2178 6070 2183
rect 6070 2178 6104 2183
rect 6104 2178 6121 2183
rect 6069 2138 6121 2178
rect 6069 2131 6070 2138
rect 6070 2131 6104 2138
rect 6104 2131 6121 2138
rect 6133 2178 6142 2183
rect 6142 2178 6176 2183
rect 6176 2178 6185 2183
rect 6133 2138 6185 2178
rect 6133 2131 6142 2138
rect 6142 2131 6176 2138
rect 6176 2131 6185 2138
rect 6197 2178 6214 2183
rect 6214 2178 6248 2183
rect 6248 2178 6249 2183
rect 6197 2138 6249 2178
rect 6197 2131 6214 2138
rect 6214 2131 6248 2138
rect 6248 2131 6249 2138
rect 6069 2104 6070 2118
rect 6070 2104 6104 2118
rect 6104 2104 6121 2118
rect 6069 2066 6121 2104
rect 6133 2104 6142 2118
rect 6142 2104 6176 2118
rect 6176 2104 6185 2118
rect 6133 2066 6185 2104
rect 6197 2104 6214 2118
rect 6214 2104 6248 2118
rect 6248 2104 6249 2118
rect 6197 2066 6249 2104
rect 6069 2030 6070 2053
rect 6070 2030 6104 2053
rect 6104 2030 6121 2053
rect 6069 2001 6121 2030
rect 6133 2030 6142 2053
rect 6142 2030 6176 2053
rect 6176 2030 6185 2053
rect 6133 2001 6185 2030
rect 6197 2030 6214 2053
rect 6214 2030 6248 2053
rect 6248 2030 6249 2053
rect 6197 2001 6249 2030
rect 6069 1956 6070 1987
rect 6070 1956 6104 1987
rect 6104 1956 6121 1987
rect 6069 1935 6121 1956
rect 6133 1956 6142 1987
rect 6142 1956 6176 1987
rect 6176 1956 6185 1987
rect 6133 1935 6185 1956
rect 6197 1956 6214 1987
rect 6214 1956 6248 1987
rect 6248 1956 6249 1987
rect 6197 1935 6249 1956
rect 6069 1916 6121 1921
rect 6069 1882 6070 1916
rect 6070 1882 6104 1916
rect 6104 1882 6121 1916
rect 6069 1869 6121 1882
rect 6133 1916 6185 1921
rect 6133 1882 6142 1916
rect 6142 1882 6176 1916
rect 6176 1882 6185 1916
rect 6133 1869 6185 1882
rect 6197 1916 6249 1921
rect 6197 1882 6214 1916
rect 6214 1882 6248 1916
rect 6248 1882 6249 1916
rect 6197 1869 6249 1882
rect 6069 1842 6121 1855
rect 6069 1808 6070 1842
rect 6070 1808 6104 1842
rect 6104 1808 6121 1842
rect 6069 1803 6121 1808
rect 6133 1842 6185 1855
rect 6133 1808 6142 1842
rect 6142 1808 6176 1842
rect 6176 1808 6185 1842
rect 6133 1803 6185 1808
rect 6197 1842 6249 1855
rect 6197 1808 6214 1842
rect 6214 1808 6248 1842
rect 6248 1808 6249 1842
rect 6197 1803 6249 1808
rect 6069 1768 6121 1789
rect 6069 1737 6070 1768
rect 6070 1737 6104 1768
rect 6104 1737 6121 1768
rect 6133 1768 6185 1789
rect 6133 1737 6142 1768
rect 6142 1737 6176 1768
rect 6176 1737 6185 1768
rect 6197 1768 6249 1789
rect 6197 1737 6214 1768
rect 6214 1737 6248 1768
rect 6248 1737 6249 1768
rect 6069 1694 6121 1723
rect 6069 1671 6070 1694
rect 6070 1671 6104 1694
rect 6104 1671 6121 1694
rect 6133 1694 6185 1723
rect 6133 1671 6142 1694
rect 6142 1671 6176 1694
rect 6176 1671 6185 1694
rect 6197 1694 6249 1723
rect 6197 1671 6214 1694
rect 6214 1671 6248 1694
rect 6248 1671 6249 1694
rect 6069 1620 6121 1657
rect 6069 1605 6070 1620
rect 6070 1605 6104 1620
rect 6104 1605 6121 1620
rect 6133 1620 6185 1657
rect 6133 1605 6142 1620
rect 6142 1605 6176 1620
rect 6176 1605 6185 1620
rect 6197 1620 6249 1657
rect 6197 1605 6214 1620
rect 6214 1605 6248 1620
rect 6248 1605 6249 1620
rect 6069 1586 6070 1591
rect 6070 1586 6104 1591
rect 6104 1586 6121 1591
rect 6069 1545 6121 1586
rect 6069 1539 6070 1545
rect 6070 1539 6104 1545
rect 6104 1539 6121 1545
rect 6133 1586 6142 1591
rect 6142 1586 6176 1591
rect 6176 1586 6185 1591
rect 6133 1545 6185 1586
rect 6133 1539 6142 1545
rect 6142 1539 6176 1545
rect 6176 1539 6185 1545
rect 6197 1586 6214 1591
rect 6214 1586 6248 1591
rect 6248 1586 6249 1591
rect 6197 1545 6249 1586
rect 6197 1539 6214 1545
rect 6214 1539 6248 1545
rect 6248 1539 6249 1545
rect 6069 1511 6070 1525
rect 6070 1511 6104 1525
rect 6104 1511 6121 1525
rect 6069 1473 6121 1511
rect 6133 1511 6142 1525
rect 6142 1511 6176 1525
rect 6176 1511 6185 1525
rect 6133 1473 6185 1511
rect 6197 1511 6214 1525
rect 6214 1511 6248 1525
rect 6248 1511 6249 1525
rect 6197 1473 6249 1511
rect 6565 4050 6617 4068
rect 6629 4062 6681 4068
rect 6629 4050 6638 4062
rect 6638 4050 6672 4062
rect 6672 4050 6681 4062
rect 6693 4050 6745 4068
rect 6565 4016 6566 4050
rect 6566 4016 6617 4050
rect 6629 4016 6681 4050
rect 6693 4016 6744 4050
rect 6744 4016 6745 4050
rect 6565 3951 6566 4003
rect 6566 3951 6617 4003
rect 6629 3951 6681 4003
rect 6693 3951 6744 4003
rect 6744 3951 6745 4003
rect 6565 3886 6566 3938
rect 6566 3886 6617 3938
rect 6629 3886 6681 3938
rect 6693 3886 6744 3938
rect 6744 3886 6745 3938
rect 6565 3821 6566 3873
rect 6566 3821 6617 3873
rect 6629 3821 6681 3873
rect 6693 3821 6744 3873
rect 6744 3821 6745 3873
rect 6565 3756 6566 3808
rect 6566 3756 6617 3808
rect 6629 3756 6681 3808
rect 6693 3756 6744 3808
rect 6744 3756 6745 3808
rect 6565 3691 6566 3743
rect 6566 3691 6617 3743
rect 6629 3691 6681 3743
rect 6693 3691 6744 3743
rect 6744 3691 6745 3743
rect 6565 3626 6566 3678
rect 6566 3626 6617 3678
rect 6629 3626 6681 3678
rect 6693 3626 6744 3678
rect 6744 3626 6745 3678
rect 6565 3561 6566 3613
rect 6566 3561 6617 3613
rect 6629 3561 6681 3613
rect 6693 3561 6744 3613
rect 6744 3561 6745 3613
rect 6565 3496 6566 3548
rect 6566 3496 6617 3548
rect 6629 3496 6681 3548
rect 6693 3496 6744 3548
rect 6744 3496 6745 3548
rect 6565 3431 6566 3483
rect 6566 3431 6617 3483
rect 6629 3431 6681 3483
rect 6693 3431 6744 3483
rect 6744 3431 6745 3483
rect 6565 3366 6566 3418
rect 6566 3366 6617 3418
rect 6629 3366 6681 3418
rect 6693 3366 6744 3418
rect 6744 3366 6745 3418
rect 6565 3301 6566 3353
rect 6566 3301 6617 3353
rect 6629 3301 6681 3353
rect 6693 3301 6744 3353
rect 6744 3301 6745 3353
rect 6565 3236 6566 3288
rect 6566 3236 6617 3288
rect 6629 3236 6681 3288
rect 6693 3236 6744 3288
rect 6744 3236 6745 3288
rect 6565 3171 6566 3223
rect 6566 3171 6617 3223
rect 6629 3171 6681 3223
rect 6693 3171 6744 3223
rect 6744 3171 6745 3223
rect 6565 3106 6566 3158
rect 6566 3106 6617 3158
rect 6629 3106 6681 3158
rect 6693 3106 6744 3158
rect 6744 3106 6745 3158
rect 6565 3080 6566 3093
rect 6566 3092 6617 3093
rect 6629 3092 6681 3093
rect 6693 3092 6744 3093
rect 6566 3080 6600 3092
rect 6600 3080 6617 3092
rect 6565 3041 6617 3080
rect 6629 3041 6681 3092
rect 6693 3080 6710 3092
rect 6710 3080 6744 3092
rect 6744 3080 6745 3093
rect 6693 3041 6745 3080
rect 6565 2976 6566 3028
rect 6566 2976 6617 3028
rect 6629 2976 6681 3028
rect 6693 2976 6744 3028
rect 6744 2976 6745 3028
rect 6565 2911 6566 2963
rect 6566 2911 6617 2963
rect 6629 2911 6681 2963
rect 6693 2911 6744 2963
rect 6744 2911 6745 2963
rect 6565 2846 6566 2898
rect 6566 2846 6617 2898
rect 6629 2846 6681 2898
rect 6693 2846 6744 2898
rect 6744 2846 6745 2898
rect 6565 2781 6566 2833
rect 6566 2781 6617 2833
rect 6629 2781 6681 2833
rect 6693 2781 6744 2833
rect 6744 2781 6745 2833
rect 6565 2716 6566 2768
rect 6566 2716 6617 2768
rect 6629 2716 6681 2768
rect 6693 2716 6744 2768
rect 6744 2716 6745 2768
rect 6565 2651 6566 2703
rect 6566 2651 6617 2703
rect 6629 2651 6681 2703
rect 6693 2651 6744 2703
rect 6744 2651 6745 2703
rect 6565 2586 6566 2638
rect 6566 2586 6617 2638
rect 6629 2586 6681 2638
rect 6693 2586 6744 2638
rect 6744 2586 6745 2638
rect 6565 2535 6617 2573
rect 6565 2521 6566 2535
rect 6566 2521 6600 2535
rect 6600 2521 6617 2535
rect 6629 2535 6681 2573
rect 6629 2521 6638 2535
rect 6638 2521 6672 2535
rect 6672 2521 6681 2535
rect 6693 2535 6745 2573
rect 6693 2521 6710 2535
rect 6710 2521 6744 2535
rect 6744 2521 6745 2535
rect 6565 2501 6566 2508
rect 6566 2501 6600 2508
rect 6600 2501 6617 2508
rect 6565 2456 6617 2501
rect 6629 2501 6638 2508
rect 6638 2501 6672 2508
rect 6672 2501 6681 2508
rect 6629 2461 6681 2501
rect 6629 2456 6638 2461
rect 6638 2456 6672 2461
rect 6672 2456 6681 2461
rect 6693 2501 6710 2508
rect 6710 2501 6744 2508
rect 6744 2501 6745 2508
rect 6693 2456 6745 2501
rect 6565 2391 6566 2443
rect 6566 2391 6617 2443
rect 6629 2391 6681 2443
rect 6693 2391 6744 2443
rect 6744 2391 6745 2443
rect 6565 2326 6566 2378
rect 6566 2326 6617 2378
rect 6629 2326 6681 2378
rect 6693 2326 6744 2378
rect 6744 2326 6745 2378
rect 6565 2261 6566 2313
rect 6566 2261 6617 2313
rect 6629 2261 6681 2313
rect 6693 2261 6744 2313
rect 6744 2261 6745 2313
rect 6565 2196 6566 2248
rect 6566 2196 6617 2248
rect 6629 2196 6681 2248
rect 6693 2196 6744 2248
rect 6744 2196 6745 2248
rect 6565 2131 6566 2183
rect 6566 2131 6617 2183
rect 6629 2131 6681 2183
rect 6693 2131 6744 2183
rect 6744 2131 6745 2183
rect 6565 2066 6566 2118
rect 6566 2066 6617 2118
rect 6629 2066 6681 2118
rect 6693 2066 6744 2118
rect 6744 2066 6745 2118
rect 6565 2001 6566 2053
rect 6566 2001 6617 2053
rect 6629 2001 6681 2053
rect 6693 2001 6744 2053
rect 6744 2001 6745 2053
rect 6565 1935 6566 1987
rect 6566 1935 6617 1987
rect 6629 1935 6681 1987
rect 6693 1935 6744 1987
rect 6744 1935 6745 1987
rect 6565 1869 6566 1921
rect 6566 1869 6617 1921
rect 6629 1869 6681 1921
rect 6693 1869 6744 1921
rect 6744 1869 6745 1921
rect 6565 1803 6566 1855
rect 6566 1803 6617 1855
rect 6629 1803 6681 1855
rect 6693 1803 6744 1855
rect 6744 1803 6745 1855
rect 6565 1737 6566 1789
rect 6566 1737 6617 1789
rect 6629 1737 6681 1789
rect 6693 1737 6744 1789
rect 6744 1737 6745 1789
rect 6565 1671 6566 1723
rect 6566 1671 6617 1723
rect 6629 1671 6681 1723
rect 6693 1671 6744 1723
rect 6744 1671 6745 1723
rect 6565 1605 6566 1657
rect 6566 1605 6617 1657
rect 6629 1605 6681 1657
rect 6693 1605 6744 1657
rect 6744 1605 6745 1657
rect 6565 1539 6566 1591
rect 6566 1539 6617 1591
rect 6629 1539 6681 1591
rect 6693 1539 6744 1591
rect 6744 1539 6745 1591
rect 6565 1479 6566 1525
rect 6566 1491 6617 1525
rect 6629 1491 6681 1525
rect 6693 1491 6744 1525
rect 6566 1479 6600 1491
rect 6600 1479 6617 1491
rect 6565 1473 6617 1479
rect 6629 1473 6681 1491
rect 6693 1479 6710 1491
rect 6710 1479 6744 1491
rect 6744 1479 6745 1525
rect 6693 1473 6745 1479
rect 7061 4062 7113 4068
rect 7061 4028 7062 4062
rect 7062 4028 7096 4062
rect 7096 4028 7113 4062
rect 7061 4016 7113 4028
rect 7125 4062 7177 4068
rect 7125 4028 7134 4062
rect 7134 4028 7168 4062
rect 7168 4028 7177 4062
rect 7125 4016 7177 4028
rect 7189 4062 7241 4068
rect 7189 4028 7206 4062
rect 7206 4028 7240 4062
rect 7240 4028 7241 4062
rect 7189 4016 7241 4028
rect 7061 3988 7113 4003
rect 7061 3954 7062 3988
rect 7062 3954 7096 3988
rect 7096 3954 7113 3988
rect 7061 3951 7113 3954
rect 7125 3988 7177 4003
rect 7125 3954 7134 3988
rect 7134 3954 7168 3988
rect 7168 3954 7177 3988
rect 7125 3951 7177 3954
rect 7189 3988 7241 4003
rect 7189 3954 7206 3988
rect 7206 3954 7240 3988
rect 7240 3954 7241 3988
rect 7189 3951 7241 3954
rect 7061 3914 7113 3938
rect 7061 3886 7062 3914
rect 7062 3886 7096 3914
rect 7096 3886 7113 3914
rect 7125 3914 7177 3938
rect 7125 3886 7134 3914
rect 7134 3886 7168 3914
rect 7168 3886 7177 3914
rect 7189 3914 7241 3938
rect 7189 3886 7206 3914
rect 7206 3886 7240 3914
rect 7240 3886 7241 3914
rect 7061 3840 7113 3873
rect 7061 3821 7062 3840
rect 7062 3821 7096 3840
rect 7096 3821 7113 3840
rect 7125 3840 7177 3873
rect 7125 3821 7134 3840
rect 7134 3821 7168 3840
rect 7168 3821 7177 3840
rect 7189 3840 7241 3873
rect 7189 3821 7206 3840
rect 7206 3821 7240 3840
rect 7240 3821 7241 3840
rect 7061 3806 7062 3808
rect 7062 3806 7096 3808
rect 7096 3806 7113 3808
rect 7061 3766 7113 3806
rect 7061 3756 7062 3766
rect 7062 3756 7096 3766
rect 7096 3756 7113 3766
rect 7125 3806 7134 3808
rect 7134 3806 7168 3808
rect 7168 3806 7177 3808
rect 7125 3766 7177 3806
rect 7125 3756 7134 3766
rect 7134 3756 7168 3766
rect 7168 3756 7177 3766
rect 7189 3806 7206 3808
rect 7206 3806 7240 3808
rect 7240 3806 7241 3808
rect 7189 3766 7241 3806
rect 7189 3756 7206 3766
rect 7206 3756 7240 3766
rect 7240 3756 7241 3766
rect 7061 3732 7062 3743
rect 7062 3732 7096 3743
rect 7096 3732 7113 3743
rect 7061 3692 7113 3732
rect 7061 3691 7062 3692
rect 7062 3691 7096 3692
rect 7096 3691 7113 3692
rect 7125 3732 7134 3743
rect 7134 3732 7168 3743
rect 7168 3732 7177 3743
rect 7125 3692 7177 3732
rect 7125 3691 7134 3692
rect 7134 3691 7168 3692
rect 7168 3691 7177 3692
rect 7189 3732 7206 3743
rect 7206 3732 7240 3743
rect 7240 3732 7241 3743
rect 7189 3692 7241 3732
rect 7189 3691 7206 3692
rect 7206 3691 7240 3692
rect 7240 3691 7241 3692
rect 7061 3658 7062 3678
rect 7062 3658 7096 3678
rect 7096 3658 7113 3678
rect 7061 3626 7113 3658
rect 7125 3658 7134 3678
rect 7134 3658 7168 3678
rect 7168 3658 7177 3678
rect 7125 3626 7177 3658
rect 7189 3658 7206 3678
rect 7206 3658 7240 3678
rect 7240 3658 7241 3678
rect 7189 3626 7241 3658
rect 7061 3584 7062 3613
rect 7062 3584 7096 3613
rect 7096 3584 7113 3613
rect 7061 3561 7113 3584
rect 7125 3584 7134 3613
rect 7134 3584 7168 3613
rect 7168 3584 7177 3613
rect 7125 3561 7177 3584
rect 7189 3584 7206 3613
rect 7206 3584 7240 3613
rect 7240 3584 7241 3613
rect 7189 3561 7241 3584
rect 7061 3544 7113 3548
rect 7061 3510 7062 3544
rect 7062 3510 7096 3544
rect 7096 3510 7113 3544
rect 7061 3496 7113 3510
rect 7125 3544 7177 3548
rect 7125 3510 7134 3544
rect 7134 3510 7168 3544
rect 7168 3510 7177 3544
rect 7125 3496 7177 3510
rect 7189 3544 7241 3548
rect 7189 3510 7206 3544
rect 7206 3510 7240 3544
rect 7240 3510 7241 3544
rect 7189 3496 7241 3510
rect 7061 3470 7113 3483
rect 7061 3436 7062 3470
rect 7062 3436 7096 3470
rect 7096 3436 7113 3470
rect 7061 3431 7113 3436
rect 7125 3470 7177 3483
rect 7125 3436 7134 3470
rect 7134 3436 7168 3470
rect 7168 3436 7177 3470
rect 7125 3431 7177 3436
rect 7189 3470 7241 3483
rect 7189 3436 7206 3470
rect 7206 3436 7240 3470
rect 7240 3436 7241 3470
rect 7189 3431 7241 3436
rect 7061 3396 7113 3418
rect 7061 3366 7062 3396
rect 7062 3366 7096 3396
rect 7096 3366 7113 3396
rect 7125 3396 7177 3418
rect 7125 3366 7134 3396
rect 7134 3366 7168 3396
rect 7168 3366 7177 3396
rect 7189 3396 7241 3418
rect 7189 3366 7206 3396
rect 7206 3366 7240 3396
rect 7240 3366 7241 3396
rect 7061 3322 7113 3353
rect 7061 3301 7062 3322
rect 7062 3301 7096 3322
rect 7096 3301 7113 3322
rect 7125 3322 7177 3353
rect 7125 3301 7134 3322
rect 7134 3301 7168 3322
rect 7168 3301 7177 3322
rect 7189 3322 7241 3353
rect 7189 3301 7206 3322
rect 7206 3301 7240 3322
rect 7240 3301 7241 3322
rect 7061 3248 7113 3288
rect 7061 3236 7062 3248
rect 7062 3236 7096 3248
rect 7096 3236 7113 3248
rect 7125 3248 7177 3288
rect 7125 3236 7134 3248
rect 7134 3236 7168 3248
rect 7168 3236 7177 3248
rect 7189 3248 7241 3288
rect 7189 3236 7206 3248
rect 7206 3236 7240 3248
rect 7240 3236 7241 3248
rect 7061 3214 7062 3223
rect 7062 3214 7096 3223
rect 7096 3214 7113 3223
rect 7061 3174 7113 3214
rect 7061 3171 7062 3174
rect 7062 3171 7096 3174
rect 7096 3171 7113 3174
rect 7125 3214 7134 3223
rect 7134 3214 7168 3223
rect 7168 3214 7177 3223
rect 7125 3174 7177 3214
rect 7125 3171 7134 3174
rect 7134 3171 7168 3174
rect 7168 3171 7177 3174
rect 7189 3214 7206 3223
rect 7206 3214 7240 3223
rect 7240 3214 7241 3223
rect 7189 3174 7241 3214
rect 7189 3171 7206 3174
rect 7206 3171 7240 3174
rect 7240 3171 7241 3174
rect 7061 3140 7062 3158
rect 7062 3140 7096 3158
rect 7096 3140 7113 3158
rect 7061 3106 7113 3140
rect 7125 3140 7134 3158
rect 7134 3140 7168 3158
rect 7168 3140 7177 3158
rect 7125 3106 7177 3140
rect 7189 3140 7206 3158
rect 7206 3140 7240 3158
rect 7240 3140 7241 3158
rect 7189 3106 7241 3140
rect 7061 3066 7062 3093
rect 7062 3066 7096 3093
rect 7096 3066 7113 3093
rect 7061 3041 7113 3066
rect 7125 3066 7134 3093
rect 7134 3066 7168 3093
rect 7168 3066 7177 3093
rect 7125 3041 7177 3066
rect 7189 3066 7206 3093
rect 7206 3066 7240 3093
rect 7240 3066 7241 3093
rect 7189 3041 7241 3066
rect 7061 3026 7113 3028
rect 7061 2992 7062 3026
rect 7062 2992 7096 3026
rect 7096 2992 7113 3026
rect 7061 2976 7113 2992
rect 7125 3026 7177 3028
rect 7125 2992 7134 3026
rect 7134 2992 7168 3026
rect 7168 2992 7177 3026
rect 7125 2976 7177 2992
rect 7189 3026 7241 3028
rect 7189 2992 7206 3026
rect 7206 2992 7240 3026
rect 7240 2992 7241 3026
rect 7189 2976 7241 2992
rect 7061 2952 7113 2963
rect 7061 2918 7062 2952
rect 7062 2918 7096 2952
rect 7096 2918 7113 2952
rect 7061 2911 7113 2918
rect 7125 2952 7177 2963
rect 7125 2918 7134 2952
rect 7134 2918 7168 2952
rect 7168 2918 7177 2952
rect 7125 2911 7177 2918
rect 7189 2952 7241 2963
rect 7189 2918 7206 2952
rect 7206 2918 7240 2952
rect 7240 2918 7241 2952
rect 7189 2911 7241 2918
rect 7061 2878 7113 2898
rect 7061 2846 7062 2878
rect 7062 2846 7096 2878
rect 7096 2846 7113 2878
rect 7125 2878 7177 2898
rect 7125 2846 7134 2878
rect 7134 2846 7168 2878
rect 7168 2846 7177 2878
rect 7189 2878 7241 2898
rect 7189 2846 7206 2878
rect 7206 2846 7240 2878
rect 7240 2846 7241 2878
rect 7061 2804 7113 2833
rect 7061 2781 7062 2804
rect 7062 2781 7096 2804
rect 7096 2781 7113 2804
rect 7125 2804 7177 2833
rect 7125 2781 7134 2804
rect 7134 2781 7168 2804
rect 7168 2781 7177 2804
rect 7189 2804 7241 2833
rect 7189 2781 7206 2804
rect 7206 2781 7240 2804
rect 7240 2781 7241 2804
rect 7061 2730 7113 2768
rect 7061 2716 7062 2730
rect 7062 2716 7096 2730
rect 7096 2716 7113 2730
rect 7125 2730 7177 2768
rect 7125 2716 7134 2730
rect 7134 2716 7168 2730
rect 7168 2716 7177 2730
rect 7189 2730 7241 2768
rect 7189 2716 7206 2730
rect 7206 2716 7240 2730
rect 7240 2716 7241 2730
rect 7061 2696 7062 2703
rect 7062 2696 7096 2703
rect 7096 2696 7113 2703
rect 7061 2656 7113 2696
rect 7061 2651 7062 2656
rect 7062 2651 7096 2656
rect 7096 2651 7113 2656
rect 7125 2696 7134 2703
rect 7134 2696 7168 2703
rect 7168 2696 7177 2703
rect 7125 2656 7177 2696
rect 7125 2651 7134 2656
rect 7134 2651 7168 2656
rect 7168 2651 7177 2656
rect 7189 2696 7206 2703
rect 7206 2696 7240 2703
rect 7240 2696 7241 2703
rect 7189 2656 7241 2696
rect 7189 2651 7206 2656
rect 7206 2651 7240 2656
rect 7240 2651 7241 2656
rect 7061 2622 7062 2638
rect 7062 2622 7096 2638
rect 7096 2622 7113 2638
rect 7061 2586 7113 2622
rect 7125 2622 7134 2638
rect 7134 2622 7168 2638
rect 7168 2622 7177 2638
rect 7125 2586 7177 2622
rect 7189 2622 7206 2638
rect 7206 2622 7240 2638
rect 7240 2622 7241 2638
rect 7189 2586 7241 2622
rect 7061 2548 7062 2573
rect 7062 2548 7096 2573
rect 7096 2548 7113 2573
rect 7061 2521 7113 2548
rect 7125 2548 7134 2573
rect 7134 2548 7168 2573
rect 7168 2548 7177 2573
rect 7125 2521 7177 2548
rect 7189 2548 7206 2573
rect 7206 2548 7240 2573
rect 7240 2548 7241 2573
rect 7189 2521 7241 2548
rect 7061 2474 7062 2508
rect 7062 2474 7096 2508
rect 7096 2474 7113 2508
rect 7061 2456 7113 2474
rect 7125 2474 7134 2508
rect 7134 2474 7168 2508
rect 7168 2474 7177 2508
rect 7125 2456 7177 2474
rect 7189 2474 7206 2508
rect 7206 2474 7240 2508
rect 7240 2474 7241 2508
rect 7189 2456 7241 2474
rect 7061 2434 7113 2443
rect 7061 2400 7062 2434
rect 7062 2400 7096 2434
rect 7096 2400 7113 2434
rect 7061 2391 7113 2400
rect 7125 2434 7177 2443
rect 7125 2400 7134 2434
rect 7134 2400 7168 2434
rect 7168 2400 7177 2434
rect 7125 2391 7177 2400
rect 7189 2434 7241 2443
rect 7189 2400 7206 2434
rect 7206 2400 7240 2434
rect 7240 2400 7241 2434
rect 7189 2391 7241 2400
rect 7061 2360 7113 2378
rect 7061 2326 7062 2360
rect 7062 2326 7096 2360
rect 7096 2326 7113 2360
rect 7125 2360 7177 2378
rect 7125 2326 7134 2360
rect 7134 2326 7168 2360
rect 7168 2326 7177 2360
rect 7189 2360 7241 2378
rect 7189 2326 7206 2360
rect 7206 2326 7240 2360
rect 7240 2326 7241 2360
rect 7061 2286 7113 2313
rect 7061 2261 7062 2286
rect 7062 2261 7096 2286
rect 7096 2261 7113 2286
rect 7125 2286 7177 2313
rect 7125 2261 7134 2286
rect 7134 2261 7168 2286
rect 7168 2261 7177 2286
rect 7189 2286 7241 2313
rect 7189 2261 7206 2286
rect 7206 2261 7240 2286
rect 7240 2261 7241 2286
rect 7061 2212 7113 2248
rect 7061 2196 7062 2212
rect 7062 2196 7096 2212
rect 7096 2196 7113 2212
rect 7125 2212 7177 2248
rect 7125 2196 7134 2212
rect 7134 2196 7168 2212
rect 7168 2196 7177 2212
rect 7189 2212 7241 2248
rect 7189 2196 7206 2212
rect 7206 2196 7240 2212
rect 7240 2196 7241 2212
rect 7061 2178 7062 2183
rect 7062 2178 7096 2183
rect 7096 2178 7113 2183
rect 7061 2138 7113 2178
rect 7061 2131 7062 2138
rect 7062 2131 7096 2138
rect 7096 2131 7113 2138
rect 7125 2178 7134 2183
rect 7134 2178 7168 2183
rect 7168 2178 7177 2183
rect 7125 2138 7177 2178
rect 7125 2131 7134 2138
rect 7134 2131 7168 2138
rect 7168 2131 7177 2138
rect 7189 2178 7206 2183
rect 7206 2178 7240 2183
rect 7240 2178 7241 2183
rect 7189 2138 7241 2178
rect 7189 2131 7206 2138
rect 7206 2131 7240 2138
rect 7240 2131 7241 2138
rect 7061 2104 7062 2118
rect 7062 2104 7096 2118
rect 7096 2104 7113 2118
rect 7061 2066 7113 2104
rect 7125 2104 7134 2118
rect 7134 2104 7168 2118
rect 7168 2104 7177 2118
rect 7125 2066 7177 2104
rect 7189 2104 7206 2118
rect 7206 2104 7240 2118
rect 7240 2104 7241 2118
rect 7189 2066 7241 2104
rect 7061 2030 7062 2053
rect 7062 2030 7096 2053
rect 7096 2030 7113 2053
rect 7061 2001 7113 2030
rect 7125 2030 7134 2053
rect 7134 2030 7168 2053
rect 7168 2030 7177 2053
rect 7125 2001 7177 2030
rect 7189 2030 7206 2053
rect 7206 2030 7240 2053
rect 7240 2030 7241 2053
rect 7189 2001 7241 2030
rect 7061 1956 7062 1987
rect 7062 1956 7096 1987
rect 7096 1956 7113 1987
rect 7061 1935 7113 1956
rect 7125 1956 7134 1987
rect 7134 1956 7168 1987
rect 7168 1956 7177 1987
rect 7125 1935 7177 1956
rect 7189 1956 7206 1987
rect 7206 1956 7240 1987
rect 7240 1956 7241 1987
rect 7189 1935 7241 1956
rect 7061 1916 7113 1921
rect 7061 1882 7062 1916
rect 7062 1882 7096 1916
rect 7096 1882 7113 1916
rect 7061 1869 7113 1882
rect 7125 1916 7177 1921
rect 7125 1882 7134 1916
rect 7134 1882 7168 1916
rect 7168 1882 7177 1916
rect 7125 1869 7177 1882
rect 7189 1916 7241 1921
rect 7189 1882 7206 1916
rect 7206 1882 7240 1916
rect 7240 1882 7241 1916
rect 7189 1869 7241 1882
rect 7061 1842 7113 1855
rect 7061 1808 7062 1842
rect 7062 1808 7096 1842
rect 7096 1808 7113 1842
rect 7061 1803 7113 1808
rect 7125 1842 7177 1855
rect 7125 1808 7134 1842
rect 7134 1808 7168 1842
rect 7168 1808 7177 1842
rect 7125 1803 7177 1808
rect 7189 1842 7241 1855
rect 7189 1808 7206 1842
rect 7206 1808 7240 1842
rect 7240 1808 7241 1842
rect 7189 1803 7241 1808
rect 7061 1768 7113 1789
rect 7061 1737 7062 1768
rect 7062 1737 7096 1768
rect 7096 1737 7113 1768
rect 7125 1768 7177 1789
rect 7125 1737 7134 1768
rect 7134 1737 7168 1768
rect 7168 1737 7177 1768
rect 7189 1768 7241 1789
rect 7189 1737 7206 1768
rect 7206 1737 7240 1768
rect 7240 1737 7241 1768
rect 7061 1694 7113 1723
rect 7061 1671 7062 1694
rect 7062 1671 7096 1694
rect 7096 1671 7113 1694
rect 7125 1694 7177 1723
rect 7125 1671 7134 1694
rect 7134 1671 7168 1694
rect 7168 1671 7177 1694
rect 7189 1694 7241 1723
rect 7189 1671 7206 1694
rect 7206 1671 7240 1694
rect 7240 1671 7241 1694
rect 7061 1620 7113 1657
rect 7061 1605 7062 1620
rect 7062 1605 7096 1620
rect 7096 1605 7113 1620
rect 7125 1620 7177 1657
rect 7125 1605 7134 1620
rect 7134 1605 7168 1620
rect 7168 1605 7177 1620
rect 7189 1620 7241 1657
rect 7189 1605 7206 1620
rect 7206 1605 7240 1620
rect 7240 1605 7241 1620
rect 7061 1586 7062 1591
rect 7062 1586 7096 1591
rect 7096 1586 7113 1591
rect 7061 1545 7113 1586
rect 7061 1539 7062 1545
rect 7062 1539 7096 1545
rect 7096 1539 7113 1545
rect 7125 1586 7134 1591
rect 7134 1586 7168 1591
rect 7168 1586 7177 1591
rect 7125 1545 7177 1586
rect 7125 1539 7134 1545
rect 7134 1539 7168 1545
rect 7168 1539 7177 1545
rect 7189 1586 7206 1591
rect 7206 1586 7240 1591
rect 7240 1586 7241 1591
rect 7189 1545 7241 1586
rect 7189 1539 7206 1545
rect 7206 1539 7240 1545
rect 7240 1539 7241 1545
rect 7061 1511 7062 1525
rect 7062 1511 7096 1525
rect 7096 1511 7113 1525
rect 7061 1473 7113 1511
rect 7125 1511 7134 1525
rect 7134 1511 7168 1525
rect 7168 1511 7177 1525
rect 7125 1473 7177 1511
rect 7189 1511 7206 1525
rect 7206 1511 7240 1525
rect 7240 1511 7241 1525
rect 7189 1473 7241 1511
rect 7557 4050 7609 4068
rect 7621 4062 7673 4068
rect 7621 4050 7630 4062
rect 7630 4050 7664 4062
rect 7664 4050 7673 4062
rect 7685 4050 7737 4068
rect 7557 4016 7558 4050
rect 7558 4016 7609 4050
rect 7621 4016 7673 4050
rect 7685 4016 7736 4050
rect 7736 4016 7737 4050
rect 7557 3951 7558 4003
rect 7558 3951 7609 4003
rect 7621 3951 7673 4003
rect 7685 3951 7736 4003
rect 7736 3951 7737 4003
rect 7557 3886 7558 3938
rect 7558 3886 7609 3938
rect 7621 3886 7673 3938
rect 7685 3886 7736 3938
rect 7736 3886 7737 3938
rect 7557 3821 7558 3873
rect 7558 3821 7609 3873
rect 7621 3821 7673 3873
rect 7685 3821 7736 3873
rect 7736 3821 7737 3873
rect 7557 3756 7558 3808
rect 7558 3756 7609 3808
rect 7621 3756 7673 3808
rect 7685 3756 7736 3808
rect 7736 3756 7737 3808
rect 7557 3691 7558 3743
rect 7558 3691 7609 3743
rect 7621 3691 7673 3743
rect 7685 3691 7736 3743
rect 7736 3691 7737 3743
rect 7557 3626 7558 3678
rect 7558 3626 7609 3678
rect 7621 3626 7673 3678
rect 7685 3626 7736 3678
rect 7736 3626 7737 3678
rect 7557 3561 7558 3613
rect 7558 3561 7609 3613
rect 7621 3561 7673 3613
rect 7685 3561 7736 3613
rect 7736 3561 7737 3613
rect 7557 3496 7558 3548
rect 7558 3496 7609 3548
rect 7621 3496 7673 3548
rect 7685 3496 7736 3548
rect 7736 3496 7737 3548
rect 7557 3431 7558 3483
rect 7558 3431 7609 3483
rect 7621 3431 7673 3483
rect 7685 3431 7736 3483
rect 7736 3431 7737 3483
rect 7557 3366 7558 3418
rect 7558 3366 7609 3418
rect 7621 3366 7673 3418
rect 7685 3366 7736 3418
rect 7736 3366 7737 3418
rect 7557 3301 7558 3353
rect 7558 3301 7609 3353
rect 7621 3301 7673 3353
rect 7685 3301 7736 3353
rect 7736 3301 7737 3353
rect 7557 3236 7558 3288
rect 7558 3236 7609 3288
rect 7621 3236 7673 3288
rect 7685 3236 7736 3288
rect 7736 3236 7737 3288
rect 7557 3171 7558 3223
rect 7558 3171 7609 3223
rect 7621 3171 7673 3223
rect 7685 3171 7736 3223
rect 7736 3171 7737 3223
rect 7557 3106 7558 3158
rect 7558 3106 7609 3158
rect 7621 3106 7673 3158
rect 7685 3106 7736 3158
rect 7736 3106 7737 3158
rect 7557 3080 7558 3093
rect 7558 3092 7609 3093
rect 7621 3092 7673 3093
rect 7685 3092 7736 3093
rect 7558 3080 7592 3092
rect 7592 3080 7609 3092
rect 7557 3041 7609 3080
rect 7621 3041 7673 3092
rect 7685 3080 7702 3092
rect 7702 3080 7736 3092
rect 7736 3080 7737 3093
rect 7685 3041 7737 3080
rect 7557 2976 7558 3028
rect 7558 2976 7609 3028
rect 7621 2976 7673 3028
rect 7685 2976 7736 3028
rect 7736 2976 7737 3028
rect 7557 2911 7558 2963
rect 7558 2911 7609 2963
rect 7621 2911 7673 2963
rect 7685 2911 7736 2963
rect 7736 2911 7737 2963
rect 7557 2846 7558 2898
rect 7558 2846 7609 2898
rect 7621 2846 7673 2898
rect 7685 2846 7736 2898
rect 7736 2846 7737 2898
rect 7557 2781 7558 2833
rect 7558 2781 7609 2833
rect 7621 2781 7673 2833
rect 7685 2781 7736 2833
rect 7736 2781 7737 2833
rect 7557 2716 7558 2768
rect 7558 2716 7609 2768
rect 7621 2716 7673 2768
rect 7685 2716 7736 2768
rect 7736 2716 7737 2768
rect 7557 2651 7558 2703
rect 7558 2651 7609 2703
rect 7621 2651 7673 2703
rect 7685 2651 7736 2703
rect 7736 2651 7737 2703
rect 7557 2586 7558 2638
rect 7558 2586 7609 2638
rect 7621 2586 7673 2638
rect 7685 2586 7736 2638
rect 7736 2586 7737 2638
rect 7557 2535 7609 2573
rect 7557 2521 7558 2535
rect 7558 2521 7592 2535
rect 7592 2521 7609 2535
rect 7621 2535 7673 2573
rect 7621 2521 7630 2535
rect 7630 2521 7664 2535
rect 7664 2521 7673 2535
rect 7685 2535 7737 2573
rect 7685 2521 7702 2535
rect 7702 2521 7736 2535
rect 7736 2521 7737 2535
rect 7557 2501 7558 2508
rect 7558 2501 7592 2508
rect 7592 2501 7609 2508
rect 7557 2456 7609 2501
rect 7621 2501 7630 2508
rect 7630 2501 7664 2508
rect 7664 2501 7673 2508
rect 7621 2461 7673 2501
rect 7621 2456 7630 2461
rect 7630 2456 7664 2461
rect 7664 2456 7673 2461
rect 7685 2501 7702 2508
rect 7702 2501 7736 2508
rect 7736 2501 7737 2508
rect 7685 2456 7737 2501
rect 7557 2391 7558 2443
rect 7558 2391 7609 2443
rect 7621 2391 7673 2443
rect 7685 2391 7736 2443
rect 7736 2391 7737 2443
rect 7557 2326 7558 2378
rect 7558 2326 7609 2378
rect 7621 2326 7673 2378
rect 7685 2326 7736 2378
rect 7736 2326 7737 2378
rect 7557 2261 7558 2313
rect 7558 2261 7609 2313
rect 7621 2261 7673 2313
rect 7685 2261 7736 2313
rect 7736 2261 7737 2313
rect 7557 2196 7558 2248
rect 7558 2196 7609 2248
rect 7621 2196 7673 2248
rect 7685 2196 7736 2248
rect 7736 2196 7737 2248
rect 7557 2131 7558 2183
rect 7558 2131 7609 2183
rect 7621 2131 7673 2183
rect 7685 2131 7736 2183
rect 7736 2131 7737 2183
rect 7557 2066 7558 2118
rect 7558 2066 7609 2118
rect 7621 2066 7673 2118
rect 7685 2066 7736 2118
rect 7736 2066 7737 2118
rect 7557 2001 7558 2053
rect 7558 2001 7609 2053
rect 7621 2001 7673 2053
rect 7685 2001 7736 2053
rect 7736 2001 7737 2053
rect 7557 1935 7558 1987
rect 7558 1935 7609 1987
rect 7621 1935 7673 1987
rect 7685 1935 7736 1987
rect 7736 1935 7737 1987
rect 7557 1869 7558 1921
rect 7558 1869 7609 1921
rect 7621 1869 7673 1921
rect 7685 1869 7736 1921
rect 7736 1869 7737 1921
rect 7557 1803 7558 1855
rect 7558 1803 7609 1855
rect 7621 1803 7673 1855
rect 7685 1803 7736 1855
rect 7736 1803 7737 1855
rect 7557 1737 7558 1789
rect 7558 1737 7609 1789
rect 7621 1737 7673 1789
rect 7685 1737 7736 1789
rect 7736 1737 7737 1789
rect 7557 1671 7558 1723
rect 7558 1671 7609 1723
rect 7621 1671 7673 1723
rect 7685 1671 7736 1723
rect 7736 1671 7737 1723
rect 7557 1605 7558 1657
rect 7558 1605 7609 1657
rect 7621 1605 7673 1657
rect 7685 1605 7736 1657
rect 7736 1605 7737 1657
rect 7557 1539 7558 1591
rect 7558 1539 7609 1591
rect 7621 1539 7673 1591
rect 7685 1539 7736 1591
rect 7736 1539 7737 1591
rect 7557 1479 7558 1525
rect 7558 1491 7609 1525
rect 7621 1491 7673 1525
rect 7685 1491 7736 1525
rect 7558 1479 7592 1491
rect 7592 1479 7609 1491
rect 7557 1473 7609 1479
rect 7621 1473 7673 1491
rect 7685 1479 7702 1491
rect 7702 1479 7736 1491
rect 7736 1479 7737 1525
rect 7685 1473 7737 1479
rect 8053 4062 8105 4068
rect 8053 4028 8054 4062
rect 8054 4028 8088 4062
rect 8088 4028 8105 4062
rect 8053 4016 8105 4028
rect 8117 4062 8169 4068
rect 8117 4028 8126 4062
rect 8126 4028 8160 4062
rect 8160 4028 8169 4062
rect 8117 4016 8169 4028
rect 8181 4062 8233 4068
rect 8181 4028 8198 4062
rect 8198 4028 8232 4062
rect 8232 4028 8233 4062
rect 8181 4016 8233 4028
rect 8053 3988 8105 4003
rect 8053 3954 8054 3988
rect 8054 3954 8088 3988
rect 8088 3954 8105 3988
rect 8053 3951 8105 3954
rect 8117 3988 8169 4003
rect 8117 3954 8126 3988
rect 8126 3954 8160 3988
rect 8160 3954 8169 3988
rect 8117 3951 8169 3954
rect 8181 3988 8233 4003
rect 8181 3954 8198 3988
rect 8198 3954 8232 3988
rect 8232 3954 8233 3988
rect 8181 3951 8233 3954
rect 8053 3914 8105 3938
rect 8053 3886 8054 3914
rect 8054 3886 8088 3914
rect 8088 3886 8105 3914
rect 8117 3914 8169 3938
rect 8117 3886 8126 3914
rect 8126 3886 8160 3914
rect 8160 3886 8169 3914
rect 8181 3914 8233 3938
rect 8181 3886 8198 3914
rect 8198 3886 8232 3914
rect 8232 3886 8233 3914
rect 8053 3840 8105 3873
rect 8053 3821 8054 3840
rect 8054 3821 8088 3840
rect 8088 3821 8105 3840
rect 8117 3840 8169 3873
rect 8117 3821 8126 3840
rect 8126 3821 8160 3840
rect 8160 3821 8169 3840
rect 8181 3840 8233 3873
rect 8181 3821 8198 3840
rect 8198 3821 8232 3840
rect 8232 3821 8233 3840
rect 8053 3806 8054 3808
rect 8054 3806 8088 3808
rect 8088 3806 8105 3808
rect 8053 3766 8105 3806
rect 8053 3756 8054 3766
rect 8054 3756 8088 3766
rect 8088 3756 8105 3766
rect 8117 3806 8126 3808
rect 8126 3806 8160 3808
rect 8160 3806 8169 3808
rect 8117 3766 8169 3806
rect 8117 3756 8126 3766
rect 8126 3756 8160 3766
rect 8160 3756 8169 3766
rect 8181 3806 8198 3808
rect 8198 3806 8232 3808
rect 8232 3806 8233 3808
rect 8181 3766 8233 3806
rect 8181 3756 8198 3766
rect 8198 3756 8232 3766
rect 8232 3756 8233 3766
rect 8053 3732 8054 3743
rect 8054 3732 8088 3743
rect 8088 3732 8105 3743
rect 8053 3692 8105 3732
rect 8053 3691 8054 3692
rect 8054 3691 8088 3692
rect 8088 3691 8105 3692
rect 8117 3732 8126 3743
rect 8126 3732 8160 3743
rect 8160 3732 8169 3743
rect 8117 3692 8169 3732
rect 8117 3691 8126 3692
rect 8126 3691 8160 3692
rect 8160 3691 8169 3692
rect 8181 3732 8198 3743
rect 8198 3732 8232 3743
rect 8232 3732 8233 3743
rect 8181 3692 8233 3732
rect 8181 3691 8198 3692
rect 8198 3691 8232 3692
rect 8232 3691 8233 3692
rect 8053 3658 8054 3678
rect 8054 3658 8088 3678
rect 8088 3658 8105 3678
rect 8053 3626 8105 3658
rect 8117 3658 8126 3678
rect 8126 3658 8160 3678
rect 8160 3658 8169 3678
rect 8117 3626 8169 3658
rect 8181 3658 8198 3678
rect 8198 3658 8232 3678
rect 8232 3658 8233 3678
rect 8181 3626 8233 3658
rect 8053 3584 8054 3613
rect 8054 3584 8088 3613
rect 8088 3584 8105 3613
rect 8053 3561 8105 3584
rect 8117 3584 8126 3613
rect 8126 3584 8160 3613
rect 8160 3584 8169 3613
rect 8117 3561 8169 3584
rect 8181 3584 8198 3613
rect 8198 3584 8232 3613
rect 8232 3584 8233 3613
rect 8181 3561 8233 3584
rect 8053 3544 8105 3548
rect 8053 3510 8054 3544
rect 8054 3510 8088 3544
rect 8088 3510 8105 3544
rect 8053 3496 8105 3510
rect 8117 3544 8169 3548
rect 8117 3510 8126 3544
rect 8126 3510 8160 3544
rect 8160 3510 8169 3544
rect 8117 3496 8169 3510
rect 8181 3544 8233 3548
rect 8181 3510 8198 3544
rect 8198 3510 8232 3544
rect 8232 3510 8233 3544
rect 8181 3496 8233 3510
rect 8053 3470 8105 3483
rect 8053 3436 8054 3470
rect 8054 3436 8088 3470
rect 8088 3436 8105 3470
rect 8053 3431 8105 3436
rect 8117 3470 8169 3483
rect 8117 3436 8126 3470
rect 8126 3436 8160 3470
rect 8160 3436 8169 3470
rect 8117 3431 8169 3436
rect 8181 3470 8233 3483
rect 8181 3436 8198 3470
rect 8198 3436 8232 3470
rect 8232 3436 8233 3470
rect 8181 3431 8233 3436
rect 8053 3396 8105 3418
rect 8053 3366 8054 3396
rect 8054 3366 8088 3396
rect 8088 3366 8105 3396
rect 8117 3396 8169 3418
rect 8117 3366 8126 3396
rect 8126 3366 8160 3396
rect 8160 3366 8169 3396
rect 8181 3396 8233 3418
rect 8181 3366 8198 3396
rect 8198 3366 8232 3396
rect 8232 3366 8233 3396
rect 8053 3322 8105 3353
rect 8053 3301 8054 3322
rect 8054 3301 8088 3322
rect 8088 3301 8105 3322
rect 8117 3322 8169 3353
rect 8117 3301 8126 3322
rect 8126 3301 8160 3322
rect 8160 3301 8169 3322
rect 8181 3322 8233 3353
rect 8181 3301 8198 3322
rect 8198 3301 8232 3322
rect 8232 3301 8233 3322
rect 8053 3248 8105 3288
rect 8053 3236 8054 3248
rect 8054 3236 8088 3248
rect 8088 3236 8105 3248
rect 8117 3248 8169 3288
rect 8117 3236 8126 3248
rect 8126 3236 8160 3248
rect 8160 3236 8169 3248
rect 8181 3248 8233 3288
rect 8181 3236 8198 3248
rect 8198 3236 8232 3248
rect 8232 3236 8233 3248
rect 8053 3214 8054 3223
rect 8054 3214 8088 3223
rect 8088 3214 8105 3223
rect 8053 3174 8105 3214
rect 8053 3171 8054 3174
rect 8054 3171 8088 3174
rect 8088 3171 8105 3174
rect 8117 3214 8126 3223
rect 8126 3214 8160 3223
rect 8160 3214 8169 3223
rect 8117 3174 8169 3214
rect 8117 3171 8126 3174
rect 8126 3171 8160 3174
rect 8160 3171 8169 3174
rect 8181 3214 8198 3223
rect 8198 3214 8232 3223
rect 8232 3214 8233 3223
rect 8181 3174 8233 3214
rect 8181 3171 8198 3174
rect 8198 3171 8232 3174
rect 8232 3171 8233 3174
rect 8053 3140 8054 3158
rect 8054 3140 8088 3158
rect 8088 3140 8105 3158
rect 8053 3106 8105 3140
rect 8117 3140 8126 3158
rect 8126 3140 8160 3158
rect 8160 3140 8169 3158
rect 8117 3106 8169 3140
rect 8181 3140 8198 3158
rect 8198 3140 8232 3158
rect 8232 3140 8233 3158
rect 8181 3106 8233 3140
rect 8053 3066 8054 3093
rect 8054 3066 8088 3093
rect 8088 3066 8105 3093
rect 8053 3041 8105 3066
rect 8117 3066 8126 3093
rect 8126 3066 8160 3093
rect 8160 3066 8169 3093
rect 8117 3041 8169 3066
rect 8181 3066 8198 3093
rect 8198 3066 8232 3093
rect 8232 3066 8233 3093
rect 8181 3041 8233 3066
rect 8053 3026 8105 3028
rect 8053 2992 8054 3026
rect 8054 2992 8088 3026
rect 8088 2992 8105 3026
rect 8053 2976 8105 2992
rect 8117 3026 8169 3028
rect 8117 2992 8126 3026
rect 8126 2992 8160 3026
rect 8160 2992 8169 3026
rect 8117 2976 8169 2992
rect 8181 3026 8233 3028
rect 8181 2992 8198 3026
rect 8198 2992 8232 3026
rect 8232 2992 8233 3026
rect 8181 2976 8233 2992
rect 8053 2952 8105 2963
rect 8053 2918 8054 2952
rect 8054 2918 8088 2952
rect 8088 2918 8105 2952
rect 8053 2911 8105 2918
rect 8117 2952 8169 2963
rect 8117 2918 8126 2952
rect 8126 2918 8160 2952
rect 8160 2918 8169 2952
rect 8117 2911 8169 2918
rect 8181 2952 8233 2963
rect 8181 2918 8198 2952
rect 8198 2918 8232 2952
rect 8232 2918 8233 2952
rect 8181 2911 8233 2918
rect 8053 2878 8105 2898
rect 8053 2846 8054 2878
rect 8054 2846 8088 2878
rect 8088 2846 8105 2878
rect 8117 2878 8169 2898
rect 8117 2846 8126 2878
rect 8126 2846 8160 2878
rect 8160 2846 8169 2878
rect 8181 2878 8233 2898
rect 8181 2846 8198 2878
rect 8198 2846 8232 2878
rect 8232 2846 8233 2878
rect 8053 2804 8105 2833
rect 8053 2781 8054 2804
rect 8054 2781 8088 2804
rect 8088 2781 8105 2804
rect 8117 2804 8169 2833
rect 8117 2781 8126 2804
rect 8126 2781 8160 2804
rect 8160 2781 8169 2804
rect 8181 2804 8233 2833
rect 8181 2781 8198 2804
rect 8198 2781 8232 2804
rect 8232 2781 8233 2804
rect 8053 2730 8105 2768
rect 8053 2716 8054 2730
rect 8054 2716 8088 2730
rect 8088 2716 8105 2730
rect 8117 2730 8169 2768
rect 8117 2716 8126 2730
rect 8126 2716 8160 2730
rect 8160 2716 8169 2730
rect 8181 2730 8233 2768
rect 8181 2716 8198 2730
rect 8198 2716 8232 2730
rect 8232 2716 8233 2730
rect 8053 2696 8054 2703
rect 8054 2696 8088 2703
rect 8088 2696 8105 2703
rect 8053 2656 8105 2696
rect 8053 2651 8054 2656
rect 8054 2651 8088 2656
rect 8088 2651 8105 2656
rect 8117 2696 8126 2703
rect 8126 2696 8160 2703
rect 8160 2696 8169 2703
rect 8117 2656 8169 2696
rect 8117 2651 8126 2656
rect 8126 2651 8160 2656
rect 8160 2651 8169 2656
rect 8181 2696 8198 2703
rect 8198 2696 8232 2703
rect 8232 2696 8233 2703
rect 8181 2656 8233 2696
rect 8181 2651 8198 2656
rect 8198 2651 8232 2656
rect 8232 2651 8233 2656
rect 8053 2622 8054 2638
rect 8054 2622 8088 2638
rect 8088 2622 8105 2638
rect 8053 2586 8105 2622
rect 8117 2622 8126 2638
rect 8126 2622 8160 2638
rect 8160 2622 8169 2638
rect 8117 2586 8169 2622
rect 8181 2622 8198 2638
rect 8198 2622 8232 2638
rect 8232 2622 8233 2638
rect 8181 2586 8233 2622
rect 8053 2548 8054 2573
rect 8054 2548 8088 2573
rect 8088 2548 8105 2573
rect 8053 2521 8105 2548
rect 8117 2548 8126 2573
rect 8126 2548 8160 2573
rect 8160 2548 8169 2573
rect 8117 2521 8169 2548
rect 8181 2548 8198 2573
rect 8198 2548 8232 2573
rect 8232 2548 8233 2573
rect 8181 2521 8233 2548
rect 8053 2474 8054 2508
rect 8054 2474 8088 2508
rect 8088 2474 8105 2508
rect 8053 2456 8105 2474
rect 8117 2474 8126 2508
rect 8126 2474 8160 2508
rect 8160 2474 8169 2508
rect 8117 2456 8169 2474
rect 8181 2474 8198 2508
rect 8198 2474 8232 2508
rect 8232 2474 8233 2508
rect 8181 2456 8233 2474
rect 8053 2434 8105 2443
rect 8053 2400 8054 2434
rect 8054 2400 8088 2434
rect 8088 2400 8105 2434
rect 8053 2391 8105 2400
rect 8117 2434 8169 2443
rect 8117 2400 8126 2434
rect 8126 2400 8160 2434
rect 8160 2400 8169 2434
rect 8117 2391 8169 2400
rect 8181 2434 8233 2443
rect 8181 2400 8198 2434
rect 8198 2400 8232 2434
rect 8232 2400 8233 2434
rect 8181 2391 8233 2400
rect 8053 2360 8105 2378
rect 8053 2326 8054 2360
rect 8054 2326 8088 2360
rect 8088 2326 8105 2360
rect 8117 2360 8169 2378
rect 8117 2326 8126 2360
rect 8126 2326 8160 2360
rect 8160 2326 8169 2360
rect 8181 2360 8233 2378
rect 8181 2326 8198 2360
rect 8198 2326 8232 2360
rect 8232 2326 8233 2360
rect 8053 2286 8105 2313
rect 8053 2261 8054 2286
rect 8054 2261 8088 2286
rect 8088 2261 8105 2286
rect 8117 2286 8169 2313
rect 8117 2261 8126 2286
rect 8126 2261 8160 2286
rect 8160 2261 8169 2286
rect 8181 2286 8233 2313
rect 8181 2261 8198 2286
rect 8198 2261 8232 2286
rect 8232 2261 8233 2286
rect 8053 2212 8105 2248
rect 8053 2196 8054 2212
rect 8054 2196 8088 2212
rect 8088 2196 8105 2212
rect 8117 2212 8169 2248
rect 8117 2196 8126 2212
rect 8126 2196 8160 2212
rect 8160 2196 8169 2212
rect 8181 2212 8233 2248
rect 8181 2196 8198 2212
rect 8198 2196 8232 2212
rect 8232 2196 8233 2212
rect 8053 2178 8054 2183
rect 8054 2178 8088 2183
rect 8088 2178 8105 2183
rect 8053 2138 8105 2178
rect 8053 2131 8054 2138
rect 8054 2131 8088 2138
rect 8088 2131 8105 2138
rect 8117 2178 8126 2183
rect 8126 2178 8160 2183
rect 8160 2178 8169 2183
rect 8117 2138 8169 2178
rect 8117 2131 8126 2138
rect 8126 2131 8160 2138
rect 8160 2131 8169 2138
rect 8181 2178 8198 2183
rect 8198 2178 8232 2183
rect 8232 2178 8233 2183
rect 8181 2138 8233 2178
rect 8181 2131 8198 2138
rect 8198 2131 8232 2138
rect 8232 2131 8233 2138
rect 8053 2104 8054 2118
rect 8054 2104 8088 2118
rect 8088 2104 8105 2118
rect 8053 2066 8105 2104
rect 8117 2104 8126 2118
rect 8126 2104 8160 2118
rect 8160 2104 8169 2118
rect 8117 2066 8169 2104
rect 8181 2104 8198 2118
rect 8198 2104 8232 2118
rect 8232 2104 8233 2118
rect 8181 2066 8233 2104
rect 8053 2030 8054 2053
rect 8054 2030 8088 2053
rect 8088 2030 8105 2053
rect 8053 2001 8105 2030
rect 8117 2030 8126 2053
rect 8126 2030 8160 2053
rect 8160 2030 8169 2053
rect 8117 2001 8169 2030
rect 8181 2030 8198 2053
rect 8198 2030 8232 2053
rect 8232 2030 8233 2053
rect 8181 2001 8233 2030
rect 8053 1956 8054 1987
rect 8054 1956 8088 1987
rect 8088 1956 8105 1987
rect 8053 1935 8105 1956
rect 8117 1956 8126 1987
rect 8126 1956 8160 1987
rect 8160 1956 8169 1987
rect 8117 1935 8169 1956
rect 8181 1956 8198 1987
rect 8198 1956 8232 1987
rect 8232 1956 8233 1987
rect 8181 1935 8233 1956
rect 8053 1916 8105 1921
rect 8053 1882 8054 1916
rect 8054 1882 8088 1916
rect 8088 1882 8105 1916
rect 8053 1869 8105 1882
rect 8117 1916 8169 1921
rect 8117 1882 8126 1916
rect 8126 1882 8160 1916
rect 8160 1882 8169 1916
rect 8117 1869 8169 1882
rect 8181 1916 8233 1921
rect 8181 1882 8198 1916
rect 8198 1882 8232 1916
rect 8232 1882 8233 1916
rect 8181 1869 8233 1882
rect 8053 1842 8105 1855
rect 8053 1808 8054 1842
rect 8054 1808 8088 1842
rect 8088 1808 8105 1842
rect 8053 1803 8105 1808
rect 8117 1842 8169 1855
rect 8117 1808 8126 1842
rect 8126 1808 8160 1842
rect 8160 1808 8169 1842
rect 8117 1803 8169 1808
rect 8181 1842 8233 1855
rect 8181 1808 8198 1842
rect 8198 1808 8232 1842
rect 8232 1808 8233 1842
rect 8181 1803 8233 1808
rect 8053 1768 8105 1789
rect 8053 1737 8054 1768
rect 8054 1737 8088 1768
rect 8088 1737 8105 1768
rect 8117 1768 8169 1789
rect 8117 1737 8126 1768
rect 8126 1737 8160 1768
rect 8160 1737 8169 1768
rect 8181 1768 8233 1789
rect 8181 1737 8198 1768
rect 8198 1737 8232 1768
rect 8232 1737 8233 1768
rect 8053 1694 8105 1723
rect 8053 1671 8054 1694
rect 8054 1671 8088 1694
rect 8088 1671 8105 1694
rect 8117 1694 8169 1723
rect 8117 1671 8126 1694
rect 8126 1671 8160 1694
rect 8160 1671 8169 1694
rect 8181 1694 8233 1723
rect 8181 1671 8198 1694
rect 8198 1671 8232 1694
rect 8232 1671 8233 1694
rect 8053 1620 8105 1657
rect 8053 1605 8054 1620
rect 8054 1605 8088 1620
rect 8088 1605 8105 1620
rect 8117 1620 8169 1657
rect 8117 1605 8126 1620
rect 8126 1605 8160 1620
rect 8160 1605 8169 1620
rect 8181 1620 8233 1657
rect 8181 1605 8198 1620
rect 8198 1605 8232 1620
rect 8232 1605 8233 1620
rect 8053 1586 8054 1591
rect 8054 1586 8088 1591
rect 8088 1586 8105 1591
rect 8053 1545 8105 1586
rect 8053 1539 8054 1545
rect 8054 1539 8088 1545
rect 8088 1539 8105 1545
rect 8117 1586 8126 1591
rect 8126 1586 8160 1591
rect 8160 1586 8169 1591
rect 8117 1545 8169 1586
rect 8117 1539 8126 1545
rect 8126 1539 8160 1545
rect 8160 1539 8169 1545
rect 8181 1586 8198 1591
rect 8198 1586 8232 1591
rect 8232 1586 8233 1591
rect 8181 1545 8233 1586
rect 8181 1539 8198 1545
rect 8198 1539 8232 1545
rect 8232 1539 8233 1545
rect 8053 1511 8054 1525
rect 8054 1511 8088 1525
rect 8088 1511 8105 1525
rect 8053 1473 8105 1511
rect 8117 1511 8126 1525
rect 8126 1511 8160 1525
rect 8160 1511 8169 1525
rect 8117 1473 8169 1511
rect 8181 1511 8198 1525
rect 8198 1511 8232 1525
rect 8232 1511 8233 1525
rect 8181 1473 8233 1511
rect 8549 4050 8601 4068
rect 8613 4062 8665 4068
rect 8613 4050 8622 4062
rect 8622 4050 8656 4062
rect 8656 4050 8665 4062
rect 8677 4050 8729 4068
rect 8549 4016 8550 4050
rect 8550 4016 8601 4050
rect 8613 4016 8665 4050
rect 8677 4016 8728 4050
rect 8728 4016 8729 4050
rect 8549 3951 8550 4003
rect 8550 3951 8601 4003
rect 8613 3951 8665 4003
rect 8677 3951 8728 4003
rect 8728 3951 8729 4003
rect 8549 3886 8550 3938
rect 8550 3886 8601 3938
rect 8613 3886 8665 3938
rect 8677 3886 8728 3938
rect 8728 3886 8729 3938
rect 8549 3821 8550 3873
rect 8550 3821 8601 3873
rect 8613 3821 8665 3873
rect 8677 3821 8728 3873
rect 8728 3821 8729 3873
rect 8549 3756 8550 3808
rect 8550 3756 8601 3808
rect 8613 3756 8665 3808
rect 8677 3756 8728 3808
rect 8728 3756 8729 3808
rect 8549 3691 8550 3743
rect 8550 3691 8601 3743
rect 8613 3691 8665 3743
rect 8677 3691 8728 3743
rect 8728 3691 8729 3743
rect 8549 3626 8550 3678
rect 8550 3626 8601 3678
rect 8613 3626 8665 3678
rect 8677 3626 8728 3678
rect 8728 3626 8729 3678
rect 8549 3561 8550 3613
rect 8550 3561 8601 3613
rect 8613 3561 8665 3613
rect 8677 3561 8728 3613
rect 8728 3561 8729 3613
rect 8549 3496 8550 3548
rect 8550 3496 8601 3548
rect 8613 3496 8665 3548
rect 8677 3496 8728 3548
rect 8728 3496 8729 3548
rect 8549 3431 8550 3483
rect 8550 3431 8601 3483
rect 8613 3431 8665 3483
rect 8677 3431 8728 3483
rect 8728 3431 8729 3483
rect 8549 3366 8550 3418
rect 8550 3366 8601 3418
rect 8613 3366 8665 3418
rect 8677 3366 8728 3418
rect 8728 3366 8729 3418
rect 8549 3301 8550 3353
rect 8550 3301 8601 3353
rect 8613 3301 8665 3353
rect 8677 3301 8728 3353
rect 8728 3301 8729 3353
rect 8549 3236 8550 3288
rect 8550 3236 8601 3288
rect 8613 3236 8665 3288
rect 8677 3236 8728 3288
rect 8728 3236 8729 3288
rect 8549 3171 8550 3223
rect 8550 3171 8601 3223
rect 8613 3171 8665 3223
rect 8677 3171 8728 3223
rect 8728 3171 8729 3223
rect 8549 3106 8550 3158
rect 8550 3106 8601 3158
rect 8613 3106 8665 3158
rect 8677 3106 8728 3158
rect 8728 3106 8729 3158
rect 8549 3080 8550 3093
rect 8550 3092 8601 3093
rect 8613 3092 8665 3093
rect 8677 3092 8728 3093
rect 8550 3080 8584 3092
rect 8584 3080 8601 3092
rect 8549 3041 8601 3080
rect 8613 3041 8665 3092
rect 8677 3080 8694 3092
rect 8694 3080 8728 3092
rect 8728 3080 8729 3093
rect 8677 3041 8729 3080
rect 8549 2976 8550 3028
rect 8550 2976 8601 3028
rect 8613 2976 8665 3028
rect 8677 2976 8728 3028
rect 8728 2976 8729 3028
rect 8549 2911 8550 2963
rect 8550 2911 8601 2963
rect 8613 2911 8665 2963
rect 8677 2911 8728 2963
rect 8728 2911 8729 2963
rect 8549 2846 8550 2898
rect 8550 2846 8601 2898
rect 8613 2846 8665 2898
rect 8677 2846 8728 2898
rect 8728 2846 8729 2898
rect 8549 2781 8550 2833
rect 8550 2781 8601 2833
rect 8613 2781 8665 2833
rect 8677 2781 8728 2833
rect 8728 2781 8729 2833
rect 8549 2716 8550 2768
rect 8550 2716 8601 2768
rect 8613 2716 8665 2768
rect 8677 2716 8728 2768
rect 8728 2716 8729 2768
rect 8549 2651 8550 2703
rect 8550 2651 8601 2703
rect 8613 2651 8665 2703
rect 8677 2651 8728 2703
rect 8728 2651 8729 2703
rect 8549 2586 8550 2638
rect 8550 2586 8601 2638
rect 8613 2586 8665 2638
rect 8677 2586 8728 2638
rect 8728 2586 8729 2638
rect 8549 2535 8601 2573
rect 8549 2521 8550 2535
rect 8550 2521 8584 2535
rect 8584 2521 8601 2535
rect 8613 2535 8665 2573
rect 8613 2521 8622 2535
rect 8622 2521 8656 2535
rect 8656 2521 8665 2535
rect 8677 2535 8729 2573
rect 8677 2521 8694 2535
rect 8694 2521 8728 2535
rect 8728 2521 8729 2535
rect 8549 2501 8550 2508
rect 8550 2501 8584 2508
rect 8584 2501 8601 2508
rect 8549 2456 8601 2501
rect 8613 2501 8622 2508
rect 8622 2501 8656 2508
rect 8656 2501 8665 2508
rect 8613 2461 8665 2501
rect 8613 2456 8622 2461
rect 8622 2456 8656 2461
rect 8656 2456 8665 2461
rect 8677 2501 8694 2508
rect 8694 2501 8728 2508
rect 8728 2501 8729 2508
rect 8677 2456 8729 2501
rect 8549 2391 8550 2443
rect 8550 2391 8601 2443
rect 8613 2391 8665 2443
rect 8677 2391 8728 2443
rect 8728 2391 8729 2443
rect 8549 2326 8550 2378
rect 8550 2326 8601 2378
rect 8613 2326 8665 2378
rect 8677 2326 8728 2378
rect 8728 2326 8729 2378
rect 8549 2261 8550 2313
rect 8550 2261 8601 2313
rect 8613 2261 8665 2313
rect 8677 2261 8728 2313
rect 8728 2261 8729 2313
rect 8549 2196 8550 2248
rect 8550 2196 8601 2248
rect 8613 2196 8665 2248
rect 8677 2196 8728 2248
rect 8728 2196 8729 2248
rect 8549 2131 8550 2183
rect 8550 2131 8601 2183
rect 8613 2131 8665 2183
rect 8677 2131 8728 2183
rect 8728 2131 8729 2183
rect 8549 2066 8550 2118
rect 8550 2066 8601 2118
rect 8613 2066 8665 2118
rect 8677 2066 8728 2118
rect 8728 2066 8729 2118
rect 8549 2001 8550 2053
rect 8550 2001 8601 2053
rect 8613 2001 8665 2053
rect 8677 2001 8728 2053
rect 8728 2001 8729 2053
rect 8549 1935 8550 1987
rect 8550 1935 8601 1987
rect 8613 1935 8665 1987
rect 8677 1935 8728 1987
rect 8728 1935 8729 1987
rect 8549 1869 8550 1921
rect 8550 1869 8601 1921
rect 8613 1869 8665 1921
rect 8677 1869 8728 1921
rect 8728 1869 8729 1921
rect 8549 1803 8550 1855
rect 8550 1803 8601 1855
rect 8613 1803 8665 1855
rect 8677 1803 8728 1855
rect 8728 1803 8729 1855
rect 8549 1737 8550 1789
rect 8550 1737 8601 1789
rect 8613 1737 8665 1789
rect 8677 1737 8728 1789
rect 8728 1737 8729 1789
rect 8549 1671 8550 1723
rect 8550 1671 8601 1723
rect 8613 1671 8665 1723
rect 8677 1671 8728 1723
rect 8728 1671 8729 1723
rect 8549 1605 8550 1657
rect 8550 1605 8601 1657
rect 8613 1605 8665 1657
rect 8677 1605 8728 1657
rect 8728 1605 8729 1657
rect 8549 1539 8550 1591
rect 8550 1539 8601 1591
rect 8613 1539 8665 1591
rect 8677 1539 8728 1591
rect 8728 1539 8729 1591
rect 8549 1479 8550 1525
rect 8550 1491 8601 1525
rect 8613 1491 8665 1525
rect 8677 1491 8728 1525
rect 8550 1479 8584 1491
rect 8584 1479 8601 1491
rect 8549 1473 8601 1479
rect 8613 1473 8665 1491
rect 8677 1479 8694 1491
rect 8694 1479 8728 1491
rect 8728 1479 8729 1525
rect 8677 1473 8729 1479
rect 9045 4062 9097 4068
rect 9045 4028 9046 4062
rect 9046 4028 9080 4062
rect 9080 4028 9097 4062
rect 9045 4016 9097 4028
rect 9109 4062 9161 4068
rect 9109 4028 9118 4062
rect 9118 4028 9152 4062
rect 9152 4028 9161 4062
rect 9109 4016 9161 4028
rect 9173 4062 9225 4068
rect 9173 4028 9190 4062
rect 9190 4028 9224 4062
rect 9224 4028 9225 4062
rect 9173 4016 9225 4028
rect 9045 3988 9097 4003
rect 9045 3954 9046 3988
rect 9046 3954 9080 3988
rect 9080 3954 9097 3988
rect 9045 3951 9097 3954
rect 9109 3988 9161 4003
rect 9109 3954 9118 3988
rect 9118 3954 9152 3988
rect 9152 3954 9161 3988
rect 9109 3951 9161 3954
rect 9173 3988 9225 4003
rect 9173 3954 9190 3988
rect 9190 3954 9224 3988
rect 9224 3954 9225 3988
rect 9173 3951 9225 3954
rect 9045 3914 9097 3938
rect 9045 3886 9046 3914
rect 9046 3886 9080 3914
rect 9080 3886 9097 3914
rect 9109 3914 9161 3938
rect 9109 3886 9118 3914
rect 9118 3886 9152 3914
rect 9152 3886 9161 3914
rect 9173 3914 9225 3938
rect 9173 3886 9190 3914
rect 9190 3886 9224 3914
rect 9224 3886 9225 3914
rect 9045 3840 9097 3873
rect 9045 3821 9046 3840
rect 9046 3821 9080 3840
rect 9080 3821 9097 3840
rect 9109 3840 9161 3873
rect 9109 3821 9118 3840
rect 9118 3821 9152 3840
rect 9152 3821 9161 3840
rect 9173 3840 9225 3873
rect 9173 3821 9190 3840
rect 9190 3821 9224 3840
rect 9224 3821 9225 3840
rect 9045 3806 9046 3808
rect 9046 3806 9080 3808
rect 9080 3806 9097 3808
rect 9045 3766 9097 3806
rect 9045 3756 9046 3766
rect 9046 3756 9080 3766
rect 9080 3756 9097 3766
rect 9109 3806 9118 3808
rect 9118 3806 9152 3808
rect 9152 3806 9161 3808
rect 9109 3766 9161 3806
rect 9109 3756 9118 3766
rect 9118 3756 9152 3766
rect 9152 3756 9161 3766
rect 9173 3806 9190 3808
rect 9190 3806 9224 3808
rect 9224 3806 9225 3808
rect 9173 3766 9225 3806
rect 9173 3756 9190 3766
rect 9190 3756 9224 3766
rect 9224 3756 9225 3766
rect 9045 3732 9046 3743
rect 9046 3732 9080 3743
rect 9080 3732 9097 3743
rect 9045 3692 9097 3732
rect 9045 3691 9046 3692
rect 9046 3691 9080 3692
rect 9080 3691 9097 3692
rect 9109 3732 9118 3743
rect 9118 3732 9152 3743
rect 9152 3732 9161 3743
rect 9109 3692 9161 3732
rect 9109 3691 9118 3692
rect 9118 3691 9152 3692
rect 9152 3691 9161 3692
rect 9173 3732 9190 3743
rect 9190 3732 9224 3743
rect 9224 3732 9225 3743
rect 9173 3692 9225 3732
rect 9173 3691 9190 3692
rect 9190 3691 9224 3692
rect 9224 3691 9225 3692
rect 9045 3658 9046 3678
rect 9046 3658 9080 3678
rect 9080 3658 9097 3678
rect 9045 3626 9097 3658
rect 9109 3658 9118 3678
rect 9118 3658 9152 3678
rect 9152 3658 9161 3678
rect 9109 3626 9161 3658
rect 9173 3658 9190 3678
rect 9190 3658 9224 3678
rect 9224 3658 9225 3678
rect 9173 3626 9225 3658
rect 9045 3584 9046 3613
rect 9046 3584 9080 3613
rect 9080 3584 9097 3613
rect 9045 3561 9097 3584
rect 9109 3584 9118 3613
rect 9118 3584 9152 3613
rect 9152 3584 9161 3613
rect 9109 3561 9161 3584
rect 9173 3584 9190 3613
rect 9190 3584 9224 3613
rect 9224 3584 9225 3613
rect 9173 3561 9225 3584
rect 9045 3544 9097 3548
rect 9045 3510 9046 3544
rect 9046 3510 9080 3544
rect 9080 3510 9097 3544
rect 9045 3496 9097 3510
rect 9109 3544 9161 3548
rect 9109 3510 9118 3544
rect 9118 3510 9152 3544
rect 9152 3510 9161 3544
rect 9109 3496 9161 3510
rect 9173 3544 9225 3548
rect 9173 3510 9190 3544
rect 9190 3510 9224 3544
rect 9224 3510 9225 3544
rect 9173 3496 9225 3510
rect 9045 3470 9097 3483
rect 9045 3436 9046 3470
rect 9046 3436 9080 3470
rect 9080 3436 9097 3470
rect 9045 3431 9097 3436
rect 9109 3470 9161 3483
rect 9109 3436 9118 3470
rect 9118 3436 9152 3470
rect 9152 3436 9161 3470
rect 9109 3431 9161 3436
rect 9173 3470 9225 3483
rect 9173 3436 9190 3470
rect 9190 3436 9224 3470
rect 9224 3436 9225 3470
rect 9173 3431 9225 3436
rect 9045 3396 9097 3418
rect 9045 3366 9046 3396
rect 9046 3366 9080 3396
rect 9080 3366 9097 3396
rect 9109 3396 9161 3418
rect 9109 3366 9118 3396
rect 9118 3366 9152 3396
rect 9152 3366 9161 3396
rect 9173 3396 9225 3418
rect 9173 3366 9190 3396
rect 9190 3366 9224 3396
rect 9224 3366 9225 3396
rect 9045 3322 9097 3353
rect 9045 3301 9046 3322
rect 9046 3301 9080 3322
rect 9080 3301 9097 3322
rect 9109 3322 9161 3353
rect 9109 3301 9118 3322
rect 9118 3301 9152 3322
rect 9152 3301 9161 3322
rect 9173 3322 9225 3353
rect 9173 3301 9190 3322
rect 9190 3301 9224 3322
rect 9224 3301 9225 3322
rect 9045 3248 9097 3288
rect 9045 3236 9046 3248
rect 9046 3236 9080 3248
rect 9080 3236 9097 3248
rect 9109 3248 9161 3288
rect 9109 3236 9118 3248
rect 9118 3236 9152 3248
rect 9152 3236 9161 3248
rect 9173 3248 9225 3288
rect 9173 3236 9190 3248
rect 9190 3236 9224 3248
rect 9224 3236 9225 3248
rect 9045 3214 9046 3223
rect 9046 3214 9080 3223
rect 9080 3214 9097 3223
rect 9045 3174 9097 3214
rect 9045 3171 9046 3174
rect 9046 3171 9080 3174
rect 9080 3171 9097 3174
rect 9109 3214 9118 3223
rect 9118 3214 9152 3223
rect 9152 3214 9161 3223
rect 9109 3174 9161 3214
rect 9109 3171 9118 3174
rect 9118 3171 9152 3174
rect 9152 3171 9161 3174
rect 9173 3214 9190 3223
rect 9190 3214 9224 3223
rect 9224 3214 9225 3223
rect 9173 3174 9225 3214
rect 9173 3171 9190 3174
rect 9190 3171 9224 3174
rect 9224 3171 9225 3174
rect 9045 3140 9046 3158
rect 9046 3140 9080 3158
rect 9080 3140 9097 3158
rect 9045 3106 9097 3140
rect 9109 3140 9118 3158
rect 9118 3140 9152 3158
rect 9152 3140 9161 3158
rect 9109 3106 9161 3140
rect 9173 3140 9190 3158
rect 9190 3140 9224 3158
rect 9224 3140 9225 3158
rect 9173 3106 9225 3140
rect 9045 3066 9046 3093
rect 9046 3066 9080 3093
rect 9080 3066 9097 3093
rect 9045 3041 9097 3066
rect 9109 3066 9118 3093
rect 9118 3066 9152 3093
rect 9152 3066 9161 3093
rect 9109 3041 9161 3066
rect 9173 3066 9190 3093
rect 9190 3066 9224 3093
rect 9224 3066 9225 3093
rect 9173 3041 9225 3066
rect 9045 3026 9097 3028
rect 9045 2992 9046 3026
rect 9046 2992 9080 3026
rect 9080 2992 9097 3026
rect 9045 2976 9097 2992
rect 9109 3026 9161 3028
rect 9109 2992 9118 3026
rect 9118 2992 9152 3026
rect 9152 2992 9161 3026
rect 9109 2976 9161 2992
rect 9173 3026 9225 3028
rect 9173 2992 9190 3026
rect 9190 2992 9224 3026
rect 9224 2992 9225 3026
rect 9173 2976 9225 2992
rect 9045 2952 9097 2963
rect 9045 2918 9046 2952
rect 9046 2918 9080 2952
rect 9080 2918 9097 2952
rect 9045 2911 9097 2918
rect 9109 2952 9161 2963
rect 9109 2918 9118 2952
rect 9118 2918 9152 2952
rect 9152 2918 9161 2952
rect 9109 2911 9161 2918
rect 9173 2952 9225 2963
rect 9173 2918 9190 2952
rect 9190 2918 9224 2952
rect 9224 2918 9225 2952
rect 9173 2911 9225 2918
rect 9045 2878 9097 2898
rect 9045 2846 9046 2878
rect 9046 2846 9080 2878
rect 9080 2846 9097 2878
rect 9109 2878 9161 2898
rect 9109 2846 9118 2878
rect 9118 2846 9152 2878
rect 9152 2846 9161 2878
rect 9173 2878 9225 2898
rect 9173 2846 9190 2878
rect 9190 2846 9224 2878
rect 9224 2846 9225 2878
rect 9045 2804 9097 2833
rect 9045 2781 9046 2804
rect 9046 2781 9080 2804
rect 9080 2781 9097 2804
rect 9109 2804 9161 2833
rect 9109 2781 9118 2804
rect 9118 2781 9152 2804
rect 9152 2781 9161 2804
rect 9173 2804 9225 2833
rect 9173 2781 9190 2804
rect 9190 2781 9224 2804
rect 9224 2781 9225 2804
rect 9045 2730 9097 2768
rect 9045 2716 9046 2730
rect 9046 2716 9080 2730
rect 9080 2716 9097 2730
rect 9109 2730 9161 2768
rect 9109 2716 9118 2730
rect 9118 2716 9152 2730
rect 9152 2716 9161 2730
rect 9173 2730 9225 2768
rect 9173 2716 9190 2730
rect 9190 2716 9224 2730
rect 9224 2716 9225 2730
rect 9045 2696 9046 2703
rect 9046 2696 9080 2703
rect 9080 2696 9097 2703
rect 9045 2656 9097 2696
rect 9045 2651 9046 2656
rect 9046 2651 9080 2656
rect 9080 2651 9097 2656
rect 9109 2696 9118 2703
rect 9118 2696 9152 2703
rect 9152 2696 9161 2703
rect 9109 2656 9161 2696
rect 9109 2651 9118 2656
rect 9118 2651 9152 2656
rect 9152 2651 9161 2656
rect 9173 2696 9190 2703
rect 9190 2696 9224 2703
rect 9224 2696 9225 2703
rect 9173 2656 9225 2696
rect 9173 2651 9190 2656
rect 9190 2651 9224 2656
rect 9224 2651 9225 2656
rect 9045 2622 9046 2638
rect 9046 2622 9080 2638
rect 9080 2622 9097 2638
rect 9045 2586 9097 2622
rect 9109 2622 9118 2638
rect 9118 2622 9152 2638
rect 9152 2622 9161 2638
rect 9109 2586 9161 2622
rect 9173 2622 9190 2638
rect 9190 2622 9224 2638
rect 9224 2622 9225 2638
rect 9173 2586 9225 2622
rect 9045 2548 9046 2573
rect 9046 2548 9080 2573
rect 9080 2548 9097 2573
rect 9045 2521 9097 2548
rect 9109 2548 9118 2573
rect 9118 2548 9152 2573
rect 9152 2548 9161 2573
rect 9109 2521 9161 2548
rect 9173 2548 9190 2573
rect 9190 2548 9224 2573
rect 9224 2548 9225 2573
rect 9173 2521 9225 2548
rect 9045 2474 9046 2508
rect 9046 2474 9080 2508
rect 9080 2474 9097 2508
rect 9045 2456 9097 2474
rect 9109 2474 9118 2508
rect 9118 2474 9152 2508
rect 9152 2474 9161 2508
rect 9109 2456 9161 2474
rect 9173 2474 9190 2508
rect 9190 2474 9224 2508
rect 9224 2474 9225 2508
rect 9173 2456 9225 2474
rect 9045 2434 9097 2443
rect 9045 2400 9046 2434
rect 9046 2400 9080 2434
rect 9080 2400 9097 2434
rect 9045 2391 9097 2400
rect 9109 2434 9161 2443
rect 9109 2400 9118 2434
rect 9118 2400 9152 2434
rect 9152 2400 9161 2434
rect 9109 2391 9161 2400
rect 9173 2434 9225 2443
rect 9173 2400 9190 2434
rect 9190 2400 9224 2434
rect 9224 2400 9225 2434
rect 9173 2391 9225 2400
rect 9045 2360 9097 2378
rect 9045 2326 9046 2360
rect 9046 2326 9080 2360
rect 9080 2326 9097 2360
rect 9109 2360 9161 2378
rect 9109 2326 9118 2360
rect 9118 2326 9152 2360
rect 9152 2326 9161 2360
rect 9173 2360 9225 2378
rect 9173 2326 9190 2360
rect 9190 2326 9224 2360
rect 9224 2326 9225 2360
rect 9045 2286 9097 2313
rect 9045 2261 9046 2286
rect 9046 2261 9080 2286
rect 9080 2261 9097 2286
rect 9109 2286 9161 2313
rect 9109 2261 9118 2286
rect 9118 2261 9152 2286
rect 9152 2261 9161 2286
rect 9173 2286 9225 2313
rect 9173 2261 9190 2286
rect 9190 2261 9224 2286
rect 9224 2261 9225 2286
rect 9045 2212 9097 2248
rect 9045 2196 9046 2212
rect 9046 2196 9080 2212
rect 9080 2196 9097 2212
rect 9109 2212 9161 2248
rect 9109 2196 9118 2212
rect 9118 2196 9152 2212
rect 9152 2196 9161 2212
rect 9173 2212 9225 2248
rect 9173 2196 9190 2212
rect 9190 2196 9224 2212
rect 9224 2196 9225 2212
rect 9045 2178 9046 2183
rect 9046 2178 9080 2183
rect 9080 2178 9097 2183
rect 9045 2138 9097 2178
rect 9045 2131 9046 2138
rect 9046 2131 9080 2138
rect 9080 2131 9097 2138
rect 9109 2178 9118 2183
rect 9118 2178 9152 2183
rect 9152 2178 9161 2183
rect 9109 2138 9161 2178
rect 9109 2131 9118 2138
rect 9118 2131 9152 2138
rect 9152 2131 9161 2138
rect 9173 2178 9190 2183
rect 9190 2178 9224 2183
rect 9224 2178 9225 2183
rect 9173 2138 9225 2178
rect 9173 2131 9190 2138
rect 9190 2131 9224 2138
rect 9224 2131 9225 2138
rect 9045 2104 9046 2118
rect 9046 2104 9080 2118
rect 9080 2104 9097 2118
rect 9045 2066 9097 2104
rect 9109 2104 9118 2118
rect 9118 2104 9152 2118
rect 9152 2104 9161 2118
rect 9109 2066 9161 2104
rect 9173 2104 9190 2118
rect 9190 2104 9224 2118
rect 9224 2104 9225 2118
rect 9173 2066 9225 2104
rect 9045 2030 9046 2053
rect 9046 2030 9080 2053
rect 9080 2030 9097 2053
rect 9045 2001 9097 2030
rect 9109 2030 9118 2053
rect 9118 2030 9152 2053
rect 9152 2030 9161 2053
rect 9109 2001 9161 2030
rect 9173 2030 9190 2053
rect 9190 2030 9224 2053
rect 9224 2030 9225 2053
rect 9173 2001 9225 2030
rect 9045 1956 9046 1987
rect 9046 1956 9080 1987
rect 9080 1956 9097 1987
rect 9045 1935 9097 1956
rect 9109 1956 9118 1987
rect 9118 1956 9152 1987
rect 9152 1956 9161 1987
rect 9109 1935 9161 1956
rect 9173 1956 9190 1987
rect 9190 1956 9224 1987
rect 9224 1956 9225 1987
rect 9173 1935 9225 1956
rect 9045 1916 9097 1921
rect 9045 1882 9046 1916
rect 9046 1882 9080 1916
rect 9080 1882 9097 1916
rect 9045 1869 9097 1882
rect 9109 1916 9161 1921
rect 9109 1882 9118 1916
rect 9118 1882 9152 1916
rect 9152 1882 9161 1916
rect 9109 1869 9161 1882
rect 9173 1916 9225 1921
rect 9173 1882 9190 1916
rect 9190 1882 9224 1916
rect 9224 1882 9225 1916
rect 9173 1869 9225 1882
rect 9045 1842 9097 1855
rect 9045 1808 9046 1842
rect 9046 1808 9080 1842
rect 9080 1808 9097 1842
rect 9045 1803 9097 1808
rect 9109 1842 9161 1855
rect 9109 1808 9118 1842
rect 9118 1808 9152 1842
rect 9152 1808 9161 1842
rect 9109 1803 9161 1808
rect 9173 1842 9225 1855
rect 9173 1808 9190 1842
rect 9190 1808 9224 1842
rect 9224 1808 9225 1842
rect 9173 1803 9225 1808
rect 9045 1768 9097 1789
rect 9045 1737 9046 1768
rect 9046 1737 9080 1768
rect 9080 1737 9097 1768
rect 9109 1768 9161 1789
rect 9109 1737 9118 1768
rect 9118 1737 9152 1768
rect 9152 1737 9161 1768
rect 9173 1768 9225 1789
rect 9173 1737 9190 1768
rect 9190 1737 9224 1768
rect 9224 1737 9225 1768
rect 9045 1694 9097 1723
rect 9045 1671 9046 1694
rect 9046 1671 9080 1694
rect 9080 1671 9097 1694
rect 9109 1694 9161 1723
rect 9109 1671 9118 1694
rect 9118 1671 9152 1694
rect 9152 1671 9161 1694
rect 9173 1694 9225 1723
rect 9173 1671 9190 1694
rect 9190 1671 9224 1694
rect 9224 1671 9225 1694
rect 9045 1620 9097 1657
rect 9045 1605 9046 1620
rect 9046 1605 9080 1620
rect 9080 1605 9097 1620
rect 9109 1620 9161 1657
rect 9109 1605 9118 1620
rect 9118 1605 9152 1620
rect 9152 1605 9161 1620
rect 9173 1620 9225 1657
rect 9173 1605 9190 1620
rect 9190 1605 9224 1620
rect 9224 1605 9225 1620
rect 9045 1586 9046 1591
rect 9046 1586 9080 1591
rect 9080 1586 9097 1591
rect 9045 1545 9097 1586
rect 9045 1539 9046 1545
rect 9046 1539 9080 1545
rect 9080 1539 9097 1545
rect 9109 1586 9118 1591
rect 9118 1586 9152 1591
rect 9152 1586 9161 1591
rect 9109 1545 9161 1586
rect 9109 1539 9118 1545
rect 9118 1539 9152 1545
rect 9152 1539 9161 1545
rect 9173 1586 9190 1591
rect 9190 1586 9224 1591
rect 9224 1586 9225 1591
rect 9173 1545 9225 1586
rect 9173 1539 9190 1545
rect 9190 1539 9224 1545
rect 9224 1539 9225 1545
rect 9045 1511 9046 1525
rect 9046 1511 9080 1525
rect 9080 1511 9097 1525
rect 9045 1473 9097 1511
rect 9109 1511 9118 1525
rect 9118 1511 9152 1525
rect 9152 1511 9161 1525
rect 9109 1473 9161 1511
rect 9173 1511 9190 1525
rect 9190 1511 9224 1525
rect 9224 1511 9225 1525
rect 9173 1473 9225 1511
rect 9541 4050 9593 4068
rect 9605 4062 9657 4068
rect 9605 4050 9614 4062
rect 9614 4050 9648 4062
rect 9648 4050 9657 4062
rect 9669 4050 9721 4068
rect 9541 4016 9542 4050
rect 9542 4016 9593 4050
rect 9605 4016 9657 4050
rect 9669 4016 9720 4050
rect 9720 4016 9721 4050
rect 9541 3951 9542 4003
rect 9542 3951 9593 4003
rect 9605 3951 9657 4003
rect 9669 3951 9720 4003
rect 9720 3951 9721 4003
rect 9541 3886 9542 3938
rect 9542 3886 9593 3938
rect 9605 3886 9657 3938
rect 9669 3886 9720 3938
rect 9720 3886 9721 3938
rect 9541 3821 9542 3873
rect 9542 3821 9593 3873
rect 9605 3821 9657 3873
rect 9669 3821 9720 3873
rect 9720 3821 9721 3873
rect 9541 3756 9542 3808
rect 9542 3756 9593 3808
rect 9605 3756 9657 3808
rect 9669 3756 9720 3808
rect 9720 3756 9721 3808
rect 9541 3691 9542 3743
rect 9542 3691 9593 3743
rect 9605 3691 9657 3743
rect 9669 3691 9720 3743
rect 9720 3691 9721 3743
rect 9541 3626 9542 3678
rect 9542 3626 9593 3678
rect 9605 3626 9657 3678
rect 9669 3626 9720 3678
rect 9720 3626 9721 3678
rect 9541 3561 9542 3613
rect 9542 3561 9593 3613
rect 9605 3561 9657 3613
rect 9669 3561 9720 3613
rect 9720 3561 9721 3613
rect 9541 3496 9542 3548
rect 9542 3496 9593 3548
rect 9605 3496 9657 3548
rect 9669 3496 9720 3548
rect 9720 3496 9721 3548
rect 9541 3431 9542 3483
rect 9542 3431 9593 3483
rect 9605 3431 9657 3483
rect 9669 3431 9720 3483
rect 9720 3431 9721 3483
rect 9541 3366 9542 3418
rect 9542 3366 9593 3418
rect 9605 3366 9657 3418
rect 9669 3366 9720 3418
rect 9720 3366 9721 3418
rect 9541 3301 9542 3353
rect 9542 3301 9593 3353
rect 9605 3301 9657 3353
rect 9669 3301 9720 3353
rect 9720 3301 9721 3353
rect 9541 3236 9542 3288
rect 9542 3236 9593 3288
rect 9605 3236 9657 3288
rect 9669 3236 9720 3288
rect 9720 3236 9721 3288
rect 9541 3171 9542 3223
rect 9542 3171 9593 3223
rect 9605 3171 9657 3223
rect 9669 3171 9720 3223
rect 9720 3171 9721 3223
rect 9541 3106 9542 3158
rect 9542 3106 9593 3158
rect 9605 3106 9657 3158
rect 9669 3106 9720 3158
rect 9720 3106 9721 3158
rect 9541 3080 9542 3093
rect 9542 3092 9593 3093
rect 9605 3092 9657 3093
rect 9669 3092 9720 3093
rect 9542 3080 9576 3092
rect 9576 3080 9593 3092
rect 9541 3041 9593 3080
rect 9605 3041 9657 3092
rect 9669 3080 9686 3092
rect 9686 3080 9720 3092
rect 9720 3080 9721 3093
rect 9669 3041 9721 3080
rect 9541 2976 9542 3028
rect 9542 2976 9593 3028
rect 9605 2976 9657 3028
rect 9669 2976 9720 3028
rect 9720 2976 9721 3028
rect 9541 2911 9542 2963
rect 9542 2911 9593 2963
rect 9605 2911 9657 2963
rect 9669 2911 9720 2963
rect 9720 2911 9721 2963
rect 9541 2846 9542 2898
rect 9542 2846 9593 2898
rect 9605 2846 9657 2898
rect 9669 2846 9720 2898
rect 9720 2846 9721 2898
rect 9541 2781 9542 2833
rect 9542 2781 9593 2833
rect 9605 2781 9657 2833
rect 9669 2781 9720 2833
rect 9720 2781 9721 2833
rect 9541 2716 9542 2768
rect 9542 2716 9593 2768
rect 9605 2716 9657 2768
rect 9669 2716 9720 2768
rect 9720 2716 9721 2768
rect 9541 2651 9542 2703
rect 9542 2651 9593 2703
rect 9605 2651 9657 2703
rect 9669 2651 9720 2703
rect 9720 2651 9721 2703
rect 9541 2586 9542 2638
rect 9542 2586 9593 2638
rect 9605 2586 9657 2638
rect 9669 2586 9720 2638
rect 9720 2586 9721 2638
rect 9541 2535 9593 2573
rect 9541 2521 9542 2535
rect 9542 2521 9576 2535
rect 9576 2521 9593 2535
rect 9605 2535 9657 2573
rect 9605 2521 9614 2535
rect 9614 2521 9648 2535
rect 9648 2521 9657 2535
rect 9669 2535 9721 2573
rect 9669 2521 9686 2535
rect 9686 2521 9720 2535
rect 9720 2521 9721 2535
rect 9541 2501 9542 2508
rect 9542 2501 9576 2508
rect 9576 2501 9593 2508
rect 9541 2456 9593 2501
rect 9605 2501 9614 2508
rect 9614 2501 9648 2508
rect 9648 2501 9657 2508
rect 9605 2461 9657 2501
rect 9605 2456 9614 2461
rect 9614 2456 9648 2461
rect 9648 2456 9657 2461
rect 9669 2501 9686 2508
rect 9686 2501 9720 2508
rect 9720 2501 9721 2508
rect 9669 2456 9721 2501
rect 9541 2391 9542 2443
rect 9542 2391 9593 2443
rect 9605 2391 9657 2443
rect 9669 2391 9720 2443
rect 9720 2391 9721 2443
rect 9541 2326 9542 2378
rect 9542 2326 9593 2378
rect 9605 2326 9657 2378
rect 9669 2326 9720 2378
rect 9720 2326 9721 2378
rect 9541 2261 9542 2313
rect 9542 2261 9593 2313
rect 9605 2261 9657 2313
rect 9669 2261 9720 2313
rect 9720 2261 9721 2313
rect 9541 2196 9542 2248
rect 9542 2196 9593 2248
rect 9605 2196 9657 2248
rect 9669 2196 9720 2248
rect 9720 2196 9721 2248
rect 9541 2131 9542 2183
rect 9542 2131 9593 2183
rect 9605 2131 9657 2183
rect 9669 2131 9720 2183
rect 9720 2131 9721 2183
rect 9541 2066 9542 2118
rect 9542 2066 9593 2118
rect 9605 2066 9657 2118
rect 9669 2066 9720 2118
rect 9720 2066 9721 2118
rect 9541 2001 9542 2053
rect 9542 2001 9593 2053
rect 9605 2001 9657 2053
rect 9669 2001 9720 2053
rect 9720 2001 9721 2053
rect 9541 1935 9542 1987
rect 9542 1935 9593 1987
rect 9605 1935 9657 1987
rect 9669 1935 9720 1987
rect 9720 1935 9721 1987
rect 9541 1869 9542 1921
rect 9542 1869 9593 1921
rect 9605 1869 9657 1921
rect 9669 1869 9720 1921
rect 9720 1869 9721 1921
rect 9541 1803 9542 1855
rect 9542 1803 9593 1855
rect 9605 1803 9657 1855
rect 9669 1803 9720 1855
rect 9720 1803 9721 1855
rect 9541 1737 9542 1789
rect 9542 1737 9593 1789
rect 9605 1737 9657 1789
rect 9669 1737 9720 1789
rect 9720 1737 9721 1789
rect 9541 1671 9542 1723
rect 9542 1671 9593 1723
rect 9605 1671 9657 1723
rect 9669 1671 9720 1723
rect 9720 1671 9721 1723
rect 9541 1605 9542 1657
rect 9542 1605 9593 1657
rect 9605 1605 9657 1657
rect 9669 1605 9720 1657
rect 9720 1605 9721 1657
rect 9541 1539 9542 1591
rect 9542 1539 9593 1591
rect 9605 1539 9657 1591
rect 9669 1539 9720 1591
rect 9720 1539 9721 1591
rect 9541 1479 9542 1525
rect 9542 1491 9593 1525
rect 9605 1491 9657 1525
rect 9669 1491 9720 1525
rect 9542 1479 9576 1491
rect 9576 1479 9593 1491
rect 9541 1473 9593 1479
rect 9605 1473 9657 1491
rect 9669 1479 9686 1491
rect 9686 1479 9720 1491
rect 9720 1479 9721 1525
rect 9669 1473 9721 1479
rect 10037 4062 10089 4068
rect 10037 4028 10038 4062
rect 10038 4028 10072 4062
rect 10072 4028 10089 4062
rect 10037 4016 10089 4028
rect 10101 4062 10153 4068
rect 10101 4028 10110 4062
rect 10110 4028 10144 4062
rect 10144 4028 10153 4062
rect 10101 4016 10153 4028
rect 10165 4062 10217 4068
rect 10165 4028 10182 4062
rect 10182 4028 10216 4062
rect 10216 4028 10217 4062
rect 10165 4016 10217 4028
rect 10037 3988 10089 4003
rect 10037 3954 10038 3988
rect 10038 3954 10072 3988
rect 10072 3954 10089 3988
rect 10037 3951 10089 3954
rect 10101 3988 10153 4003
rect 10101 3954 10110 3988
rect 10110 3954 10144 3988
rect 10144 3954 10153 3988
rect 10101 3951 10153 3954
rect 10165 3988 10217 4003
rect 10165 3954 10182 3988
rect 10182 3954 10216 3988
rect 10216 3954 10217 3988
rect 10165 3951 10217 3954
rect 10037 3914 10089 3938
rect 10037 3886 10038 3914
rect 10038 3886 10072 3914
rect 10072 3886 10089 3914
rect 10101 3914 10153 3938
rect 10101 3886 10110 3914
rect 10110 3886 10144 3914
rect 10144 3886 10153 3914
rect 10165 3914 10217 3938
rect 10165 3886 10182 3914
rect 10182 3886 10216 3914
rect 10216 3886 10217 3914
rect 10037 3840 10089 3873
rect 10037 3821 10038 3840
rect 10038 3821 10072 3840
rect 10072 3821 10089 3840
rect 10101 3840 10153 3873
rect 10101 3821 10110 3840
rect 10110 3821 10144 3840
rect 10144 3821 10153 3840
rect 10165 3840 10217 3873
rect 10165 3821 10182 3840
rect 10182 3821 10216 3840
rect 10216 3821 10217 3840
rect 10037 3806 10038 3808
rect 10038 3806 10072 3808
rect 10072 3806 10089 3808
rect 10037 3766 10089 3806
rect 10037 3756 10038 3766
rect 10038 3756 10072 3766
rect 10072 3756 10089 3766
rect 10101 3806 10110 3808
rect 10110 3806 10144 3808
rect 10144 3806 10153 3808
rect 10101 3766 10153 3806
rect 10101 3756 10110 3766
rect 10110 3756 10144 3766
rect 10144 3756 10153 3766
rect 10165 3806 10182 3808
rect 10182 3806 10216 3808
rect 10216 3806 10217 3808
rect 10165 3766 10217 3806
rect 10165 3756 10182 3766
rect 10182 3756 10216 3766
rect 10216 3756 10217 3766
rect 10037 3732 10038 3743
rect 10038 3732 10072 3743
rect 10072 3732 10089 3743
rect 10037 3692 10089 3732
rect 10037 3691 10038 3692
rect 10038 3691 10072 3692
rect 10072 3691 10089 3692
rect 10101 3732 10110 3743
rect 10110 3732 10144 3743
rect 10144 3732 10153 3743
rect 10101 3692 10153 3732
rect 10101 3691 10110 3692
rect 10110 3691 10144 3692
rect 10144 3691 10153 3692
rect 10165 3732 10182 3743
rect 10182 3732 10216 3743
rect 10216 3732 10217 3743
rect 10165 3692 10217 3732
rect 10165 3691 10182 3692
rect 10182 3691 10216 3692
rect 10216 3691 10217 3692
rect 10037 3658 10038 3678
rect 10038 3658 10072 3678
rect 10072 3658 10089 3678
rect 10037 3626 10089 3658
rect 10101 3658 10110 3678
rect 10110 3658 10144 3678
rect 10144 3658 10153 3678
rect 10101 3626 10153 3658
rect 10165 3658 10182 3678
rect 10182 3658 10216 3678
rect 10216 3658 10217 3678
rect 10165 3626 10217 3658
rect 10037 3584 10038 3613
rect 10038 3584 10072 3613
rect 10072 3584 10089 3613
rect 10037 3561 10089 3584
rect 10101 3584 10110 3613
rect 10110 3584 10144 3613
rect 10144 3584 10153 3613
rect 10101 3561 10153 3584
rect 10165 3584 10182 3613
rect 10182 3584 10216 3613
rect 10216 3584 10217 3613
rect 10165 3561 10217 3584
rect 10037 3544 10089 3548
rect 10037 3510 10038 3544
rect 10038 3510 10072 3544
rect 10072 3510 10089 3544
rect 10037 3496 10089 3510
rect 10101 3544 10153 3548
rect 10101 3510 10110 3544
rect 10110 3510 10144 3544
rect 10144 3510 10153 3544
rect 10101 3496 10153 3510
rect 10165 3544 10217 3548
rect 10165 3510 10182 3544
rect 10182 3510 10216 3544
rect 10216 3510 10217 3544
rect 10165 3496 10217 3510
rect 10037 3470 10089 3483
rect 10037 3436 10038 3470
rect 10038 3436 10072 3470
rect 10072 3436 10089 3470
rect 10037 3431 10089 3436
rect 10101 3470 10153 3483
rect 10101 3436 10110 3470
rect 10110 3436 10144 3470
rect 10144 3436 10153 3470
rect 10101 3431 10153 3436
rect 10165 3470 10217 3483
rect 10165 3436 10182 3470
rect 10182 3436 10216 3470
rect 10216 3436 10217 3470
rect 10165 3431 10217 3436
rect 10037 3396 10089 3418
rect 10037 3366 10038 3396
rect 10038 3366 10072 3396
rect 10072 3366 10089 3396
rect 10101 3396 10153 3418
rect 10101 3366 10110 3396
rect 10110 3366 10144 3396
rect 10144 3366 10153 3396
rect 10165 3396 10217 3418
rect 10165 3366 10182 3396
rect 10182 3366 10216 3396
rect 10216 3366 10217 3396
rect 10037 3322 10089 3353
rect 10037 3301 10038 3322
rect 10038 3301 10072 3322
rect 10072 3301 10089 3322
rect 10101 3322 10153 3353
rect 10101 3301 10110 3322
rect 10110 3301 10144 3322
rect 10144 3301 10153 3322
rect 10165 3322 10217 3353
rect 10165 3301 10182 3322
rect 10182 3301 10216 3322
rect 10216 3301 10217 3322
rect 10037 3248 10089 3288
rect 10037 3236 10038 3248
rect 10038 3236 10072 3248
rect 10072 3236 10089 3248
rect 10101 3248 10153 3288
rect 10101 3236 10110 3248
rect 10110 3236 10144 3248
rect 10144 3236 10153 3248
rect 10165 3248 10217 3288
rect 10165 3236 10182 3248
rect 10182 3236 10216 3248
rect 10216 3236 10217 3248
rect 10037 3214 10038 3223
rect 10038 3214 10072 3223
rect 10072 3214 10089 3223
rect 10037 3174 10089 3214
rect 10037 3171 10038 3174
rect 10038 3171 10072 3174
rect 10072 3171 10089 3174
rect 10101 3214 10110 3223
rect 10110 3214 10144 3223
rect 10144 3214 10153 3223
rect 10101 3174 10153 3214
rect 10101 3171 10110 3174
rect 10110 3171 10144 3174
rect 10144 3171 10153 3174
rect 10165 3214 10182 3223
rect 10182 3214 10216 3223
rect 10216 3214 10217 3223
rect 10165 3174 10217 3214
rect 10165 3171 10182 3174
rect 10182 3171 10216 3174
rect 10216 3171 10217 3174
rect 10037 3140 10038 3158
rect 10038 3140 10072 3158
rect 10072 3140 10089 3158
rect 10037 3106 10089 3140
rect 10101 3140 10110 3158
rect 10110 3140 10144 3158
rect 10144 3140 10153 3158
rect 10101 3106 10153 3140
rect 10165 3140 10182 3158
rect 10182 3140 10216 3158
rect 10216 3140 10217 3158
rect 10165 3106 10217 3140
rect 10037 3066 10038 3093
rect 10038 3066 10072 3093
rect 10072 3066 10089 3093
rect 10037 3041 10089 3066
rect 10101 3066 10110 3093
rect 10110 3066 10144 3093
rect 10144 3066 10153 3093
rect 10101 3041 10153 3066
rect 10165 3066 10182 3093
rect 10182 3066 10216 3093
rect 10216 3066 10217 3093
rect 10165 3041 10217 3066
rect 10037 3026 10089 3028
rect 10037 2992 10038 3026
rect 10038 2992 10072 3026
rect 10072 2992 10089 3026
rect 10037 2976 10089 2992
rect 10101 3026 10153 3028
rect 10101 2992 10110 3026
rect 10110 2992 10144 3026
rect 10144 2992 10153 3026
rect 10101 2976 10153 2992
rect 10165 3026 10217 3028
rect 10165 2992 10182 3026
rect 10182 2992 10216 3026
rect 10216 2992 10217 3026
rect 10165 2976 10217 2992
rect 10037 2952 10089 2963
rect 10037 2918 10038 2952
rect 10038 2918 10072 2952
rect 10072 2918 10089 2952
rect 10037 2911 10089 2918
rect 10101 2952 10153 2963
rect 10101 2918 10110 2952
rect 10110 2918 10144 2952
rect 10144 2918 10153 2952
rect 10101 2911 10153 2918
rect 10165 2952 10217 2963
rect 10165 2918 10182 2952
rect 10182 2918 10216 2952
rect 10216 2918 10217 2952
rect 10165 2911 10217 2918
rect 10037 2878 10089 2898
rect 10037 2846 10038 2878
rect 10038 2846 10072 2878
rect 10072 2846 10089 2878
rect 10101 2878 10153 2898
rect 10101 2846 10110 2878
rect 10110 2846 10144 2878
rect 10144 2846 10153 2878
rect 10165 2878 10217 2898
rect 10165 2846 10182 2878
rect 10182 2846 10216 2878
rect 10216 2846 10217 2878
rect 10037 2804 10089 2833
rect 10037 2781 10038 2804
rect 10038 2781 10072 2804
rect 10072 2781 10089 2804
rect 10101 2804 10153 2833
rect 10101 2781 10110 2804
rect 10110 2781 10144 2804
rect 10144 2781 10153 2804
rect 10165 2804 10217 2833
rect 10165 2781 10182 2804
rect 10182 2781 10216 2804
rect 10216 2781 10217 2804
rect 10037 2730 10089 2768
rect 10037 2716 10038 2730
rect 10038 2716 10072 2730
rect 10072 2716 10089 2730
rect 10101 2730 10153 2768
rect 10101 2716 10110 2730
rect 10110 2716 10144 2730
rect 10144 2716 10153 2730
rect 10165 2730 10217 2768
rect 10165 2716 10182 2730
rect 10182 2716 10216 2730
rect 10216 2716 10217 2730
rect 10037 2696 10038 2703
rect 10038 2696 10072 2703
rect 10072 2696 10089 2703
rect 10037 2656 10089 2696
rect 10037 2651 10038 2656
rect 10038 2651 10072 2656
rect 10072 2651 10089 2656
rect 10101 2696 10110 2703
rect 10110 2696 10144 2703
rect 10144 2696 10153 2703
rect 10101 2656 10153 2696
rect 10101 2651 10110 2656
rect 10110 2651 10144 2656
rect 10144 2651 10153 2656
rect 10165 2696 10182 2703
rect 10182 2696 10216 2703
rect 10216 2696 10217 2703
rect 10165 2656 10217 2696
rect 10165 2651 10182 2656
rect 10182 2651 10216 2656
rect 10216 2651 10217 2656
rect 10037 2622 10038 2638
rect 10038 2622 10072 2638
rect 10072 2622 10089 2638
rect 10037 2586 10089 2622
rect 10101 2622 10110 2638
rect 10110 2622 10144 2638
rect 10144 2622 10153 2638
rect 10101 2586 10153 2622
rect 10165 2622 10182 2638
rect 10182 2622 10216 2638
rect 10216 2622 10217 2638
rect 10165 2586 10217 2622
rect 10037 2548 10038 2573
rect 10038 2548 10072 2573
rect 10072 2548 10089 2573
rect 10037 2521 10089 2548
rect 10101 2548 10110 2573
rect 10110 2548 10144 2573
rect 10144 2548 10153 2573
rect 10101 2521 10153 2548
rect 10165 2548 10182 2573
rect 10182 2548 10216 2573
rect 10216 2548 10217 2573
rect 10165 2521 10217 2548
rect 10037 2474 10038 2508
rect 10038 2474 10072 2508
rect 10072 2474 10089 2508
rect 10037 2456 10089 2474
rect 10101 2474 10110 2508
rect 10110 2474 10144 2508
rect 10144 2474 10153 2508
rect 10101 2456 10153 2474
rect 10165 2474 10182 2508
rect 10182 2474 10216 2508
rect 10216 2474 10217 2508
rect 10165 2456 10217 2474
rect 10037 2434 10089 2443
rect 10037 2400 10038 2434
rect 10038 2400 10072 2434
rect 10072 2400 10089 2434
rect 10037 2391 10089 2400
rect 10101 2434 10153 2443
rect 10101 2400 10110 2434
rect 10110 2400 10144 2434
rect 10144 2400 10153 2434
rect 10101 2391 10153 2400
rect 10165 2434 10217 2443
rect 10165 2400 10182 2434
rect 10182 2400 10216 2434
rect 10216 2400 10217 2434
rect 10165 2391 10217 2400
rect 10037 2360 10089 2378
rect 10037 2326 10038 2360
rect 10038 2326 10072 2360
rect 10072 2326 10089 2360
rect 10101 2360 10153 2378
rect 10101 2326 10110 2360
rect 10110 2326 10144 2360
rect 10144 2326 10153 2360
rect 10165 2360 10217 2378
rect 10165 2326 10182 2360
rect 10182 2326 10216 2360
rect 10216 2326 10217 2360
rect 10037 2286 10089 2313
rect 10037 2261 10038 2286
rect 10038 2261 10072 2286
rect 10072 2261 10089 2286
rect 10101 2286 10153 2313
rect 10101 2261 10110 2286
rect 10110 2261 10144 2286
rect 10144 2261 10153 2286
rect 10165 2286 10217 2313
rect 10165 2261 10182 2286
rect 10182 2261 10216 2286
rect 10216 2261 10217 2286
rect 10037 2212 10089 2248
rect 10037 2196 10038 2212
rect 10038 2196 10072 2212
rect 10072 2196 10089 2212
rect 10101 2212 10153 2248
rect 10101 2196 10110 2212
rect 10110 2196 10144 2212
rect 10144 2196 10153 2212
rect 10165 2212 10217 2248
rect 10165 2196 10182 2212
rect 10182 2196 10216 2212
rect 10216 2196 10217 2212
rect 10037 2178 10038 2183
rect 10038 2178 10072 2183
rect 10072 2178 10089 2183
rect 10037 2138 10089 2178
rect 10037 2131 10038 2138
rect 10038 2131 10072 2138
rect 10072 2131 10089 2138
rect 10101 2178 10110 2183
rect 10110 2178 10144 2183
rect 10144 2178 10153 2183
rect 10101 2138 10153 2178
rect 10101 2131 10110 2138
rect 10110 2131 10144 2138
rect 10144 2131 10153 2138
rect 10165 2178 10182 2183
rect 10182 2178 10216 2183
rect 10216 2178 10217 2183
rect 10165 2138 10217 2178
rect 10165 2131 10182 2138
rect 10182 2131 10216 2138
rect 10216 2131 10217 2138
rect 10037 2104 10038 2118
rect 10038 2104 10072 2118
rect 10072 2104 10089 2118
rect 10037 2066 10089 2104
rect 10101 2104 10110 2118
rect 10110 2104 10144 2118
rect 10144 2104 10153 2118
rect 10101 2066 10153 2104
rect 10165 2104 10182 2118
rect 10182 2104 10216 2118
rect 10216 2104 10217 2118
rect 10165 2066 10217 2104
rect 10037 2030 10038 2053
rect 10038 2030 10072 2053
rect 10072 2030 10089 2053
rect 10037 2001 10089 2030
rect 10101 2030 10110 2053
rect 10110 2030 10144 2053
rect 10144 2030 10153 2053
rect 10101 2001 10153 2030
rect 10165 2030 10182 2053
rect 10182 2030 10216 2053
rect 10216 2030 10217 2053
rect 10165 2001 10217 2030
rect 10037 1956 10038 1987
rect 10038 1956 10072 1987
rect 10072 1956 10089 1987
rect 10037 1935 10089 1956
rect 10101 1956 10110 1987
rect 10110 1956 10144 1987
rect 10144 1956 10153 1987
rect 10101 1935 10153 1956
rect 10165 1956 10182 1987
rect 10182 1956 10216 1987
rect 10216 1956 10217 1987
rect 10165 1935 10217 1956
rect 10037 1916 10089 1921
rect 10037 1882 10038 1916
rect 10038 1882 10072 1916
rect 10072 1882 10089 1916
rect 10037 1869 10089 1882
rect 10101 1916 10153 1921
rect 10101 1882 10110 1916
rect 10110 1882 10144 1916
rect 10144 1882 10153 1916
rect 10101 1869 10153 1882
rect 10165 1916 10217 1921
rect 10165 1882 10182 1916
rect 10182 1882 10216 1916
rect 10216 1882 10217 1916
rect 10165 1869 10217 1882
rect 10037 1842 10089 1855
rect 10037 1808 10038 1842
rect 10038 1808 10072 1842
rect 10072 1808 10089 1842
rect 10037 1803 10089 1808
rect 10101 1842 10153 1855
rect 10101 1808 10110 1842
rect 10110 1808 10144 1842
rect 10144 1808 10153 1842
rect 10101 1803 10153 1808
rect 10165 1842 10217 1855
rect 10165 1808 10182 1842
rect 10182 1808 10216 1842
rect 10216 1808 10217 1842
rect 10165 1803 10217 1808
rect 10037 1768 10089 1789
rect 10037 1737 10038 1768
rect 10038 1737 10072 1768
rect 10072 1737 10089 1768
rect 10101 1768 10153 1789
rect 10101 1737 10110 1768
rect 10110 1737 10144 1768
rect 10144 1737 10153 1768
rect 10165 1768 10217 1789
rect 10165 1737 10182 1768
rect 10182 1737 10216 1768
rect 10216 1737 10217 1768
rect 10037 1694 10089 1723
rect 10037 1671 10038 1694
rect 10038 1671 10072 1694
rect 10072 1671 10089 1694
rect 10101 1694 10153 1723
rect 10101 1671 10110 1694
rect 10110 1671 10144 1694
rect 10144 1671 10153 1694
rect 10165 1694 10217 1723
rect 10165 1671 10182 1694
rect 10182 1671 10216 1694
rect 10216 1671 10217 1694
rect 10037 1620 10089 1657
rect 10037 1605 10038 1620
rect 10038 1605 10072 1620
rect 10072 1605 10089 1620
rect 10101 1620 10153 1657
rect 10101 1605 10110 1620
rect 10110 1605 10144 1620
rect 10144 1605 10153 1620
rect 10165 1620 10217 1657
rect 10165 1605 10182 1620
rect 10182 1605 10216 1620
rect 10216 1605 10217 1620
rect 10037 1586 10038 1591
rect 10038 1586 10072 1591
rect 10072 1586 10089 1591
rect 10037 1545 10089 1586
rect 10037 1539 10038 1545
rect 10038 1539 10072 1545
rect 10072 1539 10089 1545
rect 10101 1586 10110 1591
rect 10110 1586 10144 1591
rect 10144 1586 10153 1591
rect 10101 1545 10153 1586
rect 10101 1539 10110 1545
rect 10110 1539 10144 1545
rect 10144 1539 10153 1545
rect 10165 1586 10182 1591
rect 10182 1586 10216 1591
rect 10216 1586 10217 1591
rect 10165 1545 10217 1586
rect 10165 1539 10182 1545
rect 10182 1539 10216 1545
rect 10216 1539 10217 1545
rect 10037 1511 10038 1525
rect 10038 1511 10072 1525
rect 10072 1511 10089 1525
rect 10037 1473 10089 1511
rect 10101 1511 10110 1525
rect 10110 1511 10144 1525
rect 10144 1511 10153 1525
rect 10101 1473 10153 1511
rect 10165 1511 10182 1525
rect 10182 1511 10216 1525
rect 10216 1511 10217 1525
rect 10165 1473 10217 1511
rect 10533 4050 10585 4068
rect 10597 4062 10649 4068
rect 10597 4050 10606 4062
rect 10606 4050 10640 4062
rect 10640 4050 10649 4062
rect 10661 4050 10713 4068
rect 10533 4016 10534 4050
rect 10534 4016 10585 4050
rect 10597 4016 10649 4050
rect 10661 4016 10712 4050
rect 10712 4016 10713 4050
rect 10533 3951 10534 4003
rect 10534 3951 10585 4003
rect 10597 3951 10649 4003
rect 10661 3951 10712 4003
rect 10712 3951 10713 4003
rect 10533 3886 10534 3938
rect 10534 3886 10585 3938
rect 10597 3886 10649 3938
rect 10661 3886 10712 3938
rect 10712 3886 10713 3938
rect 10533 3821 10534 3873
rect 10534 3821 10585 3873
rect 10597 3821 10649 3873
rect 10661 3821 10712 3873
rect 10712 3821 10713 3873
rect 10533 3756 10534 3808
rect 10534 3756 10585 3808
rect 10597 3756 10649 3808
rect 10661 3756 10712 3808
rect 10712 3756 10713 3808
rect 10533 3691 10534 3743
rect 10534 3691 10585 3743
rect 10597 3691 10649 3743
rect 10661 3691 10712 3743
rect 10712 3691 10713 3743
rect 10533 3626 10534 3678
rect 10534 3626 10585 3678
rect 10597 3626 10649 3678
rect 10661 3626 10712 3678
rect 10712 3626 10713 3678
rect 10533 3561 10534 3613
rect 10534 3561 10585 3613
rect 10597 3561 10649 3613
rect 10661 3561 10712 3613
rect 10712 3561 10713 3613
rect 10533 3496 10534 3548
rect 10534 3496 10585 3548
rect 10597 3496 10649 3548
rect 10661 3496 10712 3548
rect 10712 3496 10713 3548
rect 10533 3431 10534 3483
rect 10534 3431 10585 3483
rect 10597 3431 10649 3483
rect 10661 3431 10712 3483
rect 10712 3431 10713 3483
rect 10533 3366 10534 3418
rect 10534 3366 10585 3418
rect 10597 3366 10649 3418
rect 10661 3366 10712 3418
rect 10712 3366 10713 3418
rect 10533 3301 10534 3353
rect 10534 3301 10585 3353
rect 10597 3301 10649 3353
rect 10661 3301 10712 3353
rect 10712 3301 10713 3353
rect 10533 3236 10534 3288
rect 10534 3236 10585 3288
rect 10597 3236 10649 3288
rect 10661 3236 10712 3288
rect 10712 3236 10713 3288
rect 10533 3171 10534 3223
rect 10534 3171 10585 3223
rect 10597 3171 10649 3223
rect 10661 3171 10712 3223
rect 10712 3171 10713 3223
rect 10533 3106 10534 3158
rect 10534 3106 10585 3158
rect 10597 3106 10649 3158
rect 10661 3106 10712 3158
rect 10712 3106 10713 3158
rect 10533 3080 10534 3093
rect 10534 3092 10585 3093
rect 10597 3092 10649 3093
rect 10661 3092 10712 3093
rect 10534 3080 10568 3092
rect 10568 3080 10585 3092
rect 10533 3041 10585 3080
rect 10597 3041 10649 3092
rect 10661 3080 10678 3092
rect 10678 3080 10712 3092
rect 10712 3080 10713 3093
rect 10661 3041 10713 3080
rect 10533 3003 10534 3028
rect 10534 3003 10568 3028
rect 10568 3003 10585 3028
rect 10533 2976 10585 3003
rect 10597 3003 10606 3028
rect 10606 3003 10640 3028
rect 10640 3003 10649 3028
rect 10597 2976 10649 3003
rect 10661 3003 10678 3028
rect 10678 3003 10712 3028
rect 10712 3003 10713 3028
rect 10661 2976 10713 3003
rect 10533 2954 10585 2963
rect 10533 2920 10534 2954
rect 10534 2920 10568 2954
rect 10568 2920 10585 2954
rect 10533 2911 10585 2920
rect 10597 2954 10649 2963
rect 10597 2920 10606 2954
rect 10606 2920 10640 2954
rect 10640 2920 10649 2954
rect 10597 2911 10649 2920
rect 10661 2954 10713 2963
rect 10661 2920 10678 2954
rect 10678 2920 10712 2954
rect 10712 2920 10713 2954
rect 10661 2911 10713 2920
rect 10533 2871 10585 2898
rect 10533 2846 10534 2871
rect 10534 2846 10568 2871
rect 10568 2846 10585 2871
rect 10597 2871 10649 2898
rect 10597 2846 10606 2871
rect 10606 2846 10640 2871
rect 10640 2846 10649 2871
rect 10661 2871 10713 2898
rect 10661 2846 10678 2871
rect 10678 2846 10712 2871
rect 10712 2846 10713 2871
rect 10533 2787 10585 2833
rect 10533 2781 10534 2787
rect 10534 2781 10568 2787
rect 10568 2781 10585 2787
rect 10597 2787 10649 2833
rect 10597 2781 10606 2787
rect 10606 2781 10640 2787
rect 10640 2781 10649 2787
rect 10661 2787 10713 2833
rect 10661 2781 10678 2787
rect 10678 2781 10712 2787
rect 10712 2781 10713 2787
rect 10533 2753 10534 2768
rect 10534 2753 10568 2768
rect 10568 2753 10585 2768
rect 10533 2716 10585 2753
rect 10597 2753 10606 2768
rect 10606 2753 10640 2768
rect 10640 2753 10649 2768
rect 10597 2716 10649 2753
rect 10661 2753 10678 2768
rect 10678 2753 10712 2768
rect 10712 2753 10713 2768
rect 10661 2716 10713 2753
rect 10533 2669 10534 2703
rect 10534 2669 10568 2703
rect 10568 2669 10585 2703
rect 10533 2651 10585 2669
rect 10597 2669 10606 2703
rect 10606 2669 10640 2703
rect 10640 2669 10649 2703
rect 10597 2651 10649 2669
rect 10661 2669 10678 2703
rect 10678 2669 10712 2703
rect 10712 2669 10713 2703
rect 10661 2651 10713 2669
rect 10533 2619 10585 2638
rect 10533 2586 10534 2619
rect 10534 2586 10568 2619
rect 10568 2586 10585 2619
rect 10597 2619 10649 2638
rect 10597 2586 10606 2619
rect 10606 2586 10640 2619
rect 10640 2586 10649 2619
rect 10661 2619 10713 2638
rect 10661 2586 10678 2619
rect 10678 2586 10712 2619
rect 10712 2586 10713 2619
rect 10533 2535 10585 2573
rect 10533 2521 10534 2535
rect 10534 2521 10568 2535
rect 10568 2521 10585 2535
rect 10597 2535 10649 2573
rect 10597 2521 10606 2535
rect 10606 2521 10640 2535
rect 10640 2521 10649 2535
rect 10661 2535 10713 2573
rect 10661 2521 10678 2535
rect 10678 2521 10712 2535
rect 10712 2521 10713 2535
rect 10533 2501 10534 2508
rect 10534 2501 10568 2508
rect 10568 2501 10585 2508
rect 10533 2456 10585 2501
rect 10597 2501 10606 2508
rect 10606 2501 10640 2508
rect 10640 2501 10649 2508
rect 10597 2461 10649 2501
rect 10597 2456 10606 2461
rect 10606 2456 10640 2461
rect 10640 2456 10649 2461
rect 10661 2501 10678 2508
rect 10678 2501 10712 2508
rect 10712 2501 10713 2508
rect 10661 2456 10713 2501
rect 10533 2391 10534 2443
rect 10534 2391 10585 2443
rect 10597 2391 10649 2443
rect 10661 2391 10712 2443
rect 10712 2391 10713 2443
rect 10533 2326 10534 2378
rect 10534 2326 10585 2378
rect 10597 2326 10649 2378
rect 10661 2326 10712 2378
rect 10712 2326 10713 2378
rect 10533 2261 10534 2313
rect 10534 2261 10585 2313
rect 10597 2261 10649 2313
rect 10661 2261 10712 2313
rect 10712 2261 10713 2313
rect 10533 2196 10534 2248
rect 10534 2196 10585 2248
rect 10597 2196 10649 2248
rect 10661 2196 10712 2248
rect 10712 2196 10713 2248
rect 10533 2131 10534 2183
rect 10534 2131 10585 2183
rect 10597 2131 10649 2183
rect 10661 2131 10712 2183
rect 10712 2131 10713 2183
rect 10533 2066 10534 2118
rect 10534 2066 10585 2118
rect 10597 2066 10649 2118
rect 10661 2066 10712 2118
rect 10712 2066 10713 2118
rect 10533 2001 10534 2053
rect 10534 2001 10585 2053
rect 10597 2001 10649 2053
rect 10661 2001 10712 2053
rect 10712 2001 10713 2053
rect 10533 1935 10534 1987
rect 10534 1935 10585 1987
rect 10597 1935 10649 1987
rect 10661 1935 10712 1987
rect 10712 1935 10713 1987
rect 10533 1869 10534 1921
rect 10534 1869 10585 1921
rect 10597 1869 10649 1921
rect 10661 1869 10712 1921
rect 10712 1869 10713 1921
rect 10533 1803 10534 1855
rect 10534 1803 10585 1855
rect 10597 1803 10649 1855
rect 10661 1803 10712 1855
rect 10712 1803 10713 1855
rect 10533 1737 10534 1789
rect 10534 1737 10585 1789
rect 10597 1737 10649 1789
rect 10661 1737 10712 1789
rect 10712 1737 10713 1789
rect 10533 1671 10534 1723
rect 10534 1671 10585 1723
rect 10597 1671 10649 1723
rect 10661 1671 10712 1723
rect 10712 1671 10713 1723
rect 10533 1605 10534 1657
rect 10534 1605 10585 1657
rect 10597 1605 10649 1657
rect 10661 1605 10712 1657
rect 10712 1605 10713 1657
rect 10533 1539 10534 1591
rect 10534 1539 10585 1591
rect 10597 1539 10649 1591
rect 10661 1539 10712 1591
rect 10712 1539 10713 1591
rect 10533 1479 10534 1525
rect 10534 1491 10585 1525
rect 10597 1491 10649 1525
rect 10661 1491 10712 1525
rect 10534 1479 10568 1491
rect 10568 1479 10585 1491
rect 10533 1473 10585 1479
rect 10597 1473 10649 1491
rect 10661 1479 10678 1491
rect 10678 1479 10712 1491
rect 10712 1479 10713 1525
rect 10661 1473 10713 1479
rect 11029 4062 11081 4068
rect 11029 4028 11030 4062
rect 11030 4028 11064 4062
rect 11064 4028 11081 4062
rect 11029 4016 11081 4028
rect 11093 4062 11145 4068
rect 11093 4028 11102 4062
rect 11102 4028 11136 4062
rect 11136 4028 11145 4062
rect 11093 4016 11145 4028
rect 11157 4062 11209 4068
rect 11157 4028 11174 4062
rect 11174 4028 11208 4062
rect 11208 4028 11209 4062
rect 11157 4016 11209 4028
rect 11029 3988 11081 4003
rect 11029 3954 11030 3988
rect 11030 3954 11064 3988
rect 11064 3954 11081 3988
rect 11029 3951 11081 3954
rect 11093 3988 11145 4003
rect 11093 3954 11102 3988
rect 11102 3954 11136 3988
rect 11136 3954 11145 3988
rect 11093 3951 11145 3954
rect 11157 3988 11209 4003
rect 11157 3954 11174 3988
rect 11174 3954 11208 3988
rect 11208 3954 11209 3988
rect 11157 3951 11209 3954
rect 11029 3914 11081 3938
rect 11029 3886 11030 3914
rect 11030 3886 11064 3914
rect 11064 3886 11081 3914
rect 11093 3914 11145 3938
rect 11093 3886 11102 3914
rect 11102 3886 11136 3914
rect 11136 3886 11145 3914
rect 11157 3914 11209 3938
rect 11157 3886 11174 3914
rect 11174 3886 11208 3914
rect 11208 3886 11209 3914
rect 11029 3840 11081 3873
rect 11029 3821 11030 3840
rect 11030 3821 11064 3840
rect 11064 3821 11081 3840
rect 11093 3840 11145 3873
rect 11093 3821 11102 3840
rect 11102 3821 11136 3840
rect 11136 3821 11145 3840
rect 11157 3840 11209 3873
rect 11157 3821 11174 3840
rect 11174 3821 11208 3840
rect 11208 3821 11209 3840
rect 11029 3806 11030 3808
rect 11030 3806 11064 3808
rect 11064 3806 11081 3808
rect 11029 3766 11081 3806
rect 11029 3756 11030 3766
rect 11030 3756 11064 3766
rect 11064 3756 11081 3766
rect 11093 3806 11102 3808
rect 11102 3806 11136 3808
rect 11136 3806 11145 3808
rect 11093 3766 11145 3806
rect 11093 3756 11102 3766
rect 11102 3756 11136 3766
rect 11136 3756 11145 3766
rect 11157 3806 11174 3808
rect 11174 3806 11208 3808
rect 11208 3806 11209 3808
rect 11157 3766 11209 3806
rect 11157 3756 11174 3766
rect 11174 3756 11208 3766
rect 11208 3756 11209 3766
rect 11029 3732 11030 3743
rect 11030 3732 11064 3743
rect 11064 3732 11081 3743
rect 11029 3692 11081 3732
rect 11029 3691 11030 3692
rect 11030 3691 11064 3692
rect 11064 3691 11081 3692
rect 11093 3732 11102 3743
rect 11102 3732 11136 3743
rect 11136 3732 11145 3743
rect 11093 3692 11145 3732
rect 11093 3691 11102 3692
rect 11102 3691 11136 3692
rect 11136 3691 11145 3692
rect 11157 3732 11174 3743
rect 11174 3732 11208 3743
rect 11208 3732 11209 3743
rect 11157 3692 11209 3732
rect 11157 3691 11174 3692
rect 11174 3691 11208 3692
rect 11208 3691 11209 3692
rect 11029 3658 11030 3678
rect 11030 3658 11064 3678
rect 11064 3658 11081 3678
rect 11029 3626 11081 3658
rect 11093 3658 11102 3678
rect 11102 3658 11136 3678
rect 11136 3658 11145 3678
rect 11093 3626 11145 3658
rect 11157 3658 11174 3678
rect 11174 3658 11208 3678
rect 11208 3658 11209 3678
rect 11157 3626 11209 3658
rect 11029 3584 11030 3613
rect 11030 3584 11064 3613
rect 11064 3584 11081 3613
rect 11029 3561 11081 3584
rect 11093 3584 11102 3613
rect 11102 3584 11136 3613
rect 11136 3584 11145 3613
rect 11093 3561 11145 3584
rect 11157 3584 11174 3613
rect 11174 3584 11208 3613
rect 11208 3584 11209 3613
rect 11157 3561 11209 3584
rect 11029 3544 11081 3548
rect 11029 3510 11030 3544
rect 11030 3510 11064 3544
rect 11064 3510 11081 3544
rect 11029 3496 11081 3510
rect 11093 3544 11145 3548
rect 11093 3510 11102 3544
rect 11102 3510 11136 3544
rect 11136 3510 11145 3544
rect 11093 3496 11145 3510
rect 11157 3544 11209 3548
rect 11157 3510 11174 3544
rect 11174 3510 11208 3544
rect 11208 3510 11209 3544
rect 11157 3496 11209 3510
rect 11029 3470 11081 3483
rect 11029 3436 11030 3470
rect 11030 3436 11064 3470
rect 11064 3436 11081 3470
rect 11029 3431 11081 3436
rect 11093 3470 11145 3483
rect 11093 3436 11102 3470
rect 11102 3436 11136 3470
rect 11136 3436 11145 3470
rect 11093 3431 11145 3436
rect 11157 3470 11209 3483
rect 11157 3436 11174 3470
rect 11174 3436 11208 3470
rect 11208 3436 11209 3470
rect 11157 3431 11209 3436
rect 11029 3396 11081 3418
rect 11029 3366 11030 3396
rect 11030 3366 11064 3396
rect 11064 3366 11081 3396
rect 11093 3396 11145 3418
rect 11093 3366 11102 3396
rect 11102 3366 11136 3396
rect 11136 3366 11145 3396
rect 11157 3396 11209 3418
rect 11157 3366 11174 3396
rect 11174 3366 11208 3396
rect 11208 3366 11209 3396
rect 11029 3322 11081 3353
rect 11029 3301 11030 3322
rect 11030 3301 11064 3322
rect 11064 3301 11081 3322
rect 11093 3322 11145 3353
rect 11093 3301 11102 3322
rect 11102 3301 11136 3322
rect 11136 3301 11145 3322
rect 11157 3322 11209 3353
rect 11157 3301 11174 3322
rect 11174 3301 11208 3322
rect 11208 3301 11209 3322
rect 11029 3248 11081 3288
rect 11029 3236 11030 3248
rect 11030 3236 11064 3248
rect 11064 3236 11081 3248
rect 11093 3248 11145 3288
rect 11093 3236 11102 3248
rect 11102 3236 11136 3248
rect 11136 3236 11145 3248
rect 11157 3248 11209 3288
rect 11157 3236 11174 3248
rect 11174 3236 11208 3248
rect 11208 3236 11209 3248
rect 11029 3214 11030 3223
rect 11030 3214 11064 3223
rect 11064 3214 11081 3223
rect 11029 3174 11081 3214
rect 11029 3171 11030 3174
rect 11030 3171 11064 3174
rect 11064 3171 11081 3174
rect 11093 3214 11102 3223
rect 11102 3214 11136 3223
rect 11136 3214 11145 3223
rect 11093 3174 11145 3214
rect 11093 3171 11102 3174
rect 11102 3171 11136 3174
rect 11136 3171 11145 3174
rect 11157 3214 11174 3223
rect 11174 3214 11208 3223
rect 11208 3214 11209 3223
rect 11157 3174 11209 3214
rect 11157 3171 11174 3174
rect 11174 3171 11208 3174
rect 11208 3171 11209 3174
rect 11029 3140 11030 3158
rect 11030 3140 11064 3158
rect 11064 3140 11081 3158
rect 11029 3106 11081 3140
rect 11093 3140 11102 3158
rect 11102 3140 11136 3158
rect 11136 3140 11145 3158
rect 11093 3106 11145 3140
rect 11157 3140 11174 3158
rect 11174 3140 11208 3158
rect 11208 3140 11209 3158
rect 11157 3106 11209 3140
rect 11029 3066 11030 3093
rect 11030 3066 11064 3093
rect 11064 3066 11081 3093
rect 11029 3041 11081 3066
rect 11093 3066 11102 3093
rect 11102 3066 11136 3093
rect 11136 3066 11145 3093
rect 11093 3041 11145 3066
rect 11157 3066 11174 3093
rect 11174 3066 11208 3093
rect 11208 3066 11209 3093
rect 11157 3041 11209 3066
rect 11029 3026 11081 3028
rect 11029 2992 11030 3026
rect 11030 2992 11064 3026
rect 11064 2992 11081 3026
rect 11029 2976 11081 2992
rect 11093 3026 11145 3028
rect 11093 2992 11102 3026
rect 11102 2992 11136 3026
rect 11136 2992 11145 3026
rect 11093 2976 11145 2992
rect 11157 3026 11209 3028
rect 11157 2992 11174 3026
rect 11174 2992 11208 3026
rect 11208 2992 11209 3026
rect 11157 2976 11209 2992
rect 11029 2952 11081 2963
rect 11029 2918 11030 2952
rect 11030 2918 11064 2952
rect 11064 2918 11081 2952
rect 11029 2911 11081 2918
rect 11093 2952 11145 2963
rect 11093 2918 11102 2952
rect 11102 2918 11136 2952
rect 11136 2918 11145 2952
rect 11093 2911 11145 2918
rect 11157 2952 11209 2963
rect 11157 2918 11174 2952
rect 11174 2918 11208 2952
rect 11208 2918 11209 2952
rect 11157 2911 11209 2918
rect 11029 2878 11081 2898
rect 11029 2846 11030 2878
rect 11030 2846 11064 2878
rect 11064 2846 11081 2878
rect 11093 2878 11145 2898
rect 11093 2846 11102 2878
rect 11102 2846 11136 2878
rect 11136 2846 11145 2878
rect 11157 2878 11209 2898
rect 11157 2846 11174 2878
rect 11174 2846 11208 2878
rect 11208 2846 11209 2878
rect 11029 2804 11081 2833
rect 11029 2781 11030 2804
rect 11030 2781 11064 2804
rect 11064 2781 11081 2804
rect 11093 2804 11145 2833
rect 11093 2781 11102 2804
rect 11102 2781 11136 2804
rect 11136 2781 11145 2804
rect 11157 2804 11209 2833
rect 11157 2781 11174 2804
rect 11174 2781 11208 2804
rect 11208 2781 11209 2804
rect 11029 2730 11081 2768
rect 11029 2716 11030 2730
rect 11030 2716 11064 2730
rect 11064 2716 11081 2730
rect 11093 2730 11145 2768
rect 11093 2716 11102 2730
rect 11102 2716 11136 2730
rect 11136 2716 11145 2730
rect 11157 2730 11209 2768
rect 11157 2716 11174 2730
rect 11174 2716 11208 2730
rect 11208 2716 11209 2730
rect 11029 2696 11030 2703
rect 11030 2696 11064 2703
rect 11064 2696 11081 2703
rect 11029 2656 11081 2696
rect 11029 2651 11030 2656
rect 11030 2651 11064 2656
rect 11064 2651 11081 2656
rect 11093 2696 11102 2703
rect 11102 2696 11136 2703
rect 11136 2696 11145 2703
rect 11093 2656 11145 2696
rect 11093 2651 11102 2656
rect 11102 2651 11136 2656
rect 11136 2651 11145 2656
rect 11157 2696 11174 2703
rect 11174 2696 11208 2703
rect 11208 2696 11209 2703
rect 11157 2656 11209 2696
rect 11157 2651 11174 2656
rect 11174 2651 11208 2656
rect 11208 2651 11209 2656
rect 11029 2622 11030 2638
rect 11030 2622 11064 2638
rect 11064 2622 11081 2638
rect 11029 2586 11081 2622
rect 11093 2622 11102 2638
rect 11102 2622 11136 2638
rect 11136 2622 11145 2638
rect 11093 2586 11145 2622
rect 11157 2622 11174 2638
rect 11174 2622 11208 2638
rect 11208 2622 11209 2638
rect 11157 2586 11209 2622
rect 11029 2548 11030 2573
rect 11030 2548 11064 2573
rect 11064 2548 11081 2573
rect 11029 2521 11081 2548
rect 11093 2548 11102 2573
rect 11102 2548 11136 2573
rect 11136 2548 11145 2573
rect 11093 2521 11145 2548
rect 11157 2548 11174 2573
rect 11174 2548 11208 2573
rect 11208 2548 11209 2573
rect 11157 2521 11209 2548
rect 11029 2474 11030 2508
rect 11030 2474 11064 2508
rect 11064 2474 11081 2508
rect 11029 2456 11081 2474
rect 11093 2474 11102 2508
rect 11102 2474 11136 2508
rect 11136 2474 11145 2508
rect 11093 2456 11145 2474
rect 11157 2474 11174 2508
rect 11174 2474 11208 2508
rect 11208 2474 11209 2508
rect 11157 2456 11209 2474
rect 11029 2434 11081 2443
rect 11029 2400 11030 2434
rect 11030 2400 11064 2434
rect 11064 2400 11081 2434
rect 11029 2391 11081 2400
rect 11093 2434 11145 2443
rect 11093 2400 11102 2434
rect 11102 2400 11136 2434
rect 11136 2400 11145 2434
rect 11093 2391 11145 2400
rect 11157 2434 11209 2443
rect 11157 2400 11174 2434
rect 11174 2400 11208 2434
rect 11208 2400 11209 2434
rect 11157 2391 11209 2400
rect 11029 2360 11081 2378
rect 11029 2326 11030 2360
rect 11030 2326 11064 2360
rect 11064 2326 11081 2360
rect 11093 2360 11145 2378
rect 11093 2326 11102 2360
rect 11102 2326 11136 2360
rect 11136 2326 11145 2360
rect 11157 2360 11209 2378
rect 11157 2326 11174 2360
rect 11174 2326 11208 2360
rect 11208 2326 11209 2360
rect 11029 2286 11081 2313
rect 11029 2261 11030 2286
rect 11030 2261 11064 2286
rect 11064 2261 11081 2286
rect 11093 2286 11145 2313
rect 11093 2261 11102 2286
rect 11102 2261 11136 2286
rect 11136 2261 11145 2286
rect 11157 2286 11209 2313
rect 11157 2261 11174 2286
rect 11174 2261 11208 2286
rect 11208 2261 11209 2286
rect 11029 2212 11081 2248
rect 11029 2196 11030 2212
rect 11030 2196 11064 2212
rect 11064 2196 11081 2212
rect 11093 2212 11145 2248
rect 11093 2196 11102 2212
rect 11102 2196 11136 2212
rect 11136 2196 11145 2212
rect 11157 2212 11209 2248
rect 11157 2196 11174 2212
rect 11174 2196 11208 2212
rect 11208 2196 11209 2212
rect 11029 2178 11030 2183
rect 11030 2178 11064 2183
rect 11064 2178 11081 2183
rect 11029 2138 11081 2178
rect 11029 2131 11030 2138
rect 11030 2131 11064 2138
rect 11064 2131 11081 2138
rect 11093 2178 11102 2183
rect 11102 2178 11136 2183
rect 11136 2178 11145 2183
rect 11093 2138 11145 2178
rect 11093 2131 11102 2138
rect 11102 2131 11136 2138
rect 11136 2131 11145 2138
rect 11157 2178 11174 2183
rect 11174 2178 11208 2183
rect 11208 2178 11209 2183
rect 11157 2138 11209 2178
rect 11157 2131 11174 2138
rect 11174 2131 11208 2138
rect 11208 2131 11209 2138
rect 11029 2104 11030 2118
rect 11030 2104 11064 2118
rect 11064 2104 11081 2118
rect 11029 2066 11081 2104
rect 11093 2104 11102 2118
rect 11102 2104 11136 2118
rect 11136 2104 11145 2118
rect 11093 2066 11145 2104
rect 11157 2104 11174 2118
rect 11174 2104 11208 2118
rect 11208 2104 11209 2118
rect 11157 2066 11209 2104
rect 11029 2030 11030 2053
rect 11030 2030 11064 2053
rect 11064 2030 11081 2053
rect 11029 2001 11081 2030
rect 11093 2030 11102 2053
rect 11102 2030 11136 2053
rect 11136 2030 11145 2053
rect 11093 2001 11145 2030
rect 11157 2030 11174 2053
rect 11174 2030 11208 2053
rect 11208 2030 11209 2053
rect 11157 2001 11209 2030
rect 11029 1956 11030 1987
rect 11030 1956 11064 1987
rect 11064 1956 11081 1987
rect 11029 1935 11081 1956
rect 11093 1956 11102 1987
rect 11102 1956 11136 1987
rect 11136 1956 11145 1987
rect 11093 1935 11145 1956
rect 11157 1956 11174 1987
rect 11174 1956 11208 1987
rect 11208 1956 11209 1987
rect 11157 1935 11209 1956
rect 11029 1916 11081 1921
rect 11029 1882 11030 1916
rect 11030 1882 11064 1916
rect 11064 1882 11081 1916
rect 11029 1869 11081 1882
rect 11093 1916 11145 1921
rect 11093 1882 11102 1916
rect 11102 1882 11136 1916
rect 11136 1882 11145 1916
rect 11093 1869 11145 1882
rect 11157 1916 11209 1921
rect 11157 1882 11174 1916
rect 11174 1882 11208 1916
rect 11208 1882 11209 1916
rect 11157 1869 11209 1882
rect 11029 1842 11081 1855
rect 11029 1808 11030 1842
rect 11030 1808 11064 1842
rect 11064 1808 11081 1842
rect 11029 1803 11081 1808
rect 11093 1842 11145 1855
rect 11093 1808 11102 1842
rect 11102 1808 11136 1842
rect 11136 1808 11145 1842
rect 11093 1803 11145 1808
rect 11157 1842 11209 1855
rect 11157 1808 11174 1842
rect 11174 1808 11208 1842
rect 11208 1808 11209 1842
rect 11157 1803 11209 1808
rect 11029 1768 11081 1789
rect 11029 1737 11030 1768
rect 11030 1737 11064 1768
rect 11064 1737 11081 1768
rect 11093 1768 11145 1789
rect 11093 1737 11102 1768
rect 11102 1737 11136 1768
rect 11136 1737 11145 1768
rect 11157 1768 11209 1789
rect 11157 1737 11174 1768
rect 11174 1737 11208 1768
rect 11208 1737 11209 1768
rect 11029 1694 11081 1723
rect 11029 1671 11030 1694
rect 11030 1671 11064 1694
rect 11064 1671 11081 1694
rect 11093 1694 11145 1723
rect 11093 1671 11102 1694
rect 11102 1671 11136 1694
rect 11136 1671 11145 1694
rect 11157 1694 11209 1723
rect 11157 1671 11174 1694
rect 11174 1671 11208 1694
rect 11208 1671 11209 1694
rect 11029 1620 11081 1657
rect 11029 1605 11030 1620
rect 11030 1605 11064 1620
rect 11064 1605 11081 1620
rect 11093 1620 11145 1657
rect 11093 1605 11102 1620
rect 11102 1605 11136 1620
rect 11136 1605 11145 1620
rect 11157 1620 11209 1657
rect 11157 1605 11174 1620
rect 11174 1605 11208 1620
rect 11208 1605 11209 1620
rect 11029 1586 11030 1591
rect 11030 1586 11064 1591
rect 11064 1586 11081 1591
rect 11029 1545 11081 1586
rect 11029 1539 11030 1545
rect 11030 1539 11064 1545
rect 11064 1539 11081 1545
rect 11093 1586 11102 1591
rect 11102 1586 11136 1591
rect 11136 1586 11145 1591
rect 11093 1545 11145 1586
rect 11093 1539 11102 1545
rect 11102 1539 11136 1545
rect 11136 1539 11145 1545
rect 11157 1586 11174 1591
rect 11174 1586 11208 1591
rect 11208 1586 11209 1591
rect 11157 1545 11209 1586
rect 11157 1539 11174 1545
rect 11174 1539 11208 1545
rect 11208 1539 11209 1545
rect 11029 1511 11030 1525
rect 11030 1511 11064 1525
rect 11064 1511 11081 1525
rect 11029 1473 11081 1511
rect 11093 1511 11102 1525
rect 11102 1511 11136 1525
rect 11136 1511 11145 1525
rect 11093 1473 11145 1511
rect 11157 1511 11174 1525
rect 11174 1511 11208 1525
rect 11208 1511 11209 1525
rect 11157 1473 11209 1511
rect 11525 4050 11577 4068
rect 11589 4062 11641 4068
rect 11589 4050 11598 4062
rect 11598 4050 11632 4062
rect 11632 4050 11641 4062
rect 11653 4050 11705 4068
rect 11525 4016 11526 4050
rect 11526 4016 11577 4050
rect 11589 4016 11641 4050
rect 11653 4016 11704 4050
rect 11704 4016 11705 4050
rect 11525 3951 11526 4003
rect 11526 3951 11577 4003
rect 11589 3951 11641 4003
rect 11653 3951 11704 4003
rect 11704 3951 11705 4003
rect 11525 3886 11526 3938
rect 11526 3886 11577 3938
rect 11589 3886 11641 3938
rect 11653 3886 11704 3938
rect 11704 3886 11705 3938
rect 11525 3821 11526 3873
rect 11526 3821 11577 3873
rect 11589 3821 11641 3873
rect 11653 3821 11704 3873
rect 11704 3821 11705 3873
rect 11525 3756 11526 3808
rect 11526 3756 11577 3808
rect 11589 3756 11641 3808
rect 11653 3756 11704 3808
rect 11704 3756 11705 3808
rect 11525 3691 11526 3743
rect 11526 3691 11577 3743
rect 11589 3691 11641 3743
rect 11653 3691 11704 3743
rect 11704 3691 11705 3743
rect 11525 3626 11526 3678
rect 11526 3626 11577 3678
rect 11589 3626 11641 3678
rect 11653 3626 11704 3678
rect 11704 3626 11705 3678
rect 11525 3561 11526 3613
rect 11526 3561 11577 3613
rect 11589 3561 11641 3613
rect 11653 3561 11704 3613
rect 11704 3561 11705 3613
rect 11525 3496 11526 3548
rect 11526 3496 11577 3548
rect 11589 3496 11641 3548
rect 11653 3496 11704 3548
rect 11704 3496 11705 3548
rect 11525 3431 11526 3483
rect 11526 3431 11577 3483
rect 11589 3431 11641 3483
rect 11653 3431 11704 3483
rect 11704 3431 11705 3483
rect 11525 3366 11526 3418
rect 11526 3366 11577 3418
rect 11589 3366 11641 3418
rect 11653 3366 11704 3418
rect 11704 3366 11705 3418
rect 11525 3301 11526 3353
rect 11526 3301 11577 3353
rect 11589 3301 11641 3353
rect 11653 3301 11704 3353
rect 11704 3301 11705 3353
rect 11525 3236 11526 3288
rect 11526 3236 11577 3288
rect 11589 3236 11641 3288
rect 11653 3236 11704 3288
rect 11704 3236 11705 3288
rect 11525 3171 11526 3223
rect 11526 3171 11577 3223
rect 11589 3171 11641 3223
rect 11653 3171 11704 3223
rect 11704 3171 11705 3223
rect 11525 3106 11526 3158
rect 11526 3106 11577 3158
rect 11589 3106 11641 3158
rect 11653 3106 11704 3158
rect 11704 3106 11705 3158
rect 11525 3080 11526 3093
rect 11526 3092 11577 3093
rect 11589 3092 11641 3093
rect 11653 3092 11704 3093
rect 11526 3080 11560 3092
rect 11560 3080 11577 3092
rect 11525 3041 11577 3080
rect 11589 3041 11641 3092
rect 11653 3080 11670 3092
rect 11670 3080 11704 3092
rect 11704 3080 11705 3093
rect 11653 3041 11705 3080
rect 11525 3003 11526 3028
rect 11526 3003 11560 3028
rect 11560 3003 11577 3028
rect 11525 2976 11577 3003
rect 11589 3003 11598 3028
rect 11598 3003 11632 3028
rect 11632 3003 11641 3028
rect 11589 2976 11641 3003
rect 11653 3003 11670 3028
rect 11670 3003 11704 3028
rect 11704 3003 11705 3028
rect 11653 2976 11705 3003
rect 11525 2954 11577 2963
rect 11525 2920 11526 2954
rect 11526 2920 11560 2954
rect 11560 2920 11577 2954
rect 11525 2911 11577 2920
rect 11589 2954 11641 2963
rect 11589 2920 11598 2954
rect 11598 2920 11632 2954
rect 11632 2920 11641 2954
rect 11589 2911 11641 2920
rect 11653 2954 11705 2963
rect 11653 2920 11670 2954
rect 11670 2920 11704 2954
rect 11704 2920 11705 2954
rect 11653 2911 11705 2920
rect 11525 2871 11577 2898
rect 11525 2846 11526 2871
rect 11526 2846 11560 2871
rect 11560 2846 11577 2871
rect 11589 2871 11641 2898
rect 11589 2846 11598 2871
rect 11598 2846 11632 2871
rect 11632 2846 11641 2871
rect 11653 2871 11705 2898
rect 11653 2846 11670 2871
rect 11670 2846 11704 2871
rect 11704 2846 11705 2871
rect 11525 2787 11577 2833
rect 11525 2781 11526 2787
rect 11526 2781 11560 2787
rect 11560 2781 11577 2787
rect 11589 2787 11641 2833
rect 11589 2781 11598 2787
rect 11598 2781 11632 2787
rect 11632 2781 11641 2787
rect 11653 2787 11705 2833
rect 11653 2781 11670 2787
rect 11670 2781 11704 2787
rect 11704 2781 11705 2787
rect 11525 2753 11526 2768
rect 11526 2753 11560 2768
rect 11560 2753 11577 2768
rect 11525 2716 11577 2753
rect 11589 2753 11598 2768
rect 11598 2753 11632 2768
rect 11632 2753 11641 2768
rect 11589 2716 11641 2753
rect 11653 2753 11670 2768
rect 11670 2753 11704 2768
rect 11704 2753 11705 2768
rect 11653 2716 11705 2753
rect 11525 2669 11526 2703
rect 11526 2669 11560 2703
rect 11560 2669 11577 2703
rect 11525 2651 11577 2669
rect 11589 2669 11598 2703
rect 11598 2669 11632 2703
rect 11632 2669 11641 2703
rect 11589 2651 11641 2669
rect 11653 2669 11670 2703
rect 11670 2669 11704 2703
rect 11704 2669 11705 2703
rect 11653 2651 11705 2669
rect 11525 2619 11577 2638
rect 11525 2586 11526 2619
rect 11526 2586 11560 2619
rect 11560 2586 11577 2619
rect 11589 2619 11641 2638
rect 11589 2586 11598 2619
rect 11598 2586 11632 2619
rect 11632 2586 11641 2619
rect 11653 2619 11705 2638
rect 11653 2586 11670 2619
rect 11670 2586 11704 2619
rect 11704 2586 11705 2619
rect 11525 2535 11577 2573
rect 11525 2521 11526 2535
rect 11526 2521 11560 2535
rect 11560 2521 11577 2535
rect 11589 2535 11641 2573
rect 11589 2521 11598 2535
rect 11598 2521 11632 2535
rect 11632 2521 11641 2535
rect 11653 2535 11705 2573
rect 11653 2521 11670 2535
rect 11670 2521 11704 2535
rect 11704 2521 11705 2535
rect 11525 2501 11526 2508
rect 11526 2501 11560 2508
rect 11560 2501 11577 2508
rect 11525 2456 11577 2501
rect 11589 2501 11598 2508
rect 11598 2501 11632 2508
rect 11632 2501 11641 2508
rect 11589 2461 11641 2501
rect 11589 2456 11598 2461
rect 11598 2456 11632 2461
rect 11632 2456 11641 2461
rect 11653 2501 11670 2508
rect 11670 2501 11704 2508
rect 11704 2501 11705 2508
rect 11653 2456 11705 2501
rect 11525 2391 11526 2443
rect 11526 2391 11577 2443
rect 11589 2391 11641 2443
rect 11653 2391 11704 2443
rect 11704 2391 11705 2443
rect 11525 2326 11526 2378
rect 11526 2326 11577 2378
rect 11589 2326 11641 2378
rect 11653 2326 11704 2378
rect 11704 2326 11705 2378
rect 11525 2261 11526 2313
rect 11526 2261 11577 2313
rect 11589 2261 11641 2313
rect 11653 2261 11704 2313
rect 11704 2261 11705 2313
rect 11525 2196 11526 2248
rect 11526 2196 11577 2248
rect 11589 2196 11641 2248
rect 11653 2196 11704 2248
rect 11704 2196 11705 2248
rect 11525 2131 11526 2183
rect 11526 2131 11577 2183
rect 11589 2131 11641 2183
rect 11653 2131 11704 2183
rect 11704 2131 11705 2183
rect 11525 2066 11526 2118
rect 11526 2066 11577 2118
rect 11589 2066 11641 2118
rect 11653 2066 11704 2118
rect 11704 2066 11705 2118
rect 11525 2001 11526 2053
rect 11526 2001 11577 2053
rect 11589 2001 11641 2053
rect 11653 2001 11704 2053
rect 11704 2001 11705 2053
rect 11525 1935 11526 1987
rect 11526 1935 11577 1987
rect 11589 1935 11641 1987
rect 11653 1935 11704 1987
rect 11704 1935 11705 1987
rect 11525 1869 11526 1921
rect 11526 1869 11577 1921
rect 11589 1869 11641 1921
rect 11653 1869 11704 1921
rect 11704 1869 11705 1921
rect 11525 1803 11526 1855
rect 11526 1803 11577 1855
rect 11589 1803 11641 1855
rect 11653 1803 11704 1855
rect 11704 1803 11705 1855
rect 11525 1737 11526 1789
rect 11526 1737 11577 1789
rect 11589 1737 11641 1789
rect 11653 1737 11704 1789
rect 11704 1737 11705 1789
rect 11525 1671 11526 1723
rect 11526 1671 11577 1723
rect 11589 1671 11641 1723
rect 11653 1671 11704 1723
rect 11704 1671 11705 1723
rect 11525 1605 11526 1657
rect 11526 1605 11577 1657
rect 11589 1605 11641 1657
rect 11653 1605 11704 1657
rect 11704 1605 11705 1657
rect 11525 1539 11526 1591
rect 11526 1539 11577 1591
rect 11589 1539 11641 1591
rect 11653 1539 11704 1591
rect 11704 1539 11705 1591
rect 11525 1479 11526 1525
rect 11526 1491 11577 1525
rect 11589 1491 11641 1525
rect 11653 1491 11704 1525
rect 11526 1479 11560 1491
rect 11560 1479 11577 1491
rect 11525 1473 11577 1479
rect 11589 1473 11641 1491
rect 11653 1479 11670 1491
rect 11670 1479 11704 1491
rect 11704 1479 11705 1525
rect 11653 1473 11705 1479
rect 12021 4062 12073 4068
rect 12021 4028 12022 4062
rect 12022 4028 12056 4062
rect 12056 4028 12073 4062
rect 12021 4016 12073 4028
rect 12085 4062 12137 4068
rect 12085 4028 12094 4062
rect 12094 4028 12128 4062
rect 12128 4028 12137 4062
rect 12085 4016 12137 4028
rect 12149 4062 12201 4068
rect 12149 4028 12166 4062
rect 12166 4028 12200 4062
rect 12200 4028 12201 4062
rect 12149 4016 12201 4028
rect 12021 3988 12073 4003
rect 12021 3954 12022 3988
rect 12022 3954 12056 3988
rect 12056 3954 12073 3988
rect 12021 3951 12073 3954
rect 12085 3988 12137 4003
rect 12085 3954 12094 3988
rect 12094 3954 12128 3988
rect 12128 3954 12137 3988
rect 12085 3951 12137 3954
rect 12149 3988 12201 4003
rect 12149 3954 12166 3988
rect 12166 3954 12200 3988
rect 12200 3954 12201 3988
rect 12149 3951 12201 3954
rect 12021 3914 12073 3938
rect 12021 3886 12022 3914
rect 12022 3886 12056 3914
rect 12056 3886 12073 3914
rect 12085 3914 12137 3938
rect 12085 3886 12094 3914
rect 12094 3886 12128 3914
rect 12128 3886 12137 3914
rect 12149 3914 12201 3938
rect 12149 3886 12166 3914
rect 12166 3886 12200 3914
rect 12200 3886 12201 3914
rect 12021 3840 12073 3873
rect 12021 3821 12022 3840
rect 12022 3821 12056 3840
rect 12056 3821 12073 3840
rect 12085 3840 12137 3873
rect 12085 3821 12094 3840
rect 12094 3821 12128 3840
rect 12128 3821 12137 3840
rect 12149 3840 12201 3873
rect 12149 3821 12166 3840
rect 12166 3821 12200 3840
rect 12200 3821 12201 3840
rect 12021 3806 12022 3808
rect 12022 3806 12056 3808
rect 12056 3806 12073 3808
rect 12021 3766 12073 3806
rect 12021 3756 12022 3766
rect 12022 3756 12056 3766
rect 12056 3756 12073 3766
rect 12085 3806 12094 3808
rect 12094 3806 12128 3808
rect 12128 3806 12137 3808
rect 12085 3766 12137 3806
rect 12085 3756 12094 3766
rect 12094 3756 12128 3766
rect 12128 3756 12137 3766
rect 12149 3806 12166 3808
rect 12166 3806 12200 3808
rect 12200 3806 12201 3808
rect 12149 3766 12201 3806
rect 12149 3756 12166 3766
rect 12166 3756 12200 3766
rect 12200 3756 12201 3766
rect 12021 3732 12022 3743
rect 12022 3732 12056 3743
rect 12056 3732 12073 3743
rect 12021 3692 12073 3732
rect 12021 3691 12022 3692
rect 12022 3691 12056 3692
rect 12056 3691 12073 3692
rect 12085 3732 12094 3743
rect 12094 3732 12128 3743
rect 12128 3732 12137 3743
rect 12085 3692 12137 3732
rect 12085 3691 12094 3692
rect 12094 3691 12128 3692
rect 12128 3691 12137 3692
rect 12149 3732 12166 3743
rect 12166 3732 12200 3743
rect 12200 3732 12201 3743
rect 12149 3692 12201 3732
rect 12149 3691 12166 3692
rect 12166 3691 12200 3692
rect 12200 3691 12201 3692
rect 12021 3658 12022 3678
rect 12022 3658 12056 3678
rect 12056 3658 12073 3678
rect 12021 3626 12073 3658
rect 12085 3658 12094 3678
rect 12094 3658 12128 3678
rect 12128 3658 12137 3678
rect 12085 3626 12137 3658
rect 12149 3658 12166 3678
rect 12166 3658 12200 3678
rect 12200 3658 12201 3678
rect 12149 3626 12201 3658
rect 12021 3584 12022 3613
rect 12022 3584 12056 3613
rect 12056 3584 12073 3613
rect 12021 3561 12073 3584
rect 12085 3584 12094 3613
rect 12094 3584 12128 3613
rect 12128 3584 12137 3613
rect 12085 3561 12137 3584
rect 12149 3584 12166 3613
rect 12166 3584 12200 3613
rect 12200 3584 12201 3613
rect 12149 3561 12201 3584
rect 12021 3544 12073 3548
rect 12021 3510 12022 3544
rect 12022 3510 12056 3544
rect 12056 3510 12073 3544
rect 12021 3496 12073 3510
rect 12085 3544 12137 3548
rect 12085 3510 12094 3544
rect 12094 3510 12128 3544
rect 12128 3510 12137 3544
rect 12085 3496 12137 3510
rect 12149 3544 12201 3548
rect 12149 3510 12166 3544
rect 12166 3510 12200 3544
rect 12200 3510 12201 3544
rect 12149 3496 12201 3510
rect 12021 3470 12073 3483
rect 12021 3436 12022 3470
rect 12022 3436 12056 3470
rect 12056 3436 12073 3470
rect 12021 3431 12073 3436
rect 12085 3470 12137 3483
rect 12085 3436 12094 3470
rect 12094 3436 12128 3470
rect 12128 3436 12137 3470
rect 12085 3431 12137 3436
rect 12149 3470 12201 3483
rect 12149 3436 12166 3470
rect 12166 3436 12200 3470
rect 12200 3436 12201 3470
rect 12149 3431 12201 3436
rect 12021 3396 12073 3418
rect 12021 3366 12022 3396
rect 12022 3366 12056 3396
rect 12056 3366 12073 3396
rect 12085 3396 12137 3418
rect 12085 3366 12094 3396
rect 12094 3366 12128 3396
rect 12128 3366 12137 3396
rect 12149 3396 12201 3418
rect 12149 3366 12166 3396
rect 12166 3366 12200 3396
rect 12200 3366 12201 3396
rect 12021 3322 12073 3353
rect 12021 3301 12022 3322
rect 12022 3301 12056 3322
rect 12056 3301 12073 3322
rect 12085 3322 12137 3353
rect 12085 3301 12094 3322
rect 12094 3301 12128 3322
rect 12128 3301 12137 3322
rect 12149 3322 12201 3353
rect 12149 3301 12166 3322
rect 12166 3301 12200 3322
rect 12200 3301 12201 3322
rect 12021 3248 12073 3288
rect 12021 3236 12022 3248
rect 12022 3236 12056 3248
rect 12056 3236 12073 3248
rect 12085 3248 12137 3288
rect 12085 3236 12094 3248
rect 12094 3236 12128 3248
rect 12128 3236 12137 3248
rect 12149 3248 12201 3288
rect 12149 3236 12166 3248
rect 12166 3236 12200 3248
rect 12200 3236 12201 3248
rect 12021 3214 12022 3223
rect 12022 3214 12056 3223
rect 12056 3214 12073 3223
rect 12021 3174 12073 3214
rect 12021 3171 12022 3174
rect 12022 3171 12056 3174
rect 12056 3171 12073 3174
rect 12085 3214 12094 3223
rect 12094 3214 12128 3223
rect 12128 3214 12137 3223
rect 12085 3174 12137 3214
rect 12085 3171 12094 3174
rect 12094 3171 12128 3174
rect 12128 3171 12137 3174
rect 12149 3214 12166 3223
rect 12166 3214 12200 3223
rect 12200 3214 12201 3223
rect 12149 3174 12201 3214
rect 12149 3171 12166 3174
rect 12166 3171 12200 3174
rect 12200 3171 12201 3174
rect 12021 3140 12022 3158
rect 12022 3140 12056 3158
rect 12056 3140 12073 3158
rect 12021 3106 12073 3140
rect 12085 3140 12094 3158
rect 12094 3140 12128 3158
rect 12128 3140 12137 3158
rect 12085 3106 12137 3140
rect 12149 3140 12166 3158
rect 12166 3140 12200 3158
rect 12200 3140 12201 3158
rect 12149 3106 12201 3140
rect 12021 3066 12022 3093
rect 12022 3066 12056 3093
rect 12056 3066 12073 3093
rect 12021 3041 12073 3066
rect 12085 3066 12094 3093
rect 12094 3066 12128 3093
rect 12128 3066 12137 3093
rect 12085 3041 12137 3066
rect 12149 3066 12166 3093
rect 12166 3066 12200 3093
rect 12200 3066 12201 3093
rect 12149 3041 12201 3066
rect 12021 3026 12073 3028
rect 12021 2992 12022 3026
rect 12022 2992 12056 3026
rect 12056 2992 12073 3026
rect 12021 2976 12073 2992
rect 12085 3026 12137 3028
rect 12085 2992 12094 3026
rect 12094 2992 12128 3026
rect 12128 2992 12137 3026
rect 12085 2976 12137 2992
rect 12149 3026 12201 3028
rect 12149 2992 12166 3026
rect 12166 2992 12200 3026
rect 12200 2992 12201 3026
rect 12149 2976 12201 2992
rect 12021 2952 12073 2963
rect 12021 2918 12022 2952
rect 12022 2918 12056 2952
rect 12056 2918 12073 2952
rect 12021 2911 12073 2918
rect 12085 2952 12137 2963
rect 12085 2918 12094 2952
rect 12094 2918 12128 2952
rect 12128 2918 12137 2952
rect 12085 2911 12137 2918
rect 12149 2952 12201 2963
rect 12149 2918 12166 2952
rect 12166 2918 12200 2952
rect 12200 2918 12201 2952
rect 12149 2911 12201 2918
rect 12021 2878 12073 2898
rect 12021 2846 12022 2878
rect 12022 2846 12056 2878
rect 12056 2846 12073 2878
rect 12085 2878 12137 2898
rect 12085 2846 12094 2878
rect 12094 2846 12128 2878
rect 12128 2846 12137 2878
rect 12149 2878 12201 2898
rect 12149 2846 12166 2878
rect 12166 2846 12200 2878
rect 12200 2846 12201 2878
rect 12021 2804 12073 2833
rect 12021 2781 12022 2804
rect 12022 2781 12056 2804
rect 12056 2781 12073 2804
rect 12085 2804 12137 2833
rect 12085 2781 12094 2804
rect 12094 2781 12128 2804
rect 12128 2781 12137 2804
rect 12149 2804 12201 2833
rect 12149 2781 12166 2804
rect 12166 2781 12200 2804
rect 12200 2781 12201 2804
rect 12021 2730 12073 2768
rect 12021 2716 12022 2730
rect 12022 2716 12056 2730
rect 12056 2716 12073 2730
rect 12085 2730 12137 2768
rect 12085 2716 12094 2730
rect 12094 2716 12128 2730
rect 12128 2716 12137 2730
rect 12149 2730 12201 2768
rect 12149 2716 12166 2730
rect 12166 2716 12200 2730
rect 12200 2716 12201 2730
rect 12021 2696 12022 2703
rect 12022 2696 12056 2703
rect 12056 2696 12073 2703
rect 12021 2656 12073 2696
rect 12021 2651 12022 2656
rect 12022 2651 12056 2656
rect 12056 2651 12073 2656
rect 12085 2696 12094 2703
rect 12094 2696 12128 2703
rect 12128 2696 12137 2703
rect 12085 2656 12137 2696
rect 12085 2651 12094 2656
rect 12094 2651 12128 2656
rect 12128 2651 12137 2656
rect 12149 2696 12166 2703
rect 12166 2696 12200 2703
rect 12200 2696 12201 2703
rect 12149 2656 12201 2696
rect 12149 2651 12166 2656
rect 12166 2651 12200 2656
rect 12200 2651 12201 2656
rect 12021 2622 12022 2638
rect 12022 2622 12056 2638
rect 12056 2622 12073 2638
rect 12021 2586 12073 2622
rect 12085 2622 12094 2638
rect 12094 2622 12128 2638
rect 12128 2622 12137 2638
rect 12085 2586 12137 2622
rect 12149 2622 12166 2638
rect 12166 2622 12200 2638
rect 12200 2622 12201 2638
rect 12149 2586 12201 2622
rect 12021 2548 12022 2573
rect 12022 2548 12056 2573
rect 12056 2548 12073 2573
rect 12021 2521 12073 2548
rect 12085 2548 12094 2573
rect 12094 2548 12128 2573
rect 12128 2548 12137 2573
rect 12085 2521 12137 2548
rect 12149 2548 12166 2573
rect 12166 2548 12200 2573
rect 12200 2548 12201 2573
rect 12149 2521 12201 2548
rect 12021 2474 12022 2508
rect 12022 2474 12056 2508
rect 12056 2474 12073 2508
rect 12021 2456 12073 2474
rect 12085 2474 12094 2508
rect 12094 2474 12128 2508
rect 12128 2474 12137 2508
rect 12085 2456 12137 2474
rect 12149 2474 12166 2508
rect 12166 2474 12200 2508
rect 12200 2474 12201 2508
rect 12149 2456 12201 2474
rect 12021 2434 12073 2443
rect 12021 2400 12022 2434
rect 12022 2400 12056 2434
rect 12056 2400 12073 2434
rect 12021 2391 12073 2400
rect 12085 2434 12137 2443
rect 12085 2400 12094 2434
rect 12094 2400 12128 2434
rect 12128 2400 12137 2434
rect 12085 2391 12137 2400
rect 12149 2434 12201 2443
rect 12149 2400 12166 2434
rect 12166 2400 12200 2434
rect 12200 2400 12201 2434
rect 12149 2391 12201 2400
rect 12021 2360 12073 2378
rect 12021 2326 12022 2360
rect 12022 2326 12056 2360
rect 12056 2326 12073 2360
rect 12085 2360 12137 2378
rect 12085 2326 12094 2360
rect 12094 2326 12128 2360
rect 12128 2326 12137 2360
rect 12149 2360 12201 2378
rect 12149 2326 12166 2360
rect 12166 2326 12200 2360
rect 12200 2326 12201 2360
rect 12021 2286 12073 2313
rect 12021 2261 12022 2286
rect 12022 2261 12056 2286
rect 12056 2261 12073 2286
rect 12085 2286 12137 2313
rect 12085 2261 12094 2286
rect 12094 2261 12128 2286
rect 12128 2261 12137 2286
rect 12149 2286 12201 2313
rect 12149 2261 12166 2286
rect 12166 2261 12200 2286
rect 12200 2261 12201 2286
rect 12021 2212 12073 2248
rect 12021 2196 12022 2212
rect 12022 2196 12056 2212
rect 12056 2196 12073 2212
rect 12085 2212 12137 2248
rect 12085 2196 12094 2212
rect 12094 2196 12128 2212
rect 12128 2196 12137 2212
rect 12149 2212 12201 2248
rect 12149 2196 12166 2212
rect 12166 2196 12200 2212
rect 12200 2196 12201 2212
rect 12021 2178 12022 2183
rect 12022 2178 12056 2183
rect 12056 2178 12073 2183
rect 12021 2138 12073 2178
rect 12021 2131 12022 2138
rect 12022 2131 12056 2138
rect 12056 2131 12073 2138
rect 12085 2178 12094 2183
rect 12094 2178 12128 2183
rect 12128 2178 12137 2183
rect 12085 2138 12137 2178
rect 12085 2131 12094 2138
rect 12094 2131 12128 2138
rect 12128 2131 12137 2138
rect 12149 2178 12166 2183
rect 12166 2178 12200 2183
rect 12200 2178 12201 2183
rect 12149 2138 12201 2178
rect 12149 2131 12166 2138
rect 12166 2131 12200 2138
rect 12200 2131 12201 2138
rect 12021 2104 12022 2118
rect 12022 2104 12056 2118
rect 12056 2104 12073 2118
rect 12021 2066 12073 2104
rect 12085 2104 12094 2118
rect 12094 2104 12128 2118
rect 12128 2104 12137 2118
rect 12085 2066 12137 2104
rect 12149 2104 12166 2118
rect 12166 2104 12200 2118
rect 12200 2104 12201 2118
rect 12149 2066 12201 2104
rect 12021 2030 12022 2053
rect 12022 2030 12056 2053
rect 12056 2030 12073 2053
rect 12021 2001 12073 2030
rect 12085 2030 12094 2053
rect 12094 2030 12128 2053
rect 12128 2030 12137 2053
rect 12085 2001 12137 2030
rect 12149 2030 12166 2053
rect 12166 2030 12200 2053
rect 12200 2030 12201 2053
rect 12149 2001 12201 2030
rect 12021 1956 12022 1987
rect 12022 1956 12056 1987
rect 12056 1956 12073 1987
rect 12021 1935 12073 1956
rect 12085 1956 12094 1987
rect 12094 1956 12128 1987
rect 12128 1956 12137 1987
rect 12085 1935 12137 1956
rect 12149 1956 12166 1987
rect 12166 1956 12200 1987
rect 12200 1956 12201 1987
rect 12149 1935 12201 1956
rect 12021 1916 12073 1921
rect 12021 1882 12022 1916
rect 12022 1882 12056 1916
rect 12056 1882 12073 1916
rect 12021 1869 12073 1882
rect 12085 1916 12137 1921
rect 12085 1882 12094 1916
rect 12094 1882 12128 1916
rect 12128 1882 12137 1916
rect 12085 1869 12137 1882
rect 12149 1916 12201 1921
rect 12149 1882 12166 1916
rect 12166 1882 12200 1916
rect 12200 1882 12201 1916
rect 12149 1869 12201 1882
rect 12021 1842 12073 1855
rect 12021 1808 12022 1842
rect 12022 1808 12056 1842
rect 12056 1808 12073 1842
rect 12021 1803 12073 1808
rect 12085 1842 12137 1855
rect 12085 1808 12094 1842
rect 12094 1808 12128 1842
rect 12128 1808 12137 1842
rect 12085 1803 12137 1808
rect 12149 1842 12201 1855
rect 12149 1808 12166 1842
rect 12166 1808 12200 1842
rect 12200 1808 12201 1842
rect 12149 1803 12201 1808
rect 12021 1768 12073 1789
rect 12021 1737 12022 1768
rect 12022 1737 12056 1768
rect 12056 1737 12073 1768
rect 12085 1768 12137 1789
rect 12085 1737 12094 1768
rect 12094 1737 12128 1768
rect 12128 1737 12137 1768
rect 12149 1768 12201 1789
rect 12149 1737 12166 1768
rect 12166 1737 12200 1768
rect 12200 1737 12201 1768
rect 12021 1694 12073 1723
rect 12021 1671 12022 1694
rect 12022 1671 12056 1694
rect 12056 1671 12073 1694
rect 12085 1694 12137 1723
rect 12085 1671 12094 1694
rect 12094 1671 12128 1694
rect 12128 1671 12137 1694
rect 12149 1694 12201 1723
rect 12149 1671 12166 1694
rect 12166 1671 12200 1694
rect 12200 1671 12201 1694
rect 12021 1620 12073 1657
rect 12021 1605 12022 1620
rect 12022 1605 12056 1620
rect 12056 1605 12073 1620
rect 12085 1620 12137 1657
rect 12085 1605 12094 1620
rect 12094 1605 12128 1620
rect 12128 1605 12137 1620
rect 12149 1620 12201 1657
rect 12149 1605 12166 1620
rect 12166 1605 12200 1620
rect 12200 1605 12201 1620
rect 12021 1586 12022 1591
rect 12022 1586 12056 1591
rect 12056 1586 12073 1591
rect 12021 1545 12073 1586
rect 12021 1539 12022 1545
rect 12022 1539 12056 1545
rect 12056 1539 12073 1545
rect 12085 1586 12094 1591
rect 12094 1586 12128 1591
rect 12128 1586 12137 1591
rect 12085 1545 12137 1586
rect 12085 1539 12094 1545
rect 12094 1539 12128 1545
rect 12128 1539 12137 1545
rect 12149 1586 12166 1591
rect 12166 1586 12200 1591
rect 12200 1586 12201 1591
rect 12149 1545 12201 1586
rect 12149 1539 12166 1545
rect 12166 1539 12200 1545
rect 12200 1539 12201 1545
rect 12021 1511 12022 1525
rect 12022 1511 12056 1525
rect 12056 1511 12073 1525
rect 12021 1473 12073 1511
rect 12085 1511 12094 1525
rect 12094 1511 12128 1525
rect 12128 1511 12137 1525
rect 12085 1473 12137 1511
rect 12149 1511 12166 1525
rect 12166 1511 12200 1525
rect 12200 1511 12201 1525
rect 12149 1473 12201 1511
rect 12517 4050 12569 4068
rect 12581 4062 12633 4068
rect 12581 4050 12590 4062
rect 12590 4050 12624 4062
rect 12624 4050 12633 4062
rect 12645 4050 12697 4068
rect 12517 4016 12518 4050
rect 12518 4016 12569 4050
rect 12581 4016 12633 4050
rect 12645 4016 12696 4050
rect 12696 4016 12697 4050
rect 12517 3951 12518 4003
rect 12518 3951 12569 4003
rect 12581 3951 12633 4003
rect 12645 3951 12696 4003
rect 12696 3951 12697 4003
rect 12517 3886 12518 3938
rect 12518 3886 12569 3938
rect 12581 3886 12633 3938
rect 12645 3886 12696 3938
rect 12696 3886 12697 3938
rect 12517 3821 12518 3873
rect 12518 3821 12569 3873
rect 12581 3821 12633 3873
rect 12645 3821 12696 3873
rect 12696 3821 12697 3873
rect 12517 3756 12518 3808
rect 12518 3756 12569 3808
rect 12581 3756 12633 3808
rect 12645 3756 12696 3808
rect 12696 3756 12697 3808
rect 12517 3691 12518 3743
rect 12518 3691 12569 3743
rect 12581 3691 12633 3743
rect 12645 3691 12696 3743
rect 12696 3691 12697 3743
rect 12517 3626 12518 3678
rect 12518 3626 12569 3678
rect 12581 3626 12633 3678
rect 12645 3626 12696 3678
rect 12696 3626 12697 3678
rect 12517 3561 12518 3613
rect 12518 3561 12569 3613
rect 12581 3561 12633 3613
rect 12645 3561 12696 3613
rect 12696 3561 12697 3613
rect 12517 3496 12518 3548
rect 12518 3496 12569 3548
rect 12581 3496 12633 3548
rect 12645 3496 12696 3548
rect 12696 3496 12697 3548
rect 12517 3431 12518 3483
rect 12518 3431 12569 3483
rect 12581 3431 12633 3483
rect 12645 3431 12696 3483
rect 12696 3431 12697 3483
rect 12517 3366 12518 3418
rect 12518 3366 12569 3418
rect 12581 3366 12633 3418
rect 12645 3366 12696 3418
rect 12696 3366 12697 3418
rect 12517 3301 12518 3353
rect 12518 3301 12569 3353
rect 12581 3301 12633 3353
rect 12645 3301 12696 3353
rect 12696 3301 12697 3353
rect 12517 3236 12518 3288
rect 12518 3236 12569 3288
rect 12581 3236 12633 3288
rect 12645 3236 12696 3288
rect 12696 3236 12697 3288
rect 12517 3171 12518 3223
rect 12518 3171 12569 3223
rect 12581 3171 12633 3223
rect 12645 3171 12696 3223
rect 12696 3171 12697 3223
rect 12517 3106 12518 3158
rect 12518 3106 12569 3158
rect 12581 3106 12633 3158
rect 12645 3106 12696 3158
rect 12696 3106 12697 3158
rect 12517 3080 12518 3093
rect 12518 3092 12569 3093
rect 12581 3092 12633 3093
rect 12645 3092 12696 3093
rect 12518 3080 12552 3092
rect 12552 3080 12569 3092
rect 12517 3041 12569 3080
rect 12581 3041 12633 3092
rect 12645 3080 12662 3092
rect 12662 3080 12696 3092
rect 12696 3080 12697 3093
rect 12645 3041 12697 3080
rect 12517 3004 12518 3028
rect 12518 3004 12552 3028
rect 12552 3004 12569 3028
rect 12517 2976 12569 3004
rect 12581 3004 12590 3028
rect 12590 3004 12624 3028
rect 12624 3004 12633 3028
rect 12581 2976 12633 3004
rect 12645 3004 12662 3028
rect 12662 3004 12696 3028
rect 12696 3004 12697 3028
rect 12645 2976 12697 3004
rect 12517 2955 12569 2963
rect 12517 2921 12518 2955
rect 12518 2921 12552 2955
rect 12552 2921 12569 2955
rect 12517 2911 12569 2921
rect 12581 2955 12633 2963
rect 12581 2921 12590 2955
rect 12590 2921 12624 2955
rect 12624 2921 12633 2955
rect 12581 2911 12633 2921
rect 12645 2955 12697 2963
rect 12645 2921 12662 2955
rect 12662 2921 12696 2955
rect 12696 2921 12697 2955
rect 12645 2911 12697 2921
rect 12517 2871 12569 2898
rect 12517 2846 12518 2871
rect 12518 2846 12552 2871
rect 12552 2846 12569 2871
rect 12581 2871 12633 2898
rect 12581 2846 12590 2871
rect 12590 2846 12624 2871
rect 12624 2846 12633 2871
rect 12645 2871 12697 2898
rect 12645 2846 12662 2871
rect 12662 2846 12696 2871
rect 12696 2846 12697 2871
rect 12517 2787 12569 2833
rect 12517 2781 12518 2787
rect 12518 2781 12552 2787
rect 12552 2781 12569 2787
rect 12581 2787 12633 2833
rect 12581 2781 12590 2787
rect 12590 2781 12624 2787
rect 12624 2781 12633 2787
rect 12645 2787 12697 2833
rect 12645 2781 12662 2787
rect 12662 2781 12696 2787
rect 12696 2781 12697 2787
rect 12517 2753 12518 2768
rect 12518 2753 12552 2768
rect 12552 2753 12569 2768
rect 12517 2716 12569 2753
rect 12581 2753 12590 2768
rect 12590 2753 12624 2768
rect 12624 2753 12633 2768
rect 12581 2716 12633 2753
rect 12645 2753 12662 2768
rect 12662 2753 12696 2768
rect 12696 2753 12697 2768
rect 12645 2716 12697 2753
rect 12517 2669 12518 2703
rect 12518 2669 12552 2703
rect 12552 2669 12569 2703
rect 12517 2651 12569 2669
rect 12581 2669 12590 2703
rect 12590 2669 12624 2703
rect 12624 2669 12633 2703
rect 12581 2651 12633 2669
rect 12645 2669 12662 2703
rect 12662 2669 12696 2703
rect 12696 2669 12697 2703
rect 12645 2651 12697 2669
rect 12517 2619 12569 2638
rect 12517 2586 12518 2619
rect 12518 2586 12552 2619
rect 12552 2586 12569 2619
rect 12581 2619 12633 2638
rect 12581 2586 12590 2619
rect 12590 2586 12624 2619
rect 12624 2586 12633 2619
rect 12645 2619 12697 2638
rect 12645 2586 12662 2619
rect 12662 2586 12696 2619
rect 12696 2586 12697 2619
rect 12517 2535 12569 2573
rect 12517 2521 12518 2535
rect 12518 2521 12552 2535
rect 12552 2521 12569 2535
rect 12581 2535 12633 2573
rect 12581 2521 12590 2535
rect 12590 2521 12624 2535
rect 12624 2521 12633 2535
rect 12645 2535 12697 2573
rect 12645 2521 12662 2535
rect 12662 2521 12696 2535
rect 12696 2521 12697 2535
rect 12517 2501 12518 2508
rect 12518 2501 12552 2508
rect 12552 2501 12569 2508
rect 12517 2456 12569 2501
rect 12581 2501 12590 2508
rect 12590 2501 12624 2508
rect 12624 2501 12633 2508
rect 12581 2461 12633 2501
rect 12581 2456 12590 2461
rect 12590 2456 12624 2461
rect 12624 2456 12633 2461
rect 12645 2501 12662 2508
rect 12662 2501 12696 2508
rect 12696 2501 12697 2508
rect 12645 2456 12697 2501
rect 12517 2391 12518 2443
rect 12518 2391 12569 2443
rect 12581 2391 12633 2443
rect 12645 2391 12696 2443
rect 12696 2391 12697 2443
rect 12517 2326 12518 2378
rect 12518 2326 12569 2378
rect 12581 2326 12633 2378
rect 12645 2326 12696 2378
rect 12696 2326 12697 2378
rect 12517 2261 12518 2313
rect 12518 2261 12569 2313
rect 12581 2261 12633 2313
rect 12645 2261 12696 2313
rect 12696 2261 12697 2313
rect 12517 2196 12518 2248
rect 12518 2196 12569 2248
rect 12581 2196 12633 2248
rect 12645 2196 12696 2248
rect 12696 2196 12697 2248
rect 12517 2131 12518 2183
rect 12518 2131 12569 2183
rect 12581 2131 12633 2183
rect 12645 2131 12696 2183
rect 12696 2131 12697 2183
rect 12517 2066 12518 2118
rect 12518 2066 12569 2118
rect 12581 2066 12633 2118
rect 12645 2066 12696 2118
rect 12696 2066 12697 2118
rect 12517 2001 12518 2053
rect 12518 2001 12569 2053
rect 12581 2001 12633 2053
rect 12645 2001 12696 2053
rect 12696 2001 12697 2053
rect 12517 1935 12518 1987
rect 12518 1935 12569 1987
rect 12581 1935 12633 1987
rect 12645 1935 12696 1987
rect 12696 1935 12697 1987
rect 12517 1869 12518 1921
rect 12518 1869 12569 1921
rect 12581 1869 12633 1921
rect 12645 1869 12696 1921
rect 12696 1869 12697 1921
rect 12517 1803 12518 1855
rect 12518 1803 12569 1855
rect 12581 1803 12633 1855
rect 12645 1803 12696 1855
rect 12696 1803 12697 1855
rect 12517 1737 12518 1789
rect 12518 1737 12569 1789
rect 12581 1737 12633 1789
rect 12645 1737 12696 1789
rect 12696 1737 12697 1789
rect 12517 1671 12518 1723
rect 12518 1671 12569 1723
rect 12581 1671 12633 1723
rect 12645 1671 12696 1723
rect 12696 1671 12697 1723
rect 12517 1605 12518 1657
rect 12518 1605 12569 1657
rect 12581 1605 12633 1657
rect 12645 1605 12696 1657
rect 12696 1605 12697 1657
rect 12517 1539 12518 1591
rect 12518 1539 12569 1591
rect 12581 1539 12633 1591
rect 12645 1539 12696 1591
rect 12696 1539 12697 1591
rect 12517 1479 12518 1525
rect 12518 1491 12569 1525
rect 12581 1491 12633 1525
rect 12645 1491 12696 1525
rect 12518 1479 12552 1491
rect 12552 1479 12569 1491
rect 12517 1473 12569 1479
rect 12581 1473 12633 1491
rect 12645 1479 12662 1491
rect 12662 1479 12696 1491
rect 12696 1479 12697 1525
rect 12645 1473 12697 1479
rect 13013 4062 13065 4068
rect 13013 4028 13014 4062
rect 13014 4028 13048 4062
rect 13048 4028 13065 4062
rect 13013 4016 13065 4028
rect 13077 4062 13129 4068
rect 13077 4028 13086 4062
rect 13086 4028 13120 4062
rect 13120 4028 13129 4062
rect 13077 4016 13129 4028
rect 13141 4062 13193 4068
rect 13141 4028 13158 4062
rect 13158 4028 13192 4062
rect 13192 4028 13193 4062
rect 13141 4016 13193 4028
rect 13013 3988 13065 4003
rect 13013 3954 13014 3988
rect 13014 3954 13048 3988
rect 13048 3954 13065 3988
rect 13013 3951 13065 3954
rect 13077 3988 13129 4003
rect 13077 3954 13086 3988
rect 13086 3954 13120 3988
rect 13120 3954 13129 3988
rect 13077 3951 13129 3954
rect 13141 3988 13193 4003
rect 13141 3954 13158 3988
rect 13158 3954 13192 3988
rect 13192 3954 13193 3988
rect 13141 3951 13193 3954
rect 13013 3914 13065 3938
rect 13013 3886 13014 3914
rect 13014 3886 13048 3914
rect 13048 3886 13065 3914
rect 13077 3914 13129 3938
rect 13077 3886 13086 3914
rect 13086 3886 13120 3914
rect 13120 3886 13129 3914
rect 13141 3914 13193 3938
rect 13141 3886 13158 3914
rect 13158 3886 13192 3914
rect 13192 3886 13193 3914
rect 13013 3840 13065 3873
rect 13013 3821 13014 3840
rect 13014 3821 13048 3840
rect 13048 3821 13065 3840
rect 13077 3840 13129 3873
rect 13077 3821 13086 3840
rect 13086 3821 13120 3840
rect 13120 3821 13129 3840
rect 13141 3840 13193 3873
rect 13141 3821 13158 3840
rect 13158 3821 13192 3840
rect 13192 3821 13193 3840
rect 13013 3806 13014 3808
rect 13014 3806 13048 3808
rect 13048 3806 13065 3808
rect 13013 3766 13065 3806
rect 13013 3756 13014 3766
rect 13014 3756 13048 3766
rect 13048 3756 13065 3766
rect 13077 3806 13086 3808
rect 13086 3806 13120 3808
rect 13120 3806 13129 3808
rect 13077 3766 13129 3806
rect 13077 3756 13086 3766
rect 13086 3756 13120 3766
rect 13120 3756 13129 3766
rect 13141 3806 13158 3808
rect 13158 3806 13192 3808
rect 13192 3806 13193 3808
rect 13141 3766 13193 3806
rect 13141 3756 13158 3766
rect 13158 3756 13192 3766
rect 13192 3756 13193 3766
rect 13013 3732 13014 3743
rect 13014 3732 13048 3743
rect 13048 3732 13065 3743
rect 13013 3692 13065 3732
rect 13013 3691 13014 3692
rect 13014 3691 13048 3692
rect 13048 3691 13065 3692
rect 13077 3732 13086 3743
rect 13086 3732 13120 3743
rect 13120 3732 13129 3743
rect 13077 3692 13129 3732
rect 13077 3691 13086 3692
rect 13086 3691 13120 3692
rect 13120 3691 13129 3692
rect 13141 3732 13158 3743
rect 13158 3732 13192 3743
rect 13192 3732 13193 3743
rect 13141 3692 13193 3732
rect 13141 3691 13158 3692
rect 13158 3691 13192 3692
rect 13192 3691 13193 3692
rect 13013 3658 13014 3678
rect 13014 3658 13048 3678
rect 13048 3658 13065 3678
rect 13013 3626 13065 3658
rect 13077 3658 13086 3678
rect 13086 3658 13120 3678
rect 13120 3658 13129 3678
rect 13077 3626 13129 3658
rect 13141 3658 13158 3678
rect 13158 3658 13192 3678
rect 13192 3658 13193 3678
rect 13141 3626 13193 3658
rect 13013 3584 13014 3613
rect 13014 3584 13048 3613
rect 13048 3584 13065 3613
rect 13013 3561 13065 3584
rect 13077 3584 13086 3613
rect 13086 3584 13120 3613
rect 13120 3584 13129 3613
rect 13077 3561 13129 3584
rect 13141 3584 13158 3613
rect 13158 3584 13192 3613
rect 13192 3584 13193 3613
rect 13141 3561 13193 3584
rect 13013 3544 13065 3548
rect 13013 3510 13014 3544
rect 13014 3510 13048 3544
rect 13048 3510 13065 3544
rect 13013 3496 13065 3510
rect 13077 3544 13129 3548
rect 13077 3510 13086 3544
rect 13086 3510 13120 3544
rect 13120 3510 13129 3544
rect 13077 3496 13129 3510
rect 13141 3544 13193 3548
rect 13141 3510 13158 3544
rect 13158 3510 13192 3544
rect 13192 3510 13193 3544
rect 13141 3496 13193 3510
rect 13013 3470 13065 3483
rect 13013 3436 13014 3470
rect 13014 3436 13048 3470
rect 13048 3436 13065 3470
rect 13013 3431 13065 3436
rect 13077 3470 13129 3483
rect 13077 3436 13086 3470
rect 13086 3436 13120 3470
rect 13120 3436 13129 3470
rect 13077 3431 13129 3436
rect 13141 3470 13193 3483
rect 13141 3436 13158 3470
rect 13158 3436 13192 3470
rect 13192 3436 13193 3470
rect 13141 3431 13193 3436
rect 13013 3396 13065 3418
rect 13013 3366 13014 3396
rect 13014 3366 13048 3396
rect 13048 3366 13065 3396
rect 13077 3396 13129 3418
rect 13077 3366 13086 3396
rect 13086 3366 13120 3396
rect 13120 3366 13129 3396
rect 13141 3396 13193 3418
rect 13141 3366 13158 3396
rect 13158 3366 13192 3396
rect 13192 3366 13193 3396
rect 13013 3322 13065 3353
rect 13013 3301 13014 3322
rect 13014 3301 13048 3322
rect 13048 3301 13065 3322
rect 13077 3322 13129 3353
rect 13077 3301 13086 3322
rect 13086 3301 13120 3322
rect 13120 3301 13129 3322
rect 13141 3322 13193 3353
rect 13141 3301 13158 3322
rect 13158 3301 13192 3322
rect 13192 3301 13193 3322
rect 13013 3248 13065 3288
rect 13013 3236 13014 3248
rect 13014 3236 13048 3248
rect 13048 3236 13065 3248
rect 13077 3248 13129 3288
rect 13077 3236 13086 3248
rect 13086 3236 13120 3248
rect 13120 3236 13129 3248
rect 13141 3248 13193 3288
rect 13141 3236 13158 3248
rect 13158 3236 13192 3248
rect 13192 3236 13193 3248
rect 13013 3214 13014 3223
rect 13014 3214 13048 3223
rect 13048 3214 13065 3223
rect 13013 3174 13065 3214
rect 13013 3171 13014 3174
rect 13014 3171 13048 3174
rect 13048 3171 13065 3174
rect 13077 3214 13086 3223
rect 13086 3214 13120 3223
rect 13120 3214 13129 3223
rect 13077 3174 13129 3214
rect 13077 3171 13086 3174
rect 13086 3171 13120 3174
rect 13120 3171 13129 3174
rect 13141 3214 13158 3223
rect 13158 3214 13192 3223
rect 13192 3214 13193 3223
rect 13141 3174 13193 3214
rect 13141 3171 13158 3174
rect 13158 3171 13192 3174
rect 13192 3171 13193 3174
rect 13013 3140 13014 3158
rect 13014 3140 13048 3158
rect 13048 3140 13065 3158
rect 13013 3106 13065 3140
rect 13077 3140 13086 3158
rect 13086 3140 13120 3158
rect 13120 3140 13129 3158
rect 13077 3106 13129 3140
rect 13141 3140 13158 3158
rect 13158 3140 13192 3158
rect 13192 3140 13193 3158
rect 13141 3106 13193 3140
rect 13013 3066 13014 3093
rect 13014 3066 13048 3093
rect 13048 3066 13065 3093
rect 13013 3041 13065 3066
rect 13077 3066 13086 3093
rect 13086 3066 13120 3093
rect 13120 3066 13129 3093
rect 13077 3041 13129 3066
rect 13141 3066 13158 3093
rect 13158 3066 13192 3093
rect 13192 3066 13193 3093
rect 13141 3041 13193 3066
rect 13013 3026 13065 3028
rect 13013 2992 13014 3026
rect 13014 2992 13048 3026
rect 13048 2992 13065 3026
rect 13013 2976 13065 2992
rect 13077 3026 13129 3028
rect 13077 2992 13086 3026
rect 13086 2992 13120 3026
rect 13120 2992 13129 3026
rect 13077 2976 13129 2992
rect 13141 3026 13193 3028
rect 13141 2992 13158 3026
rect 13158 2992 13192 3026
rect 13192 2992 13193 3026
rect 13141 2976 13193 2992
rect 13013 2952 13065 2963
rect 13013 2918 13014 2952
rect 13014 2918 13048 2952
rect 13048 2918 13065 2952
rect 13013 2911 13065 2918
rect 13077 2952 13129 2963
rect 13077 2918 13086 2952
rect 13086 2918 13120 2952
rect 13120 2918 13129 2952
rect 13077 2911 13129 2918
rect 13141 2952 13193 2963
rect 13141 2918 13158 2952
rect 13158 2918 13192 2952
rect 13192 2918 13193 2952
rect 13141 2911 13193 2918
rect 13013 2878 13065 2898
rect 13013 2846 13014 2878
rect 13014 2846 13048 2878
rect 13048 2846 13065 2878
rect 13077 2878 13129 2898
rect 13077 2846 13086 2878
rect 13086 2846 13120 2878
rect 13120 2846 13129 2878
rect 13141 2878 13193 2898
rect 13141 2846 13158 2878
rect 13158 2846 13192 2878
rect 13192 2846 13193 2878
rect 13013 2804 13065 2833
rect 13013 2781 13014 2804
rect 13014 2781 13048 2804
rect 13048 2781 13065 2804
rect 13077 2804 13129 2833
rect 13077 2781 13086 2804
rect 13086 2781 13120 2804
rect 13120 2781 13129 2804
rect 13141 2804 13193 2833
rect 13141 2781 13158 2804
rect 13158 2781 13192 2804
rect 13192 2781 13193 2804
rect 13013 2730 13065 2768
rect 13013 2716 13014 2730
rect 13014 2716 13048 2730
rect 13048 2716 13065 2730
rect 13077 2730 13129 2768
rect 13077 2716 13086 2730
rect 13086 2716 13120 2730
rect 13120 2716 13129 2730
rect 13141 2730 13193 2768
rect 13141 2716 13158 2730
rect 13158 2716 13192 2730
rect 13192 2716 13193 2730
rect 13013 2696 13014 2703
rect 13014 2696 13048 2703
rect 13048 2696 13065 2703
rect 13013 2656 13065 2696
rect 13013 2651 13014 2656
rect 13014 2651 13048 2656
rect 13048 2651 13065 2656
rect 13077 2696 13086 2703
rect 13086 2696 13120 2703
rect 13120 2696 13129 2703
rect 13077 2656 13129 2696
rect 13077 2651 13086 2656
rect 13086 2651 13120 2656
rect 13120 2651 13129 2656
rect 13141 2696 13158 2703
rect 13158 2696 13192 2703
rect 13192 2696 13193 2703
rect 13141 2656 13193 2696
rect 13141 2651 13158 2656
rect 13158 2651 13192 2656
rect 13192 2651 13193 2656
rect 13013 2622 13014 2638
rect 13014 2622 13048 2638
rect 13048 2622 13065 2638
rect 13013 2586 13065 2622
rect 13077 2622 13086 2638
rect 13086 2622 13120 2638
rect 13120 2622 13129 2638
rect 13077 2586 13129 2622
rect 13141 2622 13158 2638
rect 13158 2622 13192 2638
rect 13192 2622 13193 2638
rect 13141 2586 13193 2622
rect 13013 2548 13014 2573
rect 13014 2548 13048 2573
rect 13048 2548 13065 2573
rect 13013 2521 13065 2548
rect 13077 2548 13086 2573
rect 13086 2548 13120 2573
rect 13120 2548 13129 2573
rect 13077 2521 13129 2548
rect 13141 2548 13158 2573
rect 13158 2548 13192 2573
rect 13192 2548 13193 2573
rect 13141 2521 13193 2548
rect 13013 2474 13014 2508
rect 13014 2474 13048 2508
rect 13048 2474 13065 2508
rect 13013 2456 13065 2474
rect 13077 2474 13086 2508
rect 13086 2474 13120 2508
rect 13120 2474 13129 2508
rect 13077 2456 13129 2474
rect 13141 2474 13158 2508
rect 13158 2474 13192 2508
rect 13192 2474 13193 2508
rect 13141 2456 13193 2474
rect 13013 2434 13065 2443
rect 13013 2400 13014 2434
rect 13014 2400 13048 2434
rect 13048 2400 13065 2434
rect 13013 2391 13065 2400
rect 13077 2434 13129 2443
rect 13077 2400 13086 2434
rect 13086 2400 13120 2434
rect 13120 2400 13129 2434
rect 13077 2391 13129 2400
rect 13141 2434 13193 2443
rect 13141 2400 13158 2434
rect 13158 2400 13192 2434
rect 13192 2400 13193 2434
rect 13141 2391 13193 2400
rect 13013 2360 13065 2378
rect 13013 2326 13014 2360
rect 13014 2326 13048 2360
rect 13048 2326 13065 2360
rect 13077 2360 13129 2378
rect 13077 2326 13086 2360
rect 13086 2326 13120 2360
rect 13120 2326 13129 2360
rect 13141 2360 13193 2378
rect 13141 2326 13158 2360
rect 13158 2326 13192 2360
rect 13192 2326 13193 2360
rect 13013 2286 13065 2313
rect 13013 2261 13014 2286
rect 13014 2261 13048 2286
rect 13048 2261 13065 2286
rect 13077 2286 13129 2313
rect 13077 2261 13086 2286
rect 13086 2261 13120 2286
rect 13120 2261 13129 2286
rect 13141 2286 13193 2313
rect 13141 2261 13158 2286
rect 13158 2261 13192 2286
rect 13192 2261 13193 2286
rect 13013 2212 13065 2248
rect 13013 2196 13014 2212
rect 13014 2196 13048 2212
rect 13048 2196 13065 2212
rect 13077 2212 13129 2248
rect 13077 2196 13086 2212
rect 13086 2196 13120 2212
rect 13120 2196 13129 2212
rect 13141 2212 13193 2248
rect 13141 2196 13158 2212
rect 13158 2196 13192 2212
rect 13192 2196 13193 2212
rect 13013 2178 13014 2183
rect 13014 2178 13048 2183
rect 13048 2178 13065 2183
rect 13013 2138 13065 2178
rect 13013 2131 13014 2138
rect 13014 2131 13048 2138
rect 13048 2131 13065 2138
rect 13077 2178 13086 2183
rect 13086 2178 13120 2183
rect 13120 2178 13129 2183
rect 13077 2138 13129 2178
rect 13077 2131 13086 2138
rect 13086 2131 13120 2138
rect 13120 2131 13129 2138
rect 13141 2178 13158 2183
rect 13158 2178 13192 2183
rect 13192 2178 13193 2183
rect 13141 2138 13193 2178
rect 13141 2131 13158 2138
rect 13158 2131 13192 2138
rect 13192 2131 13193 2138
rect 13013 2104 13014 2118
rect 13014 2104 13048 2118
rect 13048 2104 13065 2118
rect 13013 2066 13065 2104
rect 13077 2104 13086 2118
rect 13086 2104 13120 2118
rect 13120 2104 13129 2118
rect 13077 2066 13129 2104
rect 13141 2104 13158 2118
rect 13158 2104 13192 2118
rect 13192 2104 13193 2118
rect 13141 2066 13193 2104
rect 13013 2030 13014 2053
rect 13014 2030 13048 2053
rect 13048 2030 13065 2053
rect 13013 2001 13065 2030
rect 13077 2030 13086 2053
rect 13086 2030 13120 2053
rect 13120 2030 13129 2053
rect 13077 2001 13129 2030
rect 13141 2030 13158 2053
rect 13158 2030 13192 2053
rect 13192 2030 13193 2053
rect 13141 2001 13193 2030
rect 13013 1956 13014 1987
rect 13014 1956 13048 1987
rect 13048 1956 13065 1987
rect 13013 1935 13065 1956
rect 13077 1956 13086 1987
rect 13086 1956 13120 1987
rect 13120 1956 13129 1987
rect 13077 1935 13129 1956
rect 13141 1956 13158 1987
rect 13158 1956 13192 1987
rect 13192 1956 13193 1987
rect 13141 1935 13193 1956
rect 13013 1916 13065 1921
rect 13013 1882 13014 1916
rect 13014 1882 13048 1916
rect 13048 1882 13065 1916
rect 13013 1869 13065 1882
rect 13077 1916 13129 1921
rect 13077 1882 13086 1916
rect 13086 1882 13120 1916
rect 13120 1882 13129 1916
rect 13077 1869 13129 1882
rect 13141 1916 13193 1921
rect 13141 1882 13158 1916
rect 13158 1882 13192 1916
rect 13192 1882 13193 1916
rect 13141 1869 13193 1882
rect 13013 1842 13065 1855
rect 13013 1808 13014 1842
rect 13014 1808 13048 1842
rect 13048 1808 13065 1842
rect 13013 1803 13065 1808
rect 13077 1842 13129 1855
rect 13077 1808 13086 1842
rect 13086 1808 13120 1842
rect 13120 1808 13129 1842
rect 13077 1803 13129 1808
rect 13141 1842 13193 1855
rect 13141 1808 13158 1842
rect 13158 1808 13192 1842
rect 13192 1808 13193 1842
rect 13141 1803 13193 1808
rect 13013 1768 13065 1789
rect 13013 1737 13014 1768
rect 13014 1737 13048 1768
rect 13048 1737 13065 1768
rect 13077 1768 13129 1789
rect 13077 1737 13086 1768
rect 13086 1737 13120 1768
rect 13120 1737 13129 1768
rect 13141 1768 13193 1789
rect 13141 1737 13158 1768
rect 13158 1737 13192 1768
rect 13192 1737 13193 1768
rect 13013 1694 13065 1723
rect 13013 1671 13014 1694
rect 13014 1671 13048 1694
rect 13048 1671 13065 1694
rect 13077 1694 13129 1723
rect 13077 1671 13086 1694
rect 13086 1671 13120 1694
rect 13120 1671 13129 1694
rect 13141 1694 13193 1723
rect 13141 1671 13158 1694
rect 13158 1671 13192 1694
rect 13192 1671 13193 1694
rect 13013 1620 13065 1657
rect 13013 1605 13014 1620
rect 13014 1605 13048 1620
rect 13048 1605 13065 1620
rect 13077 1620 13129 1657
rect 13077 1605 13086 1620
rect 13086 1605 13120 1620
rect 13120 1605 13129 1620
rect 13141 1620 13193 1657
rect 13141 1605 13158 1620
rect 13158 1605 13192 1620
rect 13192 1605 13193 1620
rect 13013 1586 13014 1591
rect 13014 1586 13048 1591
rect 13048 1586 13065 1591
rect 13013 1545 13065 1586
rect 13013 1539 13014 1545
rect 13014 1539 13048 1545
rect 13048 1539 13065 1545
rect 13077 1586 13086 1591
rect 13086 1586 13120 1591
rect 13120 1586 13129 1591
rect 13077 1545 13129 1586
rect 13077 1539 13086 1545
rect 13086 1539 13120 1545
rect 13120 1539 13129 1545
rect 13141 1586 13158 1591
rect 13158 1586 13192 1591
rect 13192 1586 13193 1591
rect 13141 1545 13193 1586
rect 13141 1539 13158 1545
rect 13158 1539 13192 1545
rect 13192 1539 13193 1545
rect 13013 1511 13014 1525
rect 13014 1511 13048 1525
rect 13048 1511 13065 1525
rect 13013 1473 13065 1511
rect 13077 1511 13086 1525
rect 13086 1511 13120 1525
rect 13120 1511 13129 1525
rect 13077 1473 13129 1511
rect 13141 1511 13158 1525
rect 13158 1511 13192 1525
rect 13192 1511 13193 1525
rect 13141 1473 13193 1511
rect 13509 4050 13561 4068
rect 13573 4062 13625 4068
rect 13573 4050 13582 4062
rect 13582 4050 13616 4062
rect 13616 4050 13625 4062
rect 13637 4050 13689 4068
rect 13509 4016 13510 4050
rect 13510 4016 13561 4050
rect 13573 4016 13625 4050
rect 13637 4016 13688 4050
rect 13688 4016 13689 4050
rect 13509 3951 13510 4003
rect 13510 3951 13561 4003
rect 13573 3951 13625 4003
rect 13637 3951 13688 4003
rect 13688 3951 13689 4003
rect 13509 3886 13510 3938
rect 13510 3886 13561 3938
rect 13573 3886 13625 3938
rect 13637 3886 13688 3938
rect 13688 3886 13689 3938
rect 13509 3821 13510 3873
rect 13510 3821 13561 3873
rect 13573 3821 13625 3873
rect 13637 3821 13688 3873
rect 13688 3821 13689 3873
rect 13509 3756 13510 3808
rect 13510 3756 13561 3808
rect 13573 3756 13625 3808
rect 13637 3756 13688 3808
rect 13688 3756 13689 3808
rect 13509 3691 13510 3743
rect 13510 3691 13561 3743
rect 13573 3691 13625 3743
rect 13637 3691 13688 3743
rect 13688 3691 13689 3743
rect 13509 3626 13510 3678
rect 13510 3626 13561 3678
rect 13573 3626 13625 3678
rect 13637 3626 13688 3678
rect 13688 3626 13689 3678
rect 13509 3561 13510 3613
rect 13510 3561 13561 3613
rect 13573 3561 13625 3613
rect 13637 3561 13688 3613
rect 13688 3561 13689 3613
rect 13509 3496 13510 3548
rect 13510 3496 13561 3548
rect 13573 3496 13625 3548
rect 13637 3496 13688 3548
rect 13688 3496 13689 3548
rect 13509 3431 13510 3483
rect 13510 3431 13561 3483
rect 13573 3431 13625 3483
rect 13637 3431 13688 3483
rect 13688 3431 13689 3483
rect 13509 3366 13510 3418
rect 13510 3366 13561 3418
rect 13573 3366 13625 3418
rect 13637 3366 13688 3418
rect 13688 3366 13689 3418
rect 13509 3301 13510 3353
rect 13510 3301 13561 3353
rect 13573 3301 13625 3353
rect 13637 3301 13688 3353
rect 13688 3301 13689 3353
rect 13509 3236 13510 3288
rect 13510 3236 13561 3288
rect 13573 3236 13625 3288
rect 13637 3236 13688 3288
rect 13688 3236 13689 3288
rect 13509 3171 13510 3223
rect 13510 3171 13561 3223
rect 13573 3171 13625 3223
rect 13637 3171 13688 3223
rect 13688 3171 13689 3223
rect 13509 3106 13510 3158
rect 13510 3106 13561 3158
rect 13573 3106 13625 3158
rect 13637 3106 13688 3158
rect 13688 3106 13689 3158
rect 13509 3080 13510 3093
rect 13510 3092 13561 3093
rect 13573 3092 13625 3093
rect 13637 3092 13688 3093
rect 13510 3080 13544 3092
rect 13544 3080 13561 3092
rect 13509 3041 13561 3080
rect 13573 3041 13625 3092
rect 13637 3080 13654 3092
rect 13654 3080 13688 3092
rect 13688 3080 13689 3093
rect 13637 3041 13689 3080
rect 13509 2976 13510 3028
rect 13510 2976 13561 3028
rect 13573 2976 13625 3028
rect 13637 2976 13688 3028
rect 13688 2976 13689 3028
rect 13509 2911 13510 2963
rect 13510 2911 13561 2963
rect 13573 2911 13625 2963
rect 13637 2911 13688 2963
rect 13688 2911 13689 2963
rect 13509 2846 13510 2898
rect 13510 2846 13561 2898
rect 13573 2846 13625 2898
rect 13637 2846 13688 2898
rect 13688 2846 13689 2898
rect 13509 2781 13510 2833
rect 13510 2781 13561 2833
rect 13573 2781 13625 2833
rect 13637 2781 13688 2833
rect 13688 2781 13689 2833
rect 13509 2716 13510 2768
rect 13510 2716 13561 2768
rect 13573 2716 13625 2768
rect 13637 2716 13688 2768
rect 13688 2716 13689 2768
rect 13509 2651 13510 2703
rect 13510 2651 13561 2703
rect 13573 2651 13625 2703
rect 13637 2651 13688 2703
rect 13688 2651 13689 2703
rect 13509 2586 13510 2638
rect 13510 2586 13561 2638
rect 13573 2586 13625 2638
rect 13637 2586 13688 2638
rect 13688 2586 13689 2638
rect 13509 2535 13561 2573
rect 13509 2521 13510 2535
rect 13510 2521 13544 2535
rect 13544 2521 13561 2535
rect 13573 2535 13625 2573
rect 13573 2521 13582 2535
rect 13582 2521 13616 2535
rect 13616 2521 13625 2535
rect 13637 2535 13689 2573
rect 13637 2521 13654 2535
rect 13654 2521 13688 2535
rect 13688 2521 13689 2535
rect 13509 2501 13510 2508
rect 13510 2501 13544 2508
rect 13544 2501 13561 2508
rect 13509 2456 13561 2501
rect 13573 2501 13582 2508
rect 13582 2501 13616 2508
rect 13616 2501 13625 2508
rect 13573 2461 13625 2501
rect 13573 2456 13582 2461
rect 13582 2456 13616 2461
rect 13616 2456 13625 2461
rect 13637 2501 13654 2508
rect 13654 2501 13688 2508
rect 13688 2501 13689 2508
rect 13637 2456 13689 2501
rect 13509 2391 13510 2443
rect 13510 2391 13561 2443
rect 13573 2391 13625 2443
rect 13637 2391 13688 2443
rect 13688 2391 13689 2443
rect 13509 2326 13510 2378
rect 13510 2326 13561 2378
rect 13573 2326 13625 2378
rect 13637 2326 13688 2378
rect 13688 2326 13689 2378
rect 13509 2261 13510 2313
rect 13510 2261 13561 2313
rect 13573 2261 13625 2313
rect 13637 2261 13688 2313
rect 13688 2261 13689 2313
rect 13509 2196 13510 2248
rect 13510 2196 13561 2248
rect 13573 2196 13625 2248
rect 13637 2196 13688 2248
rect 13688 2196 13689 2248
rect 13509 2131 13510 2183
rect 13510 2131 13561 2183
rect 13573 2131 13625 2183
rect 13637 2131 13688 2183
rect 13688 2131 13689 2183
rect 13509 2066 13510 2118
rect 13510 2066 13561 2118
rect 13573 2066 13625 2118
rect 13637 2066 13688 2118
rect 13688 2066 13689 2118
rect 13509 2001 13510 2053
rect 13510 2001 13561 2053
rect 13573 2001 13625 2053
rect 13637 2001 13688 2053
rect 13688 2001 13689 2053
rect 13509 1935 13510 1987
rect 13510 1935 13561 1987
rect 13573 1935 13625 1987
rect 13637 1935 13688 1987
rect 13688 1935 13689 1987
rect 13509 1869 13510 1921
rect 13510 1869 13561 1921
rect 13573 1869 13625 1921
rect 13637 1869 13688 1921
rect 13688 1869 13689 1921
rect 13509 1803 13510 1855
rect 13510 1803 13561 1855
rect 13573 1803 13625 1855
rect 13637 1803 13688 1855
rect 13688 1803 13689 1855
rect 13509 1737 13510 1789
rect 13510 1737 13561 1789
rect 13573 1737 13625 1789
rect 13637 1737 13688 1789
rect 13688 1737 13689 1789
rect 13509 1671 13510 1723
rect 13510 1671 13561 1723
rect 13573 1671 13625 1723
rect 13637 1671 13688 1723
rect 13688 1671 13689 1723
rect 13509 1605 13510 1657
rect 13510 1605 13561 1657
rect 13573 1605 13625 1657
rect 13637 1605 13688 1657
rect 13688 1605 13689 1657
rect 13509 1539 13510 1591
rect 13510 1539 13561 1591
rect 13573 1539 13625 1591
rect 13637 1539 13688 1591
rect 13688 1539 13689 1591
rect 13509 1479 13510 1525
rect 13510 1491 13561 1525
rect 13573 1491 13625 1525
rect 13637 1491 13688 1525
rect 13510 1479 13544 1491
rect 13544 1479 13561 1491
rect 13509 1473 13561 1479
rect 13573 1473 13625 1491
rect 13637 1479 13654 1491
rect 13654 1479 13688 1491
rect 13688 1479 13689 1525
rect 13637 1473 13689 1479
rect 14037 4062 14089 4068
rect 14105 4062 14157 4068
rect 14037 4016 14089 4062
rect 14105 4016 14112 4062
rect 14112 4016 14157 4062
rect 14173 4016 14225 4068
rect 14037 3951 14089 4003
rect 14105 3951 14112 4003
rect 14112 3951 14157 4003
rect 14173 3951 14225 4003
rect 14037 3886 14089 3938
rect 14105 3886 14112 3938
rect 14112 3886 14157 3938
rect 14173 3886 14225 3938
rect 14037 3821 14089 3873
rect 14105 3821 14112 3873
rect 14112 3821 14157 3873
rect 14173 3821 14225 3873
rect 14037 3756 14089 3808
rect 14105 3756 14112 3808
rect 14112 3756 14157 3808
rect 14173 3756 14225 3808
rect 14037 3691 14089 3743
rect 14105 3691 14112 3743
rect 14112 3691 14157 3743
rect 14173 3691 14225 3743
rect 14037 3626 14089 3678
rect 14105 3626 14112 3678
rect 14112 3626 14157 3678
rect 14173 3626 14225 3678
rect 14037 3561 14089 3613
rect 14105 3561 14112 3613
rect 14112 3561 14157 3613
rect 14173 3561 14225 3613
rect 14037 3496 14089 3548
rect 14105 3496 14112 3548
rect 14112 3496 14157 3548
rect 14173 3496 14225 3548
rect 14037 3431 14089 3483
rect 14105 3431 14112 3483
rect 14112 3431 14157 3483
rect 14173 3431 14225 3483
rect 14037 3366 14089 3418
rect 14105 3366 14112 3418
rect 14112 3366 14157 3418
rect 14173 3366 14225 3418
rect 14037 3301 14089 3353
rect 14105 3301 14112 3353
rect 14112 3301 14157 3353
rect 14173 3301 14225 3353
rect 14037 3236 14089 3288
rect 14105 3236 14112 3288
rect 14112 3236 14157 3288
rect 14173 3236 14225 3288
rect 14037 3171 14089 3223
rect 14105 3171 14112 3223
rect 14112 3171 14157 3223
rect 14173 3171 14225 3223
rect 14037 3106 14089 3158
rect 14105 3106 14112 3158
rect 14112 3106 14157 3158
rect 14173 3106 14225 3158
rect 14037 3041 14089 3093
rect 14105 3041 14112 3093
rect 14112 3041 14157 3093
rect 14173 3041 14225 3093
rect 14037 2976 14089 3028
rect 14105 2976 14112 3028
rect 14112 2976 14157 3028
rect 14173 2976 14225 3028
rect 14037 2911 14089 2963
rect 14105 2911 14112 2963
rect 14112 2911 14157 2963
rect 14173 2911 14225 2963
rect 14037 2846 14089 2898
rect 14105 2846 14112 2898
rect 14112 2846 14157 2898
rect 14173 2846 14225 2898
rect 14037 2781 14089 2833
rect 14105 2781 14112 2833
rect 14112 2781 14157 2833
rect 14173 2781 14225 2833
rect 14037 2732 14089 2768
rect 14105 2732 14112 2768
rect 14112 2732 14157 2768
rect 14037 2716 14089 2732
rect 14105 2716 14157 2732
rect 14173 2716 14225 2768
rect 14037 2693 14089 2703
rect 14105 2693 14157 2703
rect 14037 2659 14040 2693
rect 14040 2659 14078 2693
rect 14078 2659 14089 2693
rect 14105 2659 14112 2693
rect 14112 2659 14157 2693
rect 14037 2651 14089 2659
rect 14105 2651 14157 2659
rect 14173 2651 14225 2703
rect 14037 2620 14089 2638
rect 14105 2620 14157 2638
rect 14037 2586 14040 2620
rect 14040 2586 14078 2620
rect 14078 2586 14089 2620
rect 14105 2586 14112 2620
rect 14112 2586 14157 2620
rect 14173 2586 14225 2638
rect 14037 2547 14089 2573
rect 14105 2547 14157 2573
rect 14037 2521 14040 2547
rect 14040 2521 14078 2547
rect 14078 2521 14089 2547
rect 14105 2521 14112 2547
rect 14112 2521 14157 2547
rect 14173 2521 14225 2573
rect 14037 2474 14089 2508
rect 14105 2474 14157 2508
rect 14037 2456 14040 2474
rect 14040 2456 14078 2474
rect 14078 2456 14089 2474
rect 14105 2456 14112 2474
rect 14112 2456 14157 2474
rect 14173 2456 14225 2508
rect 14037 2440 14040 2443
rect 14040 2440 14078 2443
rect 14078 2440 14089 2443
rect 14105 2440 14112 2443
rect 14112 2440 14157 2443
rect 14037 2401 14089 2440
rect 14105 2401 14157 2440
rect 14037 2391 14040 2401
rect 14040 2391 14078 2401
rect 14078 2391 14089 2401
rect 14105 2391 14112 2401
rect 14112 2391 14157 2401
rect 14173 2391 14225 2443
rect 14037 2367 14040 2378
rect 14040 2367 14078 2378
rect 14078 2367 14089 2378
rect 14105 2367 14112 2378
rect 14112 2367 14157 2378
rect 14037 2328 14089 2367
rect 14105 2328 14157 2367
rect 14037 2326 14040 2328
rect 14040 2326 14078 2328
rect 14078 2326 14089 2328
rect 14105 2326 14112 2328
rect 14112 2326 14157 2328
rect 14173 2326 14225 2378
rect 14037 2294 14040 2313
rect 14040 2294 14078 2313
rect 14078 2294 14089 2313
rect 14105 2294 14112 2313
rect 14112 2294 14157 2313
rect 14037 2261 14089 2294
rect 14105 2261 14157 2294
rect 14173 2261 14225 2313
rect 14037 2221 14040 2248
rect 14040 2221 14078 2248
rect 14078 2221 14089 2248
rect 14105 2221 14112 2248
rect 14112 2221 14157 2248
rect 14037 2196 14089 2221
rect 14105 2196 14157 2221
rect 14173 2196 14225 2248
rect 14037 2182 14089 2183
rect 14105 2182 14157 2183
rect 14037 2148 14040 2182
rect 14040 2148 14078 2182
rect 14078 2148 14089 2182
rect 14105 2148 14112 2182
rect 14112 2148 14157 2182
rect 14037 2131 14089 2148
rect 14105 2131 14157 2148
rect 14173 2131 14225 2183
rect 14037 2109 14089 2118
rect 14105 2109 14157 2118
rect 14037 2075 14040 2109
rect 14040 2075 14078 2109
rect 14078 2075 14089 2109
rect 14105 2075 14112 2109
rect 14112 2075 14157 2109
rect 14037 2066 14089 2075
rect 14105 2066 14157 2075
rect 14173 2066 14225 2118
rect 14037 2036 14089 2053
rect 14105 2036 14157 2053
rect 14037 2002 14040 2036
rect 14040 2002 14078 2036
rect 14078 2002 14089 2036
rect 14105 2002 14112 2036
rect 14112 2002 14157 2036
rect 14037 2001 14089 2002
rect 14105 2001 14157 2002
rect 14173 2001 14225 2053
rect 14037 1963 14089 1987
rect 14105 1963 14157 1987
rect 14037 1935 14040 1963
rect 14040 1935 14078 1963
rect 14078 1935 14089 1963
rect 14105 1935 14112 1963
rect 14112 1935 14157 1963
rect 14173 1935 14225 1987
rect 14037 1890 14089 1921
rect 14105 1890 14157 1921
rect 14037 1869 14040 1890
rect 14040 1869 14078 1890
rect 14078 1869 14089 1890
rect 14105 1869 14112 1890
rect 14112 1869 14157 1890
rect 14173 1869 14225 1921
rect 14037 1817 14089 1855
rect 14105 1817 14157 1855
rect 14037 1803 14040 1817
rect 14040 1803 14078 1817
rect 14078 1803 14089 1817
rect 14105 1803 14112 1817
rect 14112 1803 14157 1817
rect 14173 1803 14225 1855
rect 14037 1783 14040 1789
rect 14040 1783 14078 1789
rect 14078 1783 14089 1789
rect 14105 1783 14112 1789
rect 14112 1783 14157 1789
rect 14037 1744 14089 1783
rect 14105 1744 14157 1783
rect 14037 1737 14040 1744
rect 14040 1737 14078 1744
rect 14078 1737 14089 1744
rect 14105 1737 14112 1744
rect 14112 1737 14157 1744
rect 14173 1737 14225 1789
rect 14037 1710 14040 1723
rect 14040 1710 14078 1723
rect 14078 1710 14089 1723
rect 14105 1710 14112 1723
rect 14112 1710 14157 1723
rect 14037 1671 14089 1710
rect 14105 1671 14157 1710
rect 14173 1671 14225 1723
rect 14037 1637 14040 1657
rect 14040 1637 14078 1657
rect 14078 1637 14089 1657
rect 14105 1637 14112 1657
rect 14112 1637 14157 1657
rect 14037 1605 14089 1637
rect 14105 1605 14157 1637
rect 14173 1605 14225 1657
rect 14037 1564 14040 1591
rect 14040 1564 14078 1591
rect 14078 1564 14089 1591
rect 14105 1564 14112 1591
rect 14112 1564 14157 1591
rect 14037 1539 14089 1564
rect 14105 1539 14157 1564
rect 14173 1539 14225 1591
rect 14037 1491 14040 1525
rect 14040 1491 14078 1525
rect 14078 1491 14089 1525
rect 14105 1491 14112 1525
rect 14112 1491 14157 1525
rect 14037 1473 14089 1491
rect 14105 1473 14157 1491
rect 14173 1473 14225 1525
rect 14400 4044 14452 4068
rect 14488 4052 14510 4068
rect 14510 4052 14540 4068
rect 14576 4052 14582 4068
rect 14582 4052 14616 4068
rect 14616 4052 14628 4068
rect 14400 4016 14431 4044
rect 14431 4016 14452 4044
rect 14488 4016 14540 4052
rect 14576 4016 14628 4052
rect 14400 3971 14452 4003
rect 14488 3979 14510 4003
rect 14510 3979 14540 4003
rect 14576 3979 14582 4003
rect 14582 3979 14616 4003
rect 14616 3979 14628 4003
rect 14400 3951 14431 3971
rect 14431 3951 14452 3971
rect 14488 3951 14540 3979
rect 14576 3951 14628 3979
rect 14400 3937 14431 3938
rect 14431 3937 14452 3938
rect 14400 3898 14452 3937
rect 14488 3906 14510 3938
rect 14510 3906 14540 3938
rect 14576 3906 14582 3938
rect 14582 3906 14616 3938
rect 14616 3906 14628 3938
rect 14400 3886 14431 3898
rect 14431 3886 14452 3898
rect 14488 3886 14540 3906
rect 14576 3886 14628 3906
rect 14400 3864 14431 3873
rect 14431 3864 14452 3873
rect 14488 3867 14540 3873
rect 14576 3867 14628 3873
rect 14400 3825 14452 3864
rect 14488 3833 14510 3867
rect 14510 3833 14540 3867
rect 14576 3833 14582 3867
rect 14582 3833 14616 3867
rect 14616 3833 14628 3867
rect 14400 3821 14431 3825
rect 14431 3821 14452 3825
rect 14488 3821 14540 3833
rect 14576 3821 14628 3833
rect 14400 3791 14431 3808
rect 14431 3791 14452 3808
rect 14488 3794 14540 3808
rect 14576 3794 14628 3808
rect 14400 3756 14452 3791
rect 14488 3760 14510 3794
rect 14510 3760 14540 3794
rect 14576 3760 14582 3794
rect 14582 3760 14616 3794
rect 14616 3760 14628 3794
rect 14488 3756 14540 3760
rect 14576 3756 14628 3760
rect 14400 3718 14431 3743
rect 14431 3718 14452 3743
rect 14488 3721 14540 3743
rect 14576 3721 14628 3743
rect 14400 3691 14452 3718
rect 14488 3691 14510 3721
rect 14510 3691 14540 3721
rect 14576 3691 14582 3721
rect 14582 3691 14616 3721
rect 14616 3691 14628 3721
rect 14400 3645 14431 3678
rect 14431 3645 14452 3678
rect 14488 3648 14540 3678
rect 14576 3648 14628 3678
rect 14400 3626 14452 3645
rect 14488 3626 14510 3648
rect 14510 3626 14540 3648
rect 14576 3626 14582 3648
rect 14582 3626 14616 3648
rect 14616 3626 14628 3648
rect 14400 3606 14452 3613
rect 14400 3572 14431 3606
rect 14431 3572 14452 3606
rect 14488 3575 14540 3613
rect 14576 3575 14628 3613
rect 14400 3561 14452 3572
rect 14488 3561 14510 3575
rect 14510 3561 14540 3575
rect 14576 3561 14582 3575
rect 14582 3561 14616 3575
rect 14616 3561 14628 3575
rect 14400 3533 14452 3548
rect 14488 3541 14510 3548
rect 14510 3541 14540 3548
rect 14576 3541 14582 3548
rect 14582 3541 14616 3548
rect 14616 3541 14628 3548
rect 14400 3499 14431 3533
rect 14431 3499 14452 3533
rect 14488 3502 14540 3541
rect 14576 3502 14628 3541
rect 14400 3496 14452 3499
rect 14488 3496 14510 3502
rect 14510 3496 14540 3502
rect 14576 3496 14582 3502
rect 14582 3496 14616 3502
rect 14616 3496 14628 3502
rect 14400 3460 14452 3483
rect 14488 3468 14510 3483
rect 14510 3468 14540 3483
rect 14576 3468 14582 3483
rect 14582 3468 14616 3483
rect 14616 3468 14628 3483
rect 14400 3431 14431 3460
rect 14431 3431 14452 3460
rect 14488 3431 14540 3468
rect 14576 3431 14628 3468
rect 14400 3387 14452 3418
rect 14488 3395 14510 3418
rect 14510 3395 14540 3418
rect 14576 3395 14582 3418
rect 14582 3395 14616 3418
rect 14616 3395 14628 3418
rect 14400 3366 14431 3387
rect 14431 3366 14452 3387
rect 14488 3366 14540 3395
rect 14576 3366 14628 3395
rect 14400 3314 14452 3353
rect 14488 3322 14510 3353
rect 14510 3322 14540 3353
rect 14576 3322 14582 3353
rect 14582 3322 14616 3353
rect 14616 3322 14628 3353
rect 14400 3301 14431 3314
rect 14431 3301 14452 3314
rect 14488 3301 14540 3322
rect 14576 3301 14628 3322
rect 14400 3280 14431 3288
rect 14431 3280 14452 3288
rect 14488 3283 14540 3288
rect 14576 3283 14628 3288
rect 14400 3241 14452 3280
rect 14488 3249 14510 3283
rect 14510 3249 14540 3283
rect 14576 3249 14582 3283
rect 14582 3249 14616 3283
rect 14616 3249 14628 3283
rect 14400 3236 14431 3241
rect 14431 3236 14452 3241
rect 14488 3236 14540 3249
rect 14576 3236 14628 3249
rect 14400 3207 14431 3223
rect 14431 3207 14452 3223
rect 14488 3210 14540 3223
rect 14576 3210 14628 3223
rect 14400 3171 14452 3207
rect 14488 3176 14510 3210
rect 14510 3176 14540 3210
rect 14576 3176 14582 3210
rect 14582 3176 14616 3210
rect 14616 3176 14628 3210
rect 14488 3171 14540 3176
rect 14576 3171 14628 3176
rect 14400 3134 14431 3158
rect 14431 3134 14452 3158
rect 14488 3137 14540 3158
rect 14576 3137 14628 3158
rect 14400 3106 14452 3134
rect 14488 3106 14510 3137
rect 14510 3106 14540 3137
rect 14576 3106 14582 3137
rect 14582 3106 14616 3137
rect 14616 3106 14628 3137
rect 14400 3061 14431 3093
rect 14431 3061 14452 3093
rect 14488 3064 14540 3093
rect 14576 3064 14628 3093
rect 14400 3041 14452 3061
rect 14488 3041 14510 3064
rect 14510 3041 14540 3064
rect 14576 3041 14582 3064
rect 14582 3041 14616 3064
rect 14616 3041 14628 3064
rect 14400 3022 14452 3028
rect 14400 2988 14431 3022
rect 14431 2988 14452 3022
rect 14488 2991 14540 3028
rect 14576 2991 14628 3028
rect 14400 2976 14452 2988
rect 14488 2976 14510 2991
rect 14510 2976 14540 2991
rect 14576 2976 14582 2991
rect 14582 2976 14616 2991
rect 14616 2976 14628 2991
rect 14400 2949 14452 2963
rect 14488 2957 14510 2963
rect 14510 2957 14540 2963
rect 14576 2957 14582 2963
rect 14582 2957 14616 2963
rect 14616 2957 14628 2963
rect 14400 2915 14431 2949
rect 14431 2915 14452 2949
rect 14488 2918 14540 2957
rect 14576 2918 14628 2957
rect 14400 2911 14452 2915
rect 14488 2911 14510 2918
rect 14510 2911 14540 2918
rect 14576 2911 14582 2918
rect 14582 2911 14616 2918
rect 14616 2911 14628 2918
rect 14400 2876 14452 2898
rect 14488 2884 14510 2898
rect 14510 2884 14540 2898
rect 14576 2884 14582 2898
rect 14582 2884 14616 2898
rect 14616 2884 14628 2898
rect 14400 2846 14431 2876
rect 14431 2846 14452 2876
rect 14488 2846 14540 2884
rect 14576 2846 14628 2884
rect 14400 2803 14452 2833
rect 14488 2811 14510 2833
rect 14510 2811 14540 2833
rect 14576 2811 14582 2833
rect 14582 2811 14616 2833
rect 14616 2811 14628 2833
rect 14400 2781 14431 2803
rect 14431 2781 14452 2803
rect 14488 2781 14540 2811
rect 14576 2781 14628 2811
rect 14400 2730 14452 2768
rect 14488 2738 14510 2768
rect 14510 2738 14540 2768
rect 14576 2738 14582 2768
rect 14582 2738 14616 2768
rect 14616 2738 14628 2768
rect 14400 2716 14431 2730
rect 14431 2716 14452 2730
rect 14488 2716 14540 2738
rect 14576 2716 14628 2738
rect 14400 2696 14431 2703
rect 14431 2696 14452 2703
rect 14488 2699 14540 2703
rect 14576 2699 14628 2703
rect 14400 2657 14452 2696
rect 14488 2665 14510 2699
rect 14510 2665 14540 2699
rect 14576 2665 14582 2699
rect 14582 2665 14616 2699
rect 14616 2665 14628 2699
rect 14400 2651 14431 2657
rect 14431 2651 14452 2657
rect 14488 2651 14540 2665
rect 14576 2651 14628 2665
rect 14400 2623 14431 2638
rect 14431 2623 14452 2638
rect 14488 2626 14540 2638
rect 14576 2626 14628 2638
rect 14400 2586 14452 2623
rect 14488 2592 14510 2626
rect 14510 2592 14540 2626
rect 14576 2592 14582 2626
rect 14582 2592 14616 2626
rect 14616 2592 14628 2626
rect 14488 2586 14540 2592
rect 14576 2586 14628 2592
rect 14400 2550 14431 2573
rect 14431 2550 14452 2573
rect 14488 2553 14540 2573
rect 14576 2553 14628 2573
rect 14400 2521 14452 2550
rect 14488 2521 14510 2553
rect 14510 2521 14540 2553
rect 14576 2521 14582 2553
rect 14582 2521 14616 2553
rect 14616 2521 14628 2553
rect 14400 2477 14431 2508
rect 14431 2477 14452 2508
rect 14488 2480 14540 2508
rect 14576 2480 14628 2508
rect 14400 2456 14452 2477
rect 14488 2456 14510 2480
rect 14510 2456 14540 2480
rect 14576 2456 14582 2480
rect 14582 2456 14616 2480
rect 14616 2456 14628 2480
rect 14400 2438 14452 2443
rect 14400 2404 14431 2438
rect 14431 2404 14452 2438
rect 14488 2407 14540 2443
rect 14576 2407 14628 2443
rect 14400 2391 14452 2404
rect 14488 2391 14510 2407
rect 14510 2391 14540 2407
rect 14576 2391 14582 2407
rect 14582 2391 14616 2407
rect 14616 2391 14628 2407
rect 14400 2365 14452 2378
rect 14488 2373 14510 2378
rect 14510 2373 14540 2378
rect 14576 2373 14582 2378
rect 14582 2373 14616 2378
rect 14616 2373 14628 2378
rect 14400 2331 14431 2365
rect 14431 2331 14452 2365
rect 14488 2334 14540 2373
rect 14576 2334 14628 2373
rect 14400 2326 14452 2331
rect 14488 2326 14510 2334
rect 14510 2326 14540 2334
rect 14576 2326 14582 2334
rect 14582 2326 14616 2334
rect 14616 2326 14628 2334
rect 14400 2292 14452 2313
rect 14488 2300 14510 2313
rect 14510 2300 14540 2313
rect 14576 2300 14582 2313
rect 14582 2300 14616 2313
rect 14616 2300 14628 2313
rect 14400 2261 14431 2292
rect 14431 2261 14452 2292
rect 14488 2261 14540 2300
rect 14576 2261 14628 2300
rect 14400 2219 14452 2248
rect 14488 2226 14510 2248
rect 14510 2226 14540 2248
rect 14576 2226 14582 2248
rect 14582 2226 14616 2248
rect 14616 2226 14628 2248
rect 14400 2196 14431 2219
rect 14431 2196 14452 2219
rect 14488 2196 14540 2226
rect 14576 2196 14628 2226
rect 14400 2146 14452 2183
rect 14488 2152 14510 2183
rect 14510 2152 14540 2183
rect 14576 2152 14582 2183
rect 14582 2152 14616 2183
rect 14616 2152 14628 2183
rect 14400 2131 14431 2146
rect 14431 2131 14452 2146
rect 14488 2131 14540 2152
rect 14576 2131 14628 2152
rect 14400 2112 14431 2118
rect 14431 2112 14452 2118
rect 14488 2112 14540 2118
rect 14576 2112 14628 2118
rect 14400 2073 14452 2112
rect 14488 2078 14510 2112
rect 14510 2078 14540 2112
rect 14576 2078 14582 2112
rect 14582 2078 14616 2112
rect 14616 2078 14628 2112
rect 14400 2066 14431 2073
rect 14431 2066 14452 2073
rect 14488 2066 14540 2078
rect 14576 2066 14628 2078
rect 14400 2039 14431 2053
rect 14431 2039 14452 2053
rect 14400 2001 14452 2039
rect 14488 2038 14540 2053
rect 14576 2038 14628 2053
rect 14488 2004 14510 2038
rect 14510 2004 14540 2038
rect 14576 2004 14582 2038
rect 14582 2004 14616 2038
rect 14616 2004 14628 2038
rect 14488 2001 14540 2004
rect 14576 2001 14628 2004
rect 14400 1966 14431 1987
rect 14431 1966 14452 1987
rect 14400 1935 14452 1966
rect 14488 1964 14540 1987
rect 14576 1964 14628 1987
rect 14488 1935 14510 1964
rect 14510 1935 14540 1964
rect 14576 1935 14582 1964
rect 14582 1935 14616 1964
rect 14616 1935 14628 1964
rect 14400 1893 14431 1921
rect 14431 1893 14452 1921
rect 14400 1869 14452 1893
rect 14488 1890 14540 1921
rect 14576 1890 14628 1921
rect 14488 1869 14510 1890
rect 14510 1869 14540 1890
rect 14576 1869 14582 1890
rect 14582 1869 14616 1890
rect 14616 1869 14628 1890
rect 14400 1854 14452 1855
rect 14400 1820 14431 1854
rect 14431 1820 14452 1854
rect 14400 1803 14452 1820
rect 14488 1816 14540 1855
rect 14576 1816 14628 1855
rect 14488 1803 14510 1816
rect 14510 1803 14540 1816
rect 14576 1803 14582 1816
rect 14582 1803 14616 1816
rect 14616 1803 14628 1816
rect 14400 1781 14452 1789
rect 14488 1782 14510 1789
rect 14510 1782 14540 1789
rect 14576 1782 14582 1789
rect 14582 1782 14616 1789
rect 14616 1782 14628 1789
rect 14400 1747 14431 1781
rect 14431 1747 14452 1781
rect 14400 1737 14452 1747
rect 14488 1742 14540 1782
rect 14576 1742 14628 1782
rect 14488 1737 14510 1742
rect 14510 1737 14540 1742
rect 14576 1737 14582 1742
rect 14582 1737 14616 1742
rect 14616 1737 14628 1742
rect 14400 1708 14452 1723
rect 14488 1708 14510 1723
rect 14510 1708 14540 1723
rect 14576 1708 14582 1723
rect 14582 1708 14616 1723
rect 14616 1708 14628 1723
rect 14400 1674 14431 1708
rect 14431 1674 14452 1708
rect 14400 1671 14452 1674
rect 14488 1671 14540 1708
rect 14576 1671 14628 1708
rect 14400 1635 14452 1657
rect 14400 1605 14431 1635
rect 14431 1605 14452 1635
rect 14488 1634 14510 1657
rect 14510 1634 14540 1657
rect 14576 1634 14582 1657
rect 14582 1634 14616 1657
rect 14616 1634 14628 1657
rect 14488 1605 14540 1634
rect 14576 1605 14628 1634
rect 14400 1562 14452 1591
rect 14400 1539 14431 1562
rect 14431 1539 14452 1562
rect 14488 1560 14510 1591
rect 14510 1560 14540 1591
rect 14576 1560 14582 1591
rect 14582 1560 14616 1591
rect 14616 1560 14628 1591
rect 14488 1539 14540 1560
rect 14576 1539 14628 1560
rect 14400 1489 14452 1525
rect 14488 1520 14540 1525
rect 14576 1520 14628 1525
rect 14400 1473 14431 1489
rect 14431 1473 14452 1489
rect 14488 1486 14510 1520
rect 14510 1486 14540 1520
rect 14576 1486 14582 1520
rect 14582 1486 14616 1520
rect 14616 1486 14628 1520
rect 14488 1473 14540 1486
rect 14576 1473 14628 1486
<< metal2 >>
rect 575 4068 803 4074
rect 627 4016 663 4068
rect 715 4016 751 4068
rect 575 4003 803 4016
rect 627 3951 663 4003
rect 715 3951 751 4003
rect 575 3938 803 3951
rect 627 3886 663 3938
rect 715 3886 751 3938
rect 575 3873 803 3886
rect 627 3821 663 3873
rect 715 3821 751 3873
rect 575 3808 803 3821
rect 627 3756 663 3808
rect 715 3756 751 3808
rect 575 3743 803 3756
rect 627 3691 663 3743
rect 715 3691 751 3743
rect 575 3678 803 3691
rect 627 3626 663 3678
rect 715 3626 751 3678
rect 575 3613 803 3626
rect 627 3561 663 3613
rect 715 3561 751 3613
rect 575 3548 803 3561
rect 627 3496 663 3548
rect 715 3496 751 3548
rect 575 3483 803 3496
rect 627 3431 663 3483
rect 715 3431 751 3483
rect 575 3418 803 3431
rect 627 3366 663 3418
rect 715 3366 751 3418
rect 575 3353 803 3366
rect 627 3301 663 3353
rect 715 3301 751 3353
rect 575 3288 803 3301
rect 627 3236 663 3288
rect 715 3236 751 3288
rect 575 3223 803 3236
rect 627 3171 663 3223
rect 715 3171 751 3223
rect 575 3158 803 3171
rect 627 3106 663 3158
rect 715 3106 751 3158
rect 575 3093 803 3106
rect 627 3041 663 3093
rect 715 3041 751 3093
rect 575 3028 803 3041
rect 627 2976 663 3028
rect 715 2976 751 3028
rect 575 2963 803 2976
rect 627 2911 663 2963
rect 715 2911 751 2963
rect 575 2898 803 2911
rect 627 2846 663 2898
rect 715 2846 751 2898
rect 575 2833 803 2846
rect 627 2781 663 2833
rect 715 2781 751 2833
rect 575 2768 803 2781
rect 627 2716 663 2768
rect 715 2716 751 2768
rect 575 2703 803 2716
rect 627 2651 663 2703
rect 715 2651 751 2703
rect 575 2638 803 2651
rect 627 2586 663 2638
rect 715 2586 751 2638
rect 575 2573 803 2586
rect 627 2521 663 2573
rect 715 2521 751 2573
rect 575 2508 803 2521
rect 627 2456 663 2508
rect 715 2456 751 2508
rect 575 2443 803 2456
rect 627 2391 663 2443
rect 715 2391 751 2443
rect 575 2378 803 2391
rect 627 2326 663 2378
rect 715 2326 751 2378
rect 575 2313 803 2326
rect 627 2261 663 2313
rect 715 2261 751 2313
rect 575 2248 803 2261
rect 627 2196 663 2248
rect 715 2196 751 2248
rect 575 2183 803 2196
rect 627 2131 663 2183
rect 715 2131 751 2183
rect 575 2118 803 2131
rect 627 2066 663 2118
rect 715 2066 751 2118
rect 575 2053 803 2066
rect 627 2001 663 2053
rect 715 2001 751 2053
rect 575 1987 803 2001
rect 627 1935 663 1987
rect 715 1935 751 1987
rect 575 1921 803 1935
rect 627 1869 663 1921
rect 715 1869 751 1921
rect 575 1855 803 1869
rect 627 1803 663 1855
rect 715 1803 751 1855
rect 575 1789 803 1803
rect 627 1737 663 1789
rect 715 1737 751 1789
rect 575 1723 803 1737
rect 627 1671 663 1723
rect 715 1671 751 1723
rect 575 1657 803 1671
rect 627 1605 663 1657
rect 715 1605 751 1657
rect 575 1591 803 1605
rect 627 1539 663 1591
rect 715 1539 751 1591
rect 575 1525 803 1539
rect 627 1473 663 1525
rect 715 1473 751 1525
rect 575 1467 803 1473
rect 1104 4068 1294 4074
rect 1104 4016 1109 4068
rect 1161 4016 1173 4068
rect 1225 4016 1237 4068
rect 1289 4016 1294 4068
rect 1104 4003 1294 4016
rect 1104 3951 1109 4003
rect 1161 3951 1173 4003
rect 1225 3951 1237 4003
rect 1289 3951 1294 4003
rect 1104 3938 1294 3951
rect 1104 3886 1109 3938
rect 1161 3886 1173 3938
rect 1225 3886 1237 3938
rect 1289 3886 1294 3938
rect 1104 3873 1294 3886
rect 1104 3821 1109 3873
rect 1161 3821 1173 3873
rect 1225 3821 1237 3873
rect 1289 3821 1294 3873
rect 1104 3808 1294 3821
rect 1104 3756 1109 3808
rect 1161 3756 1173 3808
rect 1225 3756 1237 3808
rect 1289 3756 1294 3808
rect 1104 3743 1294 3756
rect 1104 3691 1109 3743
rect 1161 3691 1173 3743
rect 1225 3691 1237 3743
rect 1289 3691 1294 3743
rect 1104 3678 1294 3691
rect 1104 3626 1109 3678
rect 1161 3626 1173 3678
rect 1225 3626 1237 3678
rect 1289 3626 1294 3678
rect 1104 3613 1294 3626
rect 1104 3561 1109 3613
rect 1161 3561 1173 3613
rect 1225 3561 1237 3613
rect 1289 3561 1294 3613
rect 1104 3548 1294 3561
rect 1104 3496 1109 3548
rect 1161 3496 1173 3548
rect 1225 3496 1237 3548
rect 1289 3496 1294 3548
rect 1104 3483 1294 3496
rect 1104 3431 1109 3483
rect 1161 3431 1173 3483
rect 1225 3431 1237 3483
rect 1289 3431 1294 3483
rect 1104 3418 1294 3431
rect 1104 3366 1109 3418
rect 1161 3366 1173 3418
rect 1225 3366 1237 3418
rect 1289 3366 1294 3418
rect 1104 3353 1294 3366
rect 1104 3301 1109 3353
rect 1161 3301 1173 3353
rect 1225 3301 1237 3353
rect 1289 3301 1294 3353
rect 1104 3288 1294 3301
rect 1104 3236 1109 3288
rect 1161 3236 1173 3288
rect 1225 3236 1237 3288
rect 1289 3236 1294 3288
rect 1104 3223 1294 3236
rect 1104 3171 1109 3223
rect 1161 3171 1173 3223
rect 1225 3171 1237 3223
rect 1289 3171 1294 3223
rect 1104 3158 1294 3171
rect 1104 3106 1109 3158
rect 1161 3106 1173 3158
rect 1225 3106 1237 3158
rect 1289 3106 1294 3158
rect 1104 3093 1294 3106
rect 1104 3041 1109 3093
rect 1161 3041 1173 3093
rect 1225 3041 1237 3093
rect 1289 3041 1294 3093
rect 1104 3028 1294 3041
rect 1104 2976 1109 3028
rect 1161 2976 1173 3028
rect 1225 2976 1237 3028
rect 1289 2976 1294 3028
rect 1104 2963 1294 2976
rect 1104 2911 1109 2963
rect 1161 2911 1173 2963
rect 1225 2911 1237 2963
rect 1289 2911 1294 2963
rect 1104 2898 1294 2911
rect 1104 2846 1109 2898
rect 1161 2846 1173 2898
rect 1225 2846 1237 2898
rect 1289 2846 1294 2898
rect 1104 2833 1294 2846
rect 1104 2781 1109 2833
rect 1161 2781 1173 2833
rect 1225 2781 1237 2833
rect 1289 2781 1294 2833
rect 1104 2768 1294 2781
rect 1104 2716 1109 2768
rect 1161 2716 1173 2768
rect 1225 2716 1237 2768
rect 1289 2716 1294 2768
rect 1104 2703 1294 2716
rect 1104 2651 1109 2703
rect 1161 2651 1173 2703
rect 1225 2651 1237 2703
rect 1289 2651 1294 2703
rect 1104 2638 1294 2651
rect 1104 2586 1109 2638
rect 1161 2586 1173 2638
rect 1225 2586 1237 2638
rect 1289 2586 1294 2638
rect 1104 2573 1294 2586
rect 1104 2521 1109 2573
rect 1161 2521 1173 2573
rect 1225 2521 1237 2573
rect 1289 2521 1294 2573
rect 1104 2508 1294 2521
rect 1104 2456 1109 2508
rect 1161 2456 1173 2508
rect 1225 2456 1237 2508
rect 1289 2456 1294 2508
rect 1104 2443 1294 2456
rect 1104 2391 1109 2443
rect 1161 2391 1173 2443
rect 1225 2391 1237 2443
rect 1289 2391 1294 2443
rect 1104 2378 1294 2391
rect 1104 2326 1109 2378
rect 1161 2326 1173 2378
rect 1225 2326 1237 2378
rect 1289 2326 1294 2378
rect 1104 2313 1294 2326
rect 1104 2261 1109 2313
rect 1161 2261 1173 2313
rect 1225 2261 1237 2313
rect 1289 2261 1294 2313
rect 1104 2248 1294 2261
rect 1104 2196 1109 2248
rect 1161 2196 1173 2248
rect 1225 2196 1237 2248
rect 1289 2196 1294 2248
rect 1104 2183 1294 2196
rect 1104 2131 1109 2183
rect 1161 2131 1173 2183
rect 1225 2131 1237 2183
rect 1289 2131 1294 2183
rect 1104 2118 1294 2131
rect 1104 2066 1109 2118
rect 1161 2066 1173 2118
rect 1225 2066 1237 2118
rect 1289 2066 1294 2118
rect 1104 2053 1294 2066
rect 1104 2001 1109 2053
rect 1161 2001 1173 2053
rect 1225 2001 1237 2053
rect 1289 2001 1294 2053
rect 1104 1987 1294 2001
rect 1104 1935 1109 1987
rect 1161 1935 1173 1987
rect 1225 1935 1237 1987
rect 1289 1935 1294 1987
rect 1104 1921 1294 1935
rect 1104 1869 1109 1921
rect 1161 1869 1173 1921
rect 1225 1869 1237 1921
rect 1289 1869 1294 1921
rect 1104 1855 1294 1869
rect 1104 1803 1109 1855
rect 1161 1803 1173 1855
rect 1225 1803 1237 1855
rect 1289 1803 1294 1855
rect 1104 1789 1294 1803
rect 1104 1737 1109 1789
rect 1161 1737 1173 1789
rect 1225 1737 1237 1789
rect 1289 1737 1294 1789
rect 1104 1723 1294 1737
rect 1104 1671 1109 1723
rect 1161 1671 1173 1723
rect 1225 1671 1237 1723
rect 1289 1671 1294 1723
rect 1104 1657 1294 1671
rect 1104 1605 1109 1657
rect 1161 1605 1173 1657
rect 1225 1605 1237 1657
rect 1289 1605 1294 1657
rect 1104 1591 1294 1605
rect 1104 1539 1109 1591
rect 1161 1539 1173 1591
rect 1225 1539 1237 1591
rect 1289 1539 1294 1591
rect 1104 1525 1294 1539
rect 1104 1473 1109 1525
rect 1161 1473 1173 1525
rect 1225 1473 1237 1525
rect 1289 1473 1294 1525
rect 1104 1467 1294 1473
rect 1600 4068 1790 4074
rect 1600 4016 1605 4068
rect 1657 4016 1669 4068
rect 1721 4016 1733 4068
rect 1785 4016 1790 4068
rect 1600 4003 1790 4016
rect 1600 3951 1605 4003
rect 1657 3951 1669 4003
rect 1721 3951 1733 4003
rect 1785 3951 1790 4003
rect 1600 3938 1790 3951
rect 1600 3886 1605 3938
rect 1657 3886 1669 3938
rect 1721 3886 1733 3938
rect 1785 3886 1790 3938
rect 1600 3873 1790 3886
rect 1600 3821 1605 3873
rect 1657 3821 1669 3873
rect 1721 3821 1733 3873
rect 1785 3821 1790 3873
rect 1600 3808 1790 3821
rect 1600 3756 1605 3808
rect 1657 3756 1669 3808
rect 1721 3756 1733 3808
rect 1785 3756 1790 3808
rect 1600 3743 1790 3756
rect 1600 3691 1605 3743
rect 1657 3691 1669 3743
rect 1721 3691 1733 3743
rect 1785 3691 1790 3743
rect 1600 3678 1790 3691
rect 1600 3626 1605 3678
rect 1657 3626 1669 3678
rect 1721 3626 1733 3678
rect 1785 3626 1790 3678
rect 1600 3613 1790 3626
rect 1600 3561 1605 3613
rect 1657 3561 1669 3613
rect 1721 3561 1733 3613
rect 1785 3561 1790 3613
rect 1600 3548 1790 3561
rect 1600 3496 1605 3548
rect 1657 3496 1669 3548
rect 1721 3496 1733 3548
rect 1785 3496 1790 3548
rect 1600 3483 1790 3496
rect 1600 3431 1605 3483
rect 1657 3431 1669 3483
rect 1721 3431 1733 3483
rect 1785 3431 1790 3483
rect 1600 3418 1790 3431
rect 1600 3366 1605 3418
rect 1657 3366 1669 3418
rect 1721 3366 1733 3418
rect 1785 3366 1790 3418
rect 1600 3353 1790 3366
rect 1600 3301 1605 3353
rect 1657 3301 1669 3353
rect 1721 3301 1733 3353
rect 1785 3301 1790 3353
rect 1600 3288 1790 3301
rect 1600 3236 1605 3288
rect 1657 3236 1669 3288
rect 1721 3236 1733 3288
rect 1785 3236 1790 3288
rect 1600 3223 1790 3236
rect 1600 3171 1605 3223
rect 1657 3171 1669 3223
rect 1721 3171 1733 3223
rect 1785 3171 1790 3223
rect 1600 3158 1790 3171
rect 1600 3106 1605 3158
rect 1657 3106 1669 3158
rect 1721 3106 1733 3158
rect 1785 3106 1790 3158
rect 1600 3093 1790 3106
rect 1600 3041 1605 3093
rect 1657 3041 1669 3093
rect 1721 3041 1733 3093
rect 1785 3041 1790 3093
rect 1600 3028 1790 3041
rect 1600 2976 1605 3028
rect 1657 2976 1669 3028
rect 1721 2976 1733 3028
rect 1785 2976 1790 3028
rect 1600 2963 1790 2976
rect 1600 2911 1605 2963
rect 1657 2911 1669 2963
rect 1721 2911 1733 2963
rect 1785 2911 1790 2963
rect 1600 2898 1790 2911
rect 1600 2846 1605 2898
rect 1657 2846 1669 2898
rect 1721 2846 1733 2898
rect 1785 2846 1790 2898
rect 1600 2833 1790 2846
rect 1600 2781 1605 2833
rect 1657 2781 1669 2833
rect 1721 2781 1733 2833
rect 1785 2781 1790 2833
rect 1600 2768 1790 2781
rect 1600 2716 1605 2768
rect 1657 2716 1669 2768
rect 1721 2716 1733 2768
rect 1785 2716 1790 2768
rect 1600 2703 1790 2716
rect 1600 2651 1605 2703
rect 1657 2651 1669 2703
rect 1721 2651 1733 2703
rect 1785 2651 1790 2703
rect 1600 2638 1790 2651
rect 1600 2586 1605 2638
rect 1657 2586 1669 2638
rect 1721 2586 1733 2638
rect 1785 2586 1790 2638
rect 1600 2573 1790 2586
rect 1600 2521 1605 2573
rect 1657 2521 1669 2573
rect 1721 2521 1733 2573
rect 1785 2521 1790 2573
rect 1600 2508 1790 2521
rect 1600 2456 1605 2508
rect 1657 2456 1669 2508
rect 1721 2456 1733 2508
rect 1785 2456 1790 2508
rect 1600 2443 1790 2456
rect 1600 2391 1605 2443
rect 1657 2391 1669 2443
rect 1721 2391 1733 2443
rect 1785 2391 1790 2443
rect 1600 2378 1790 2391
rect 1600 2326 1605 2378
rect 1657 2326 1669 2378
rect 1721 2326 1733 2378
rect 1785 2326 1790 2378
rect 1600 2313 1790 2326
rect 1600 2261 1605 2313
rect 1657 2261 1669 2313
rect 1721 2261 1733 2313
rect 1785 2261 1790 2313
rect 1600 2248 1790 2261
rect 1600 2196 1605 2248
rect 1657 2196 1669 2248
rect 1721 2196 1733 2248
rect 1785 2196 1790 2248
rect 1600 2183 1790 2196
rect 1600 2131 1605 2183
rect 1657 2131 1669 2183
rect 1721 2131 1733 2183
rect 1785 2131 1790 2183
rect 1600 2118 1790 2131
rect 1600 2066 1605 2118
rect 1657 2066 1669 2118
rect 1721 2066 1733 2118
rect 1785 2066 1790 2118
rect 1600 2053 1790 2066
rect 1600 2001 1605 2053
rect 1657 2001 1669 2053
rect 1721 2001 1733 2053
rect 1785 2001 1790 2053
rect 1600 1987 1790 2001
rect 1600 1935 1605 1987
rect 1657 1935 1669 1987
rect 1721 1935 1733 1987
rect 1785 1935 1790 1987
rect 1600 1921 1790 1935
rect 1600 1869 1605 1921
rect 1657 1869 1669 1921
rect 1721 1869 1733 1921
rect 1785 1869 1790 1921
rect 1600 1855 1790 1869
rect 1600 1803 1605 1855
rect 1657 1803 1669 1855
rect 1721 1803 1733 1855
rect 1785 1803 1790 1855
rect 1600 1789 1790 1803
rect 1600 1737 1605 1789
rect 1657 1737 1669 1789
rect 1721 1737 1733 1789
rect 1785 1737 1790 1789
rect 1600 1723 1790 1737
rect 1600 1671 1605 1723
rect 1657 1671 1669 1723
rect 1721 1671 1733 1723
rect 1785 1671 1790 1723
rect 1600 1657 1790 1671
rect 1600 1605 1605 1657
rect 1657 1605 1669 1657
rect 1721 1605 1733 1657
rect 1785 1605 1790 1657
rect 1600 1591 1790 1605
rect 1600 1539 1605 1591
rect 1657 1539 1669 1591
rect 1721 1539 1733 1591
rect 1785 1539 1790 1591
rect 1600 1525 1790 1539
rect 1600 1473 1605 1525
rect 1657 1473 1669 1525
rect 1721 1473 1733 1525
rect 1785 1473 1790 1525
rect 1600 1467 1790 1473
rect 2096 4068 2286 4074
rect 2096 4016 2101 4068
rect 2153 4016 2165 4068
rect 2217 4016 2229 4068
rect 2281 4016 2286 4068
rect 2096 4003 2286 4016
rect 2096 3951 2101 4003
rect 2153 3951 2165 4003
rect 2217 3951 2229 4003
rect 2281 3951 2286 4003
rect 2096 3938 2286 3951
rect 2096 3886 2101 3938
rect 2153 3886 2165 3938
rect 2217 3886 2229 3938
rect 2281 3886 2286 3938
rect 2096 3873 2286 3886
rect 2096 3821 2101 3873
rect 2153 3821 2165 3873
rect 2217 3821 2229 3873
rect 2281 3821 2286 3873
rect 2096 3808 2286 3821
rect 2096 3756 2101 3808
rect 2153 3756 2165 3808
rect 2217 3756 2229 3808
rect 2281 3756 2286 3808
rect 2096 3743 2286 3756
rect 2096 3691 2101 3743
rect 2153 3691 2165 3743
rect 2217 3691 2229 3743
rect 2281 3691 2286 3743
rect 2096 3678 2286 3691
rect 2096 3626 2101 3678
rect 2153 3626 2165 3678
rect 2217 3626 2229 3678
rect 2281 3626 2286 3678
rect 2096 3613 2286 3626
rect 2096 3561 2101 3613
rect 2153 3561 2165 3613
rect 2217 3561 2229 3613
rect 2281 3561 2286 3613
rect 2096 3548 2286 3561
rect 2096 3496 2101 3548
rect 2153 3496 2165 3548
rect 2217 3496 2229 3548
rect 2281 3496 2286 3548
rect 2096 3483 2286 3496
rect 2096 3431 2101 3483
rect 2153 3431 2165 3483
rect 2217 3431 2229 3483
rect 2281 3431 2286 3483
rect 2096 3418 2286 3431
rect 2096 3366 2101 3418
rect 2153 3366 2165 3418
rect 2217 3366 2229 3418
rect 2281 3366 2286 3418
rect 2096 3353 2286 3366
rect 2096 3301 2101 3353
rect 2153 3301 2165 3353
rect 2217 3301 2229 3353
rect 2281 3301 2286 3353
rect 2096 3288 2286 3301
rect 2096 3236 2101 3288
rect 2153 3236 2165 3288
rect 2217 3236 2229 3288
rect 2281 3236 2286 3288
rect 2096 3223 2286 3236
rect 2096 3171 2101 3223
rect 2153 3171 2165 3223
rect 2217 3171 2229 3223
rect 2281 3171 2286 3223
rect 2096 3158 2286 3171
rect 2096 3106 2101 3158
rect 2153 3106 2165 3158
rect 2217 3106 2229 3158
rect 2281 3106 2286 3158
rect 2096 3093 2286 3106
rect 2096 3041 2101 3093
rect 2153 3041 2165 3093
rect 2217 3041 2229 3093
rect 2281 3041 2286 3093
rect 2096 3028 2286 3041
rect 2096 2976 2101 3028
rect 2153 2976 2165 3028
rect 2217 2976 2229 3028
rect 2281 2976 2286 3028
rect 2096 2963 2286 2976
rect 2096 2911 2101 2963
rect 2153 2911 2165 2963
rect 2217 2911 2229 2963
rect 2281 2911 2286 2963
rect 2096 2898 2286 2911
rect 2096 2846 2101 2898
rect 2153 2846 2165 2898
rect 2217 2846 2229 2898
rect 2281 2846 2286 2898
rect 2096 2833 2286 2846
rect 2096 2781 2101 2833
rect 2153 2781 2165 2833
rect 2217 2781 2229 2833
rect 2281 2781 2286 2833
rect 2096 2768 2286 2781
rect 2096 2716 2101 2768
rect 2153 2716 2165 2768
rect 2217 2716 2229 2768
rect 2281 2716 2286 2768
rect 2096 2703 2286 2716
rect 2096 2651 2101 2703
rect 2153 2651 2165 2703
rect 2217 2651 2229 2703
rect 2281 2651 2286 2703
rect 2096 2638 2286 2651
rect 2096 2586 2101 2638
rect 2153 2586 2165 2638
rect 2217 2586 2229 2638
rect 2281 2586 2286 2638
rect 2096 2573 2286 2586
rect 2096 2521 2101 2573
rect 2153 2521 2165 2573
rect 2217 2521 2229 2573
rect 2281 2521 2286 2573
rect 2096 2508 2286 2521
rect 2096 2456 2101 2508
rect 2153 2456 2165 2508
rect 2217 2456 2229 2508
rect 2281 2456 2286 2508
rect 2096 2443 2286 2456
rect 2096 2391 2101 2443
rect 2153 2391 2165 2443
rect 2217 2391 2229 2443
rect 2281 2391 2286 2443
rect 2096 2378 2286 2391
rect 2096 2326 2101 2378
rect 2153 2326 2165 2378
rect 2217 2326 2229 2378
rect 2281 2326 2286 2378
rect 2096 2313 2286 2326
rect 2096 2261 2101 2313
rect 2153 2261 2165 2313
rect 2217 2261 2229 2313
rect 2281 2261 2286 2313
rect 2096 2248 2286 2261
rect 2096 2196 2101 2248
rect 2153 2196 2165 2248
rect 2217 2196 2229 2248
rect 2281 2196 2286 2248
rect 2096 2183 2286 2196
rect 2096 2131 2101 2183
rect 2153 2131 2165 2183
rect 2217 2131 2229 2183
rect 2281 2131 2286 2183
rect 2096 2118 2286 2131
rect 2096 2066 2101 2118
rect 2153 2066 2165 2118
rect 2217 2066 2229 2118
rect 2281 2066 2286 2118
rect 2096 2053 2286 2066
rect 2096 2001 2101 2053
rect 2153 2001 2165 2053
rect 2217 2001 2229 2053
rect 2281 2001 2286 2053
rect 2096 1987 2286 2001
rect 2096 1935 2101 1987
rect 2153 1935 2165 1987
rect 2217 1935 2229 1987
rect 2281 1935 2286 1987
rect 2096 1921 2286 1935
rect 2096 1869 2101 1921
rect 2153 1869 2165 1921
rect 2217 1869 2229 1921
rect 2281 1869 2286 1921
rect 2096 1855 2286 1869
rect 2096 1803 2101 1855
rect 2153 1803 2165 1855
rect 2217 1803 2229 1855
rect 2281 1803 2286 1855
rect 2096 1789 2286 1803
rect 2096 1737 2101 1789
rect 2153 1737 2165 1789
rect 2217 1737 2229 1789
rect 2281 1737 2286 1789
rect 2096 1723 2286 1737
rect 2096 1671 2101 1723
rect 2153 1671 2165 1723
rect 2217 1671 2229 1723
rect 2281 1671 2286 1723
rect 2096 1657 2286 1671
rect 2096 1605 2101 1657
rect 2153 1605 2165 1657
rect 2217 1605 2229 1657
rect 2281 1605 2286 1657
rect 2096 1591 2286 1605
rect 2096 1539 2101 1591
rect 2153 1539 2165 1591
rect 2217 1539 2229 1591
rect 2281 1539 2286 1591
rect 2096 1525 2286 1539
rect 2096 1473 2101 1525
rect 2153 1473 2165 1525
rect 2217 1473 2229 1525
rect 2281 1473 2286 1525
rect 2096 1467 2286 1473
rect 2592 4068 2782 4074
rect 2592 4016 2597 4068
rect 2649 4016 2661 4068
rect 2713 4016 2725 4068
rect 2777 4016 2782 4068
rect 2592 4003 2782 4016
rect 2592 3951 2597 4003
rect 2649 3951 2661 4003
rect 2713 3951 2725 4003
rect 2777 3951 2782 4003
rect 2592 3938 2782 3951
rect 2592 3886 2597 3938
rect 2649 3886 2661 3938
rect 2713 3886 2725 3938
rect 2777 3886 2782 3938
rect 2592 3873 2782 3886
rect 2592 3821 2597 3873
rect 2649 3821 2661 3873
rect 2713 3821 2725 3873
rect 2777 3821 2782 3873
rect 2592 3808 2782 3821
rect 2592 3756 2597 3808
rect 2649 3756 2661 3808
rect 2713 3756 2725 3808
rect 2777 3756 2782 3808
rect 2592 3743 2782 3756
rect 2592 3691 2597 3743
rect 2649 3691 2661 3743
rect 2713 3691 2725 3743
rect 2777 3691 2782 3743
rect 2592 3678 2782 3691
rect 2592 3626 2597 3678
rect 2649 3626 2661 3678
rect 2713 3626 2725 3678
rect 2777 3626 2782 3678
rect 2592 3613 2782 3626
rect 2592 3561 2597 3613
rect 2649 3561 2661 3613
rect 2713 3561 2725 3613
rect 2777 3561 2782 3613
rect 2592 3548 2782 3561
rect 2592 3496 2597 3548
rect 2649 3496 2661 3548
rect 2713 3496 2725 3548
rect 2777 3496 2782 3548
rect 2592 3483 2782 3496
rect 2592 3431 2597 3483
rect 2649 3431 2661 3483
rect 2713 3431 2725 3483
rect 2777 3431 2782 3483
rect 2592 3418 2782 3431
rect 2592 3366 2597 3418
rect 2649 3366 2661 3418
rect 2713 3366 2725 3418
rect 2777 3366 2782 3418
rect 2592 3353 2782 3366
rect 2592 3301 2597 3353
rect 2649 3301 2661 3353
rect 2713 3301 2725 3353
rect 2777 3301 2782 3353
rect 2592 3288 2782 3301
rect 2592 3236 2597 3288
rect 2649 3236 2661 3288
rect 2713 3236 2725 3288
rect 2777 3236 2782 3288
rect 2592 3223 2782 3236
rect 2592 3171 2597 3223
rect 2649 3171 2661 3223
rect 2713 3171 2725 3223
rect 2777 3171 2782 3223
rect 2592 3158 2782 3171
rect 2592 3106 2597 3158
rect 2649 3106 2661 3158
rect 2713 3106 2725 3158
rect 2777 3106 2782 3158
rect 2592 3093 2782 3106
rect 2592 3041 2597 3093
rect 2649 3041 2661 3093
rect 2713 3041 2725 3093
rect 2777 3041 2782 3093
rect 2592 3028 2782 3041
rect 2592 2976 2597 3028
rect 2649 2976 2661 3028
rect 2713 2976 2725 3028
rect 2777 2976 2782 3028
rect 2592 2963 2782 2976
rect 2592 2911 2597 2963
rect 2649 2911 2661 2963
rect 2713 2911 2725 2963
rect 2777 2911 2782 2963
rect 2592 2898 2782 2911
rect 2592 2846 2597 2898
rect 2649 2846 2661 2898
rect 2713 2846 2725 2898
rect 2777 2846 2782 2898
rect 2592 2833 2782 2846
rect 2592 2781 2597 2833
rect 2649 2781 2661 2833
rect 2713 2781 2725 2833
rect 2777 2781 2782 2833
rect 2592 2768 2782 2781
rect 2592 2716 2597 2768
rect 2649 2716 2661 2768
rect 2713 2716 2725 2768
rect 2777 2716 2782 2768
rect 2592 2703 2782 2716
rect 2592 2651 2597 2703
rect 2649 2651 2661 2703
rect 2713 2651 2725 2703
rect 2777 2651 2782 2703
rect 2592 2638 2782 2651
rect 2592 2586 2597 2638
rect 2649 2586 2661 2638
rect 2713 2586 2725 2638
rect 2777 2586 2782 2638
rect 2592 2573 2782 2586
rect 2592 2521 2597 2573
rect 2649 2521 2661 2573
rect 2713 2521 2725 2573
rect 2777 2521 2782 2573
rect 2592 2508 2782 2521
rect 2592 2456 2597 2508
rect 2649 2456 2661 2508
rect 2713 2456 2725 2508
rect 2777 2456 2782 2508
rect 2592 2443 2782 2456
rect 2592 2391 2597 2443
rect 2649 2391 2661 2443
rect 2713 2391 2725 2443
rect 2777 2391 2782 2443
rect 2592 2378 2782 2391
rect 2592 2326 2597 2378
rect 2649 2326 2661 2378
rect 2713 2326 2725 2378
rect 2777 2326 2782 2378
rect 2592 2313 2782 2326
rect 2592 2261 2597 2313
rect 2649 2261 2661 2313
rect 2713 2261 2725 2313
rect 2777 2261 2782 2313
rect 2592 2248 2782 2261
rect 2592 2196 2597 2248
rect 2649 2196 2661 2248
rect 2713 2196 2725 2248
rect 2777 2196 2782 2248
rect 2592 2183 2782 2196
rect 2592 2131 2597 2183
rect 2649 2131 2661 2183
rect 2713 2131 2725 2183
rect 2777 2131 2782 2183
rect 2592 2118 2782 2131
rect 2592 2066 2597 2118
rect 2649 2066 2661 2118
rect 2713 2066 2725 2118
rect 2777 2066 2782 2118
rect 2592 2053 2782 2066
rect 2592 2001 2597 2053
rect 2649 2001 2661 2053
rect 2713 2001 2725 2053
rect 2777 2001 2782 2053
rect 2592 1987 2782 2001
rect 2592 1935 2597 1987
rect 2649 1935 2661 1987
rect 2713 1935 2725 1987
rect 2777 1935 2782 1987
rect 2592 1921 2782 1935
rect 2592 1869 2597 1921
rect 2649 1869 2661 1921
rect 2713 1869 2725 1921
rect 2777 1869 2782 1921
rect 2592 1855 2782 1869
rect 2592 1803 2597 1855
rect 2649 1803 2661 1855
rect 2713 1803 2725 1855
rect 2777 1803 2782 1855
rect 2592 1789 2782 1803
rect 2592 1737 2597 1789
rect 2649 1737 2661 1789
rect 2713 1737 2725 1789
rect 2777 1737 2782 1789
rect 2592 1723 2782 1737
rect 2592 1671 2597 1723
rect 2649 1671 2661 1723
rect 2713 1671 2725 1723
rect 2777 1671 2782 1723
rect 2592 1657 2782 1671
rect 2592 1605 2597 1657
rect 2649 1605 2661 1657
rect 2713 1605 2725 1657
rect 2777 1605 2782 1657
rect 2592 1591 2782 1605
rect 2592 1539 2597 1591
rect 2649 1539 2661 1591
rect 2713 1539 2725 1591
rect 2777 1539 2782 1591
rect 2592 1525 2782 1539
rect 2592 1473 2597 1525
rect 2649 1473 2661 1525
rect 2713 1473 2725 1525
rect 2777 1473 2782 1525
rect 2592 1467 2782 1473
rect 3088 4068 3278 4074
rect 3088 4016 3093 4068
rect 3145 4016 3157 4068
rect 3209 4016 3221 4068
rect 3273 4016 3278 4068
rect 3088 4003 3278 4016
rect 3088 3951 3093 4003
rect 3145 3951 3157 4003
rect 3209 3951 3221 4003
rect 3273 3951 3278 4003
rect 3088 3938 3278 3951
rect 3088 3886 3093 3938
rect 3145 3886 3157 3938
rect 3209 3886 3221 3938
rect 3273 3886 3278 3938
rect 3088 3873 3278 3886
rect 3088 3821 3093 3873
rect 3145 3821 3157 3873
rect 3209 3821 3221 3873
rect 3273 3821 3278 3873
rect 3088 3808 3278 3821
rect 3088 3756 3093 3808
rect 3145 3756 3157 3808
rect 3209 3756 3221 3808
rect 3273 3756 3278 3808
rect 3088 3743 3278 3756
rect 3088 3691 3093 3743
rect 3145 3691 3157 3743
rect 3209 3691 3221 3743
rect 3273 3691 3278 3743
rect 3088 3678 3278 3691
rect 3088 3626 3093 3678
rect 3145 3626 3157 3678
rect 3209 3626 3221 3678
rect 3273 3626 3278 3678
rect 3088 3613 3278 3626
rect 3088 3561 3093 3613
rect 3145 3561 3157 3613
rect 3209 3561 3221 3613
rect 3273 3561 3278 3613
rect 3088 3548 3278 3561
rect 3088 3496 3093 3548
rect 3145 3496 3157 3548
rect 3209 3496 3221 3548
rect 3273 3496 3278 3548
rect 3088 3483 3278 3496
rect 3088 3431 3093 3483
rect 3145 3431 3157 3483
rect 3209 3431 3221 3483
rect 3273 3431 3278 3483
rect 3088 3418 3278 3431
rect 3088 3366 3093 3418
rect 3145 3366 3157 3418
rect 3209 3366 3221 3418
rect 3273 3366 3278 3418
rect 3088 3353 3278 3366
rect 3088 3301 3093 3353
rect 3145 3301 3157 3353
rect 3209 3301 3221 3353
rect 3273 3301 3278 3353
rect 3088 3288 3278 3301
rect 3088 3236 3093 3288
rect 3145 3236 3157 3288
rect 3209 3236 3221 3288
rect 3273 3236 3278 3288
rect 3088 3223 3278 3236
rect 3088 3171 3093 3223
rect 3145 3171 3157 3223
rect 3209 3171 3221 3223
rect 3273 3171 3278 3223
rect 3088 3158 3278 3171
rect 3088 3106 3093 3158
rect 3145 3106 3157 3158
rect 3209 3106 3221 3158
rect 3273 3106 3278 3158
rect 3088 3093 3278 3106
rect 3088 3041 3093 3093
rect 3145 3041 3157 3093
rect 3209 3041 3221 3093
rect 3273 3041 3278 3093
rect 3088 3028 3278 3041
rect 3088 2976 3093 3028
rect 3145 2976 3157 3028
rect 3209 2976 3221 3028
rect 3273 2976 3278 3028
rect 3088 2963 3278 2976
rect 3088 2911 3093 2963
rect 3145 2911 3157 2963
rect 3209 2911 3221 2963
rect 3273 2911 3278 2963
rect 3088 2898 3278 2911
rect 3088 2846 3093 2898
rect 3145 2846 3157 2898
rect 3209 2846 3221 2898
rect 3273 2846 3278 2898
rect 3088 2833 3278 2846
rect 3088 2781 3093 2833
rect 3145 2781 3157 2833
rect 3209 2781 3221 2833
rect 3273 2781 3278 2833
rect 3088 2768 3278 2781
rect 3088 2716 3093 2768
rect 3145 2716 3157 2768
rect 3209 2716 3221 2768
rect 3273 2716 3278 2768
rect 3088 2703 3278 2716
rect 3088 2651 3093 2703
rect 3145 2651 3157 2703
rect 3209 2651 3221 2703
rect 3273 2651 3278 2703
rect 3088 2638 3278 2651
rect 3088 2586 3093 2638
rect 3145 2586 3157 2638
rect 3209 2586 3221 2638
rect 3273 2586 3278 2638
rect 3088 2573 3278 2586
rect 3088 2521 3093 2573
rect 3145 2521 3157 2573
rect 3209 2521 3221 2573
rect 3273 2521 3278 2573
rect 3088 2508 3278 2521
rect 3088 2456 3093 2508
rect 3145 2456 3157 2508
rect 3209 2456 3221 2508
rect 3273 2456 3278 2508
rect 3088 2443 3278 2456
rect 3088 2391 3093 2443
rect 3145 2391 3157 2443
rect 3209 2391 3221 2443
rect 3273 2391 3278 2443
rect 3088 2378 3278 2391
rect 3088 2326 3093 2378
rect 3145 2326 3157 2378
rect 3209 2326 3221 2378
rect 3273 2326 3278 2378
rect 3088 2313 3278 2326
rect 3088 2261 3093 2313
rect 3145 2261 3157 2313
rect 3209 2261 3221 2313
rect 3273 2261 3278 2313
rect 3088 2248 3278 2261
rect 3088 2196 3093 2248
rect 3145 2196 3157 2248
rect 3209 2196 3221 2248
rect 3273 2196 3278 2248
rect 3088 2183 3278 2196
rect 3088 2131 3093 2183
rect 3145 2131 3157 2183
rect 3209 2131 3221 2183
rect 3273 2131 3278 2183
rect 3088 2118 3278 2131
rect 3088 2066 3093 2118
rect 3145 2066 3157 2118
rect 3209 2066 3221 2118
rect 3273 2066 3278 2118
rect 3088 2053 3278 2066
rect 3088 2001 3093 2053
rect 3145 2001 3157 2053
rect 3209 2001 3221 2053
rect 3273 2001 3278 2053
rect 3088 1987 3278 2001
rect 3088 1935 3093 1987
rect 3145 1935 3157 1987
rect 3209 1935 3221 1987
rect 3273 1935 3278 1987
rect 3088 1921 3278 1935
rect 3088 1869 3093 1921
rect 3145 1869 3157 1921
rect 3209 1869 3221 1921
rect 3273 1869 3278 1921
rect 3088 1855 3278 1869
rect 3088 1803 3093 1855
rect 3145 1803 3157 1855
rect 3209 1803 3221 1855
rect 3273 1803 3278 1855
rect 3088 1789 3278 1803
rect 3088 1737 3093 1789
rect 3145 1737 3157 1789
rect 3209 1737 3221 1789
rect 3273 1737 3278 1789
rect 3088 1723 3278 1737
rect 3088 1671 3093 1723
rect 3145 1671 3157 1723
rect 3209 1671 3221 1723
rect 3273 1671 3278 1723
rect 3088 1657 3278 1671
rect 3088 1605 3093 1657
rect 3145 1605 3157 1657
rect 3209 1605 3221 1657
rect 3273 1605 3278 1657
rect 3088 1591 3278 1605
rect 3088 1539 3093 1591
rect 3145 1539 3157 1591
rect 3209 1539 3221 1591
rect 3273 1539 3278 1591
rect 3088 1525 3278 1539
rect 3088 1473 3093 1525
rect 3145 1473 3157 1525
rect 3209 1473 3221 1525
rect 3273 1473 3278 1525
rect 3088 1467 3278 1473
rect 3584 4068 3774 4074
rect 3584 4016 3589 4068
rect 3641 4016 3653 4068
rect 3705 4016 3717 4068
rect 3769 4016 3774 4068
rect 3584 4003 3774 4016
rect 3584 3951 3589 4003
rect 3641 3951 3653 4003
rect 3705 3951 3717 4003
rect 3769 3951 3774 4003
rect 3584 3938 3774 3951
rect 3584 3886 3589 3938
rect 3641 3886 3653 3938
rect 3705 3886 3717 3938
rect 3769 3886 3774 3938
rect 3584 3873 3774 3886
rect 3584 3821 3589 3873
rect 3641 3821 3653 3873
rect 3705 3821 3717 3873
rect 3769 3821 3774 3873
rect 3584 3808 3774 3821
rect 3584 3756 3589 3808
rect 3641 3756 3653 3808
rect 3705 3756 3717 3808
rect 3769 3756 3774 3808
rect 3584 3743 3774 3756
rect 3584 3691 3589 3743
rect 3641 3691 3653 3743
rect 3705 3691 3717 3743
rect 3769 3691 3774 3743
rect 3584 3678 3774 3691
rect 3584 3626 3589 3678
rect 3641 3626 3653 3678
rect 3705 3626 3717 3678
rect 3769 3626 3774 3678
rect 3584 3613 3774 3626
rect 3584 3561 3589 3613
rect 3641 3561 3653 3613
rect 3705 3561 3717 3613
rect 3769 3561 3774 3613
rect 3584 3548 3774 3561
rect 3584 3496 3589 3548
rect 3641 3496 3653 3548
rect 3705 3496 3717 3548
rect 3769 3496 3774 3548
rect 3584 3483 3774 3496
rect 3584 3431 3589 3483
rect 3641 3431 3653 3483
rect 3705 3431 3717 3483
rect 3769 3431 3774 3483
rect 3584 3418 3774 3431
rect 3584 3366 3589 3418
rect 3641 3366 3653 3418
rect 3705 3366 3717 3418
rect 3769 3366 3774 3418
rect 3584 3353 3774 3366
rect 3584 3301 3589 3353
rect 3641 3301 3653 3353
rect 3705 3301 3717 3353
rect 3769 3301 3774 3353
rect 3584 3288 3774 3301
rect 3584 3236 3589 3288
rect 3641 3236 3653 3288
rect 3705 3236 3717 3288
rect 3769 3236 3774 3288
rect 3584 3223 3774 3236
rect 3584 3171 3589 3223
rect 3641 3171 3653 3223
rect 3705 3171 3717 3223
rect 3769 3171 3774 3223
rect 3584 3158 3774 3171
rect 3584 3106 3589 3158
rect 3641 3106 3653 3158
rect 3705 3106 3717 3158
rect 3769 3106 3774 3158
rect 3584 3093 3774 3106
rect 3584 3041 3589 3093
rect 3641 3041 3653 3093
rect 3705 3041 3717 3093
rect 3769 3041 3774 3093
rect 3584 3028 3774 3041
rect 3584 2976 3589 3028
rect 3641 2976 3653 3028
rect 3705 2976 3717 3028
rect 3769 2976 3774 3028
rect 3584 2963 3774 2976
rect 3584 2911 3589 2963
rect 3641 2911 3653 2963
rect 3705 2911 3717 2963
rect 3769 2911 3774 2963
rect 3584 2898 3774 2911
rect 3584 2846 3589 2898
rect 3641 2846 3653 2898
rect 3705 2846 3717 2898
rect 3769 2846 3774 2898
rect 3584 2833 3774 2846
rect 3584 2781 3589 2833
rect 3641 2781 3653 2833
rect 3705 2781 3717 2833
rect 3769 2781 3774 2833
rect 3584 2768 3774 2781
rect 3584 2716 3589 2768
rect 3641 2716 3653 2768
rect 3705 2716 3717 2768
rect 3769 2716 3774 2768
rect 3584 2703 3774 2716
rect 3584 2651 3589 2703
rect 3641 2651 3653 2703
rect 3705 2651 3717 2703
rect 3769 2651 3774 2703
rect 3584 2638 3774 2651
rect 3584 2586 3589 2638
rect 3641 2586 3653 2638
rect 3705 2586 3717 2638
rect 3769 2586 3774 2638
rect 3584 2573 3774 2586
rect 3584 2521 3589 2573
rect 3641 2521 3653 2573
rect 3705 2521 3717 2573
rect 3769 2521 3774 2573
rect 3584 2508 3774 2521
rect 3584 2456 3589 2508
rect 3641 2456 3653 2508
rect 3705 2456 3717 2508
rect 3769 2456 3774 2508
rect 3584 2443 3774 2456
rect 3584 2391 3589 2443
rect 3641 2391 3653 2443
rect 3705 2391 3717 2443
rect 3769 2391 3774 2443
rect 3584 2378 3774 2391
rect 3584 2326 3589 2378
rect 3641 2326 3653 2378
rect 3705 2326 3717 2378
rect 3769 2326 3774 2378
rect 3584 2313 3774 2326
rect 3584 2261 3589 2313
rect 3641 2261 3653 2313
rect 3705 2261 3717 2313
rect 3769 2261 3774 2313
rect 3584 2248 3774 2261
rect 3584 2196 3589 2248
rect 3641 2196 3653 2248
rect 3705 2196 3717 2248
rect 3769 2196 3774 2248
rect 3584 2183 3774 2196
rect 3584 2131 3589 2183
rect 3641 2131 3653 2183
rect 3705 2131 3717 2183
rect 3769 2131 3774 2183
rect 3584 2118 3774 2131
rect 3584 2066 3589 2118
rect 3641 2066 3653 2118
rect 3705 2066 3717 2118
rect 3769 2066 3774 2118
rect 3584 2053 3774 2066
rect 3584 2001 3589 2053
rect 3641 2001 3653 2053
rect 3705 2001 3717 2053
rect 3769 2001 3774 2053
rect 3584 1987 3774 2001
rect 3584 1935 3589 1987
rect 3641 1935 3653 1987
rect 3705 1935 3717 1987
rect 3769 1935 3774 1987
rect 3584 1921 3774 1935
rect 3584 1869 3589 1921
rect 3641 1869 3653 1921
rect 3705 1869 3717 1921
rect 3769 1869 3774 1921
rect 3584 1855 3774 1869
rect 3584 1803 3589 1855
rect 3641 1803 3653 1855
rect 3705 1803 3717 1855
rect 3769 1803 3774 1855
rect 3584 1789 3774 1803
rect 3584 1737 3589 1789
rect 3641 1737 3653 1789
rect 3705 1737 3717 1789
rect 3769 1737 3774 1789
rect 3584 1723 3774 1737
rect 3584 1671 3589 1723
rect 3641 1671 3653 1723
rect 3705 1671 3717 1723
rect 3769 1671 3774 1723
rect 3584 1657 3774 1671
rect 3584 1605 3589 1657
rect 3641 1605 3653 1657
rect 3705 1605 3717 1657
rect 3769 1605 3774 1657
rect 3584 1591 3774 1605
rect 3584 1539 3589 1591
rect 3641 1539 3653 1591
rect 3705 1539 3717 1591
rect 3769 1539 3774 1591
rect 3584 1525 3774 1539
rect 3584 1473 3589 1525
rect 3641 1473 3653 1525
rect 3705 1473 3717 1525
rect 3769 1473 3774 1525
rect 3584 1467 3774 1473
rect 4080 4068 4270 4074
rect 4080 4016 4085 4068
rect 4137 4016 4149 4068
rect 4201 4016 4213 4068
rect 4265 4016 4270 4068
rect 4080 4003 4270 4016
rect 4080 3951 4085 4003
rect 4137 3951 4149 4003
rect 4201 3951 4213 4003
rect 4265 3951 4270 4003
rect 4080 3938 4270 3951
rect 4080 3886 4085 3938
rect 4137 3886 4149 3938
rect 4201 3886 4213 3938
rect 4265 3886 4270 3938
rect 4080 3873 4270 3886
rect 4080 3821 4085 3873
rect 4137 3821 4149 3873
rect 4201 3821 4213 3873
rect 4265 3821 4270 3873
rect 4080 3808 4270 3821
rect 4080 3756 4085 3808
rect 4137 3756 4149 3808
rect 4201 3756 4213 3808
rect 4265 3756 4270 3808
rect 4080 3743 4270 3756
rect 4080 3691 4085 3743
rect 4137 3691 4149 3743
rect 4201 3691 4213 3743
rect 4265 3691 4270 3743
rect 4080 3678 4270 3691
rect 4080 3626 4085 3678
rect 4137 3626 4149 3678
rect 4201 3626 4213 3678
rect 4265 3626 4270 3678
rect 4080 3613 4270 3626
rect 4080 3561 4085 3613
rect 4137 3561 4149 3613
rect 4201 3561 4213 3613
rect 4265 3561 4270 3613
rect 4080 3548 4270 3561
rect 4080 3496 4085 3548
rect 4137 3496 4149 3548
rect 4201 3496 4213 3548
rect 4265 3496 4270 3548
rect 4080 3483 4270 3496
rect 4080 3431 4085 3483
rect 4137 3431 4149 3483
rect 4201 3431 4213 3483
rect 4265 3431 4270 3483
rect 4080 3418 4270 3431
rect 4080 3366 4085 3418
rect 4137 3366 4149 3418
rect 4201 3366 4213 3418
rect 4265 3366 4270 3418
rect 4080 3353 4270 3366
rect 4080 3301 4085 3353
rect 4137 3301 4149 3353
rect 4201 3301 4213 3353
rect 4265 3301 4270 3353
rect 4080 3288 4270 3301
rect 4080 3236 4085 3288
rect 4137 3236 4149 3288
rect 4201 3236 4213 3288
rect 4265 3236 4270 3288
rect 4080 3223 4270 3236
rect 4080 3171 4085 3223
rect 4137 3171 4149 3223
rect 4201 3171 4213 3223
rect 4265 3171 4270 3223
rect 4080 3158 4270 3171
rect 4080 3106 4085 3158
rect 4137 3106 4149 3158
rect 4201 3106 4213 3158
rect 4265 3106 4270 3158
rect 4080 3093 4270 3106
rect 4080 3041 4085 3093
rect 4137 3041 4149 3093
rect 4201 3041 4213 3093
rect 4265 3041 4270 3093
rect 4080 3028 4270 3041
rect 4080 2976 4085 3028
rect 4137 2976 4149 3028
rect 4201 2976 4213 3028
rect 4265 2976 4270 3028
rect 4080 2963 4270 2976
rect 4080 2911 4085 2963
rect 4137 2911 4149 2963
rect 4201 2911 4213 2963
rect 4265 2911 4270 2963
rect 4080 2898 4270 2911
rect 4080 2846 4085 2898
rect 4137 2846 4149 2898
rect 4201 2846 4213 2898
rect 4265 2846 4270 2898
rect 4080 2833 4270 2846
rect 4080 2781 4085 2833
rect 4137 2781 4149 2833
rect 4201 2781 4213 2833
rect 4265 2781 4270 2833
rect 4080 2768 4270 2781
rect 4080 2716 4085 2768
rect 4137 2716 4149 2768
rect 4201 2716 4213 2768
rect 4265 2716 4270 2768
rect 4080 2703 4270 2716
rect 4080 2651 4085 2703
rect 4137 2651 4149 2703
rect 4201 2651 4213 2703
rect 4265 2651 4270 2703
rect 4080 2638 4270 2651
rect 4080 2586 4085 2638
rect 4137 2586 4149 2638
rect 4201 2586 4213 2638
rect 4265 2586 4270 2638
rect 4080 2573 4270 2586
rect 4080 2521 4085 2573
rect 4137 2521 4149 2573
rect 4201 2521 4213 2573
rect 4265 2521 4270 2573
rect 4080 2508 4270 2521
rect 4080 2456 4085 2508
rect 4137 2456 4149 2508
rect 4201 2456 4213 2508
rect 4265 2456 4270 2508
rect 4080 2443 4270 2456
rect 4080 2391 4085 2443
rect 4137 2391 4149 2443
rect 4201 2391 4213 2443
rect 4265 2391 4270 2443
rect 4080 2378 4270 2391
rect 4080 2326 4085 2378
rect 4137 2326 4149 2378
rect 4201 2326 4213 2378
rect 4265 2326 4270 2378
rect 4080 2313 4270 2326
rect 4080 2261 4085 2313
rect 4137 2261 4149 2313
rect 4201 2261 4213 2313
rect 4265 2261 4270 2313
rect 4080 2248 4270 2261
rect 4080 2196 4085 2248
rect 4137 2196 4149 2248
rect 4201 2196 4213 2248
rect 4265 2196 4270 2248
rect 4080 2183 4270 2196
rect 4080 2131 4085 2183
rect 4137 2131 4149 2183
rect 4201 2131 4213 2183
rect 4265 2131 4270 2183
rect 4080 2118 4270 2131
rect 4080 2066 4085 2118
rect 4137 2066 4149 2118
rect 4201 2066 4213 2118
rect 4265 2066 4270 2118
rect 4080 2053 4270 2066
rect 4080 2001 4085 2053
rect 4137 2001 4149 2053
rect 4201 2001 4213 2053
rect 4265 2001 4270 2053
rect 4080 1987 4270 2001
rect 4080 1935 4085 1987
rect 4137 1935 4149 1987
rect 4201 1935 4213 1987
rect 4265 1935 4270 1987
rect 4080 1921 4270 1935
rect 4080 1869 4085 1921
rect 4137 1869 4149 1921
rect 4201 1869 4213 1921
rect 4265 1869 4270 1921
rect 4080 1855 4270 1869
rect 4080 1803 4085 1855
rect 4137 1803 4149 1855
rect 4201 1803 4213 1855
rect 4265 1803 4270 1855
rect 4080 1789 4270 1803
rect 4080 1737 4085 1789
rect 4137 1737 4149 1789
rect 4201 1737 4213 1789
rect 4265 1737 4270 1789
rect 4080 1723 4270 1737
rect 4080 1671 4085 1723
rect 4137 1671 4149 1723
rect 4201 1671 4213 1723
rect 4265 1671 4270 1723
rect 4080 1657 4270 1671
rect 4080 1605 4085 1657
rect 4137 1605 4149 1657
rect 4201 1605 4213 1657
rect 4265 1605 4270 1657
rect 4080 1591 4270 1605
rect 4080 1539 4085 1591
rect 4137 1539 4149 1591
rect 4201 1539 4213 1591
rect 4265 1539 4270 1591
rect 4080 1525 4270 1539
rect 4080 1473 4085 1525
rect 4137 1473 4149 1525
rect 4201 1473 4213 1525
rect 4265 1473 4270 1525
rect 4080 1467 4270 1473
rect 4576 4068 4766 4074
rect 4576 4016 4581 4068
rect 4633 4016 4645 4068
rect 4697 4016 4709 4068
rect 4761 4016 4766 4068
rect 4576 4003 4766 4016
rect 4576 3951 4581 4003
rect 4633 3951 4645 4003
rect 4697 3951 4709 4003
rect 4761 3951 4766 4003
rect 4576 3938 4766 3951
rect 4576 3886 4581 3938
rect 4633 3886 4645 3938
rect 4697 3886 4709 3938
rect 4761 3886 4766 3938
rect 4576 3873 4766 3886
rect 4576 3821 4581 3873
rect 4633 3821 4645 3873
rect 4697 3821 4709 3873
rect 4761 3821 4766 3873
rect 4576 3808 4766 3821
rect 4576 3756 4581 3808
rect 4633 3756 4645 3808
rect 4697 3756 4709 3808
rect 4761 3756 4766 3808
rect 4576 3743 4766 3756
rect 4576 3691 4581 3743
rect 4633 3691 4645 3743
rect 4697 3691 4709 3743
rect 4761 3691 4766 3743
rect 4576 3678 4766 3691
rect 4576 3626 4581 3678
rect 4633 3626 4645 3678
rect 4697 3626 4709 3678
rect 4761 3626 4766 3678
rect 4576 3613 4766 3626
rect 4576 3561 4581 3613
rect 4633 3561 4645 3613
rect 4697 3561 4709 3613
rect 4761 3561 4766 3613
rect 4576 3548 4766 3561
rect 4576 3496 4581 3548
rect 4633 3496 4645 3548
rect 4697 3496 4709 3548
rect 4761 3496 4766 3548
rect 4576 3483 4766 3496
rect 4576 3431 4581 3483
rect 4633 3431 4645 3483
rect 4697 3431 4709 3483
rect 4761 3431 4766 3483
rect 4576 3418 4766 3431
rect 4576 3366 4581 3418
rect 4633 3366 4645 3418
rect 4697 3366 4709 3418
rect 4761 3366 4766 3418
rect 4576 3353 4766 3366
rect 4576 3301 4581 3353
rect 4633 3301 4645 3353
rect 4697 3301 4709 3353
rect 4761 3301 4766 3353
rect 4576 3288 4766 3301
rect 4576 3236 4581 3288
rect 4633 3236 4645 3288
rect 4697 3236 4709 3288
rect 4761 3236 4766 3288
rect 4576 3223 4766 3236
rect 4576 3171 4581 3223
rect 4633 3171 4645 3223
rect 4697 3171 4709 3223
rect 4761 3171 4766 3223
rect 4576 3158 4766 3171
rect 4576 3106 4581 3158
rect 4633 3106 4645 3158
rect 4697 3106 4709 3158
rect 4761 3106 4766 3158
rect 4576 3093 4766 3106
rect 4576 3041 4581 3093
rect 4633 3041 4645 3093
rect 4697 3041 4709 3093
rect 4761 3041 4766 3093
rect 4576 3028 4766 3041
rect 4576 2976 4581 3028
rect 4633 2976 4645 3028
rect 4697 2976 4709 3028
rect 4761 2976 4766 3028
rect 4576 2963 4766 2976
rect 4576 2911 4581 2963
rect 4633 2911 4645 2963
rect 4697 2911 4709 2963
rect 4761 2911 4766 2963
rect 4576 2898 4766 2911
rect 4576 2846 4581 2898
rect 4633 2846 4645 2898
rect 4697 2846 4709 2898
rect 4761 2846 4766 2898
rect 4576 2833 4766 2846
rect 4576 2781 4581 2833
rect 4633 2781 4645 2833
rect 4697 2781 4709 2833
rect 4761 2781 4766 2833
rect 4576 2768 4766 2781
rect 4576 2716 4581 2768
rect 4633 2716 4645 2768
rect 4697 2716 4709 2768
rect 4761 2716 4766 2768
rect 4576 2703 4766 2716
rect 4576 2651 4581 2703
rect 4633 2651 4645 2703
rect 4697 2651 4709 2703
rect 4761 2651 4766 2703
rect 4576 2638 4766 2651
rect 4576 2586 4581 2638
rect 4633 2586 4645 2638
rect 4697 2586 4709 2638
rect 4761 2586 4766 2638
rect 4576 2573 4766 2586
rect 4576 2521 4581 2573
rect 4633 2521 4645 2573
rect 4697 2521 4709 2573
rect 4761 2521 4766 2573
rect 4576 2508 4766 2521
rect 4576 2456 4581 2508
rect 4633 2456 4645 2508
rect 4697 2456 4709 2508
rect 4761 2456 4766 2508
rect 4576 2443 4766 2456
rect 4576 2391 4581 2443
rect 4633 2391 4645 2443
rect 4697 2391 4709 2443
rect 4761 2391 4766 2443
rect 4576 2378 4766 2391
rect 4576 2326 4581 2378
rect 4633 2326 4645 2378
rect 4697 2326 4709 2378
rect 4761 2326 4766 2378
rect 4576 2313 4766 2326
rect 4576 2261 4581 2313
rect 4633 2261 4645 2313
rect 4697 2261 4709 2313
rect 4761 2261 4766 2313
rect 4576 2248 4766 2261
rect 4576 2196 4581 2248
rect 4633 2196 4645 2248
rect 4697 2196 4709 2248
rect 4761 2196 4766 2248
rect 4576 2183 4766 2196
rect 4576 2131 4581 2183
rect 4633 2131 4645 2183
rect 4697 2131 4709 2183
rect 4761 2131 4766 2183
rect 4576 2118 4766 2131
rect 4576 2066 4581 2118
rect 4633 2066 4645 2118
rect 4697 2066 4709 2118
rect 4761 2066 4766 2118
rect 4576 2053 4766 2066
rect 4576 2001 4581 2053
rect 4633 2001 4645 2053
rect 4697 2001 4709 2053
rect 4761 2001 4766 2053
rect 4576 1987 4766 2001
rect 4576 1935 4581 1987
rect 4633 1935 4645 1987
rect 4697 1935 4709 1987
rect 4761 1935 4766 1987
rect 4576 1921 4766 1935
rect 4576 1869 4581 1921
rect 4633 1869 4645 1921
rect 4697 1869 4709 1921
rect 4761 1869 4766 1921
rect 4576 1855 4766 1869
rect 4576 1803 4581 1855
rect 4633 1803 4645 1855
rect 4697 1803 4709 1855
rect 4761 1803 4766 1855
rect 4576 1789 4766 1803
rect 4576 1737 4581 1789
rect 4633 1737 4645 1789
rect 4697 1737 4709 1789
rect 4761 1737 4766 1789
rect 4576 1723 4766 1737
rect 4576 1671 4581 1723
rect 4633 1671 4645 1723
rect 4697 1671 4709 1723
rect 4761 1671 4766 1723
rect 4576 1657 4766 1671
rect 4576 1605 4581 1657
rect 4633 1605 4645 1657
rect 4697 1605 4709 1657
rect 4761 1605 4766 1657
rect 4576 1591 4766 1605
rect 4576 1539 4581 1591
rect 4633 1539 4645 1591
rect 4697 1539 4709 1591
rect 4761 1539 4766 1591
rect 4576 1525 4766 1539
rect 4576 1473 4581 1525
rect 4633 1473 4645 1525
rect 4697 1473 4709 1525
rect 4761 1473 4766 1525
rect 4576 1467 4766 1473
rect 5072 4068 5262 4074
rect 5072 4016 5077 4068
rect 5129 4016 5141 4068
rect 5193 4016 5205 4068
rect 5257 4016 5262 4068
rect 5072 4003 5262 4016
rect 5072 3951 5077 4003
rect 5129 3951 5141 4003
rect 5193 3951 5205 4003
rect 5257 3951 5262 4003
rect 5072 3938 5262 3951
rect 5072 3886 5077 3938
rect 5129 3886 5141 3938
rect 5193 3886 5205 3938
rect 5257 3886 5262 3938
rect 5072 3873 5262 3886
rect 5072 3821 5077 3873
rect 5129 3821 5141 3873
rect 5193 3821 5205 3873
rect 5257 3821 5262 3873
rect 5072 3808 5262 3821
rect 5072 3756 5077 3808
rect 5129 3756 5141 3808
rect 5193 3756 5205 3808
rect 5257 3756 5262 3808
rect 5072 3743 5262 3756
rect 5072 3691 5077 3743
rect 5129 3691 5141 3743
rect 5193 3691 5205 3743
rect 5257 3691 5262 3743
rect 5072 3678 5262 3691
rect 5072 3626 5077 3678
rect 5129 3626 5141 3678
rect 5193 3626 5205 3678
rect 5257 3626 5262 3678
rect 5072 3613 5262 3626
rect 5072 3561 5077 3613
rect 5129 3561 5141 3613
rect 5193 3561 5205 3613
rect 5257 3561 5262 3613
rect 5072 3548 5262 3561
rect 5072 3496 5077 3548
rect 5129 3496 5141 3548
rect 5193 3496 5205 3548
rect 5257 3496 5262 3548
rect 5072 3483 5262 3496
rect 5072 3431 5077 3483
rect 5129 3431 5141 3483
rect 5193 3431 5205 3483
rect 5257 3431 5262 3483
rect 5072 3418 5262 3431
rect 5072 3366 5077 3418
rect 5129 3366 5141 3418
rect 5193 3366 5205 3418
rect 5257 3366 5262 3418
rect 5072 3353 5262 3366
rect 5072 3301 5077 3353
rect 5129 3301 5141 3353
rect 5193 3301 5205 3353
rect 5257 3301 5262 3353
rect 5072 3288 5262 3301
rect 5072 3236 5077 3288
rect 5129 3236 5141 3288
rect 5193 3236 5205 3288
rect 5257 3236 5262 3288
rect 5072 3223 5262 3236
rect 5072 3171 5077 3223
rect 5129 3171 5141 3223
rect 5193 3171 5205 3223
rect 5257 3171 5262 3223
rect 5072 3158 5262 3171
rect 5072 3106 5077 3158
rect 5129 3106 5141 3158
rect 5193 3106 5205 3158
rect 5257 3106 5262 3158
rect 5072 3093 5262 3106
rect 5072 3041 5077 3093
rect 5129 3041 5141 3093
rect 5193 3041 5205 3093
rect 5257 3041 5262 3093
rect 5072 3028 5262 3041
rect 5072 2976 5077 3028
rect 5129 2976 5141 3028
rect 5193 2976 5205 3028
rect 5257 2976 5262 3028
rect 5072 2963 5262 2976
rect 5072 2911 5077 2963
rect 5129 2911 5141 2963
rect 5193 2911 5205 2963
rect 5257 2911 5262 2963
rect 5072 2898 5262 2911
rect 5072 2846 5077 2898
rect 5129 2846 5141 2898
rect 5193 2846 5205 2898
rect 5257 2846 5262 2898
rect 5072 2833 5262 2846
rect 5072 2781 5077 2833
rect 5129 2781 5141 2833
rect 5193 2781 5205 2833
rect 5257 2781 5262 2833
rect 5072 2768 5262 2781
rect 5072 2716 5077 2768
rect 5129 2716 5141 2768
rect 5193 2716 5205 2768
rect 5257 2716 5262 2768
rect 5072 2703 5262 2716
rect 5072 2651 5077 2703
rect 5129 2651 5141 2703
rect 5193 2651 5205 2703
rect 5257 2651 5262 2703
rect 5072 2638 5262 2651
rect 5072 2586 5077 2638
rect 5129 2586 5141 2638
rect 5193 2586 5205 2638
rect 5257 2586 5262 2638
rect 5072 2573 5262 2586
rect 5072 2521 5077 2573
rect 5129 2521 5141 2573
rect 5193 2521 5205 2573
rect 5257 2521 5262 2573
rect 5072 2508 5262 2521
rect 5072 2456 5077 2508
rect 5129 2456 5141 2508
rect 5193 2456 5205 2508
rect 5257 2456 5262 2508
rect 5072 2443 5262 2456
rect 5072 2391 5077 2443
rect 5129 2391 5141 2443
rect 5193 2391 5205 2443
rect 5257 2391 5262 2443
rect 5072 2378 5262 2391
rect 5072 2326 5077 2378
rect 5129 2326 5141 2378
rect 5193 2326 5205 2378
rect 5257 2326 5262 2378
rect 5072 2313 5262 2326
rect 5072 2261 5077 2313
rect 5129 2261 5141 2313
rect 5193 2261 5205 2313
rect 5257 2261 5262 2313
rect 5072 2248 5262 2261
rect 5072 2196 5077 2248
rect 5129 2196 5141 2248
rect 5193 2196 5205 2248
rect 5257 2196 5262 2248
rect 5072 2183 5262 2196
rect 5072 2131 5077 2183
rect 5129 2131 5141 2183
rect 5193 2131 5205 2183
rect 5257 2131 5262 2183
rect 5072 2118 5262 2131
rect 5072 2066 5077 2118
rect 5129 2066 5141 2118
rect 5193 2066 5205 2118
rect 5257 2066 5262 2118
rect 5072 2053 5262 2066
rect 5072 2001 5077 2053
rect 5129 2001 5141 2053
rect 5193 2001 5205 2053
rect 5257 2001 5262 2053
rect 5072 1987 5262 2001
rect 5072 1935 5077 1987
rect 5129 1935 5141 1987
rect 5193 1935 5205 1987
rect 5257 1935 5262 1987
rect 5072 1921 5262 1935
rect 5072 1869 5077 1921
rect 5129 1869 5141 1921
rect 5193 1869 5205 1921
rect 5257 1869 5262 1921
rect 5072 1855 5262 1869
rect 5072 1803 5077 1855
rect 5129 1803 5141 1855
rect 5193 1803 5205 1855
rect 5257 1803 5262 1855
rect 5072 1789 5262 1803
rect 5072 1737 5077 1789
rect 5129 1737 5141 1789
rect 5193 1737 5205 1789
rect 5257 1737 5262 1789
rect 5072 1723 5262 1737
rect 5072 1671 5077 1723
rect 5129 1671 5141 1723
rect 5193 1671 5205 1723
rect 5257 1671 5262 1723
rect 5072 1657 5262 1671
rect 5072 1605 5077 1657
rect 5129 1605 5141 1657
rect 5193 1605 5205 1657
rect 5257 1605 5262 1657
rect 5072 1591 5262 1605
rect 5072 1539 5077 1591
rect 5129 1539 5141 1591
rect 5193 1539 5205 1591
rect 5257 1539 5262 1591
rect 5072 1525 5262 1539
rect 5072 1473 5077 1525
rect 5129 1473 5141 1525
rect 5193 1473 5205 1525
rect 5257 1473 5262 1525
rect 5072 1467 5262 1473
rect 5568 4068 5758 4074
rect 5568 4016 5573 4068
rect 5625 4016 5637 4068
rect 5689 4016 5701 4068
rect 5753 4016 5758 4068
rect 5568 4003 5758 4016
rect 5568 3951 5573 4003
rect 5625 3951 5637 4003
rect 5689 3951 5701 4003
rect 5753 3951 5758 4003
rect 5568 3938 5758 3951
rect 5568 3886 5573 3938
rect 5625 3886 5637 3938
rect 5689 3886 5701 3938
rect 5753 3886 5758 3938
rect 5568 3873 5758 3886
rect 5568 3821 5573 3873
rect 5625 3821 5637 3873
rect 5689 3821 5701 3873
rect 5753 3821 5758 3873
rect 5568 3808 5758 3821
rect 5568 3756 5573 3808
rect 5625 3756 5637 3808
rect 5689 3756 5701 3808
rect 5753 3756 5758 3808
rect 5568 3743 5758 3756
rect 5568 3691 5573 3743
rect 5625 3691 5637 3743
rect 5689 3691 5701 3743
rect 5753 3691 5758 3743
rect 5568 3678 5758 3691
rect 5568 3626 5573 3678
rect 5625 3626 5637 3678
rect 5689 3626 5701 3678
rect 5753 3626 5758 3678
rect 5568 3613 5758 3626
rect 5568 3561 5573 3613
rect 5625 3561 5637 3613
rect 5689 3561 5701 3613
rect 5753 3561 5758 3613
rect 5568 3548 5758 3561
rect 5568 3496 5573 3548
rect 5625 3496 5637 3548
rect 5689 3496 5701 3548
rect 5753 3496 5758 3548
rect 5568 3483 5758 3496
rect 5568 3431 5573 3483
rect 5625 3431 5637 3483
rect 5689 3431 5701 3483
rect 5753 3431 5758 3483
rect 5568 3418 5758 3431
rect 5568 3366 5573 3418
rect 5625 3366 5637 3418
rect 5689 3366 5701 3418
rect 5753 3366 5758 3418
rect 5568 3353 5758 3366
rect 5568 3301 5573 3353
rect 5625 3301 5637 3353
rect 5689 3301 5701 3353
rect 5753 3301 5758 3353
rect 5568 3288 5758 3301
rect 5568 3236 5573 3288
rect 5625 3236 5637 3288
rect 5689 3236 5701 3288
rect 5753 3236 5758 3288
rect 5568 3223 5758 3236
rect 5568 3171 5573 3223
rect 5625 3171 5637 3223
rect 5689 3171 5701 3223
rect 5753 3171 5758 3223
rect 5568 3158 5758 3171
rect 5568 3106 5573 3158
rect 5625 3106 5637 3158
rect 5689 3106 5701 3158
rect 5753 3106 5758 3158
rect 5568 3093 5758 3106
rect 5568 3041 5573 3093
rect 5625 3041 5637 3093
rect 5689 3041 5701 3093
rect 5753 3041 5758 3093
rect 5568 3028 5758 3041
rect 5568 2976 5573 3028
rect 5625 2976 5637 3028
rect 5689 2976 5701 3028
rect 5753 2976 5758 3028
rect 5568 2963 5758 2976
rect 5568 2911 5573 2963
rect 5625 2911 5637 2963
rect 5689 2911 5701 2963
rect 5753 2911 5758 2963
rect 5568 2898 5758 2911
rect 5568 2846 5573 2898
rect 5625 2846 5637 2898
rect 5689 2846 5701 2898
rect 5753 2846 5758 2898
rect 5568 2833 5758 2846
rect 5568 2781 5573 2833
rect 5625 2781 5637 2833
rect 5689 2781 5701 2833
rect 5753 2781 5758 2833
rect 5568 2768 5758 2781
rect 5568 2716 5573 2768
rect 5625 2716 5637 2768
rect 5689 2716 5701 2768
rect 5753 2716 5758 2768
rect 5568 2703 5758 2716
rect 5568 2651 5573 2703
rect 5625 2651 5637 2703
rect 5689 2651 5701 2703
rect 5753 2651 5758 2703
rect 5568 2638 5758 2651
rect 5568 2586 5573 2638
rect 5625 2586 5637 2638
rect 5689 2586 5701 2638
rect 5753 2586 5758 2638
rect 5568 2573 5758 2586
rect 5568 2521 5573 2573
rect 5625 2521 5637 2573
rect 5689 2521 5701 2573
rect 5753 2521 5758 2573
rect 5568 2508 5758 2521
rect 5568 2456 5573 2508
rect 5625 2456 5637 2508
rect 5689 2456 5701 2508
rect 5753 2456 5758 2508
rect 5568 2443 5758 2456
rect 5568 2391 5573 2443
rect 5625 2391 5637 2443
rect 5689 2391 5701 2443
rect 5753 2391 5758 2443
rect 5568 2378 5758 2391
rect 5568 2326 5573 2378
rect 5625 2326 5637 2378
rect 5689 2326 5701 2378
rect 5753 2326 5758 2378
rect 5568 2313 5758 2326
rect 5568 2261 5573 2313
rect 5625 2261 5637 2313
rect 5689 2261 5701 2313
rect 5753 2261 5758 2313
rect 5568 2248 5758 2261
rect 5568 2196 5573 2248
rect 5625 2196 5637 2248
rect 5689 2196 5701 2248
rect 5753 2196 5758 2248
rect 5568 2183 5758 2196
rect 5568 2131 5573 2183
rect 5625 2131 5637 2183
rect 5689 2131 5701 2183
rect 5753 2131 5758 2183
rect 5568 2118 5758 2131
rect 5568 2066 5573 2118
rect 5625 2066 5637 2118
rect 5689 2066 5701 2118
rect 5753 2066 5758 2118
rect 5568 2053 5758 2066
rect 5568 2001 5573 2053
rect 5625 2001 5637 2053
rect 5689 2001 5701 2053
rect 5753 2001 5758 2053
rect 5568 1987 5758 2001
rect 5568 1935 5573 1987
rect 5625 1935 5637 1987
rect 5689 1935 5701 1987
rect 5753 1935 5758 1987
rect 5568 1921 5758 1935
rect 5568 1869 5573 1921
rect 5625 1869 5637 1921
rect 5689 1869 5701 1921
rect 5753 1869 5758 1921
rect 5568 1855 5758 1869
rect 5568 1803 5573 1855
rect 5625 1803 5637 1855
rect 5689 1803 5701 1855
rect 5753 1803 5758 1855
rect 5568 1789 5758 1803
rect 5568 1737 5573 1789
rect 5625 1737 5637 1789
rect 5689 1737 5701 1789
rect 5753 1737 5758 1789
rect 5568 1723 5758 1737
rect 5568 1671 5573 1723
rect 5625 1671 5637 1723
rect 5689 1671 5701 1723
rect 5753 1671 5758 1723
rect 5568 1657 5758 1671
rect 5568 1605 5573 1657
rect 5625 1605 5637 1657
rect 5689 1605 5701 1657
rect 5753 1605 5758 1657
rect 5568 1591 5758 1605
rect 5568 1539 5573 1591
rect 5625 1539 5637 1591
rect 5689 1539 5701 1591
rect 5753 1539 5758 1591
rect 5568 1525 5758 1539
rect 5568 1473 5573 1525
rect 5625 1473 5637 1525
rect 5689 1473 5701 1525
rect 5753 1473 5758 1525
rect 5568 1467 5758 1473
rect 6064 4068 6254 4074
rect 6064 4016 6069 4068
rect 6121 4016 6133 4068
rect 6185 4016 6197 4068
rect 6249 4016 6254 4068
rect 6064 4003 6254 4016
rect 6064 3951 6069 4003
rect 6121 3951 6133 4003
rect 6185 3951 6197 4003
rect 6249 3951 6254 4003
rect 6064 3938 6254 3951
rect 6064 3886 6069 3938
rect 6121 3886 6133 3938
rect 6185 3886 6197 3938
rect 6249 3886 6254 3938
rect 6064 3873 6254 3886
rect 6064 3821 6069 3873
rect 6121 3821 6133 3873
rect 6185 3821 6197 3873
rect 6249 3821 6254 3873
rect 6064 3808 6254 3821
rect 6064 3756 6069 3808
rect 6121 3756 6133 3808
rect 6185 3756 6197 3808
rect 6249 3756 6254 3808
rect 6064 3743 6254 3756
rect 6064 3691 6069 3743
rect 6121 3691 6133 3743
rect 6185 3691 6197 3743
rect 6249 3691 6254 3743
rect 6064 3678 6254 3691
rect 6064 3626 6069 3678
rect 6121 3626 6133 3678
rect 6185 3626 6197 3678
rect 6249 3626 6254 3678
rect 6064 3613 6254 3626
rect 6064 3561 6069 3613
rect 6121 3561 6133 3613
rect 6185 3561 6197 3613
rect 6249 3561 6254 3613
rect 6064 3548 6254 3561
rect 6064 3496 6069 3548
rect 6121 3496 6133 3548
rect 6185 3496 6197 3548
rect 6249 3496 6254 3548
rect 6064 3483 6254 3496
rect 6064 3431 6069 3483
rect 6121 3431 6133 3483
rect 6185 3431 6197 3483
rect 6249 3431 6254 3483
rect 6064 3418 6254 3431
rect 6064 3366 6069 3418
rect 6121 3366 6133 3418
rect 6185 3366 6197 3418
rect 6249 3366 6254 3418
rect 6064 3353 6254 3366
rect 6064 3301 6069 3353
rect 6121 3301 6133 3353
rect 6185 3301 6197 3353
rect 6249 3301 6254 3353
rect 6064 3288 6254 3301
rect 6064 3236 6069 3288
rect 6121 3236 6133 3288
rect 6185 3236 6197 3288
rect 6249 3236 6254 3288
rect 6064 3223 6254 3236
rect 6064 3171 6069 3223
rect 6121 3171 6133 3223
rect 6185 3171 6197 3223
rect 6249 3171 6254 3223
rect 6064 3158 6254 3171
rect 6064 3106 6069 3158
rect 6121 3106 6133 3158
rect 6185 3106 6197 3158
rect 6249 3106 6254 3158
rect 6064 3093 6254 3106
rect 6064 3041 6069 3093
rect 6121 3041 6133 3093
rect 6185 3041 6197 3093
rect 6249 3041 6254 3093
rect 6064 3028 6254 3041
rect 6064 2976 6069 3028
rect 6121 2976 6133 3028
rect 6185 2976 6197 3028
rect 6249 2976 6254 3028
rect 6064 2963 6254 2976
rect 6064 2911 6069 2963
rect 6121 2911 6133 2963
rect 6185 2911 6197 2963
rect 6249 2911 6254 2963
rect 6064 2898 6254 2911
rect 6064 2846 6069 2898
rect 6121 2846 6133 2898
rect 6185 2846 6197 2898
rect 6249 2846 6254 2898
rect 6064 2833 6254 2846
rect 6064 2781 6069 2833
rect 6121 2781 6133 2833
rect 6185 2781 6197 2833
rect 6249 2781 6254 2833
rect 6064 2768 6254 2781
rect 6064 2716 6069 2768
rect 6121 2716 6133 2768
rect 6185 2716 6197 2768
rect 6249 2716 6254 2768
rect 6064 2703 6254 2716
rect 6064 2651 6069 2703
rect 6121 2651 6133 2703
rect 6185 2651 6197 2703
rect 6249 2651 6254 2703
rect 6064 2638 6254 2651
rect 6064 2586 6069 2638
rect 6121 2586 6133 2638
rect 6185 2586 6197 2638
rect 6249 2586 6254 2638
rect 6064 2573 6254 2586
rect 6064 2521 6069 2573
rect 6121 2521 6133 2573
rect 6185 2521 6197 2573
rect 6249 2521 6254 2573
rect 6064 2508 6254 2521
rect 6064 2456 6069 2508
rect 6121 2456 6133 2508
rect 6185 2456 6197 2508
rect 6249 2456 6254 2508
rect 6064 2443 6254 2456
rect 6064 2391 6069 2443
rect 6121 2391 6133 2443
rect 6185 2391 6197 2443
rect 6249 2391 6254 2443
rect 6064 2378 6254 2391
rect 6064 2326 6069 2378
rect 6121 2326 6133 2378
rect 6185 2326 6197 2378
rect 6249 2326 6254 2378
rect 6064 2313 6254 2326
rect 6064 2261 6069 2313
rect 6121 2261 6133 2313
rect 6185 2261 6197 2313
rect 6249 2261 6254 2313
rect 6064 2248 6254 2261
rect 6064 2196 6069 2248
rect 6121 2196 6133 2248
rect 6185 2196 6197 2248
rect 6249 2196 6254 2248
rect 6064 2183 6254 2196
rect 6064 2131 6069 2183
rect 6121 2131 6133 2183
rect 6185 2131 6197 2183
rect 6249 2131 6254 2183
rect 6064 2118 6254 2131
rect 6064 2066 6069 2118
rect 6121 2066 6133 2118
rect 6185 2066 6197 2118
rect 6249 2066 6254 2118
rect 6064 2053 6254 2066
rect 6064 2001 6069 2053
rect 6121 2001 6133 2053
rect 6185 2001 6197 2053
rect 6249 2001 6254 2053
rect 6064 1987 6254 2001
rect 6064 1935 6069 1987
rect 6121 1935 6133 1987
rect 6185 1935 6197 1987
rect 6249 1935 6254 1987
rect 6064 1921 6254 1935
rect 6064 1869 6069 1921
rect 6121 1869 6133 1921
rect 6185 1869 6197 1921
rect 6249 1869 6254 1921
rect 6064 1855 6254 1869
rect 6064 1803 6069 1855
rect 6121 1803 6133 1855
rect 6185 1803 6197 1855
rect 6249 1803 6254 1855
rect 6064 1789 6254 1803
rect 6064 1737 6069 1789
rect 6121 1737 6133 1789
rect 6185 1737 6197 1789
rect 6249 1737 6254 1789
rect 6064 1723 6254 1737
rect 6064 1671 6069 1723
rect 6121 1671 6133 1723
rect 6185 1671 6197 1723
rect 6249 1671 6254 1723
rect 6064 1657 6254 1671
rect 6064 1605 6069 1657
rect 6121 1605 6133 1657
rect 6185 1605 6197 1657
rect 6249 1605 6254 1657
rect 6064 1591 6254 1605
rect 6064 1539 6069 1591
rect 6121 1539 6133 1591
rect 6185 1539 6197 1591
rect 6249 1539 6254 1591
rect 6064 1525 6254 1539
rect 6064 1473 6069 1525
rect 6121 1473 6133 1525
rect 6185 1473 6197 1525
rect 6249 1473 6254 1525
rect 6064 1467 6254 1473
rect 6560 4068 6750 4074
rect 6560 4016 6565 4068
rect 6617 4016 6629 4068
rect 6681 4016 6693 4068
rect 6745 4016 6750 4068
rect 6560 4003 6750 4016
rect 6560 3951 6565 4003
rect 6617 3951 6629 4003
rect 6681 3951 6693 4003
rect 6745 3951 6750 4003
rect 6560 3938 6750 3951
rect 6560 3886 6565 3938
rect 6617 3886 6629 3938
rect 6681 3886 6693 3938
rect 6745 3886 6750 3938
rect 6560 3873 6750 3886
rect 6560 3821 6565 3873
rect 6617 3821 6629 3873
rect 6681 3821 6693 3873
rect 6745 3821 6750 3873
rect 6560 3808 6750 3821
rect 6560 3756 6565 3808
rect 6617 3756 6629 3808
rect 6681 3756 6693 3808
rect 6745 3756 6750 3808
rect 6560 3743 6750 3756
rect 6560 3691 6565 3743
rect 6617 3691 6629 3743
rect 6681 3691 6693 3743
rect 6745 3691 6750 3743
rect 6560 3678 6750 3691
rect 6560 3626 6565 3678
rect 6617 3626 6629 3678
rect 6681 3626 6693 3678
rect 6745 3626 6750 3678
rect 6560 3613 6750 3626
rect 6560 3561 6565 3613
rect 6617 3561 6629 3613
rect 6681 3561 6693 3613
rect 6745 3561 6750 3613
rect 6560 3548 6750 3561
rect 6560 3496 6565 3548
rect 6617 3496 6629 3548
rect 6681 3496 6693 3548
rect 6745 3496 6750 3548
rect 6560 3483 6750 3496
rect 6560 3431 6565 3483
rect 6617 3431 6629 3483
rect 6681 3431 6693 3483
rect 6745 3431 6750 3483
rect 6560 3418 6750 3431
rect 6560 3366 6565 3418
rect 6617 3366 6629 3418
rect 6681 3366 6693 3418
rect 6745 3366 6750 3418
rect 6560 3353 6750 3366
rect 6560 3301 6565 3353
rect 6617 3301 6629 3353
rect 6681 3301 6693 3353
rect 6745 3301 6750 3353
rect 6560 3288 6750 3301
rect 6560 3236 6565 3288
rect 6617 3236 6629 3288
rect 6681 3236 6693 3288
rect 6745 3236 6750 3288
rect 6560 3223 6750 3236
rect 6560 3171 6565 3223
rect 6617 3171 6629 3223
rect 6681 3171 6693 3223
rect 6745 3171 6750 3223
rect 6560 3158 6750 3171
rect 6560 3106 6565 3158
rect 6617 3106 6629 3158
rect 6681 3106 6693 3158
rect 6745 3106 6750 3158
rect 6560 3093 6750 3106
rect 6560 3041 6565 3093
rect 6617 3041 6629 3093
rect 6681 3041 6693 3093
rect 6745 3041 6750 3093
rect 6560 3028 6750 3041
rect 6560 2976 6565 3028
rect 6617 2976 6629 3028
rect 6681 2976 6693 3028
rect 6745 2976 6750 3028
rect 6560 2963 6750 2976
rect 6560 2911 6565 2963
rect 6617 2911 6629 2963
rect 6681 2911 6693 2963
rect 6745 2911 6750 2963
rect 6560 2898 6750 2911
rect 6560 2846 6565 2898
rect 6617 2846 6629 2898
rect 6681 2846 6693 2898
rect 6745 2846 6750 2898
rect 6560 2833 6750 2846
rect 6560 2781 6565 2833
rect 6617 2781 6629 2833
rect 6681 2781 6693 2833
rect 6745 2781 6750 2833
rect 6560 2768 6750 2781
rect 6560 2716 6565 2768
rect 6617 2716 6629 2768
rect 6681 2716 6693 2768
rect 6745 2716 6750 2768
rect 6560 2703 6750 2716
rect 6560 2651 6565 2703
rect 6617 2651 6629 2703
rect 6681 2651 6693 2703
rect 6745 2651 6750 2703
rect 6560 2638 6750 2651
rect 6560 2586 6565 2638
rect 6617 2586 6629 2638
rect 6681 2586 6693 2638
rect 6745 2586 6750 2638
rect 6560 2573 6750 2586
rect 6560 2521 6565 2573
rect 6617 2521 6629 2573
rect 6681 2521 6693 2573
rect 6745 2521 6750 2573
rect 6560 2508 6750 2521
rect 6560 2456 6565 2508
rect 6617 2456 6629 2508
rect 6681 2456 6693 2508
rect 6745 2456 6750 2508
rect 6560 2443 6750 2456
rect 6560 2391 6565 2443
rect 6617 2391 6629 2443
rect 6681 2391 6693 2443
rect 6745 2391 6750 2443
rect 6560 2378 6750 2391
rect 6560 2326 6565 2378
rect 6617 2326 6629 2378
rect 6681 2326 6693 2378
rect 6745 2326 6750 2378
rect 6560 2313 6750 2326
rect 6560 2261 6565 2313
rect 6617 2261 6629 2313
rect 6681 2261 6693 2313
rect 6745 2261 6750 2313
rect 6560 2248 6750 2261
rect 6560 2196 6565 2248
rect 6617 2196 6629 2248
rect 6681 2196 6693 2248
rect 6745 2196 6750 2248
rect 6560 2183 6750 2196
rect 6560 2131 6565 2183
rect 6617 2131 6629 2183
rect 6681 2131 6693 2183
rect 6745 2131 6750 2183
rect 6560 2118 6750 2131
rect 6560 2066 6565 2118
rect 6617 2066 6629 2118
rect 6681 2066 6693 2118
rect 6745 2066 6750 2118
rect 6560 2053 6750 2066
rect 6560 2001 6565 2053
rect 6617 2001 6629 2053
rect 6681 2001 6693 2053
rect 6745 2001 6750 2053
rect 6560 1987 6750 2001
rect 6560 1935 6565 1987
rect 6617 1935 6629 1987
rect 6681 1935 6693 1987
rect 6745 1935 6750 1987
rect 6560 1921 6750 1935
rect 6560 1869 6565 1921
rect 6617 1869 6629 1921
rect 6681 1869 6693 1921
rect 6745 1869 6750 1921
rect 6560 1855 6750 1869
rect 6560 1803 6565 1855
rect 6617 1803 6629 1855
rect 6681 1803 6693 1855
rect 6745 1803 6750 1855
rect 6560 1789 6750 1803
rect 6560 1737 6565 1789
rect 6617 1737 6629 1789
rect 6681 1737 6693 1789
rect 6745 1737 6750 1789
rect 6560 1723 6750 1737
rect 6560 1671 6565 1723
rect 6617 1671 6629 1723
rect 6681 1671 6693 1723
rect 6745 1671 6750 1723
rect 6560 1657 6750 1671
rect 6560 1605 6565 1657
rect 6617 1605 6629 1657
rect 6681 1605 6693 1657
rect 6745 1605 6750 1657
rect 6560 1591 6750 1605
rect 6560 1539 6565 1591
rect 6617 1539 6629 1591
rect 6681 1539 6693 1591
rect 6745 1539 6750 1591
rect 6560 1525 6750 1539
rect 6560 1473 6565 1525
rect 6617 1473 6629 1525
rect 6681 1473 6693 1525
rect 6745 1473 6750 1525
rect 6560 1467 6750 1473
rect 7056 4068 7246 4074
rect 7056 4016 7061 4068
rect 7113 4016 7125 4068
rect 7177 4016 7189 4068
rect 7241 4016 7246 4068
rect 7056 4003 7246 4016
rect 7056 3951 7061 4003
rect 7113 3951 7125 4003
rect 7177 3951 7189 4003
rect 7241 3951 7246 4003
rect 7056 3938 7246 3951
rect 7056 3886 7061 3938
rect 7113 3886 7125 3938
rect 7177 3886 7189 3938
rect 7241 3886 7246 3938
rect 7056 3873 7246 3886
rect 7056 3821 7061 3873
rect 7113 3821 7125 3873
rect 7177 3821 7189 3873
rect 7241 3821 7246 3873
rect 7056 3808 7246 3821
rect 7056 3756 7061 3808
rect 7113 3756 7125 3808
rect 7177 3756 7189 3808
rect 7241 3756 7246 3808
rect 7056 3743 7246 3756
rect 7056 3691 7061 3743
rect 7113 3691 7125 3743
rect 7177 3691 7189 3743
rect 7241 3691 7246 3743
rect 7056 3678 7246 3691
rect 7056 3626 7061 3678
rect 7113 3626 7125 3678
rect 7177 3626 7189 3678
rect 7241 3626 7246 3678
rect 7056 3613 7246 3626
rect 7056 3561 7061 3613
rect 7113 3561 7125 3613
rect 7177 3561 7189 3613
rect 7241 3561 7246 3613
rect 7056 3548 7246 3561
rect 7056 3496 7061 3548
rect 7113 3496 7125 3548
rect 7177 3496 7189 3548
rect 7241 3496 7246 3548
rect 7056 3483 7246 3496
rect 7056 3431 7061 3483
rect 7113 3431 7125 3483
rect 7177 3431 7189 3483
rect 7241 3431 7246 3483
rect 7056 3418 7246 3431
rect 7056 3366 7061 3418
rect 7113 3366 7125 3418
rect 7177 3366 7189 3418
rect 7241 3366 7246 3418
rect 7056 3353 7246 3366
rect 7056 3301 7061 3353
rect 7113 3301 7125 3353
rect 7177 3301 7189 3353
rect 7241 3301 7246 3353
rect 7056 3288 7246 3301
rect 7056 3236 7061 3288
rect 7113 3236 7125 3288
rect 7177 3236 7189 3288
rect 7241 3236 7246 3288
rect 7056 3223 7246 3236
rect 7056 3171 7061 3223
rect 7113 3171 7125 3223
rect 7177 3171 7189 3223
rect 7241 3171 7246 3223
rect 7056 3158 7246 3171
rect 7056 3106 7061 3158
rect 7113 3106 7125 3158
rect 7177 3106 7189 3158
rect 7241 3106 7246 3158
rect 7056 3093 7246 3106
rect 7056 3041 7061 3093
rect 7113 3041 7125 3093
rect 7177 3041 7189 3093
rect 7241 3041 7246 3093
rect 7056 3028 7246 3041
rect 7056 2976 7061 3028
rect 7113 2976 7125 3028
rect 7177 2976 7189 3028
rect 7241 2976 7246 3028
rect 7056 2963 7246 2976
rect 7056 2911 7061 2963
rect 7113 2911 7125 2963
rect 7177 2911 7189 2963
rect 7241 2911 7246 2963
rect 7056 2898 7246 2911
rect 7056 2846 7061 2898
rect 7113 2846 7125 2898
rect 7177 2846 7189 2898
rect 7241 2846 7246 2898
rect 7056 2833 7246 2846
rect 7056 2781 7061 2833
rect 7113 2781 7125 2833
rect 7177 2781 7189 2833
rect 7241 2781 7246 2833
rect 7056 2768 7246 2781
rect 7056 2716 7061 2768
rect 7113 2716 7125 2768
rect 7177 2716 7189 2768
rect 7241 2716 7246 2768
rect 7056 2703 7246 2716
rect 7056 2651 7061 2703
rect 7113 2651 7125 2703
rect 7177 2651 7189 2703
rect 7241 2651 7246 2703
rect 7056 2638 7246 2651
rect 7056 2586 7061 2638
rect 7113 2586 7125 2638
rect 7177 2586 7189 2638
rect 7241 2586 7246 2638
rect 7056 2573 7246 2586
rect 7056 2521 7061 2573
rect 7113 2521 7125 2573
rect 7177 2521 7189 2573
rect 7241 2521 7246 2573
rect 7056 2508 7246 2521
rect 7056 2456 7061 2508
rect 7113 2456 7125 2508
rect 7177 2456 7189 2508
rect 7241 2456 7246 2508
rect 7056 2443 7246 2456
rect 7056 2391 7061 2443
rect 7113 2391 7125 2443
rect 7177 2391 7189 2443
rect 7241 2391 7246 2443
rect 7056 2378 7246 2391
rect 7056 2326 7061 2378
rect 7113 2326 7125 2378
rect 7177 2326 7189 2378
rect 7241 2326 7246 2378
rect 7056 2313 7246 2326
rect 7056 2261 7061 2313
rect 7113 2261 7125 2313
rect 7177 2261 7189 2313
rect 7241 2261 7246 2313
rect 7056 2248 7246 2261
rect 7056 2196 7061 2248
rect 7113 2196 7125 2248
rect 7177 2196 7189 2248
rect 7241 2196 7246 2248
rect 7056 2183 7246 2196
rect 7056 2131 7061 2183
rect 7113 2131 7125 2183
rect 7177 2131 7189 2183
rect 7241 2131 7246 2183
rect 7056 2118 7246 2131
rect 7056 2066 7061 2118
rect 7113 2066 7125 2118
rect 7177 2066 7189 2118
rect 7241 2066 7246 2118
rect 7056 2053 7246 2066
rect 7056 2001 7061 2053
rect 7113 2001 7125 2053
rect 7177 2001 7189 2053
rect 7241 2001 7246 2053
rect 7056 1987 7246 2001
rect 7056 1935 7061 1987
rect 7113 1935 7125 1987
rect 7177 1935 7189 1987
rect 7241 1935 7246 1987
rect 7056 1921 7246 1935
rect 7056 1869 7061 1921
rect 7113 1869 7125 1921
rect 7177 1869 7189 1921
rect 7241 1869 7246 1921
rect 7056 1855 7246 1869
rect 7056 1803 7061 1855
rect 7113 1803 7125 1855
rect 7177 1803 7189 1855
rect 7241 1803 7246 1855
rect 7056 1789 7246 1803
rect 7056 1737 7061 1789
rect 7113 1737 7125 1789
rect 7177 1737 7189 1789
rect 7241 1737 7246 1789
rect 7056 1723 7246 1737
rect 7056 1671 7061 1723
rect 7113 1671 7125 1723
rect 7177 1671 7189 1723
rect 7241 1671 7246 1723
rect 7056 1657 7246 1671
rect 7056 1605 7061 1657
rect 7113 1605 7125 1657
rect 7177 1605 7189 1657
rect 7241 1605 7246 1657
rect 7056 1591 7246 1605
rect 7056 1539 7061 1591
rect 7113 1539 7125 1591
rect 7177 1539 7189 1591
rect 7241 1539 7246 1591
rect 7056 1525 7246 1539
rect 7056 1473 7061 1525
rect 7113 1473 7125 1525
rect 7177 1473 7189 1525
rect 7241 1473 7246 1525
rect 7056 1467 7246 1473
rect 7552 4068 7742 4074
rect 7552 4016 7557 4068
rect 7609 4016 7621 4068
rect 7673 4016 7685 4068
rect 7737 4016 7742 4068
rect 7552 4003 7742 4016
rect 7552 3951 7557 4003
rect 7609 3951 7621 4003
rect 7673 3951 7685 4003
rect 7737 3951 7742 4003
rect 7552 3938 7742 3951
rect 7552 3886 7557 3938
rect 7609 3886 7621 3938
rect 7673 3886 7685 3938
rect 7737 3886 7742 3938
rect 7552 3873 7742 3886
rect 7552 3821 7557 3873
rect 7609 3821 7621 3873
rect 7673 3821 7685 3873
rect 7737 3821 7742 3873
rect 7552 3808 7742 3821
rect 7552 3756 7557 3808
rect 7609 3756 7621 3808
rect 7673 3756 7685 3808
rect 7737 3756 7742 3808
rect 7552 3743 7742 3756
rect 7552 3691 7557 3743
rect 7609 3691 7621 3743
rect 7673 3691 7685 3743
rect 7737 3691 7742 3743
rect 7552 3678 7742 3691
rect 7552 3626 7557 3678
rect 7609 3626 7621 3678
rect 7673 3626 7685 3678
rect 7737 3626 7742 3678
rect 7552 3613 7742 3626
rect 7552 3561 7557 3613
rect 7609 3561 7621 3613
rect 7673 3561 7685 3613
rect 7737 3561 7742 3613
rect 7552 3548 7742 3561
rect 7552 3496 7557 3548
rect 7609 3496 7621 3548
rect 7673 3496 7685 3548
rect 7737 3496 7742 3548
rect 7552 3483 7742 3496
rect 7552 3431 7557 3483
rect 7609 3431 7621 3483
rect 7673 3431 7685 3483
rect 7737 3431 7742 3483
rect 7552 3418 7742 3431
rect 7552 3366 7557 3418
rect 7609 3366 7621 3418
rect 7673 3366 7685 3418
rect 7737 3366 7742 3418
rect 7552 3353 7742 3366
rect 7552 3301 7557 3353
rect 7609 3301 7621 3353
rect 7673 3301 7685 3353
rect 7737 3301 7742 3353
rect 7552 3288 7742 3301
rect 7552 3236 7557 3288
rect 7609 3236 7621 3288
rect 7673 3236 7685 3288
rect 7737 3236 7742 3288
rect 7552 3223 7742 3236
rect 7552 3171 7557 3223
rect 7609 3171 7621 3223
rect 7673 3171 7685 3223
rect 7737 3171 7742 3223
rect 7552 3158 7742 3171
rect 7552 3106 7557 3158
rect 7609 3106 7621 3158
rect 7673 3106 7685 3158
rect 7737 3106 7742 3158
rect 7552 3093 7742 3106
rect 7552 3041 7557 3093
rect 7609 3041 7621 3093
rect 7673 3041 7685 3093
rect 7737 3041 7742 3093
rect 7552 3028 7742 3041
rect 7552 2976 7557 3028
rect 7609 2976 7621 3028
rect 7673 2976 7685 3028
rect 7737 2976 7742 3028
rect 7552 2963 7742 2976
rect 7552 2911 7557 2963
rect 7609 2911 7621 2963
rect 7673 2911 7685 2963
rect 7737 2911 7742 2963
rect 7552 2898 7742 2911
rect 7552 2846 7557 2898
rect 7609 2846 7621 2898
rect 7673 2846 7685 2898
rect 7737 2846 7742 2898
rect 7552 2833 7742 2846
rect 7552 2781 7557 2833
rect 7609 2781 7621 2833
rect 7673 2781 7685 2833
rect 7737 2781 7742 2833
rect 7552 2768 7742 2781
rect 7552 2716 7557 2768
rect 7609 2716 7621 2768
rect 7673 2716 7685 2768
rect 7737 2716 7742 2768
rect 7552 2703 7742 2716
rect 7552 2651 7557 2703
rect 7609 2651 7621 2703
rect 7673 2651 7685 2703
rect 7737 2651 7742 2703
rect 7552 2638 7742 2651
rect 7552 2586 7557 2638
rect 7609 2586 7621 2638
rect 7673 2586 7685 2638
rect 7737 2586 7742 2638
rect 7552 2573 7742 2586
rect 7552 2521 7557 2573
rect 7609 2521 7621 2573
rect 7673 2521 7685 2573
rect 7737 2521 7742 2573
rect 7552 2508 7742 2521
rect 7552 2456 7557 2508
rect 7609 2456 7621 2508
rect 7673 2456 7685 2508
rect 7737 2456 7742 2508
rect 7552 2443 7742 2456
rect 7552 2391 7557 2443
rect 7609 2391 7621 2443
rect 7673 2391 7685 2443
rect 7737 2391 7742 2443
rect 7552 2378 7742 2391
rect 7552 2326 7557 2378
rect 7609 2326 7621 2378
rect 7673 2326 7685 2378
rect 7737 2326 7742 2378
rect 7552 2313 7742 2326
rect 7552 2261 7557 2313
rect 7609 2261 7621 2313
rect 7673 2261 7685 2313
rect 7737 2261 7742 2313
rect 7552 2248 7742 2261
rect 7552 2196 7557 2248
rect 7609 2196 7621 2248
rect 7673 2196 7685 2248
rect 7737 2196 7742 2248
rect 7552 2183 7742 2196
rect 7552 2131 7557 2183
rect 7609 2131 7621 2183
rect 7673 2131 7685 2183
rect 7737 2131 7742 2183
rect 7552 2118 7742 2131
rect 7552 2066 7557 2118
rect 7609 2066 7621 2118
rect 7673 2066 7685 2118
rect 7737 2066 7742 2118
rect 7552 2053 7742 2066
rect 7552 2001 7557 2053
rect 7609 2001 7621 2053
rect 7673 2001 7685 2053
rect 7737 2001 7742 2053
rect 7552 1987 7742 2001
rect 7552 1935 7557 1987
rect 7609 1935 7621 1987
rect 7673 1935 7685 1987
rect 7737 1935 7742 1987
rect 7552 1921 7742 1935
rect 7552 1869 7557 1921
rect 7609 1869 7621 1921
rect 7673 1869 7685 1921
rect 7737 1869 7742 1921
rect 7552 1855 7742 1869
rect 7552 1803 7557 1855
rect 7609 1803 7621 1855
rect 7673 1803 7685 1855
rect 7737 1803 7742 1855
rect 7552 1789 7742 1803
rect 7552 1737 7557 1789
rect 7609 1737 7621 1789
rect 7673 1737 7685 1789
rect 7737 1737 7742 1789
rect 7552 1723 7742 1737
rect 7552 1671 7557 1723
rect 7609 1671 7621 1723
rect 7673 1671 7685 1723
rect 7737 1671 7742 1723
rect 7552 1657 7742 1671
rect 7552 1605 7557 1657
rect 7609 1605 7621 1657
rect 7673 1605 7685 1657
rect 7737 1605 7742 1657
rect 7552 1591 7742 1605
rect 7552 1539 7557 1591
rect 7609 1539 7621 1591
rect 7673 1539 7685 1591
rect 7737 1539 7742 1591
rect 7552 1525 7742 1539
rect 7552 1473 7557 1525
rect 7609 1473 7621 1525
rect 7673 1473 7685 1525
rect 7737 1473 7742 1525
rect 7552 1467 7742 1473
rect 8048 4068 8238 4074
rect 8048 4016 8053 4068
rect 8105 4016 8117 4068
rect 8169 4016 8181 4068
rect 8233 4016 8238 4068
rect 8048 4003 8238 4016
rect 8048 3951 8053 4003
rect 8105 3951 8117 4003
rect 8169 3951 8181 4003
rect 8233 3951 8238 4003
rect 8048 3938 8238 3951
rect 8048 3886 8053 3938
rect 8105 3886 8117 3938
rect 8169 3886 8181 3938
rect 8233 3886 8238 3938
rect 8048 3873 8238 3886
rect 8048 3821 8053 3873
rect 8105 3821 8117 3873
rect 8169 3821 8181 3873
rect 8233 3821 8238 3873
rect 8048 3808 8238 3821
rect 8048 3756 8053 3808
rect 8105 3756 8117 3808
rect 8169 3756 8181 3808
rect 8233 3756 8238 3808
rect 8048 3743 8238 3756
rect 8048 3691 8053 3743
rect 8105 3691 8117 3743
rect 8169 3691 8181 3743
rect 8233 3691 8238 3743
rect 8048 3678 8238 3691
rect 8048 3626 8053 3678
rect 8105 3626 8117 3678
rect 8169 3626 8181 3678
rect 8233 3626 8238 3678
rect 8048 3613 8238 3626
rect 8048 3561 8053 3613
rect 8105 3561 8117 3613
rect 8169 3561 8181 3613
rect 8233 3561 8238 3613
rect 8048 3548 8238 3561
rect 8048 3496 8053 3548
rect 8105 3496 8117 3548
rect 8169 3496 8181 3548
rect 8233 3496 8238 3548
rect 8048 3483 8238 3496
rect 8048 3431 8053 3483
rect 8105 3431 8117 3483
rect 8169 3431 8181 3483
rect 8233 3431 8238 3483
rect 8048 3418 8238 3431
rect 8048 3366 8053 3418
rect 8105 3366 8117 3418
rect 8169 3366 8181 3418
rect 8233 3366 8238 3418
rect 8048 3353 8238 3366
rect 8048 3301 8053 3353
rect 8105 3301 8117 3353
rect 8169 3301 8181 3353
rect 8233 3301 8238 3353
rect 8048 3288 8238 3301
rect 8048 3236 8053 3288
rect 8105 3236 8117 3288
rect 8169 3236 8181 3288
rect 8233 3236 8238 3288
rect 8048 3223 8238 3236
rect 8048 3171 8053 3223
rect 8105 3171 8117 3223
rect 8169 3171 8181 3223
rect 8233 3171 8238 3223
rect 8048 3158 8238 3171
rect 8048 3106 8053 3158
rect 8105 3106 8117 3158
rect 8169 3106 8181 3158
rect 8233 3106 8238 3158
rect 8048 3093 8238 3106
rect 8048 3041 8053 3093
rect 8105 3041 8117 3093
rect 8169 3041 8181 3093
rect 8233 3041 8238 3093
rect 8048 3028 8238 3041
rect 8048 2976 8053 3028
rect 8105 2976 8117 3028
rect 8169 2976 8181 3028
rect 8233 2976 8238 3028
rect 8048 2963 8238 2976
rect 8048 2911 8053 2963
rect 8105 2911 8117 2963
rect 8169 2911 8181 2963
rect 8233 2911 8238 2963
rect 8048 2898 8238 2911
rect 8048 2846 8053 2898
rect 8105 2846 8117 2898
rect 8169 2846 8181 2898
rect 8233 2846 8238 2898
rect 8048 2833 8238 2846
rect 8048 2781 8053 2833
rect 8105 2781 8117 2833
rect 8169 2781 8181 2833
rect 8233 2781 8238 2833
rect 8048 2768 8238 2781
rect 8048 2716 8053 2768
rect 8105 2716 8117 2768
rect 8169 2716 8181 2768
rect 8233 2716 8238 2768
rect 8048 2703 8238 2716
rect 8048 2651 8053 2703
rect 8105 2651 8117 2703
rect 8169 2651 8181 2703
rect 8233 2651 8238 2703
rect 8048 2638 8238 2651
rect 8048 2586 8053 2638
rect 8105 2586 8117 2638
rect 8169 2586 8181 2638
rect 8233 2586 8238 2638
rect 8048 2573 8238 2586
rect 8048 2521 8053 2573
rect 8105 2521 8117 2573
rect 8169 2521 8181 2573
rect 8233 2521 8238 2573
rect 8048 2508 8238 2521
rect 8048 2456 8053 2508
rect 8105 2456 8117 2508
rect 8169 2456 8181 2508
rect 8233 2456 8238 2508
rect 8048 2443 8238 2456
rect 8048 2391 8053 2443
rect 8105 2391 8117 2443
rect 8169 2391 8181 2443
rect 8233 2391 8238 2443
rect 8048 2378 8238 2391
rect 8048 2326 8053 2378
rect 8105 2326 8117 2378
rect 8169 2326 8181 2378
rect 8233 2326 8238 2378
rect 8048 2313 8238 2326
rect 8048 2261 8053 2313
rect 8105 2261 8117 2313
rect 8169 2261 8181 2313
rect 8233 2261 8238 2313
rect 8048 2248 8238 2261
rect 8048 2196 8053 2248
rect 8105 2196 8117 2248
rect 8169 2196 8181 2248
rect 8233 2196 8238 2248
rect 8048 2183 8238 2196
rect 8048 2131 8053 2183
rect 8105 2131 8117 2183
rect 8169 2131 8181 2183
rect 8233 2131 8238 2183
rect 8048 2118 8238 2131
rect 8048 2066 8053 2118
rect 8105 2066 8117 2118
rect 8169 2066 8181 2118
rect 8233 2066 8238 2118
rect 8048 2053 8238 2066
rect 8048 2001 8053 2053
rect 8105 2001 8117 2053
rect 8169 2001 8181 2053
rect 8233 2001 8238 2053
rect 8048 1987 8238 2001
rect 8048 1935 8053 1987
rect 8105 1935 8117 1987
rect 8169 1935 8181 1987
rect 8233 1935 8238 1987
rect 8048 1921 8238 1935
rect 8048 1869 8053 1921
rect 8105 1869 8117 1921
rect 8169 1869 8181 1921
rect 8233 1869 8238 1921
rect 8048 1855 8238 1869
rect 8048 1803 8053 1855
rect 8105 1803 8117 1855
rect 8169 1803 8181 1855
rect 8233 1803 8238 1855
rect 8048 1789 8238 1803
rect 8048 1737 8053 1789
rect 8105 1737 8117 1789
rect 8169 1737 8181 1789
rect 8233 1737 8238 1789
rect 8048 1723 8238 1737
rect 8048 1671 8053 1723
rect 8105 1671 8117 1723
rect 8169 1671 8181 1723
rect 8233 1671 8238 1723
rect 8048 1657 8238 1671
rect 8048 1605 8053 1657
rect 8105 1605 8117 1657
rect 8169 1605 8181 1657
rect 8233 1605 8238 1657
rect 8048 1591 8238 1605
rect 8048 1539 8053 1591
rect 8105 1539 8117 1591
rect 8169 1539 8181 1591
rect 8233 1539 8238 1591
rect 8048 1525 8238 1539
rect 8048 1473 8053 1525
rect 8105 1473 8117 1525
rect 8169 1473 8181 1525
rect 8233 1473 8238 1525
rect 8048 1467 8238 1473
rect 8544 4068 8734 4074
rect 8544 4016 8549 4068
rect 8601 4016 8613 4068
rect 8665 4016 8677 4068
rect 8729 4016 8734 4068
rect 8544 4003 8734 4016
rect 8544 3951 8549 4003
rect 8601 3951 8613 4003
rect 8665 3951 8677 4003
rect 8729 3951 8734 4003
rect 8544 3938 8734 3951
rect 8544 3886 8549 3938
rect 8601 3886 8613 3938
rect 8665 3886 8677 3938
rect 8729 3886 8734 3938
rect 8544 3873 8734 3886
rect 8544 3821 8549 3873
rect 8601 3821 8613 3873
rect 8665 3821 8677 3873
rect 8729 3821 8734 3873
rect 8544 3808 8734 3821
rect 8544 3756 8549 3808
rect 8601 3756 8613 3808
rect 8665 3756 8677 3808
rect 8729 3756 8734 3808
rect 8544 3743 8734 3756
rect 8544 3691 8549 3743
rect 8601 3691 8613 3743
rect 8665 3691 8677 3743
rect 8729 3691 8734 3743
rect 8544 3678 8734 3691
rect 8544 3626 8549 3678
rect 8601 3626 8613 3678
rect 8665 3626 8677 3678
rect 8729 3626 8734 3678
rect 8544 3613 8734 3626
rect 8544 3561 8549 3613
rect 8601 3561 8613 3613
rect 8665 3561 8677 3613
rect 8729 3561 8734 3613
rect 8544 3548 8734 3561
rect 8544 3496 8549 3548
rect 8601 3496 8613 3548
rect 8665 3496 8677 3548
rect 8729 3496 8734 3548
rect 8544 3483 8734 3496
rect 8544 3431 8549 3483
rect 8601 3431 8613 3483
rect 8665 3431 8677 3483
rect 8729 3431 8734 3483
rect 8544 3418 8734 3431
rect 8544 3366 8549 3418
rect 8601 3366 8613 3418
rect 8665 3366 8677 3418
rect 8729 3366 8734 3418
rect 8544 3353 8734 3366
rect 8544 3301 8549 3353
rect 8601 3301 8613 3353
rect 8665 3301 8677 3353
rect 8729 3301 8734 3353
rect 8544 3288 8734 3301
rect 8544 3236 8549 3288
rect 8601 3236 8613 3288
rect 8665 3236 8677 3288
rect 8729 3236 8734 3288
rect 8544 3223 8734 3236
rect 8544 3171 8549 3223
rect 8601 3171 8613 3223
rect 8665 3171 8677 3223
rect 8729 3171 8734 3223
rect 8544 3158 8734 3171
rect 8544 3106 8549 3158
rect 8601 3106 8613 3158
rect 8665 3106 8677 3158
rect 8729 3106 8734 3158
rect 8544 3093 8734 3106
rect 8544 3041 8549 3093
rect 8601 3041 8613 3093
rect 8665 3041 8677 3093
rect 8729 3041 8734 3093
rect 8544 3028 8734 3041
rect 8544 2976 8549 3028
rect 8601 2976 8613 3028
rect 8665 2976 8677 3028
rect 8729 2976 8734 3028
rect 8544 2963 8734 2976
rect 8544 2911 8549 2963
rect 8601 2911 8613 2963
rect 8665 2911 8677 2963
rect 8729 2911 8734 2963
rect 8544 2898 8734 2911
rect 8544 2846 8549 2898
rect 8601 2846 8613 2898
rect 8665 2846 8677 2898
rect 8729 2846 8734 2898
rect 8544 2833 8734 2846
rect 8544 2781 8549 2833
rect 8601 2781 8613 2833
rect 8665 2781 8677 2833
rect 8729 2781 8734 2833
rect 8544 2768 8734 2781
rect 8544 2716 8549 2768
rect 8601 2716 8613 2768
rect 8665 2716 8677 2768
rect 8729 2716 8734 2768
rect 8544 2703 8734 2716
rect 8544 2651 8549 2703
rect 8601 2651 8613 2703
rect 8665 2651 8677 2703
rect 8729 2651 8734 2703
rect 8544 2638 8734 2651
rect 8544 2586 8549 2638
rect 8601 2586 8613 2638
rect 8665 2586 8677 2638
rect 8729 2586 8734 2638
rect 8544 2573 8734 2586
rect 8544 2521 8549 2573
rect 8601 2521 8613 2573
rect 8665 2521 8677 2573
rect 8729 2521 8734 2573
rect 8544 2508 8734 2521
rect 8544 2456 8549 2508
rect 8601 2456 8613 2508
rect 8665 2456 8677 2508
rect 8729 2456 8734 2508
rect 8544 2443 8734 2456
rect 8544 2391 8549 2443
rect 8601 2391 8613 2443
rect 8665 2391 8677 2443
rect 8729 2391 8734 2443
rect 8544 2378 8734 2391
rect 8544 2326 8549 2378
rect 8601 2326 8613 2378
rect 8665 2326 8677 2378
rect 8729 2326 8734 2378
rect 8544 2313 8734 2326
rect 8544 2261 8549 2313
rect 8601 2261 8613 2313
rect 8665 2261 8677 2313
rect 8729 2261 8734 2313
rect 8544 2248 8734 2261
rect 8544 2196 8549 2248
rect 8601 2196 8613 2248
rect 8665 2196 8677 2248
rect 8729 2196 8734 2248
rect 8544 2183 8734 2196
rect 8544 2131 8549 2183
rect 8601 2131 8613 2183
rect 8665 2131 8677 2183
rect 8729 2131 8734 2183
rect 8544 2118 8734 2131
rect 8544 2066 8549 2118
rect 8601 2066 8613 2118
rect 8665 2066 8677 2118
rect 8729 2066 8734 2118
rect 8544 2053 8734 2066
rect 8544 2001 8549 2053
rect 8601 2001 8613 2053
rect 8665 2001 8677 2053
rect 8729 2001 8734 2053
rect 8544 1987 8734 2001
rect 8544 1935 8549 1987
rect 8601 1935 8613 1987
rect 8665 1935 8677 1987
rect 8729 1935 8734 1987
rect 8544 1921 8734 1935
rect 8544 1869 8549 1921
rect 8601 1869 8613 1921
rect 8665 1869 8677 1921
rect 8729 1869 8734 1921
rect 8544 1855 8734 1869
rect 8544 1803 8549 1855
rect 8601 1803 8613 1855
rect 8665 1803 8677 1855
rect 8729 1803 8734 1855
rect 8544 1789 8734 1803
rect 8544 1737 8549 1789
rect 8601 1737 8613 1789
rect 8665 1737 8677 1789
rect 8729 1737 8734 1789
rect 8544 1723 8734 1737
rect 8544 1671 8549 1723
rect 8601 1671 8613 1723
rect 8665 1671 8677 1723
rect 8729 1671 8734 1723
rect 8544 1657 8734 1671
rect 8544 1605 8549 1657
rect 8601 1605 8613 1657
rect 8665 1605 8677 1657
rect 8729 1605 8734 1657
rect 8544 1591 8734 1605
rect 8544 1539 8549 1591
rect 8601 1539 8613 1591
rect 8665 1539 8677 1591
rect 8729 1539 8734 1591
rect 8544 1525 8734 1539
rect 8544 1473 8549 1525
rect 8601 1473 8613 1525
rect 8665 1473 8677 1525
rect 8729 1473 8734 1525
rect 8544 1467 8734 1473
rect 9040 4068 9230 4074
rect 9040 4016 9045 4068
rect 9097 4016 9109 4068
rect 9161 4016 9173 4068
rect 9225 4016 9230 4068
rect 9040 4003 9230 4016
rect 9040 3951 9045 4003
rect 9097 3951 9109 4003
rect 9161 3951 9173 4003
rect 9225 3951 9230 4003
rect 9040 3938 9230 3951
rect 9040 3886 9045 3938
rect 9097 3886 9109 3938
rect 9161 3886 9173 3938
rect 9225 3886 9230 3938
rect 9040 3873 9230 3886
rect 9040 3821 9045 3873
rect 9097 3821 9109 3873
rect 9161 3821 9173 3873
rect 9225 3821 9230 3873
rect 9040 3808 9230 3821
rect 9040 3756 9045 3808
rect 9097 3756 9109 3808
rect 9161 3756 9173 3808
rect 9225 3756 9230 3808
rect 9040 3743 9230 3756
rect 9040 3691 9045 3743
rect 9097 3691 9109 3743
rect 9161 3691 9173 3743
rect 9225 3691 9230 3743
rect 9040 3678 9230 3691
rect 9040 3626 9045 3678
rect 9097 3626 9109 3678
rect 9161 3626 9173 3678
rect 9225 3626 9230 3678
rect 9040 3613 9230 3626
rect 9040 3561 9045 3613
rect 9097 3561 9109 3613
rect 9161 3561 9173 3613
rect 9225 3561 9230 3613
rect 9040 3548 9230 3561
rect 9040 3496 9045 3548
rect 9097 3496 9109 3548
rect 9161 3496 9173 3548
rect 9225 3496 9230 3548
rect 9040 3483 9230 3496
rect 9040 3431 9045 3483
rect 9097 3431 9109 3483
rect 9161 3431 9173 3483
rect 9225 3431 9230 3483
rect 9040 3418 9230 3431
rect 9040 3366 9045 3418
rect 9097 3366 9109 3418
rect 9161 3366 9173 3418
rect 9225 3366 9230 3418
rect 9040 3353 9230 3366
rect 9040 3301 9045 3353
rect 9097 3301 9109 3353
rect 9161 3301 9173 3353
rect 9225 3301 9230 3353
rect 9040 3288 9230 3301
rect 9040 3236 9045 3288
rect 9097 3236 9109 3288
rect 9161 3236 9173 3288
rect 9225 3236 9230 3288
rect 9040 3223 9230 3236
rect 9040 3171 9045 3223
rect 9097 3171 9109 3223
rect 9161 3171 9173 3223
rect 9225 3171 9230 3223
rect 9040 3158 9230 3171
rect 9040 3106 9045 3158
rect 9097 3106 9109 3158
rect 9161 3106 9173 3158
rect 9225 3106 9230 3158
rect 9040 3093 9230 3106
rect 9040 3041 9045 3093
rect 9097 3041 9109 3093
rect 9161 3041 9173 3093
rect 9225 3041 9230 3093
rect 9040 3028 9230 3041
rect 9040 2976 9045 3028
rect 9097 2976 9109 3028
rect 9161 2976 9173 3028
rect 9225 2976 9230 3028
rect 9040 2963 9230 2976
rect 9040 2911 9045 2963
rect 9097 2911 9109 2963
rect 9161 2911 9173 2963
rect 9225 2911 9230 2963
rect 9040 2898 9230 2911
rect 9040 2846 9045 2898
rect 9097 2846 9109 2898
rect 9161 2846 9173 2898
rect 9225 2846 9230 2898
rect 9040 2833 9230 2846
rect 9040 2781 9045 2833
rect 9097 2781 9109 2833
rect 9161 2781 9173 2833
rect 9225 2781 9230 2833
rect 9040 2768 9230 2781
rect 9040 2716 9045 2768
rect 9097 2716 9109 2768
rect 9161 2716 9173 2768
rect 9225 2716 9230 2768
rect 9040 2703 9230 2716
rect 9040 2651 9045 2703
rect 9097 2651 9109 2703
rect 9161 2651 9173 2703
rect 9225 2651 9230 2703
rect 9040 2638 9230 2651
rect 9040 2586 9045 2638
rect 9097 2586 9109 2638
rect 9161 2586 9173 2638
rect 9225 2586 9230 2638
rect 9040 2573 9230 2586
rect 9040 2521 9045 2573
rect 9097 2521 9109 2573
rect 9161 2521 9173 2573
rect 9225 2521 9230 2573
rect 9040 2508 9230 2521
rect 9040 2456 9045 2508
rect 9097 2456 9109 2508
rect 9161 2456 9173 2508
rect 9225 2456 9230 2508
rect 9040 2443 9230 2456
rect 9040 2391 9045 2443
rect 9097 2391 9109 2443
rect 9161 2391 9173 2443
rect 9225 2391 9230 2443
rect 9040 2378 9230 2391
rect 9040 2326 9045 2378
rect 9097 2326 9109 2378
rect 9161 2326 9173 2378
rect 9225 2326 9230 2378
rect 9040 2313 9230 2326
rect 9040 2261 9045 2313
rect 9097 2261 9109 2313
rect 9161 2261 9173 2313
rect 9225 2261 9230 2313
rect 9040 2248 9230 2261
rect 9040 2196 9045 2248
rect 9097 2196 9109 2248
rect 9161 2196 9173 2248
rect 9225 2196 9230 2248
rect 9040 2183 9230 2196
rect 9040 2131 9045 2183
rect 9097 2131 9109 2183
rect 9161 2131 9173 2183
rect 9225 2131 9230 2183
rect 9040 2118 9230 2131
rect 9040 2066 9045 2118
rect 9097 2066 9109 2118
rect 9161 2066 9173 2118
rect 9225 2066 9230 2118
rect 9040 2053 9230 2066
rect 9040 2001 9045 2053
rect 9097 2001 9109 2053
rect 9161 2001 9173 2053
rect 9225 2001 9230 2053
rect 9040 1987 9230 2001
rect 9040 1935 9045 1987
rect 9097 1935 9109 1987
rect 9161 1935 9173 1987
rect 9225 1935 9230 1987
rect 9040 1921 9230 1935
rect 9040 1869 9045 1921
rect 9097 1869 9109 1921
rect 9161 1869 9173 1921
rect 9225 1869 9230 1921
rect 9040 1855 9230 1869
rect 9040 1803 9045 1855
rect 9097 1803 9109 1855
rect 9161 1803 9173 1855
rect 9225 1803 9230 1855
rect 9040 1789 9230 1803
rect 9040 1737 9045 1789
rect 9097 1737 9109 1789
rect 9161 1737 9173 1789
rect 9225 1737 9230 1789
rect 9040 1723 9230 1737
rect 9040 1671 9045 1723
rect 9097 1671 9109 1723
rect 9161 1671 9173 1723
rect 9225 1671 9230 1723
rect 9040 1657 9230 1671
rect 9040 1605 9045 1657
rect 9097 1605 9109 1657
rect 9161 1605 9173 1657
rect 9225 1605 9230 1657
rect 9040 1591 9230 1605
rect 9040 1539 9045 1591
rect 9097 1539 9109 1591
rect 9161 1539 9173 1591
rect 9225 1539 9230 1591
rect 9040 1525 9230 1539
rect 9040 1473 9045 1525
rect 9097 1473 9109 1525
rect 9161 1473 9173 1525
rect 9225 1473 9230 1525
rect 9040 1467 9230 1473
rect 9536 4068 9726 4074
rect 9536 4016 9541 4068
rect 9593 4016 9605 4068
rect 9657 4016 9669 4068
rect 9721 4016 9726 4068
rect 9536 4003 9726 4016
rect 9536 3951 9541 4003
rect 9593 3951 9605 4003
rect 9657 3951 9669 4003
rect 9721 3951 9726 4003
rect 9536 3938 9726 3951
rect 9536 3886 9541 3938
rect 9593 3886 9605 3938
rect 9657 3886 9669 3938
rect 9721 3886 9726 3938
rect 9536 3873 9726 3886
rect 9536 3821 9541 3873
rect 9593 3821 9605 3873
rect 9657 3821 9669 3873
rect 9721 3821 9726 3873
rect 9536 3808 9726 3821
rect 9536 3756 9541 3808
rect 9593 3756 9605 3808
rect 9657 3756 9669 3808
rect 9721 3756 9726 3808
rect 9536 3743 9726 3756
rect 9536 3691 9541 3743
rect 9593 3691 9605 3743
rect 9657 3691 9669 3743
rect 9721 3691 9726 3743
rect 9536 3678 9726 3691
rect 9536 3626 9541 3678
rect 9593 3626 9605 3678
rect 9657 3626 9669 3678
rect 9721 3626 9726 3678
rect 9536 3613 9726 3626
rect 9536 3561 9541 3613
rect 9593 3561 9605 3613
rect 9657 3561 9669 3613
rect 9721 3561 9726 3613
rect 9536 3548 9726 3561
rect 9536 3496 9541 3548
rect 9593 3496 9605 3548
rect 9657 3496 9669 3548
rect 9721 3496 9726 3548
rect 9536 3483 9726 3496
rect 9536 3431 9541 3483
rect 9593 3431 9605 3483
rect 9657 3431 9669 3483
rect 9721 3431 9726 3483
rect 9536 3418 9726 3431
rect 9536 3366 9541 3418
rect 9593 3366 9605 3418
rect 9657 3366 9669 3418
rect 9721 3366 9726 3418
rect 9536 3353 9726 3366
rect 9536 3301 9541 3353
rect 9593 3301 9605 3353
rect 9657 3301 9669 3353
rect 9721 3301 9726 3353
rect 9536 3288 9726 3301
rect 9536 3236 9541 3288
rect 9593 3236 9605 3288
rect 9657 3236 9669 3288
rect 9721 3236 9726 3288
rect 9536 3223 9726 3236
rect 9536 3171 9541 3223
rect 9593 3171 9605 3223
rect 9657 3171 9669 3223
rect 9721 3171 9726 3223
rect 9536 3158 9726 3171
rect 9536 3106 9541 3158
rect 9593 3106 9605 3158
rect 9657 3106 9669 3158
rect 9721 3106 9726 3158
rect 9536 3093 9726 3106
rect 9536 3041 9541 3093
rect 9593 3041 9605 3093
rect 9657 3041 9669 3093
rect 9721 3041 9726 3093
rect 9536 3028 9726 3041
rect 9536 2976 9541 3028
rect 9593 2976 9605 3028
rect 9657 2976 9669 3028
rect 9721 2976 9726 3028
rect 9536 2963 9726 2976
rect 9536 2911 9541 2963
rect 9593 2911 9605 2963
rect 9657 2911 9669 2963
rect 9721 2911 9726 2963
rect 9536 2898 9726 2911
rect 9536 2846 9541 2898
rect 9593 2846 9605 2898
rect 9657 2846 9669 2898
rect 9721 2846 9726 2898
rect 9536 2833 9726 2846
rect 9536 2781 9541 2833
rect 9593 2781 9605 2833
rect 9657 2781 9669 2833
rect 9721 2781 9726 2833
rect 9536 2768 9726 2781
rect 9536 2716 9541 2768
rect 9593 2716 9605 2768
rect 9657 2716 9669 2768
rect 9721 2716 9726 2768
rect 9536 2703 9726 2716
rect 9536 2651 9541 2703
rect 9593 2651 9605 2703
rect 9657 2651 9669 2703
rect 9721 2651 9726 2703
rect 9536 2638 9726 2651
rect 9536 2586 9541 2638
rect 9593 2586 9605 2638
rect 9657 2586 9669 2638
rect 9721 2586 9726 2638
rect 9536 2573 9726 2586
rect 9536 2521 9541 2573
rect 9593 2521 9605 2573
rect 9657 2521 9669 2573
rect 9721 2521 9726 2573
rect 9536 2508 9726 2521
rect 9536 2456 9541 2508
rect 9593 2456 9605 2508
rect 9657 2456 9669 2508
rect 9721 2456 9726 2508
rect 9536 2443 9726 2456
rect 9536 2391 9541 2443
rect 9593 2391 9605 2443
rect 9657 2391 9669 2443
rect 9721 2391 9726 2443
rect 9536 2378 9726 2391
rect 9536 2326 9541 2378
rect 9593 2326 9605 2378
rect 9657 2326 9669 2378
rect 9721 2326 9726 2378
rect 9536 2313 9726 2326
rect 9536 2261 9541 2313
rect 9593 2261 9605 2313
rect 9657 2261 9669 2313
rect 9721 2261 9726 2313
rect 9536 2248 9726 2261
rect 9536 2196 9541 2248
rect 9593 2196 9605 2248
rect 9657 2196 9669 2248
rect 9721 2196 9726 2248
rect 9536 2183 9726 2196
rect 9536 2131 9541 2183
rect 9593 2131 9605 2183
rect 9657 2131 9669 2183
rect 9721 2131 9726 2183
rect 9536 2118 9726 2131
rect 9536 2066 9541 2118
rect 9593 2066 9605 2118
rect 9657 2066 9669 2118
rect 9721 2066 9726 2118
rect 9536 2053 9726 2066
rect 9536 2001 9541 2053
rect 9593 2001 9605 2053
rect 9657 2001 9669 2053
rect 9721 2001 9726 2053
rect 9536 1987 9726 2001
rect 9536 1935 9541 1987
rect 9593 1935 9605 1987
rect 9657 1935 9669 1987
rect 9721 1935 9726 1987
rect 9536 1921 9726 1935
rect 9536 1869 9541 1921
rect 9593 1869 9605 1921
rect 9657 1869 9669 1921
rect 9721 1869 9726 1921
rect 9536 1855 9726 1869
rect 9536 1803 9541 1855
rect 9593 1803 9605 1855
rect 9657 1803 9669 1855
rect 9721 1803 9726 1855
rect 9536 1789 9726 1803
rect 9536 1737 9541 1789
rect 9593 1737 9605 1789
rect 9657 1737 9669 1789
rect 9721 1737 9726 1789
rect 9536 1723 9726 1737
rect 9536 1671 9541 1723
rect 9593 1671 9605 1723
rect 9657 1671 9669 1723
rect 9721 1671 9726 1723
rect 9536 1657 9726 1671
rect 9536 1605 9541 1657
rect 9593 1605 9605 1657
rect 9657 1605 9669 1657
rect 9721 1605 9726 1657
rect 9536 1591 9726 1605
rect 9536 1539 9541 1591
rect 9593 1539 9605 1591
rect 9657 1539 9669 1591
rect 9721 1539 9726 1591
rect 9536 1525 9726 1539
rect 9536 1473 9541 1525
rect 9593 1473 9605 1525
rect 9657 1473 9669 1525
rect 9721 1473 9726 1525
rect 9536 1467 9726 1473
rect 10032 4068 10222 4074
rect 10032 4016 10037 4068
rect 10089 4016 10101 4068
rect 10153 4016 10165 4068
rect 10217 4016 10222 4068
rect 10032 4003 10222 4016
rect 10032 3951 10037 4003
rect 10089 3951 10101 4003
rect 10153 3951 10165 4003
rect 10217 3951 10222 4003
rect 10032 3938 10222 3951
rect 10032 3886 10037 3938
rect 10089 3886 10101 3938
rect 10153 3886 10165 3938
rect 10217 3886 10222 3938
rect 10032 3873 10222 3886
rect 10032 3821 10037 3873
rect 10089 3821 10101 3873
rect 10153 3821 10165 3873
rect 10217 3821 10222 3873
rect 10032 3808 10222 3821
rect 10032 3756 10037 3808
rect 10089 3756 10101 3808
rect 10153 3756 10165 3808
rect 10217 3756 10222 3808
rect 10032 3743 10222 3756
rect 10032 3691 10037 3743
rect 10089 3691 10101 3743
rect 10153 3691 10165 3743
rect 10217 3691 10222 3743
rect 10032 3678 10222 3691
rect 10032 3626 10037 3678
rect 10089 3626 10101 3678
rect 10153 3626 10165 3678
rect 10217 3626 10222 3678
rect 10032 3613 10222 3626
rect 10032 3561 10037 3613
rect 10089 3561 10101 3613
rect 10153 3561 10165 3613
rect 10217 3561 10222 3613
rect 10032 3548 10222 3561
rect 10032 3496 10037 3548
rect 10089 3496 10101 3548
rect 10153 3496 10165 3548
rect 10217 3496 10222 3548
rect 10032 3483 10222 3496
rect 10032 3431 10037 3483
rect 10089 3431 10101 3483
rect 10153 3431 10165 3483
rect 10217 3431 10222 3483
rect 10032 3418 10222 3431
rect 10032 3366 10037 3418
rect 10089 3366 10101 3418
rect 10153 3366 10165 3418
rect 10217 3366 10222 3418
rect 10032 3353 10222 3366
rect 10032 3301 10037 3353
rect 10089 3301 10101 3353
rect 10153 3301 10165 3353
rect 10217 3301 10222 3353
rect 10032 3288 10222 3301
rect 10032 3236 10037 3288
rect 10089 3236 10101 3288
rect 10153 3236 10165 3288
rect 10217 3236 10222 3288
rect 10032 3223 10222 3236
rect 10032 3171 10037 3223
rect 10089 3171 10101 3223
rect 10153 3171 10165 3223
rect 10217 3171 10222 3223
rect 10032 3158 10222 3171
rect 10032 3106 10037 3158
rect 10089 3106 10101 3158
rect 10153 3106 10165 3158
rect 10217 3106 10222 3158
rect 10032 3093 10222 3106
rect 10032 3041 10037 3093
rect 10089 3041 10101 3093
rect 10153 3041 10165 3093
rect 10217 3041 10222 3093
rect 10032 3028 10222 3041
rect 10032 2976 10037 3028
rect 10089 2976 10101 3028
rect 10153 2976 10165 3028
rect 10217 2976 10222 3028
rect 10032 2963 10222 2976
rect 10032 2911 10037 2963
rect 10089 2911 10101 2963
rect 10153 2911 10165 2963
rect 10217 2911 10222 2963
rect 10032 2898 10222 2911
rect 10032 2846 10037 2898
rect 10089 2846 10101 2898
rect 10153 2846 10165 2898
rect 10217 2846 10222 2898
rect 10032 2833 10222 2846
rect 10032 2781 10037 2833
rect 10089 2781 10101 2833
rect 10153 2781 10165 2833
rect 10217 2781 10222 2833
rect 10032 2768 10222 2781
rect 10032 2716 10037 2768
rect 10089 2716 10101 2768
rect 10153 2716 10165 2768
rect 10217 2716 10222 2768
rect 10032 2703 10222 2716
rect 10032 2651 10037 2703
rect 10089 2651 10101 2703
rect 10153 2651 10165 2703
rect 10217 2651 10222 2703
rect 10032 2638 10222 2651
rect 10032 2586 10037 2638
rect 10089 2586 10101 2638
rect 10153 2586 10165 2638
rect 10217 2586 10222 2638
rect 10032 2573 10222 2586
rect 10032 2521 10037 2573
rect 10089 2521 10101 2573
rect 10153 2521 10165 2573
rect 10217 2521 10222 2573
rect 10032 2508 10222 2521
rect 10032 2456 10037 2508
rect 10089 2456 10101 2508
rect 10153 2456 10165 2508
rect 10217 2456 10222 2508
rect 10032 2443 10222 2456
rect 10032 2391 10037 2443
rect 10089 2391 10101 2443
rect 10153 2391 10165 2443
rect 10217 2391 10222 2443
rect 10032 2378 10222 2391
rect 10032 2326 10037 2378
rect 10089 2326 10101 2378
rect 10153 2326 10165 2378
rect 10217 2326 10222 2378
rect 10032 2313 10222 2326
rect 10032 2261 10037 2313
rect 10089 2261 10101 2313
rect 10153 2261 10165 2313
rect 10217 2261 10222 2313
rect 10032 2248 10222 2261
rect 10032 2196 10037 2248
rect 10089 2196 10101 2248
rect 10153 2196 10165 2248
rect 10217 2196 10222 2248
rect 10032 2183 10222 2196
rect 10032 2131 10037 2183
rect 10089 2131 10101 2183
rect 10153 2131 10165 2183
rect 10217 2131 10222 2183
rect 10032 2118 10222 2131
rect 10032 2066 10037 2118
rect 10089 2066 10101 2118
rect 10153 2066 10165 2118
rect 10217 2066 10222 2118
rect 10032 2053 10222 2066
rect 10032 2001 10037 2053
rect 10089 2001 10101 2053
rect 10153 2001 10165 2053
rect 10217 2001 10222 2053
rect 10032 1987 10222 2001
rect 10032 1935 10037 1987
rect 10089 1935 10101 1987
rect 10153 1935 10165 1987
rect 10217 1935 10222 1987
rect 10032 1921 10222 1935
rect 10032 1869 10037 1921
rect 10089 1869 10101 1921
rect 10153 1869 10165 1921
rect 10217 1869 10222 1921
rect 10032 1855 10222 1869
rect 10032 1803 10037 1855
rect 10089 1803 10101 1855
rect 10153 1803 10165 1855
rect 10217 1803 10222 1855
rect 10032 1789 10222 1803
rect 10032 1737 10037 1789
rect 10089 1737 10101 1789
rect 10153 1737 10165 1789
rect 10217 1737 10222 1789
rect 10032 1723 10222 1737
rect 10032 1671 10037 1723
rect 10089 1671 10101 1723
rect 10153 1671 10165 1723
rect 10217 1671 10222 1723
rect 10032 1657 10222 1671
rect 10032 1605 10037 1657
rect 10089 1605 10101 1657
rect 10153 1605 10165 1657
rect 10217 1605 10222 1657
rect 10032 1591 10222 1605
rect 10032 1539 10037 1591
rect 10089 1539 10101 1591
rect 10153 1539 10165 1591
rect 10217 1539 10222 1591
rect 10032 1525 10222 1539
rect 10032 1473 10037 1525
rect 10089 1473 10101 1525
rect 10153 1473 10165 1525
rect 10217 1473 10222 1525
rect 10032 1467 10222 1473
rect 10528 4068 10718 4074
rect 10528 4016 10533 4068
rect 10585 4016 10597 4068
rect 10649 4016 10661 4068
rect 10713 4016 10718 4068
rect 10528 4003 10718 4016
rect 10528 3951 10533 4003
rect 10585 3951 10597 4003
rect 10649 3951 10661 4003
rect 10713 3951 10718 4003
rect 10528 3938 10718 3951
rect 10528 3886 10533 3938
rect 10585 3886 10597 3938
rect 10649 3886 10661 3938
rect 10713 3886 10718 3938
rect 10528 3873 10718 3886
rect 10528 3821 10533 3873
rect 10585 3821 10597 3873
rect 10649 3821 10661 3873
rect 10713 3821 10718 3873
rect 10528 3808 10718 3821
rect 10528 3756 10533 3808
rect 10585 3756 10597 3808
rect 10649 3756 10661 3808
rect 10713 3756 10718 3808
rect 10528 3743 10718 3756
rect 10528 3691 10533 3743
rect 10585 3691 10597 3743
rect 10649 3691 10661 3743
rect 10713 3691 10718 3743
rect 10528 3678 10718 3691
rect 10528 3626 10533 3678
rect 10585 3626 10597 3678
rect 10649 3626 10661 3678
rect 10713 3626 10718 3678
rect 10528 3613 10718 3626
rect 10528 3561 10533 3613
rect 10585 3561 10597 3613
rect 10649 3561 10661 3613
rect 10713 3561 10718 3613
rect 10528 3548 10718 3561
rect 10528 3496 10533 3548
rect 10585 3496 10597 3548
rect 10649 3496 10661 3548
rect 10713 3496 10718 3548
rect 10528 3483 10718 3496
rect 10528 3431 10533 3483
rect 10585 3431 10597 3483
rect 10649 3431 10661 3483
rect 10713 3431 10718 3483
rect 10528 3418 10718 3431
rect 10528 3366 10533 3418
rect 10585 3366 10597 3418
rect 10649 3366 10661 3418
rect 10713 3366 10718 3418
rect 10528 3353 10718 3366
rect 10528 3301 10533 3353
rect 10585 3301 10597 3353
rect 10649 3301 10661 3353
rect 10713 3301 10718 3353
rect 10528 3288 10718 3301
rect 10528 3236 10533 3288
rect 10585 3236 10597 3288
rect 10649 3236 10661 3288
rect 10713 3236 10718 3288
rect 10528 3223 10718 3236
rect 10528 3171 10533 3223
rect 10585 3171 10597 3223
rect 10649 3171 10661 3223
rect 10713 3171 10718 3223
rect 10528 3158 10718 3171
rect 10528 3106 10533 3158
rect 10585 3106 10597 3158
rect 10649 3106 10661 3158
rect 10713 3106 10718 3158
rect 10528 3093 10718 3106
rect 10528 3041 10533 3093
rect 10585 3041 10597 3093
rect 10649 3041 10661 3093
rect 10713 3041 10718 3093
rect 10528 3028 10718 3041
rect 10528 2976 10533 3028
rect 10585 2976 10597 3028
rect 10649 2976 10661 3028
rect 10713 2976 10718 3028
rect 10528 2963 10718 2976
rect 10528 2911 10533 2963
rect 10585 2911 10597 2963
rect 10649 2911 10661 2963
rect 10713 2911 10718 2963
rect 10528 2898 10718 2911
rect 10528 2846 10533 2898
rect 10585 2846 10597 2898
rect 10649 2846 10661 2898
rect 10713 2846 10718 2898
rect 10528 2833 10718 2846
rect 10528 2781 10533 2833
rect 10585 2781 10597 2833
rect 10649 2781 10661 2833
rect 10713 2781 10718 2833
rect 10528 2768 10718 2781
rect 10528 2716 10533 2768
rect 10585 2716 10597 2768
rect 10649 2716 10661 2768
rect 10713 2716 10718 2768
rect 10528 2703 10718 2716
rect 10528 2651 10533 2703
rect 10585 2651 10597 2703
rect 10649 2651 10661 2703
rect 10713 2651 10718 2703
rect 10528 2638 10718 2651
rect 10528 2586 10533 2638
rect 10585 2586 10597 2638
rect 10649 2586 10661 2638
rect 10713 2586 10718 2638
rect 10528 2573 10718 2586
rect 10528 2521 10533 2573
rect 10585 2521 10597 2573
rect 10649 2521 10661 2573
rect 10713 2521 10718 2573
rect 10528 2508 10718 2521
rect 10528 2456 10533 2508
rect 10585 2456 10597 2508
rect 10649 2456 10661 2508
rect 10713 2456 10718 2508
rect 10528 2443 10718 2456
rect 10528 2391 10533 2443
rect 10585 2391 10597 2443
rect 10649 2391 10661 2443
rect 10713 2391 10718 2443
rect 10528 2378 10718 2391
rect 10528 2326 10533 2378
rect 10585 2326 10597 2378
rect 10649 2326 10661 2378
rect 10713 2326 10718 2378
rect 10528 2313 10718 2326
rect 10528 2261 10533 2313
rect 10585 2261 10597 2313
rect 10649 2261 10661 2313
rect 10713 2261 10718 2313
rect 10528 2248 10718 2261
rect 10528 2196 10533 2248
rect 10585 2196 10597 2248
rect 10649 2196 10661 2248
rect 10713 2196 10718 2248
rect 10528 2183 10718 2196
rect 10528 2131 10533 2183
rect 10585 2131 10597 2183
rect 10649 2131 10661 2183
rect 10713 2131 10718 2183
rect 10528 2118 10718 2131
rect 10528 2066 10533 2118
rect 10585 2066 10597 2118
rect 10649 2066 10661 2118
rect 10713 2066 10718 2118
rect 10528 2053 10718 2066
rect 10528 2001 10533 2053
rect 10585 2001 10597 2053
rect 10649 2001 10661 2053
rect 10713 2001 10718 2053
rect 10528 1987 10718 2001
rect 10528 1935 10533 1987
rect 10585 1935 10597 1987
rect 10649 1935 10661 1987
rect 10713 1935 10718 1987
rect 10528 1921 10718 1935
rect 10528 1869 10533 1921
rect 10585 1869 10597 1921
rect 10649 1869 10661 1921
rect 10713 1869 10718 1921
rect 10528 1855 10718 1869
rect 10528 1803 10533 1855
rect 10585 1803 10597 1855
rect 10649 1803 10661 1855
rect 10713 1803 10718 1855
rect 10528 1789 10718 1803
rect 10528 1737 10533 1789
rect 10585 1737 10597 1789
rect 10649 1737 10661 1789
rect 10713 1737 10718 1789
rect 10528 1723 10718 1737
rect 10528 1671 10533 1723
rect 10585 1671 10597 1723
rect 10649 1671 10661 1723
rect 10713 1671 10718 1723
rect 10528 1657 10718 1671
rect 10528 1605 10533 1657
rect 10585 1605 10597 1657
rect 10649 1605 10661 1657
rect 10713 1605 10718 1657
rect 10528 1591 10718 1605
rect 10528 1539 10533 1591
rect 10585 1539 10597 1591
rect 10649 1539 10661 1591
rect 10713 1539 10718 1591
rect 10528 1525 10718 1539
rect 10528 1473 10533 1525
rect 10585 1473 10597 1525
rect 10649 1473 10661 1525
rect 10713 1473 10718 1525
rect 10528 1467 10718 1473
rect 11024 4068 11214 4074
rect 11024 4016 11029 4068
rect 11081 4016 11093 4068
rect 11145 4016 11157 4068
rect 11209 4016 11214 4068
rect 11024 4003 11214 4016
rect 11024 3951 11029 4003
rect 11081 3951 11093 4003
rect 11145 3951 11157 4003
rect 11209 3951 11214 4003
rect 11024 3938 11214 3951
rect 11024 3886 11029 3938
rect 11081 3886 11093 3938
rect 11145 3886 11157 3938
rect 11209 3886 11214 3938
rect 11024 3873 11214 3886
rect 11024 3821 11029 3873
rect 11081 3821 11093 3873
rect 11145 3821 11157 3873
rect 11209 3821 11214 3873
rect 11024 3808 11214 3821
rect 11024 3756 11029 3808
rect 11081 3756 11093 3808
rect 11145 3756 11157 3808
rect 11209 3756 11214 3808
rect 11024 3743 11214 3756
rect 11024 3691 11029 3743
rect 11081 3691 11093 3743
rect 11145 3691 11157 3743
rect 11209 3691 11214 3743
rect 11024 3678 11214 3691
rect 11024 3626 11029 3678
rect 11081 3626 11093 3678
rect 11145 3626 11157 3678
rect 11209 3626 11214 3678
rect 11024 3613 11214 3626
rect 11024 3561 11029 3613
rect 11081 3561 11093 3613
rect 11145 3561 11157 3613
rect 11209 3561 11214 3613
rect 11024 3548 11214 3561
rect 11024 3496 11029 3548
rect 11081 3496 11093 3548
rect 11145 3496 11157 3548
rect 11209 3496 11214 3548
rect 11024 3483 11214 3496
rect 11024 3431 11029 3483
rect 11081 3431 11093 3483
rect 11145 3431 11157 3483
rect 11209 3431 11214 3483
rect 11024 3418 11214 3431
rect 11024 3366 11029 3418
rect 11081 3366 11093 3418
rect 11145 3366 11157 3418
rect 11209 3366 11214 3418
rect 11024 3353 11214 3366
rect 11024 3301 11029 3353
rect 11081 3301 11093 3353
rect 11145 3301 11157 3353
rect 11209 3301 11214 3353
rect 11024 3288 11214 3301
rect 11024 3236 11029 3288
rect 11081 3236 11093 3288
rect 11145 3236 11157 3288
rect 11209 3236 11214 3288
rect 11024 3223 11214 3236
rect 11024 3171 11029 3223
rect 11081 3171 11093 3223
rect 11145 3171 11157 3223
rect 11209 3171 11214 3223
rect 11024 3158 11214 3171
rect 11024 3106 11029 3158
rect 11081 3106 11093 3158
rect 11145 3106 11157 3158
rect 11209 3106 11214 3158
rect 11024 3093 11214 3106
rect 11024 3041 11029 3093
rect 11081 3041 11093 3093
rect 11145 3041 11157 3093
rect 11209 3041 11214 3093
rect 11024 3028 11214 3041
rect 11024 2976 11029 3028
rect 11081 2976 11093 3028
rect 11145 2976 11157 3028
rect 11209 2976 11214 3028
rect 11024 2963 11214 2976
rect 11024 2911 11029 2963
rect 11081 2911 11093 2963
rect 11145 2911 11157 2963
rect 11209 2911 11214 2963
rect 11024 2898 11214 2911
rect 11024 2846 11029 2898
rect 11081 2846 11093 2898
rect 11145 2846 11157 2898
rect 11209 2846 11214 2898
rect 11024 2833 11214 2846
rect 11024 2781 11029 2833
rect 11081 2781 11093 2833
rect 11145 2781 11157 2833
rect 11209 2781 11214 2833
rect 11024 2768 11214 2781
rect 11024 2716 11029 2768
rect 11081 2716 11093 2768
rect 11145 2716 11157 2768
rect 11209 2716 11214 2768
rect 11024 2703 11214 2716
rect 11024 2651 11029 2703
rect 11081 2651 11093 2703
rect 11145 2651 11157 2703
rect 11209 2651 11214 2703
rect 11024 2638 11214 2651
rect 11024 2586 11029 2638
rect 11081 2586 11093 2638
rect 11145 2586 11157 2638
rect 11209 2586 11214 2638
rect 11024 2573 11214 2586
rect 11024 2521 11029 2573
rect 11081 2521 11093 2573
rect 11145 2521 11157 2573
rect 11209 2521 11214 2573
rect 11024 2508 11214 2521
rect 11024 2456 11029 2508
rect 11081 2456 11093 2508
rect 11145 2456 11157 2508
rect 11209 2456 11214 2508
rect 11024 2443 11214 2456
rect 11024 2391 11029 2443
rect 11081 2391 11093 2443
rect 11145 2391 11157 2443
rect 11209 2391 11214 2443
rect 11024 2378 11214 2391
rect 11024 2326 11029 2378
rect 11081 2326 11093 2378
rect 11145 2326 11157 2378
rect 11209 2326 11214 2378
rect 11024 2313 11214 2326
rect 11024 2261 11029 2313
rect 11081 2261 11093 2313
rect 11145 2261 11157 2313
rect 11209 2261 11214 2313
rect 11024 2248 11214 2261
rect 11024 2196 11029 2248
rect 11081 2196 11093 2248
rect 11145 2196 11157 2248
rect 11209 2196 11214 2248
rect 11024 2183 11214 2196
rect 11024 2131 11029 2183
rect 11081 2131 11093 2183
rect 11145 2131 11157 2183
rect 11209 2131 11214 2183
rect 11024 2118 11214 2131
rect 11024 2066 11029 2118
rect 11081 2066 11093 2118
rect 11145 2066 11157 2118
rect 11209 2066 11214 2118
rect 11024 2053 11214 2066
rect 11024 2001 11029 2053
rect 11081 2001 11093 2053
rect 11145 2001 11157 2053
rect 11209 2001 11214 2053
rect 11024 1987 11214 2001
rect 11024 1935 11029 1987
rect 11081 1935 11093 1987
rect 11145 1935 11157 1987
rect 11209 1935 11214 1987
rect 11024 1921 11214 1935
rect 11024 1869 11029 1921
rect 11081 1869 11093 1921
rect 11145 1869 11157 1921
rect 11209 1869 11214 1921
rect 11024 1855 11214 1869
rect 11024 1803 11029 1855
rect 11081 1803 11093 1855
rect 11145 1803 11157 1855
rect 11209 1803 11214 1855
rect 11024 1789 11214 1803
rect 11024 1737 11029 1789
rect 11081 1737 11093 1789
rect 11145 1737 11157 1789
rect 11209 1737 11214 1789
rect 11024 1723 11214 1737
rect 11024 1671 11029 1723
rect 11081 1671 11093 1723
rect 11145 1671 11157 1723
rect 11209 1671 11214 1723
rect 11024 1657 11214 1671
rect 11024 1605 11029 1657
rect 11081 1605 11093 1657
rect 11145 1605 11157 1657
rect 11209 1605 11214 1657
rect 11024 1591 11214 1605
rect 11024 1539 11029 1591
rect 11081 1539 11093 1591
rect 11145 1539 11157 1591
rect 11209 1539 11214 1591
rect 11024 1525 11214 1539
rect 11024 1473 11029 1525
rect 11081 1473 11093 1525
rect 11145 1473 11157 1525
rect 11209 1473 11214 1525
rect 11024 1467 11214 1473
rect 11520 4068 11710 4074
rect 11520 4016 11525 4068
rect 11577 4016 11589 4068
rect 11641 4016 11653 4068
rect 11705 4016 11710 4068
rect 11520 4003 11710 4016
rect 11520 3951 11525 4003
rect 11577 3951 11589 4003
rect 11641 3951 11653 4003
rect 11705 3951 11710 4003
rect 11520 3938 11710 3951
rect 11520 3886 11525 3938
rect 11577 3886 11589 3938
rect 11641 3886 11653 3938
rect 11705 3886 11710 3938
rect 11520 3873 11710 3886
rect 11520 3821 11525 3873
rect 11577 3821 11589 3873
rect 11641 3821 11653 3873
rect 11705 3821 11710 3873
rect 11520 3808 11710 3821
rect 11520 3756 11525 3808
rect 11577 3756 11589 3808
rect 11641 3756 11653 3808
rect 11705 3756 11710 3808
rect 11520 3743 11710 3756
rect 11520 3691 11525 3743
rect 11577 3691 11589 3743
rect 11641 3691 11653 3743
rect 11705 3691 11710 3743
rect 11520 3678 11710 3691
rect 11520 3626 11525 3678
rect 11577 3626 11589 3678
rect 11641 3626 11653 3678
rect 11705 3626 11710 3678
rect 11520 3613 11710 3626
rect 11520 3561 11525 3613
rect 11577 3561 11589 3613
rect 11641 3561 11653 3613
rect 11705 3561 11710 3613
rect 11520 3548 11710 3561
rect 11520 3496 11525 3548
rect 11577 3496 11589 3548
rect 11641 3496 11653 3548
rect 11705 3496 11710 3548
rect 11520 3483 11710 3496
rect 11520 3431 11525 3483
rect 11577 3431 11589 3483
rect 11641 3431 11653 3483
rect 11705 3431 11710 3483
rect 11520 3418 11710 3431
rect 11520 3366 11525 3418
rect 11577 3366 11589 3418
rect 11641 3366 11653 3418
rect 11705 3366 11710 3418
rect 11520 3353 11710 3366
rect 11520 3301 11525 3353
rect 11577 3301 11589 3353
rect 11641 3301 11653 3353
rect 11705 3301 11710 3353
rect 11520 3288 11710 3301
rect 11520 3236 11525 3288
rect 11577 3236 11589 3288
rect 11641 3236 11653 3288
rect 11705 3236 11710 3288
rect 11520 3223 11710 3236
rect 11520 3171 11525 3223
rect 11577 3171 11589 3223
rect 11641 3171 11653 3223
rect 11705 3171 11710 3223
rect 11520 3158 11710 3171
rect 11520 3106 11525 3158
rect 11577 3106 11589 3158
rect 11641 3106 11653 3158
rect 11705 3106 11710 3158
rect 11520 3093 11710 3106
rect 11520 3041 11525 3093
rect 11577 3041 11589 3093
rect 11641 3041 11653 3093
rect 11705 3041 11710 3093
rect 11520 3028 11710 3041
rect 11520 2976 11525 3028
rect 11577 2976 11589 3028
rect 11641 2976 11653 3028
rect 11705 2976 11710 3028
rect 11520 2963 11710 2976
rect 11520 2911 11525 2963
rect 11577 2911 11589 2963
rect 11641 2911 11653 2963
rect 11705 2911 11710 2963
rect 11520 2898 11710 2911
rect 11520 2846 11525 2898
rect 11577 2846 11589 2898
rect 11641 2846 11653 2898
rect 11705 2846 11710 2898
rect 11520 2833 11710 2846
rect 11520 2781 11525 2833
rect 11577 2781 11589 2833
rect 11641 2781 11653 2833
rect 11705 2781 11710 2833
rect 11520 2768 11710 2781
rect 11520 2716 11525 2768
rect 11577 2716 11589 2768
rect 11641 2716 11653 2768
rect 11705 2716 11710 2768
rect 11520 2703 11710 2716
rect 11520 2651 11525 2703
rect 11577 2651 11589 2703
rect 11641 2651 11653 2703
rect 11705 2651 11710 2703
rect 11520 2638 11710 2651
rect 11520 2586 11525 2638
rect 11577 2586 11589 2638
rect 11641 2586 11653 2638
rect 11705 2586 11710 2638
rect 11520 2573 11710 2586
rect 11520 2521 11525 2573
rect 11577 2521 11589 2573
rect 11641 2521 11653 2573
rect 11705 2521 11710 2573
rect 11520 2508 11710 2521
rect 11520 2456 11525 2508
rect 11577 2456 11589 2508
rect 11641 2456 11653 2508
rect 11705 2456 11710 2508
rect 11520 2443 11710 2456
rect 11520 2391 11525 2443
rect 11577 2391 11589 2443
rect 11641 2391 11653 2443
rect 11705 2391 11710 2443
rect 11520 2378 11710 2391
rect 11520 2326 11525 2378
rect 11577 2326 11589 2378
rect 11641 2326 11653 2378
rect 11705 2326 11710 2378
rect 11520 2313 11710 2326
rect 11520 2261 11525 2313
rect 11577 2261 11589 2313
rect 11641 2261 11653 2313
rect 11705 2261 11710 2313
rect 11520 2248 11710 2261
rect 11520 2196 11525 2248
rect 11577 2196 11589 2248
rect 11641 2196 11653 2248
rect 11705 2196 11710 2248
rect 11520 2183 11710 2196
rect 11520 2131 11525 2183
rect 11577 2131 11589 2183
rect 11641 2131 11653 2183
rect 11705 2131 11710 2183
rect 11520 2118 11710 2131
rect 11520 2066 11525 2118
rect 11577 2066 11589 2118
rect 11641 2066 11653 2118
rect 11705 2066 11710 2118
rect 11520 2053 11710 2066
rect 11520 2001 11525 2053
rect 11577 2001 11589 2053
rect 11641 2001 11653 2053
rect 11705 2001 11710 2053
rect 11520 1987 11710 2001
rect 11520 1935 11525 1987
rect 11577 1935 11589 1987
rect 11641 1935 11653 1987
rect 11705 1935 11710 1987
rect 11520 1921 11710 1935
rect 11520 1869 11525 1921
rect 11577 1869 11589 1921
rect 11641 1869 11653 1921
rect 11705 1869 11710 1921
rect 11520 1855 11710 1869
rect 11520 1803 11525 1855
rect 11577 1803 11589 1855
rect 11641 1803 11653 1855
rect 11705 1803 11710 1855
rect 11520 1789 11710 1803
rect 11520 1737 11525 1789
rect 11577 1737 11589 1789
rect 11641 1737 11653 1789
rect 11705 1737 11710 1789
rect 11520 1723 11710 1737
rect 11520 1671 11525 1723
rect 11577 1671 11589 1723
rect 11641 1671 11653 1723
rect 11705 1671 11710 1723
rect 11520 1657 11710 1671
rect 11520 1605 11525 1657
rect 11577 1605 11589 1657
rect 11641 1605 11653 1657
rect 11705 1605 11710 1657
rect 11520 1591 11710 1605
rect 11520 1539 11525 1591
rect 11577 1539 11589 1591
rect 11641 1539 11653 1591
rect 11705 1539 11710 1591
rect 11520 1525 11710 1539
rect 11520 1473 11525 1525
rect 11577 1473 11589 1525
rect 11641 1473 11653 1525
rect 11705 1473 11710 1525
rect 11520 1467 11710 1473
rect 12016 4068 12206 4074
rect 12016 4016 12021 4068
rect 12073 4016 12085 4068
rect 12137 4016 12149 4068
rect 12201 4016 12206 4068
rect 12016 4003 12206 4016
rect 12016 3951 12021 4003
rect 12073 3951 12085 4003
rect 12137 3951 12149 4003
rect 12201 3951 12206 4003
rect 12016 3938 12206 3951
rect 12016 3886 12021 3938
rect 12073 3886 12085 3938
rect 12137 3886 12149 3938
rect 12201 3886 12206 3938
rect 12016 3873 12206 3886
rect 12016 3821 12021 3873
rect 12073 3821 12085 3873
rect 12137 3821 12149 3873
rect 12201 3821 12206 3873
rect 12016 3808 12206 3821
rect 12016 3756 12021 3808
rect 12073 3756 12085 3808
rect 12137 3756 12149 3808
rect 12201 3756 12206 3808
rect 12016 3743 12206 3756
rect 12016 3691 12021 3743
rect 12073 3691 12085 3743
rect 12137 3691 12149 3743
rect 12201 3691 12206 3743
rect 12016 3678 12206 3691
rect 12016 3626 12021 3678
rect 12073 3626 12085 3678
rect 12137 3626 12149 3678
rect 12201 3626 12206 3678
rect 12016 3613 12206 3626
rect 12016 3561 12021 3613
rect 12073 3561 12085 3613
rect 12137 3561 12149 3613
rect 12201 3561 12206 3613
rect 12016 3548 12206 3561
rect 12016 3496 12021 3548
rect 12073 3496 12085 3548
rect 12137 3496 12149 3548
rect 12201 3496 12206 3548
rect 12016 3483 12206 3496
rect 12016 3431 12021 3483
rect 12073 3431 12085 3483
rect 12137 3431 12149 3483
rect 12201 3431 12206 3483
rect 12016 3418 12206 3431
rect 12016 3366 12021 3418
rect 12073 3366 12085 3418
rect 12137 3366 12149 3418
rect 12201 3366 12206 3418
rect 12016 3353 12206 3366
rect 12016 3301 12021 3353
rect 12073 3301 12085 3353
rect 12137 3301 12149 3353
rect 12201 3301 12206 3353
rect 12016 3288 12206 3301
rect 12016 3236 12021 3288
rect 12073 3236 12085 3288
rect 12137 3236 12149 3288
rect 12201 3236 12206 3288
rect 12016 3223 12206 3236
rect 12016 3171 12021 3223
rect 12073 3171 12085 3223
rect 12137 3171 12149 3223
rect 12201 3171 12206 3223
rect 12016 3158 12206 3171
rect 12016 3106 12021 3158
rect 12073 3106 12085 3158
rect 12137 3106 12149 3158
rect 12201 3106 12206 3158
rect 12016 3093 12206 3106
rect 12016 3041 12021 3093
rect 12073 3041 12085 3093
rect 12137 3041 12149 3093
rect 12201 3041 12206 3093
rect 12016 3028 12206 3041
rect 12016 2976 12021 3028
rect 12073 2976 12085 3028
rect 12137 2976 12149 3028
rect 12201 2976 12206 3028
rect 12016 2963 12206 2976
rect 12016 2911 12021 2963
rect 12073 2911 12085 2963
rect 12137 2911 12149 2963
rect 12201 2911 12206 2963
rect 12016 2898 12206 2911
rect 12016 2846 12021 2898
rect 12073 2846 12085 2898
rect 12137 2846 12149 2898
rect 12201 2846 12206 2898
rect 12016 2833 12206 2846
rect 12016 2781 12021 2833
rect 12073 2781 12085 2833
rect 12137 2781 12149 2833
rect 12201 2781 12206 2833
rect 12016 2768 12206 2781
rect 12016 2716 12021 2768
rect 12073 2716 12085 2768
rect 12137 2716 12149 2768
rect 12201 2716 12206 2768
rect 12016 2703 12206 2716
rect 12016 2651 12021 2703
rect 12073 2651 12085 2703
rect 12137 2651 12149 2703
rect 12201 2651 12206 2703
rect 12016 2638 12206 2651
rect 12016 2586 12021 2638
rect 12073 2586 12085 2638
rect 12137 2586 12149 2638
rect 12201 2586 12206 2638
rect 12016 2573 12206 2586
rect 12016 2521 12021 2573
rect 12073 2521 12085 2573
rect 12137 2521 12149 2573
rect 12201 2521 12206 2573
rect 12016 2508 12206 2521
rect 12016 2456 12021 2508
rect 12073 2456 12085 2508
rect 12137 2456 12149 2508
rect 12201 2456 12206 2508
rect 12016 2443 12206 2456
rect 12016 2391 12021 2443
rect 12073 2391 12085 2443
rect 12137 2391 12149 2443
rect 12201 2391 12206 2443
rect 12016 2378 12206 2391
rect 12016 2326 12021 2378
rect 12073 2326 12085 2378
rect 12137 2326 12149 2378
rect 12201 2326 12206 2378
rect 12016 2313 12206 2326
rect 12016 2261 12021 2313
rect 12073 2261 12085 2313
rect 12137 2261 12149 2313
rect 12201 2261 12206 2313
rect 12016 2248 12206 2261
rect 12016 2196 12021 2248
rect 12073 2196 12085 2248
rect 12137 2196 12149 2248
rect 12201 2196 12206 2248
rect 12016 2183 12206 2196
rect 12016 2131 12021 2183
rect 12073 2131 12085 2183
rect 12137 2131 12149 2183
rect 12201 2131 12206 2183
rect 12016 2118 12206 2131
rect 12016 2066 12021 2118
rect 12073 2066 12085 2118
rect 12137 2066 12149 2118
rect 12201 2066 12206 2118
rect 12016 2053 12206 2066
rect 12016 2001 12021 2053
rect 12073 2001 12085 2053
rect 12137 2001 12149 2053
rect 12201 2001 12206 2053
rect 12016 1987 12206 2001
rect 12016 1935 12021 1987
rect 12073 1935 12085 1987
rect 12137 1935 12149 1987
rect 12201 1935 12206 1987
rect 12016 1921 12206 1935
rect 12016 1869 12021 1921
rect 12073 1869 12085 1921
rect 12137 1869 12149 1921
rect 12201 1869 12206 1921
rect 12016 1855 12206 1869
rect 12016 1803 12021 1855
rect 12073 1803 12085 1855
rect 12137 1803 12149 1855
rect 12201 1803 12206 1855
rect 12016 1789 12206 1803
rect 12016 1737 12021 1789
rect 12073 1737 12085 1789
rect 12137 1737 12149 1789
rect 12201 1737 12206 1789
rect 12016 1723 12206 1737
rect 12016 1671 12021 1723
rect 12073 1671 12085 1723
rect 12137 1671 12149 1723
rect 12201 1671 12206 1723
rect 12016 1657 12206 1671
rect 12016 1605 12021 1657
rect 12073 1605 12085 1657
rect 12137 1605 12149 1657
rect 12201 1605 12206 1657
rect 12016 1591 12206 1605
rect 12016 1539 12021 1591
rect 12073 1539 12085 1591
rect 12137 1539 12149 1591
rect 12201 1539 12206 1591
rect 12016 1525 12206 1539
rect 12016 1473 12021 1525
rect 12073 1473 12085 1525
rect 12137 1473 12149 1525
rect 12201 1473 12206 1525
rect 12016 1467 12206 1473
rect 12512 4068 12702 4074
rect 12512 4016 12517 4068
rect 12569 4016 12581 4068
rect 12633 4016 12645 4068
rect 12697 4016 12702 4068
rect 12512 4003 12702 4016
rect 12512 3951 12517 4003
rect 12569 3951 12581 4003
rect 12633 3951 12645 4003
rect 12697 3951 12702 4003
rect 12512 3938 12702 3951
rect 12512 3886 12517 3938
rect 12569 3886 12581 3938
rect 12633 3886 12645 3938
rect 12697 3886 12702 3938
rect 12512 3873 12702 3886
rect 12512 3821 12517 3873
rect 12569 3821 12581 3873
rect 12633 3821 12645 3873
rect 12697 3821 12702 3873
rect 12512 3808 12702 3821
rect 12512 3756 12517 3808
rect 12569 3756 12581 3808
rect 12633 3756 12645 3808
rect 12697 3756 12702 3808
rect 12512 3743 12702 3756
rect 12512 3691 12517 3743
rect 12569 3691 12581 3743
rect 12633 3691 12645 3743
rect 12697 3691 12702 3743
rect 12512 3678 12702 3691
rect 12512 3626 12517 3678
rect 12569 3626 12581 3678
rect 12633 3626 12645 3678
rect 12697 3626 12702 3678
rect 12512 3613 12702 3626
rect 12512 3561 12517 3613
rect 12569 3561 12581 3613
rect 12633 3561 12645 3613
rect 12697 3561 12702 3613
rect 12512 3548 12702 3561
rect 12512 3496 12517 3548
rect 12569 3496 12581 3548
rect 12633 3496 12645 3548
rect 12697 3496 12702 3548
rect 12512 3483 12702 3496
rect 12512 3431 12517 3483
rect 12569 3431 12581 3483
rect 12633 3431 12645 3483
rect 12697 3431 12702 3483
rect 12512 3418 12702 3431
rect 12512 3366 12517 3418
rect 12569 3366 12581 3418
rect 12633 3366 12645 3418
rect 12697 3366 12702 3418
rect 12512 3353 12702 3366
rect 12512 3301 12517 3353
rect 12569 3301 12581 3353
rect 12633 3301 12645 3353
rect 12697 3301 12702 3353
rect 12512 3288 12702 3301
rect 12512 3236 12517 3288
rect 12569 3236 12581 3288
rect 12633 3236 12645 3288
rect 12697 3236 12702 3288
rect 12512 3223 12702 3236
rect 12512 3171 12517 3223
rect 12569 3171 12581 3223
rect 12633 3171 12645 3223
rect 12697 3171 12702 3223
rect 12512 3158 12702 3171
rect 12512 3106 12517 3158
rect 12569 3106 12581 3158
rect 12633 3106 12645 3158
rect 12697 3106 12702 3158
rect 12512 3093 12702 3106
rect 12512 3041 12517 3093
rect 12569 3041 12581 3093
rect 12633 3041 12645 3093
rect 12697 3041 12702 3093
rect 12512 3028 12702 3041
rect 12512 2976 12517 3028
rect 12569 2976 12581 3028
rect 12633 2976 12645 3028
rect 12697 2976 12702 3028
rect 12512 2963 12702 2976
rect 12512 2911 12517 2963
rect 12569 2911 12581 2963
rect 12633 2911 12645 2963
rect 12697 2911 12702 2963
rect 12512 2898 12702 2911
rect 12512 2846 12517 2898
rect 12569 2846 12581 2898
rect 12633 2846 12645 2898
rect 12697 2846 12702 2898
rect 12512 2833 12702 2846
rect 12512 2781 12517 2833
rect 12569 2781 12581 2833
rect 12633 2781 12645 2833
rect 12697 2781 12702 2833
rect 12512 2768 12702 2781
rect 12512 2716 12517 2768
rect 12569 2716 12581 2768
rect 12633 2716 12645 2768
rect 12697 2716 12702 2768
rect 12512 2703 12702 2716
rect 12512 2651 12517 2703
rect 12569 2651 12581 2703
rect 12633 2651 12645 2703
rect 12697 2651 12702 2703
rect 12512 2638 12702 2651
rect 12512 2586 12517 2638
rect 12569 2586 12581 2638
rect 12633 2586 12645 2638
rect 12697 2586 12702 2638
rect 12512 2573 12702 2586
rect 12512 2521 12517 2573
rect 12569 2521 12581 2573
rect 12633 2521 12645 2573
rect 12697 2521 12702 2573
rect 12512 2508 12702 2521
rect 12512 2456 12517 2508
rect 12569 2456 12581 2508
rect 12633 2456 12645 2508
rect 12697 2456 12702 2508
rect 12512 2443 12702 2456
rect 12512 2391 12517 2443
rect 12569 2391 12581 2443
rect 12633 2391 12645 2443
rect 12697 2391 12702 2443
rect 12512 2378 12702 2391
rect 12512 2326 12517 2378
rect 12569 2326 12581 2378
rect 12633 2326 12645 2378
rect 12697 2326 12702 2378
rect 12512 2313 12702 2326
rect 12512 2261 12517 2313
rect 12569 2261 12581 2313
rect 12633 2261 12645 2313
rect 12697 2261 12702 2313
rect 12512 2248 12702 2261
rect 12512 2196 12517 2248
rect 12569 2196 12581 2248
rect 12633 2196 12645 2248
rect 12697 2196 12702 2248
rect 12512 2183 12702 2196
rect 12512 2131 12517 2183
rect 12569 2131 12581 2183
rect 12633 2131 12645 2183
rect 12697 2131 12702 2183
rect 12512 2118 12702 2131
rect 12512 2066 12517 2118
rect 12569 2066 12581 2118
rect 12633 2066 12645 2118
rect 12697 2066 12702 2118
rect 12512 2053 12702 2066
rect 12512 2001 12517 2053
rect 12569 2001 12581 2053
rect 12633 2001 12645 2053
rect 12697 2001 12702 2053
rect 12512 1987 12702 2001
rect 12512 1935 12517 1987
rect 12569 1935 12581 1987
rect 12633 1935 12645 1987
rect 12697 1935 12702 1987
rect 12512 1921 12702 1935
rect 12512 1869 12517 1921
rect 12569 1869 12581 1921
rect 12633 1869 12645 1921
rect 12697 1869 12702 1921
rect 12512 1855 12702 1869
rect 12512 1803 12517 1855
rect 12569 1803 12581 1855
rect 12633 1803 12645 1855
rect 12697 1803 12702 1855
rect 12512 1789 12702 1803
rect 12512 1737 12517 1789
rect 12569 1737 12581 1789
rect 12633 1737 12645 1789
rect 12697 1737 12702 1789
rect 12512 1723 12702 1737
rect 12512 1671 12517 1723
rect 12569 1671 12581 1723
rect 12633 1671 12645 1723
rect 12697 1671 12702 1723
rect 12512 1657 12702 1671
rect 12512 1605 12517 1657
rect 12569 1605 12581 1657
rect 12633 1605 12645 1657
rect 12697 1605 12702 1657
rect 12512 1591 12702 1605
rect 12512 1539 12517 1591
rect 12569 1539 12581 1591
rect 12633 1539 12645 1591
rect 12697 1539 12702 1591
rect 12512 1525 12702 1539
rect 12512 1473 12517 1525
rect 12569 1473 12581 1525
rect 12633 1473 12645 1525
rect 12697 1473 12702 1525
rect 12512 1467 12702 1473
rect 13008 4068 13198 4074
rect 13008 4016 13013 4068
rect 13065 4016 13077 4068
rect 13129 4016 13141 4068
rect 13193 4016 13198 4068
rect 13008 4003 13198 4016
rect 13008 3951 13013 4003
rect 13065 3951 13077 4003
rect 13129 3951 13141 4003
rect 13193 3951 13198 4003
rect 13008 3938 13198 3951
rect 13008 3886 13013 3938
rect 13065 3886 13077 3938
rect 13129 3886 13141 3938
rect 13193 3886 13198 3938
rect 13008 3873 13198 3886
rect 13008 3821 13013 3873
rect 13065 3821 13077 3873
rect 13129 3821 13141 3873
rect 13193 3821 13198 3873
rect 13008 3808 13198 3821
rect 13008 3756 13013 3808
rect 13065 3756 13077 3808
rect 13129 3756 13141 3808
rect 13193 3756 13198 3808
rect 13008 3743 13198 3756
rect 13008 3691 13013 3743
rect 13065 3691 13077 3743
rect 13129 3691 13141 3743
rect 13193 3691 13198 3743
rect 13008 3678 13198 3691
rect 13008 3626 13013 3678
rect 13065 3626 13077 3678
rect 13129 3626 13141 3678
rect 13193 3626 13198 3678
rect 13008 3613 13198 3626
rect 13008 3561 13013 3613
rect 13065 3561 13077 3613
rect 13129 3561 13141 3613
rect 13193 3561 13198 3613
rect 13008 3548 13198 3561
rect 13008 3496 13013 3548
rect 13065 3496 13077 3548
rect 13129 3496 13141 3548
rect 13193 3496 13198 3548
rect 13008 3483 13198 3496
rect 13008 3431 13013 3483
rect 13065 3431 13077 3483
rect 13129 3431 13141 3483
rect 13193 3431 13198 3483
rect 13008 3418 13198 3431
rect 13008 3366 13013 3418
rect 13065 3366 13077 3418
rect 13129 3366 13141 3418
rect 13193 3366 13198 3418
rect 13008 3353 13198 3366
rect 13008 3301 13013 3353
rect 13065 3301 13077 3353
rect 13129 3301 13141 3353
rect 13193 3301 13198 3353
rect 13008 3288 13198 3301
rect 13008 3236 13013 3288
rect 13065 3236 13077 3288
rect 13129 3236 13141 3288
rect 13193 3236 13198 3288
rect 13008 3223 13198 3236
rect 13008 3171 13013 3223
rect 13065 3171 13077 3223
rect 13129 3171 13141 3223
rect 13193 3171 13198 3223
rect 13008 3158 13198 3171
rect 13008 3106 13013 3158
rect 13065 3106 13077 3158
rect 13129 3106 13141 3158
rect 13193 3106 13198 3158
rect 13008 3093 13198 3106
rect 13008 3041 13013 3093
rect 13065 3041 13077 3093
rect 13129 3041 13141 3093
rect 13193 3041 13198 3093
rect 13008 3028 13198 3041
rect 13008 2976 13013 3028
rect 13065 2976 13077 3028
rect 13129 2976 13141 3028
rect 13193 2976 13198 3028
rect 13008 2963 13198 2976
rect 13008 2911 13013 2963
rect 13065 2911 13077 2963
rect 13129 2911 13141 2963
rect 13193 2911 13198 2963
rect 13008 2898 13198 2911
rect 13008 2846 13013 2898
rect 13065 2846 13077 2898
rect 13129 2846 13141 2898
rect 13193 2846 13198 2898
rect 13008 2833 13198 2846
rect 13008 2781 13013 2833
rect 13065 2781 13077 2833
rect 13129 2781 13141 2833
rect 13193 2781 13198 2833
rect 13008 2768 13198 2781
rect 13008 2716 13013 2768
rect 13065 2716 13077 2768
rect 13129 2716 13141 2768
rect 13193 2716 13198 2768
rect 13008 2703 13198 2716
rect 13008 2651 13013 2703
rect 13065 2651 13077 2703
rect 13129 2651 13141 2703
rect 13193 2651 13198 2703
rect 13008 2638 13198 2651
rect 13008 2586 13013 2638
rect 13065 2586 13077 2638
rect 13129 2586 13141 2638
rect 13193 2586 13198 2638
rect 13008 2573 13198 2586
rect 13008 2521 13013 2573
rect 13065 2521 13077 2573
rect 13129 2521 13141 2573
rect 13193 2521 13198 2573
rect 13008 2508 13198 2521
rect 13008 2456 13013 2508
rect 13065 2456 13077 2508
rect 13129 2456 13141 2508
rect 13193 2456 13198 2508
rect 13008 2443 13198 2456
rect 13008 2391 13013 2443
rect 13065 2391 13077 2443
rect 13129 2391 13141 2443
rect 13193 2391 13198 2443
rect 13008 2378 13198 2391
rect 13008 2326 13013 2378
rect 13065 2326 13077 2378
rect 13129 2326 13141 2378
rect 13193 2326 13198 2378
rect 13008 2313 13198 2326
rect 13008 2261 13013 2313
rect 13065 2261 13077 2313
rect 13129 2261 13141 2313
rect 13193 2261 13198 2313
rect 13008 2248 13198 2261
rect 13008 2196 13013 2248
rect 13065 2196 13077 2248
rect 13129 2196 13141 2248
rect 13193 2196 13198 2248
rect 13008 2183 13198 2196
rect 13008 2131 13013 2183
rect 13065 2131 13077 2183
rect 13129 2131 13141 2183
rect 13193 2131 13198 2183
rect 13008 2118 13198 2131
rect 13008 2066 13013 2118
rect 13065 2066 13077 2118
rect 13129 2066 13141 2118
rect 13193 2066 13198 2118
rect 13008 2053 13198 2066
rect 13008 2001 13013 2053
rect 13065 2001 13077 2053
rect 13129 2001 13141 2053
rect 13193 2001 13198 2053
rect 13008 1987 13198 2001
rect 13008 1935 13013 1987
rect 13065 1935 13077 1987
rect 13129 1935 13141 1987
rect 13193 1935 13198 1987
rect 13008 1921 13198 1935
rect 13008 1869 13013 1921
rect 13065 1869 13077 1921
rect 13129 1869 13141 1921
rect 13193 1869 13198 1921
rect 13008 1855 13198 1869
rect 13008 1803 13013 1855
rect 13065 1803 13077 1855
rect 13129 1803 13141 1855
rect 13193 1803 13198 1855
rect 13008 1789 13198 1803
rect 13008 1737 13013 1789
rect 13065 1737 13077 1789
rect 13129 1737 13141 1789
rect 13193 1737 13198 1789
rect 13008 1723 13198 1737
rect 13008 1671 13013 1723
rect 13065 1671 13077 1723
rect 13129 1671 13141 1723
rect 13193 1671 13198 1723
rect 13008 1657 13198 1671
rect 13008 1605 13013 1657
rect 13065 1605 13077 1657
rect 13129 1605 13141 1657
rect 13193 1605 13198 1657
rect 13008 1591 13198 1605
rect 13008 1539 13013 1591
rect 13065 1539 13077 1591
rect 13129 1539 13141 1591
rect 13193 1539 13198 1591
rect 13008 1525 13198 1539
rect 13008 1473 13013 1525
rect 13065 1473 13077 1525
rect 13129 1473 13141 1525
rect 13193 1473 13198 1525
rect 13008 1467 13198 1473
rect 13504 4068 13694 4074
rect 13504 4016 13509 4068
rect 13561 4016 13573 4068
rect 13625 4016 13637 4068
rect 13689 4016 13694 4068
rect 13504 4003 13694 4016
rect 13504 3951 13509 4003
rect 13561 3951 13573 4003
rect 13625 3951 13637 4003
rect 13689 3951 13694 4003
rect 13504 3938 13694 3951
rect 13504 3886 13509 3938
rect 13561 3886 13573 3938
rect 13625 3886 13637 3938
rect 13689 3886 13694 3938
rect 13504 3873 13694 3886
rect 13504 3821 13509 3873
rect 13561 3821 13573 3873
rect 13625 3821 13637 3873
rect 13689 3821 13694 3873
rect 13504 3808 13694 3821
rect 13504 3756 13509 3808
rect 13561 3756 13573 3808
rect 13625 3756 13637 3808
rect 13689 3756 13694 3808
rect 13504 3743 13694 3756
rect 13504 3691 13509 3743
rect 13561 3691 13573 3743
rect 13625 3691 13637 3743
rect 13689 3691 13694 3743
rect 13504 3678 13694 3691
rect 13504 3626 13509 3678
rect 13561 3626 13573 3678
rect 13625 3626 13637 3678
rect 13689 3626 13694 3678
rect 13504 3613 13694 3626
rect 13504 3561 13509 3613
rect 13561 3561 13573 3613
rect 13625 3561 13637 3613
rect 13689 3561 13694 3613
rect 13504 3548 13694 3561
rect 13504 3496 13509 3548
rect 13561 3496 13573 3548
rect 13625 3496 13637 3548
rect 13689 3496 13694 3548
rect 13504 3483 13694 3496
rect 13504 3431 13509 3483
rect 13561 3431 13573 3483
rect 13625 3431 13637 3483
rect 13689 3431 13694 3483
rect 13504 3418 13694 3431
rect 13504 3366 13509 3418
rect 13561 3366 13573 3418
rect 13625 3366 13637 3418
rect 13689 3366 13694 3418
rect 13504 3353 13694 3366
rect 13504 3301 13509 3353
rect 13561 3301 13573 3353
rect 13625 3301 13637 3353
rect 13689 3301 13694 3353
rect 13504 3288 13694 3301
rect 13504 3236 13509 3288
rect 13561 3236 13573 3288
rect 13625 3236 13637 3288
rect 13689 3236 13694 3288
rect 13504 3223 13694 3236
rect 13504 3171 13509 3223
rect 13561 3171 13573 3223
rect 13625 3171 13637 3223
rect 13689 3171 13694 3223
rect 13504 3158 13694 3171
rect 13504 3106 13509 3158
rect 13561 3106 13573 3158
rect 13625 3106 13637 3158
rect 13689 3106 13694 3158
rect 13504 3093 13694 3106
rect 13504 3041 13509 3093
rect 13561 3041 13573 3093
rect 13625 3041 13637 3093
rect 13689 3041 13694 3093
rect 13504 3028 13694 3041
rect 13504 2976 13509 3028
rect 13561 2976 13573 3028
rect 13625 2976 13637 3028
rect 13689 2976 13694 3028
rect 13504 2963 13694 2976
rect 13504 2911 13509 2963
rect 13561 2911 13573 2963
rect 13625 2911 13637 2963
rect 13689 2911 13694 2963
rect 13504 2898 13694 2911
rect 13504 2846 13509 2898
rect 13561 2846 13573 2898
rect 13625 2846 13637 2898
rect 13689 2846 13694 2898
rect 13504 2833 13694 2846
rect 13504 2781 13509 2833
rect 13561 2781 13573 2833
rect 13625 2781 13637 2833
rect 13689 2781 13694 2833
rect 13504 2768 13694 2781
rect 13504 2716 13509 2768
rect 13561 2716 13573 2768
rect 13625 2716 13637 2768
rect 13689 2716 13694 2768
rect 13504 2703 13694 2716
rect 13504 2651 13509 2703
rect 13561 2651 13573 2703
rect 13625 2651 13637 2703
rect 13689 2651 13694 2703
rect 13504 2638 13694 2651
rect 13504 2586 13509 2638
rect 13561 2586 13573 2638
rect 13625 2586 13637 2638
rect 13689 2586 13694 2638
rect 13504 2573 13694 2586
rect 13504 2521 13509 2573
rect 13561 2521 13573 2573
rect 13625 2521 13637 2573
rect 13689 2521 13694 2573
rect 13504 2508 13694 2521
rect 13504 2456 13509 2508
rect 13561 2456 13573 2508
rect 13625 2456 13637 2508
rect 13689 2456 13694 2508
rect 13504 2443 13694 2456
rect 13504 2391 13509 2443
rect 13561 2391 13573 2443
rect 13625 2391 13637 2443
rect 13689 2391 13694 2443
rect 13504 2378 13694 2391
rect 13504 2326 13509 2378
rect 13561 2326 13573 2378
rect 13625 2326 13637 2378
rect 13689 2326 13694 2378
rect 13504 2313 13694 2326
rect 13504 2261 13509 2313
rect 13561 2261 13573 2313
rect 13625 2261 13637 2313
rect 13689 2261 13694 2313
rect 13504 2248 13694 2261
rect 13504 2196 13509 2248
rect 13561 2196 13573 2248
rect 13625 2196 13637 2248
rect 13689 2196 13694 2248
rect 13504 2183 13694 2196
rect 13504 2131 13509 2183
rect 13561 2131 13573 2183
rect 13625 2131 13637 2183
rect 13689 2131 13694 2183
rect 13504 2118 13694 2131
rect 13504 2066 13509 2118
rect 13561 2066 13573 2118
rect 13625 2066 13637 2118
rect 13689 2066 13694 2118
rect 13504 2053 13694 2066
rect 13504 2001 13509 2053
rect 13561 2001 13573 2053
rect 13625 2001 13637 2053
rect 13689 2001 13694 2053
rect 13504 1987 13694 2001
rect 13504 1935 13509 1987
rect 13561 1935 13573 1987
rect 13625 1935 13637 1987
rect 13689 1935 13694 1987
rect 13504 1921 13694 1935
rect 13504 1869 13509 1921
rect 13561 1869 13573 1921
rect 13625 1869 13637 1921
rect 13689 1869 13694 1921
rect 13504 1855 13694 1869
rect 13504 1803 13509 1855
rect 13561 1803 13573 1855
rect 13625 1803 13637 1855
rect 13689 1803 13694 1855
rect 13504 1789 13694 1803
rect 13504 1737 13509 1789
rect 13561 1737 13573 1789
rect 13625 1737 13637 1789
rect 13689 1737 13694 1789
rect 13504 1723 13694 1737
rect 13504 1671 13509 1723
rect 13561 1671 13573 1723
rect 13625 1671 13637 1723
rect 13689 1671 13694 1723
rect 13504 1657 13694 1671
rect 13504 1605 13509 1657
rect 13561 1605 13573 1657
rect 13625 1605 13637 1657
rect 13689 1605 13694 1657
rect 13504 1591 13694 1605
rect 13504 1539 13509 1591
rect 13561 1539 13573 1591
rect 13625 1539 13637 1591
rect 13689 1539 13694 1591
rect 13504 1525 13694 1539
rect 13504 1473 13509 1525
rect 13561 1473 13573 1525
rect 13625 1473 13637 1525
rect 13689 1473 13694 1525
rect 13504 1467 13694 1473
rect 14036 4068 14226 4074
rect 14036 4016 14037 4068
rect 14089 4016 14105 4068
rect 14157 4016 14173 4068
rect 14225 4016 14226 4068
rect 14036 4003 14226 4016
rect 14036 3951 14037 4003
rect 14089 3951 14105 4003
rect 14157 3951 14173 4003
rect 14225 3951 14226 4003
rect 14036 3938 14226 3951
rect 14036 3886 14037 3938
rect 14089 3886 14105 3938
rect 14157 3886 14173 3938
rect 14225 3886 14226 3938
rect 14036 3873 14226 3886
rect 14036 3821 14037 3873
rect 14089 3821 14105 3873
rect 14157 3821 14173 3873
rect 14225 3821 14226 3873
rect 14036 3808 14226 3821
rect 14036 3756 14037 3808
rect 14089 3756 14105 3808
rect 14157 3756 14173 3808
rect 14225 3756 14226 3808
rect 14036 3743 14226 3756
rect 14036 3691 14037 3743
rect 14089 3691 14105 3743
rect 14157 3691 14173 3743
rect 14225 3691 14226 3743
rect 14036 3678 14226 3691
rect 14036 3626 14037 3678
rect 14089 3626 14105 3678
rect 14157 3626 14173 3678
rect 14225 3626 14226 3678
rect 14036 3613 14226 3626
rect 14036 3561 14037 3613
rect 14089 3561 14105 3613
rect 14157 3561 14173 3613
rect 14225 3561 14226 3613
rect 14036 3548 14226 3561
rect 14036 3496 14037 3548
rect 14089 3496 14105 3548
rect 14157 3496 14173 3548
rect 14225 3496 14226 3548
rect 14036 3483 14226 3496
rect 14036 3431 14037 3483
rect 14089 3431 14105 3483
rect 14157 3431 14173 3483
rect 14225 3431 14226 3483
rect 14036 3418 14226 3431
rect 14036 3366 14037 3418
rect 14089 3366 14105 3418
rect 14157 3366 14173 3418
rect 14225 3366 14226 3418
rect 14036 3353 14226 3366
rect 14036 3301 14037 3353
rect 14089 3301 14105 3353
rect 14157 3301 14173 3353
rect 14225 3301 14226 3353
rect 14036 3288 14226 3301
rect 14036 3236 14037 3288
rect 14089 3236 14105 3288
rect 14157 3236 14173 3288
rect 14225 3236 14226 3288
rect 14036 3223 14226 3236
rect 14036 3171 14037 3223
rect 14089 3171 14105 3223
rect 14157 3171 14173 3223
rect 14225 3171 14226 3223
rect 14036 3158 14226 3171
rect 14036 3106 14037 3158
rect 14089 3106 14105 3158
rect 14157 3106 14173 3158
rect 14225 3106 14226 3158
rect 14036 3093 14226 3106
rect 14036 3041 14037 3093
rect 14089 3041 14105 3093
rect 14157 3041 14173 3093
rect 14225 3041 14226 3093
rect 14036 3028 14226 3041
rect 14036 2976 14037 3028
rect 14089 2976 14105 3028
rect 14157 2976 14173 3028
rect 14225 2976 14226 3028
rect 14036 2963 14226 2976
rect 14036 2911 14037 2963
rect 14089 2911 14105 2963
rect 14157 2911 14173 2963
rect 14225 2911 14226 2963
rect 14036 2898 14226 2911
rect 14036 2846 14037 2898
rect 14089 2846 14105 2898
rect 14157 2846 14173 2898
rect 14225 2846 14226 2898
rect 14036 2833 14226 2846
rect 14036 2781 14037 2833
rect 14089 2781 14105 2833
rect 14157 2781 14173 2833
rect 14225 2781 14226 2833
rect 14036 2768 14226 2781
rect 14036 2716 14037 2768
rect 14089 2716 14105 2768
rect 14157 2716 14173 2768
rect 14225 2716 14226 2768
rect 14036 2703 14226 2716
rect 14036 2651 14037 2703
rect 14089 2651 14105 2703
rect 14157 2651 14173 2703
rect 14225 2651 14226 2703
rect 14036 2638 14226 2651
rect 14036 2586 14037 2638
rect 14089 2586 14105 2638
rect 14157 2586 14173 2638
rect 14225 2586 14226 2638
rect 14036 2573 14226 2586
rect 14036 2521 14037 2573
rect 14089 2521 14105 2573
rect 14157 2521 14173 2573
rect 14225 2521 14226 2573
rect 14036 2508 14226 2521
rect 14036 2456 14037 2508
rect 14089 2456 14105 2508
rect 14157 2456 14173 2508
rect 14225 2456 14226 2508
rect 14036 2443 14226 2456
rect 14036 2391 14037 2443
rect 14089 2391 14105 2443
rect 14157 2391 14173 2443
rect 14225 2391 14226 2443
rect 14036 2378 14226 2391
rect 14036 2326 14037 2378
rect 14089 2326 14105 2378
rect 14157 2326 14173 2378
rect 14225 2326 14226 2378
rect 14036 2313 14226 2326
rect 14036 2261 14037 2313
rect 14089 2261 14105 2313
rect 14157 2261 14173 2313
rect 14225 2261 14226 2313
rect 14036 2248 14226 2261
rect 14036 2196 14037 2248
rect 14089 2196 14105 2248
rect 14157 2196 14173 2248
rect 14225 2196 14226 2248
rect 14036 2183 14226 2196
rect 14036 2131 14037 2183
rect 14089 2131 14105 2183
rect 14157 2131 14173 2183
rect 14225 2131 14226 2183
rect 14036 2118 14226 2131
rect 14036 2066 14037 2118
rect 14089 2066 14105 2118
rect 14157 2066 14173 2118
rect 14225 2066 14226 2118
rect 14036 2053 14226 2066
rect 14036 2001 14037 2053
rect 14089 2001 14105 2053
rect 14157 2001 14173 2053
rect 14225 2001 14226 2053
rect 14036 1987 14226 2001
rect 14036 1935 14037 1987
rect 14089 1935 14105 1987
rect 14157 1935 14173 1987
rect 14225 1935 14226 1987
rect 14036 1921 14226 1935
rect 14036 1869 14037 1921
rect 14089 1869 14105 1921
rect 14157 1869 14173 1921
rect 14225 1869 14226 1921
rect 14036 1855 14226 1869
rect 14036 1803 14037 1855
rect 14089 1803 14105 1855
rect 14157 1803 14173 1855
rect 14225 1803 14226 1855
rect 14036 1789 14226 1803
rect 14036 1737 14037 1789
rect 14089 1737 14105 1789
rect 14157 1737 14173 1789
rect 14225 1737 14226 1789
rect 14036 1723 14226 1737
rect 14036 1671 14037 1723
rect 14089 1671 14105 1723
rect 14157 1671 14173 1723
rect 14225 1671 14226 1723
rect 14036 1657 14226 1671
rect 14036 1605 14037 1657
rect 14089 1605 14105 1657
rect 14157 1605 14173 1657
rect 14225 1605 14226 1657
rect 14036 1591 14226 1605
rect 14036 1539 14037 1591
rect 14089 1539 14105 1591
rect 14157 1539 14173 1591
rect 14225 1539 14226 1591
rect 14036 1525 14226 1539
rect 14036 1473 14037 1525
rect 14089 1473 14105 1525
rect 14157 1473 14173 1525
rect 14225 1473 14226 1525
rect 14036 1467 14226 1473
rect 14400 4068 14628 4074
rect 14452 4016 14488 4068
rect 14540 4016 14576 4068
rect 14400 4003 14628 4016
rect 14452 3951 14488 4003
rect 14540 3951 14576 4003
rect 14400 3938 14628 3951
rect 14452 3886 14488 3938
rect 14540 3886 14576 3938
rect 14400 3873 14628 3886
rect 14452 3821 14488 3873
rect 14540 3821 14576 3873
rect 14400 3808 14628 3821
rect 14452 3756 14488 3808
rect 14540 3756 14576 3808
rect 14400 3743 14628 3756
rect 14452 3691 14488 3743
rect 14540 3691 14576 3743
rect 14400 3678 14628 3691
rect 14452 3626 14488 3678
rect 14540 3626 14576 3678
rect 14400 3613 14628 3626
rect 14452 3561 14488 3613
rect 14540 3561 14576 3613
rect 14400 3548 14628 3561
rect 14452 3496 14488 3548
rect 14540 3496 14576 3548
rect 14400 3483 14628 3496
rect 14452 3431 14488 3483
rect 14540 3431 14576 3483
rect 14400 3418 14628 3431
rect 14452 3366 14488 3418
rect 14540 3366 14576 3418
rect 14400 3353 14628 3366
rect 14452 3301 14488 3353
rect 14540 3301 14576 3353
rect 14400 3288 14628 3301
rect 14452 3236 14488 3288
rect 14540 3236 14576 3288
rect 14400 3223 14628 3236
rect 14452 3171 14488 3223
rect 14540 3171 14576 3223
rect 14400 3158 14628 3171
rect 14452 3106 14488 3158
rect 14540 3106 14576 3158
rect 14400 3093 14628 3106
rect 14452 3041 14488 3093
rect 14540 3041 14576 3093
rect 14400 3028 14628 3041
rect 14452 2976 14488 3028
rect 14540 2976 14576 3028
rect 14400 2963 14628 2976
rect 14452 2911 14488 2963
rect 14540 2911 14576 2963
rect 14400 2898 14628 2911
rect 14452 2846 14488 2898
rect 14540 2846 14576 2898
rect 14400 2833 14628 2846
rect 14452 2781 14488 2833
rect 14540 2781 14576 2833
rect 14400 2768 14628 2781
rect 14452 2716 14488 2768
rect 14540 2716 14576 2768
rect 14400 2703 14628 2716
rect 14452 2651 14488 2703
rect 14540 2651 14576 2703
rect 14400 2638 14628 2651
rect 14452 2586 14488 2638
rect 14540 2586 14576 2638
rect 14400 2573 14628 2586
rect 14452 2521 14488 2573
rect 14540 2521 14576 2573
rect 14400 2508 14628 2521
rect 14452 2456 14488 2508
rect 14540 2456 14576 2508
rect 14400 2443 14628 2456
rect 14452 2391 14488 2443
rect 14540 2391 14576 2443
rect 14400 2378 14628 2391
rect 14452 2326 14488 2378
rect 14540 2326 14576 2378
rect 14400 2313 14628 2326
rect 14452 2261 14488 2313
rect 14540 2261 14576 2313
rect 14400 2248 14628 2261
rect 14452 2196 14488 2248
rect 14540 2196 14576 2248
rect 14400 2183 14628 2196
rect 14452 2131 14488 2183
rect 14540 2131 14576 2183
rect 14400 2118 14628 2131
rect 14452 2066 14488 2118
rect 14540 2066 14576 2118
rect 14400 2053 14628 2066
rect 14452 2001 14488 2053
rect 14540 2001 14576 2053
rect 14400 1987 14628 2001
rect 14452 1935 14488 1987
rect 14540 1935 14576 1987
rect 14400 1921 14628 1935
rect 14452 1869 14488 1921
rect 14540 1869 14576 1921
rect 14400 1855 14628 1869
rect 14452 1803 14488 1855
rect 14540 1803 14576 1855
rect 14400 1789 14628 1803
rect 14452 1737 14488 1789
rect 14540 1737 14576 1789
rect 14400 1723 14628 1737
rect 14452 1671 14488 1723
rect 14540 1671 14576 1723
rect 14400 1657 14628 1671
rect 14452 1605 14488 1657
rect 14540 1605 14576 1657
rect 14400 1591 14628 1605
rect 14452 1539 14488 1591
rect 14540 1539 14576 1591
rect 14400 1525 14628 1539
rect 14452 1473 14488 1525
rect 14540 1473 14576 1525
rect 14400 1467 14628 1473
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_0
timestamp 1644511149
transform 1 0 14031 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_1
timestamp 1644511149
transform 1 0 14031 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_2
timestamp 1644511149
transform 1 0 8079 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_3
timestamp 1644511149
transform 1 0 9071 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_4
timestamp 1644511149
transform 1 0 10063 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_5
timestamp 1644511149
transform 1 0 11055 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_6
timestamp 1644511149
transform 1 0 12047 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_7
timestamp 1644511149
transform 1 0 13039 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_8
timestamp 1644511149
transform 1 0 8151 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_9
timestamp 1644511149
transform 1 0 9143 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_10
timestamp 1644511149
transform 1 0 10135 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_11
timestamp 1644511149
transform 1 0 11127 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_12
timestamp 1644511149
transform 1 0 12119 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_13
timestamp 1644511149
transform 1 0 13111 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_14
timestamp 1644511149
transform 1 0 13111 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_15
timestamp 1644511149
transform 1 0 12119 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_16
timestamp 1644511149
transform 1 0 11127 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_17
timestamp 1644511149
transform 1 0 10135 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_18
timestamp 1644511149
transform 1 0 9143 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_19
timestamp 1644511149
transform 1 0 8151 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_20
timestamp 1644511149
transform 1 0 13039 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_21
timestamp 1644511149
transform 1 0 12047 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_22
timestamp 1644511149
transform 1 0 11055 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_23
timestamp 1644511149
transform 1 0 10063 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_24
timestamp 1644511149
transform 1 0 9071 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_25
timestamp 1644511149
transform 1 0 8079 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_26
timestamp 1644511149
transform 1 0 1135 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_27
timestamp 1644511149
transform 1 0 1207 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_28
timestamp 1644511149
transform 1 0 2199 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_29
timestamp 1644511149
transform 1 0 2127 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_30
timestamp 1644511149
transform 1 0 1135 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_31
timestamp 1644511149
transform 1 0 1207 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_32
timestamp 1644511149
transform 1 0 2199 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_33
timestamp 1644511149
transform 1 0 2127 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_34
timestamp 1644511149
transform 1 0 3119 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_35
timestamp 1644511149
transform 1 0 4111 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_36
timestamp 1644511149
transform 1 0 5103 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_37
timestamp 1644511149
transform 1 0 6095 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_38
timestamp 1644511149
transform 1 0 7087 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_39
timestamp 1644511149
transform 1 0 3191 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_40
timestamp 1644511149
transform 1 0 4183 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_41
timestamp 1644511149
transform 1 0 5175 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_42
timestamp 1644511149
transform 1 0 6167 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_43
timestamp 1644511149
transform 1 0 7159 0 -1 2457
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_44
timestamp 1644511149
transform 1 0 7159 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_45
timestamp 1644511149
transform 1 0 6167 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_46
timestamp 1644511149
transform 1 0 5175 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_47
timestamp 1644511149
transform 1 0 4183 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_48
timestamp 1644511149
transform 1 0 3191 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_49
timestamp 1644511149
transform 1 0 7087 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_50
timestamp 1644511149
transform 1 0 6095 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_51
timestamp 1644511149
transform 1 0 5103 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_52
timestamp 1644511149
transform 1 0 4111 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808378  sky130_fd_pr__hvdfl1sd2__example_55959141808378_53
timestamp 1644511149
transform 1 0 3119 0 -1 4058
box 0 0 1 1
use sky130_fd_pr__nfet_01v8__example_55959141808645  sky130_fd_pr__nfet_01v8__example_55959141808645_0
timestamp 1644511149
transform 1 0 924 0 -1 2457
box -139 0 145 500
use sky130_fd_pr__nfet_01v8__example_55959141808647  sky130_fd_pr__nfet_01v8__example_55959141808647_0
timestamp 1644511149
transform 1 0 924 0 -1 4058
box -139 0 145 500
use sky130_fd_pr__nfet_01v8__example_55959141808647  sky130_fd_pr__nfet_01v8__example_55959141808647_1
timestamp 1644511149
transform -1 0 14298 0 -1 2457
box -139 0 145 500
use sky130_fd_pr__nfet_01v8__example_55959141808647  sky130_fd_pr__nfet_01v8__example_55959141808647_2
timestamp 1644511149
transform -1 0 14298 0 -1 4058
box -139 0 145 500
use sky130_fd_pr__nfet_01v8__example_55959141808648  sky130_fd_pr__nfet_01v8__example_55959141808648_0
timestamp 1644511149
transform 1 0 1916 0 -1 4058
box -25 0 12049 500
use sky130_fd_pr__nfet_01v8__example_55959141808650  sky130_fd_pr__nfet_01v8__example_55959141808650_0
timestamp 1644511149
transform -1 0 1474 0 -1 2457
box -221 0 145 500
use sky130_fd_pr__nfet_01v8__example_55959141808650  sky130_fd_pr__nfet_01v8__example_55959141808650_1
timestamp 1644511149
transform -1 0 1474 0 -1 4058
box -221 0 145 500
use sky130_fd_pr__nfet_01v8__example_55959141808651  sky130_fd_pr__nfet_01v8__example_55959141808651_0
timestamp 1644511149
transform 1 0 1916 0 -1 2457
box -25 0 12049 500
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_0
timestamp 1644511149
transform 1 0 14238 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_1
timestamp 1644511149
transform 1 0 12888 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_2
timestamp 1644511149
transform 1 0 13880 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_3
timestamp 1644511149
transform 1 0 13318 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_4
timestamp 1644511149
transform 1 0 12326 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_5
timestamp 1644511149
transform 1 0 11334 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_6
timestamp 1644511149
transform 1 0 10342 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_7
timestamp 1644511149
transform 1 0 9350 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_8
timestamp 1644511149
transform 1 0 8358 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_9
timestamp 1644511149
transform 1 0 7366 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_10
timestamp 1644511149
transform 1 0 6374 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_11
timestamp 1644511149
transform 1 0 5382 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_12
timestamp 1644511149
transform 1 0 8920 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_13
timestamp 1644511149
transform 1 0 7928 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_14
timestamp 1644511149
transform 1 0 6921 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_15
timestamp 1644511149
transform 1 0 5944 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_16
timestamp 1644511149
transform 1 0 4952 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_17
timestamp 1644511149
transform 1 0 3960 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_18
timestamp 1644511149
transform 1 0 2968 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_19
timestamp 1644511149
transform 1 0 1976 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_20
timestamp 1644511149
transform 1 0 984 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_21
timestamp 1644511149
transform 1 0 3398 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_22
timestamp 1644511149
transform 1 0 2406 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_23
timestamp 1644511149
transform 1 0 1414 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_24
timestamp 1644511149
transform 1 0 11896 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_25
timestamp 1644511149
transform 1 0 10904 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_26
timestamp 1644511149
transform 1 0 9912 0 1 4441
box 0 0 1 1
use sky130_fd_pr__via_l1m1_centered__example_559591418084  sky130_fd_pr__via_l1m1_centered__example_559591418084_27
timestamp 1644511149
transform 1 0 4390 0 1 4441
box 0 0 1 1
<< labels >>
flabel metal1 s 13239 5295 13646 5426 0 FreeSans 2000 0 0 0 VCC_IO
port 1 nsew
<< properties >>
string GDS_END 29749066
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 28946698
<< end >>
