magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< pwell >>
rect 467 350 491 401
<< locali >>
rect 0 902 876 918
rect 0 868 97 902
rect 131 868 169 902
rect 203 868 241 902
rect 275 868 313 902
rect 347 868 385 902
rect 419 868 457 902
rect 491 868 529 902
rect 563 868 601 902
rect 635 868 673 902
rect 707 868 745 902
rect 779 868 876 902
rect 0 836 876 868
rect 0 802 16 836
rect 50 802 826 836
rect 860 802 876 836
rect 0 764 876 802
rect 0 730 16 764
rect 50 730 826 764
rect 860 730 876 764
rect 0 692 876 730
rect 0 658 16 692
rect 50 658 826 692
rect 860 658 876 692
rect 0 620 876 658
rect 0 586 16 620
rect 50 586 826 620
rect 860 586 876 620
rect 0 548 876 586
rect 0 514 16 548
rect 50 514 826 548
rect 860 514 876 548
rect 0 476 876 514
rect 0 442 16 476
rect 50 442 826 476
rect 860 442 876 476
rect 0 404 876 442
rect 0 370 16 404
rect 50 370 826 404
rect 860 370 876 404
rect 0 332 876 370
rect 0 298 16 332
rect 50 298 826 332
rect 860 298 876 332
rect 0 260 876 298
rect 0 226 16 260
rect 50 226 826 260
rect 860 226 876 260
rect 0 188 876 226
rect 0 154 16 188
rect 50 154 826 188
rect 860 154 876 188
rect 0 116 876 154
rect 0 82 16 116
rect 50 82 826 116
rect 860 82 876 116
rect 0 50 876 82
rect 0 16 97 50
rect 131 16 169 50
rect 203 16 241 50
rect 275 16 313 50
rect 347 16 385 50
rect 419 16 457 50
rect 491 16 529 50
rect 563 16 601 50
rect 635 16 673 50
rect 707 16 745 50
rect 779 16 876 50
rect 0 0 876 16
<< viali >>
rect 97 868 131 902
rect 169 868 203 902
rect 241 868 275 902
rect 313 868 347 902
rect 385 868 419 902
rect 457 868 491 902
rect 529 868 563 902
rect 601 868 635 902
rect 673 868 707 902
rect 745 868 779 902
rect 16 802 50 836
rect 826 802 860 836
rect 16 730 50 764
rect 826 730 860 764
rect 16 658 50 692
rect 826 658 860 692
rect 16 586 50 620
rect 826 586 860 620
rect 16 514 50 548
rect 826 514 860 548
rect 16 442 50 476
rect 826 442 860 476
rect 16 370 50 404
rect 826 370 860 404
rect 16 298 50 332
rect 826 298 860 332
rect 16 226 50 260
rect 826 226 860 260
rect 16 154 50 188
rect 826 154 860 188
rect 16 82 50 116
rect 826 82 860 116
rect 97 16 131 50
rect 169 16 203 50
rect 241 16 275 50
rect 313 16 347 50
rect 385 16 419 50
rect 457 16 491 50
rect 529 16 563 50
rect 601 16 635 50
rect 673 16 707 50
rect 745 16 779 50
<< metal1 >>
rect 0 911 876 918
rect 0 859 52 911
rect 104 902 116 911
rect 168 902 180 911
rect 232 902 244 911
rect 168 868 169 902
rect 232 868 241 902
rect 104 859 116 868
rect 168 859 180 868
rect 232 859 244 868
rect 296 859 308 911
rect 360 902 516 911
rect 360 868 385 902
rect 419 868 457 902
rect 491 868 516 902
rect 360 859 516 868
rect 568 859 580 911
rect 632 902 644 911
rect 696 902 708 911
rect 760 902 772 911
rect 635 868 644 902
rect 707 868 708 902
rect 632 859 644 868
rect 696 859 708 868
rect 760 859 772 868
rect 824 859 876 911
rect 0 852 876 859
rect 0 842 66 852
rect 0 790 7 842
rect 59 790 66 842
rect 0 778 66 790
rect 0 726 7 778
rect 59 726 66 778
rect 0 714 66 726
rect 0 662 7 714
rect 59 662 66 714
rect 0 658 16 662
rect 50 658 66 662
rect 0 650 66 658
rect 0 598 7 650
rect 59 598 66 650
rect 0 586 16 598
rect 50 586 66 598
rect 0 534 7 586
rect 59 534 66 586
rect 0 514 16 534
rect 50 514 66 534
rect 0 476 66 514
rect 0 442 16 476
rect 50 442 66 476
rect 0 404 66 442
rect 0 384 16 404
rect 50 384 66 404
rect 0 332 7 384
rect 59 332 66 384
rect 0 320 16 332
rect 50 320 66 332
rect 0 268 7 320
rect 59 268 66 320
rect 0 260 66 268
rect 0 256 16 260
rect 50 256 66 260
rect 0 204 7 256
rect 59 204 66 256
rect 0 192 66 204
rect 0 140 7 192
rect 59 140 66 192
rect 0 128 66 140
rect 0 76 7 128
rect 59 76 66 128
rect 113 491 141 824
rect 169 519 197 852
rect 225 491 253 824
rect 281 519 309 852
rect 337 491 365 824
rect 411 818 465 824
rect 411 766 412 818
rect 464 766 465 818
rect 411 754 465 766
rect 411 702 412 754
rect 464 702 465 754
rect 411 690 465 702
rect 411 638 412 690
rect 464 638 465 690
rect 411 626 465 638
rect 411 574 412 626
rect 464 574 465 626
rect 411 562 465 574
rect 411 510 412 562
rect 464 510 465 562
rect 411 491 465 510
rect 511 491 539 824
rect 567 519 595 852
rect 623 491 651 824
rect 679 519 707 852
rect 810 842 876 852
rect 735 491 763 824
rect 113 485 763 491
rect 113 433 119 485
rect 171 433 183 485
rect 235 433 247 485
rect 299 433 311 485
rect 363 433 513 485
rect 565 433 577 485
rect 629 433 641 485
rect 693 433 705 485
rect 757 433 763 485
rect 113 427 763 433
rect 113 94 141 427
rect 0 66 66 76
rect 169 66 197 399
rect 225 94 253 427
rect 281 66 309 399
rect 337 94 365 427
rect 411 408 465 427
rect 411 356 412 408
rect 464 356 465 408
rect 411 344 465 356
rect 411 292 412 344
rect 464 292 465 344
rect 411 280 465 292
rect 411 228 412 280
rect 464 228 465 280
rect 411 216 465 228
rect 411 164 412 216
rect 464 164 465 216
rect 411 152 465 164
rect 411 100 412 152
rect 464 100 465 152
rect 411 94 465 100
rect 511 94 539 427
rect 567 66 595 399
rect 623 94 651 427
rect 679 66 707 399
rect 735 94 763 427
rect 810 790 817 842
rect 869 790 876 842
rect 810 778 876 790
rect 810 726 817 778
rect 869 726 876 778
rect 810 714 876 726
rect 810 662 817 714
rect 869 662 876 714
rect 810 658 826 662
rect 860 658 876 662
rect 810 650 876 658
rect 810 598 817 650
rect 869 598 876 650
rect 810 586 826 598
rect 860 586 876 598
rect 810 534 817 586
rect 869 534 876 586
rect 810 514 826 534
rect 860 514 876 534
rect 810 476 876 514
rect 810 442 826 476
rect 860 442 876 476
rect 810 404 876 442
rect 810 384 826 404
rect 860 384 876 404
rect 810 332 817 384
rect 869 332 876 384
rect 810 320 826 332
rect 860 320 876 332
rect 810 268 817 320
rect 869 268 876 320
rect 810 260 876 268
rect 810 256 826 260
rect 860 256 876 260
rect 810 204 817 256
rect 869 204 876 256
rect 810 192 876 204
rect 810 140 817 192
rect 869 140 876 192
rect 810 128 876 140
rect 810 76 817 128
rect 869 76 876 128
rect 810 66 876 76
rect 0 59 876 66
rect 0 7 52 59
rect 104 50 116 59
rect 168 50 180 59
rect 232 50 244 59
rect 168 16 169 50
rect 232 16 241 50
rect 104 7 116 16
rect 168 7 180 16
rect 232 7 244 16
rect 296 7 308 59
rect 360 50 516 59
rect 360 16 385 50
rect 419 16 457 50
rect 491 16 516 50
rect 360 7 516 16
rect 568 7 580 59
rect 632 50 644 59
rect 696 50 708 59
rect 760 50 772 59
rect 635 16 644 50
rect 707 16 708 50
rect 632 7 644 16
rect 696 7 708 16
rect 760 7 772 16
rect 824 7 876 59
rect 0 0 876 7
<< via1 >>
rect 52 902 104 911
rect 116 902 168 911
rect 180 902 232 911
rect 244 902 296 911
rect 52 868 97 902
rect 97 868 104 902
rect 116 868 131 902
rect 131 868 168 902
rect 180 868 203 902
rect 203 868 232 902
rect 244 868 275 902
rect 275 868 296 902
rect 52 859 104 868
rect 116 859 168 868
rect 180 859 232 868
rect 244 859 296 868
rect 308 902 360 911
rect 516 902 568 911
rect 308 868 313 902
rect 313 868 347 902
rect 347 868 360 902
rect 516 868 529 902
rect 529 868 563 902
rect 563 868 568 902
rect 308 859 360 868
rect 516 859 568 868
rect 580 902 632 911
rect 644 902 696 911
rect 708 902 760 911
rect 772 902 824 911
rect 580 868 601 902
rect 601 868 632 902
rect 644 868 673 902
rect 673 868 696 902
rect 708 868 745 902
rect 745 868 760 902
rect 772 868 779 902
rect 779 868 824 902
rect 580 859 632 868
rect 644 859 696 868
rect 708 859 760 868
rect 772 859 824 868
rect 7 836 59 842
rect 7 802 16 836
rect 16 802 50 836
rect 50 802 59 836
rect 7 790 59 802
rect 7 764 59 778
rect 7 730 16 764
rect 16 730 50 764
rect 50 730 59 764
rect 7 726 59 730
rect 7 692 59 714
rect 7 662 16 692
rect 16 662 50 692
rect 50 662 59 692
rect 7 620 59 650
rect 7 598 16 620
rect 16 598 50 620
rect 50 598 59 620
rect 7 548 59 586
rect 7 534 16 548
rect 16 534 50 548
rect 50 534 59 548
rect 7 370 16 384
rect 16 370 50 384
rect 50 370 59 384
rect 7 332 59 370
rect 7 298 16 320
rect 16 298 50 320
rect 50 298 59 320
rect 7 268 59 298
rect 7 226 16 256
rect 16 226 50 256
rect 50 226 59 256
rect 7 204 59 226
rect 7 188 59 192
rect 7 154 16 188
rect 16 154 50 188
rect 50 154 59 188
rect 7 140 59 154
rect 7 116 59 128
rect 7 82 16 116
rect 16 82 50 116
rect 50 82 59 116
rect 7 76 59 82
rect 412 766 464 818
rect 412 702 464 754
rect 412 638 464 690
rect 412 574 464 626
rect 412 510 464 562
rect 119 433 171 485
rect 183 433 235 485
rect 247 433 299 485
rect 311 433 363 485
rect 513 433 565 485
rect 577 433 629 485
rect 641 433 693 485
rect 705 433 757 485
rect 412 356 464 408
rect 412 292 464 344
rect 412 228 464 280
rect 412 164 464 216
rect 412 100 464 152
rect 817 836 869 842
rect 817 802 826 836
rect 826 802 860 836
rect 860 802 869 836
rect 817 790 869 802
rect 817 764 869 778
rect 817 730 826 764
rect 826 730 860 764
rect 860 730 869 764
rect 817 726 869 730
rect 817 692 869 714
rect 817 662 826 692
rect 826 662 860 692
rect 860 662 869 692
rect 817 620 869 650
rect 817 598 826 620
rect 826 598 860 620
rect 860 598 869 620
rect 817 548 869 586
rect 817 534 826 548
rect 826 534 860 548
rect 860 534 869 548
rect 817 370 826 384
rect 826 370 860 384
rect 860 370 869 384
rect 817 332 869 370
rect 817 298 826 320
rect 826 298 860 320
rect 860 298 869 320
rect 817 268 869 298
rect 817 226 826 256
rect 826 226 860 256
rect 860 226 869 256
rect 817 204 869 226
rect 817 188 869 192
rect 817 154 826 188
rect 826 154 860 188
rect 860 154 869 188
rect 817 140 869 154
rect 817 116 869 128
rect 817 82 826 116
rect 826 82 860 116
rect 860 82 869 116
rect 817 76 869 82
rect 52 50 104 59
rect 116 50 168 59
rect 180 50 232 59
rect 244 50 296 59
rect 52 16 97 50
rect 97 16 104 50
rect 116 16 131 50
rect 131 16 168 50
rect 180 16 203 50
rect 203 16 232 50
rect 244 16 275 50
rect 275 16 296 50
rect 52 7 104 16
rect 116 7 168 16
rect 180 7 232 16
rect 244 7 296 16
rect 308 50 360 59
rect 516 50 568 59
rect 308 16 313 50
rect 313 16 347 50
rect 347 16 360 50
rect 516 16 529 50
rect 529 16 563 50
rect 563 16 568 50
rect 308 7 360 16
rect 516 7 568 16
rect 580 50 632 59
rect 644 50 696 59
rect 708 50 760 59
rect 772 50 824 59
rect 580 16 601 50
rect 601 16 632 50
rect 644 16 673 50
rect 673 16 696 50
rect 708 16 745 50
rect 745 16 760 50
rect 772 16 779 50
rect 779 16 824 50
rect 580 7 632 16
rect 644 7 696 16
rect 708 7 760 16
rect 772 7 824 16
<< metal2 >>
rect 0 913 383 918
rect 0 911 78 913
rect 134 911 158 913
rect 214 911 238 913
rect 294 911 318 913
rect 0 859 52 911
rect 232 859 238 911
rect 296 859 308 911
rect 0 857 78 859
rect 134 857 158 859
rect 214 857 238 859
rect 294 857 318 859
rect 374 857 383 913
rect 0 852 383 857
rect 0 842 66 852
rect 0 819 7 842
rect 59 819 66 842
rect 411 824 465 918
rect 493 913 876 918
rect 493 857 502 913
rect 558 911 582 913
rect 638 911 662 913
rect 718 911 742 913
rect 798 911 876 913
rect 568 859 580 911
rect 638 859 644 911
rect 824 859 876 911
rect 558 857 582 859
rect 638 857 662 859
rect 718 857 742 859
rect 798 857 876 859
rect 493 852 876 857
rect 810 842 876 852
rect 0 763 5 819
rect 61 768 66 819
rect 94 818 782 824
rect 94 796 412 818
rect 61 763 382 768
rect 0 739 7 763
rect 59 740 382 763
rect 410 766 412 796
rect 464 796 782 818
rect 810 819 817 842
rect 869 819 876 842
rect 464 766 466 796
rect 810 768 815 819
rect 410 754 466 766
rect 59 739 66 740
rect 0 683 5 739
rect 61 683 66 739
rect 410 727 412 754
rect 464 727 466 754
rect 494 763 815 768
rect 871 763 876 819
rect 494 740 817 763
rect 94 684 410 712
rect 810 739 817 740
rect 869 739 876 763
rect 0 662 7 683
rect 59 662 66 683
rect 0 659 66 662
rect 0 603 5 659
rect 61 656 66 659
rect 466 684 782 712
rect 61 628 382 656
rect 410 647 412 671
rect 464 647 466 671
rect 810 683 815 739
rect 871 683 876 739
rect 810 662 817 683
rect 869 662 876 683
rect 810 659 876 662
rect 810 656 815 659
rect 61 603 66 628
rect 0 598 7 603
rect 59 598 66 603
rect 494 628 815 656
rect 0 586 66 598
rect 0 579 7 586
rect 59 579 66 586
rect 0 523 5 579
rect 61 544 66 579
rect 94 591 410 600
rect 810 603 815 628
rect 871 603 876 659
rect 466 591 782 600
rect 94 574 412 591
rect 464 574 782 591
rect 94 572 782 574
rect 810 598 817 603
rect 869 598 876 603
rect 810 586 876 598
rect 810 579 817 586
rect 869 579 876 586
rect 410 567 466 572
rect 61 523 382 544
rect 0 516 382 523
rect 0 514 66 516
rect 810 544 815 579
rect 494 523 815 544
rect 871 523 876 579
rect 494 516 876 523
rect 810 514 876 516
rect 410 510 412 511
rect 464 510 466 511
rect 410 487 466 510
rect 74 486 170 487
rect 0 485 170 486
rect 226 485 250 487
rect 306 485 330 487
rect 0 433 119 485
rect 235 433 247 485
rect 306 433 311 485
rect 0 432 170 433
rect 74 431 170 432
rect 226 431 250 433
rect 306 431 330 433
rect 386 431 410 487
rect 466 431 490 487
rect 546 485 570 487
rect 626 485 650 487
rect 706 486 802 487
rect 706 485 876 486
rect 565 433 570 485
rect 629 433 641 485
rect 757 433 876 485
rect 546 431 570 433
rect 626 431 650 433
rect 706 432 876 433
rect 706 431 802 432
rect 410 408 466 431
rect 410 407 412 408
rect 464 407 466 408
rect 0 402 66 404
rect 0 395 382 402
rect 0 339 5 395
rect 61 374 382 395
rect 61 339 66 374
rect 810 402 876 404
rect 494 395 876 402
rect 494 374 815 395
rect 410 346 466 351
rect 0 332 7 339
rect 59 332 66 339
rect 0 320 66 332
rect 0 315 7 320
rect 59 315 66 320
rect 94 344 782 346
rect 94 327 412 344
rect 464 327 782 344
rect 94 318 410 327
rect 0 259 5 315
rect 61 290 66 315
rect 466 318 782 327
rect 810 339 815 374
rect 871 339 876 395
rect 810 332 817 339
rect 869 332 876 339
rect 810 320 876 332
rect 61 262 382 290
rect 810 315 817 320
rect 869 315 876 320
rect 810 290 815 315
rect 61 259 66 262
rect 0 256 66 259
rect 0 235 7 256
rect 59 235 66 256
rect 0 179 5 235
rect 61 179 66 235
rect 410 247 412 271
rect 464 247 466 271
rect 494 262 815 290
rect 94 206 410 234
rect 810 259 815 262
rect 871 259 876 315
rect 810 256 876 259
rect 810 235 817 256
rect 869 235 876 256
rect 0 155 7 179
rect 59 178 66 179
rect 466 206 782 234
rect 59 155 382 178
rect 0 99 5 155
rect 61 150 382 155
rect 410 164 412 191
rect 464 164 466 191
rect 810 179 815 235
rect 871 179 876 235
rect 810 178 817 179
rect 410 152 466 164
rect 61 99 66 150
rect 410 122 412 152
rect 0 76 7 99
rect 59 76 66 99
rect 94 100 412 122
rect 464 122 466 152
rect 494 155 817 178
rect 869 155 876 179
rect 494 150 815 155
rect 464 100 782 122
rect 94 94 782 100
rect 810 99 815 150
rect 871 99 876 155
rect 0 66 66 76
rect 0 61 383 66
rect 0 59 78 61
rect 134 59 158 61
rect 214 59 238 61
rect 294 59 318 61
rect 0 7 52 59
rect 232 7 238 59
rect 296 7 308 59
rect 0 5 78 7
rect 134 5 158 7
rect 214 5 238 7
rect 294 5 318 7
rect 374 5 383 61
rect 0 0 383 5
rect 411 0 465 94
rect 810 76 817 99
rect 869 76 876 99
rect 810 66 876 76
rect 493 61 876 66
rect 493 5 502 61
rect 558 59 582 61
rect 638 59 662 61
rect 718 59 742 61
rect 798 59 876 61
rect 568 7 580 59
rect 638 7 644 59
rect 824 7 876 59
rect 558 5 582 7
rect 638 5 662 7
rect 718 5 742 7
rect 798 5 876 7
rect 493 0 876 5
<< via2 >>
rect 78 911 134 913
rect 158 911 214 913
rect 238 911 294 913
rect 318 911 374 913
rect 78 859 104 911
rect 104 859 116 911
rect 116 859 134 911
rect 158 859 168 911
rect 168 859 180 911
rect 180 859 214 911
rect 238 859 244 911
rect 244 859 294 911
rect 318 859 360 911
rect 360 859 374 911
rect 78 857 134 859
rect 158 857 214 859
rect 238 857 294 859
rect 318 857 374 859
rect 502 911 558 913
rect 582 911 638 913
rect 662 911 718 913
rect 742 911 798 913
rect 502 859 516 911
rect 516 859 558 911
rect 582 859 632 911
rect 632 859 638 911
rect 662 859 696 911
rect 696 859 708 911
rect 708 859 718 911
rect 742 859 760 911
rect 760 859 772 911
rect 772 859 798 911
rect 502 857 558 859
rect 582 857 638 859
rect 662 857 718 859
rect 742 857 798 859
rect 5 790 7 819
rect 7 790 59 819
rect 59 790 61 819
rect 5 778 61 790
rect 5 763 7 778
rect 7 763 59 778
rect 59 763 61 778
rect 815 790 817 819
rect 817 790 869 819
rect 869 790 871 819
rect 815 778 871 790
rect 5 726 7 739
rect 7 726 59 739
rect 59 726 61 739
rect 5 714 61 726
rect 5 683 7 714
rect 7 683 59 714
rect 59 683 61 714
rect 815 763 817 778
rect 817 763 869 778
rect 869 763 871 778
rect 410 702 412 727
rect 412 702 464 727
rect 464 702 466 727
rect 410 690 466 702
rect 5 650 61 659
rect 410 671 412 690
rect 412 671 464 690
rect 464 671 466 690
rect 5 603 7 650
rect 7 603 59 650
rect 59 603 61 650
rect 815 726 817 739
rect 817 726 869 739
rect 869 726 871 739
rect 815 714 871 726
rect 815 683 817 714
rect 817 683 869 714
rect 869 683 871 714
rect 410 638 412 647
rect 412 638 464 647
rect 464 638 466 647
rect 410 626 466 638
rect 815 650 871 659
rect 5 534 7 579
rect 7 534 59 579
rect 59 534 61 579
rect 410 591 412 626
rect 412 591 464 626
rect 464 591 466 626
rect 815 603 817 650
rect 817 603 869 650
rect 869 603 871 650
rect 410 562 466 567
rect 5 523 61 534
rect 410 511 412 562
rect 412 511 464 562
rect 464 511 466 562
rect 815 534 817 579
rect 817 534 869 579
rect 869 534 871 579
rect 815 523 871 534
rect 170 485 226 487
rect 250 485 306 487
rect 330 485 386 487
rect 170 433 171 485
rect 171 433 183 485
rect 183 433 226 485
rect 250 433 299 485
rect 299 433 306 485
rect 330 433 363 485
rect 363 433 386 485
rect 170 431 226 433
rect 250 431 306 433
rect 330 431 386 433
rect 410 431 466 487
rect 490 485 546 487
rect 570 485 626 487
rect 650 485 706 487
rect 490 433 513 485
rect 513 433 546 485
rect 570 433 577 485
rect 577 433 626 485
rect 650 433 693 485
rect 693 433 705 485
rect 705 433 706 485
rect 490 431 546 433
rect 570 431 626 433
rect 650 431 706 433
rect 5 384 61 395
rect 5 339 7 384
rect 7 339 59 384
rect 59 339 61 384
rect 410 356 412 407
rect 412 356 464 407
rect 464 356 466 407
rect 815 384 871 395
rect 410 351 466 356
rect 5 268 7 315
rect 7 268 59 315
rect 59 268 61 315
rect 410 292 412 327
rect 412 292 464 327
rect 464 292 466 327
rect 815 339 817 384
rect 817 339 869 384
rect 869 339 871 384
rect 5 259 61 268
rect 410 280 466 292
rect 410 271 412 280
rect 412 271 464 280
rect 464 271 466 280
rect 5 204 7 235
rect 7 204 59 235
rect 59 204 61 235
rect 5 192 61 204
rect 5 179 7 192
rect 7 179 59 192
rect 59 179 61 192
rect 815 268 817 315
rect 817 268 869 315
rect 869 268 871 315
rect 410 228 412 247
rect 412 228 464 247
rect 464 228 466 247
rect 815 259 871 268
rect 410 216 466 228
rect 410 191 412 216
rect 412 191 464 216
rect 464 191 466 216
rect 5 140 7 155
rect 7 140 59 155
rect 59 140 61 155
rect 815 204 817 235
rect 817 204 869 235
rect 869 204 871 235
rect 815 192 871 204
rect 815 179 817 192
rect 817 179 869 192
rect 869 179 871 192
rect 5 128 61 140
rect 5 99 7 128
rect 7 99 59 128
rect 59 99 61 128
rect 815 140 817 155
rect 817 140 869 155
rect 869 140 871 155
rect 815 128 871 140
rect 815 99 817 128
rect 817 99 869 128
rect 869 99 871 128
rect 78 59 134 61
rect 158 59 214 61
rect 238 59 294 61
rect 318 59 374 61
rect 78 7 104 59
rect 104 7 116 59
rect 116 7 134 59
rect 158 7 168 59
rect 168 7 180 59
rect 180 7 214 59
rect 238 7 244 59
rect 244 7 294 59
rect 318 7 360 59
rect 360 7 374 59
rect 78 5 134 7
rect 158 5 214 7
rect 238 5 294 7
rect 318 5 374 7
rect 502 59 558 61
rect 582 59 638 61
rect 662 59 718 61
rect 742 59 798 61
rect 502 7 516 59
rect 516 7 558 59
rect 582 7 632 59
rect 632 7 638 59
rect 662 7 696 59
rect 696 7 708 59
rect 708 7 718 59
rect 742 7 760 59
rect 760 7 772 59
rect 772 7 798 59
rect 502 5 558 7
rect 582 5 638 7
rect 662 5 718 7
rect 742 5 798 7
<< metal3 >>
rect 0 913 876 918
rect 0 857 78 913
rect 134 857 158 913
rect 214 857 238 913
rect 294 857 318 913
rect 374 857 502 913
rect 558 857 582 913
rect 638 857 662 913
rect 718 857 742 913
rect 798 857 876 913
rect 0 852 876 857
rect 0 819 66 852
rect 0 763 5 819
rect 61 763 66 819
rect 0 739 66 763
rect 0 683 5 739
rect 61 683 66 739
rect 0 659 66 683
rect 0 603 5 659
rect 61 603 66 659
rect 0 579 66 603
rect 0 523 5 579
rect 61 523 66 579
rect 0 395 66 523
rect 0 339 5 395
rect 61 339 66 395
rect 0 315 66 339
rect 0 259 5 315
rect 61 259 66 315
rect 0 235 66 259
rect 0 179 5 235
rect 61 179 66 235
rect 0 155 66 179
rect 0 99 5 155
rect 61 99 66 155
rect 126 492 186 792
rect 246 552 306 852
rect 405 727 471 792
rect 405 671 410 727
rect 466 671 471 727
rect 405 647 471 671
rect 405 591 410 647
rect 466 591 471 647
rect 405 567 471 591
rect 405 511 410 567
rect 466 511 471 567
rect 570 552 630 852
rect 810 819 876 852
rect 405 492 471 511
rect 690 492 750 792
rect 126 487 750 492
rect 126 431 170 487
rect 226 431 250 487
rect 306 431 330 487
rect 386 431 410 487
rect 466 431 490 487
rect 546 431 570 487
rect 626 431 650 487
rect 706 431 750 487
rect 126 426 750 431
rect 126 126 186 426
rect 405 407 471 426
rect 0 66 66 99
rect 246 66 306 366
rect 405 351 410 407
rect 466 351 471 407
rect 405 327 471 351
rect 405 271 410 327
rect 466 271 471 327
rect 405 247 471 271
rect 405 191 410 247
rect 466 191 471 247
rect 405 126 471 191
rect 570 66 630 366
rect 690 126 750 426
rect 810 763 815 819
rect 871 763 876 819
rect 810 739 876 763
rect 810 683 815 739
rect 871 683 876 739
rect 810 659 876 683
rect 810 603 815 659
rect 871 603 876 659
rect 810 579 876 603
rect 810 523 815 579
rect 871 523 876 579
rect 810 395 876 523
rect 810 339 815 395
rect 871 339 876 395
rect 810 315 876 339
rect 810 259 815 315
rect 871 259 876 315
rect 810 235 876 259
rect 810 179 815 235
rect 871 179 876 235
rect 810 155 876 179
rect 810 99 815 155
rect 871 99 876 155
rect 810 66 876 99
rect 0 61 876 66
rect 0 5 78 61
rect 134 5 158 61
rect 214 5 238 61
rect 294 5 318 61
rect 374 5 502 61
rect 558 5 582 61
rect 638 5 662 61
rect 718 5 742 61
rect 798 5 876 61
rect 0 0 876 5
<< labels >>
flabel metal2 s 292 870 319 897 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 421 868 451 900 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 467 350 491 401 0 FreeSans 200 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 74038
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 59990
<< end >>
