magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 19 21 917 203
rect 29 -17 63 21
<< scnmos >>
rect 102 47 132 177
rect 188 47 218 177
rect 397 47 427 177
rect 483 47 513 177
rect 588 47 618 177
rect 685 47 715 177
rect 793 47 823 177
<< scpmoshvt >>
rect 86 297 116 497
rect 172 297 202 497
rect 397 297 427 497
rect 469 297 499 497
rect 577 297 607 497
rect 685 297 715 497
rect 793 297 823 497
<< ndiff >>
rect 45 161 102 177
rect 45 127 53 161
rect 87 127 102 161
rect 45 93 102 127
rect 45 59 53 93
rect 87 59 102 93
rect 45 47 102 59
rect 132 169 188 177
rect 132 135 143 169
rect 177 135 188 169
rect 132 101 188 135
rect 132 67 143 101
rect 177 67 188 101
rect 132 47 188 67
rect 218 157 397 177
rect 218 123 229 157
rect 263 123 397 157
rect 218 89 397 123
rect 218 55 229 89
rect 263 55 352 89
rect 386 55 397 89
rect 218 47 397 55
rect 427 101 483 177
rect 427 67 438 101
rect 472 67 483 101
rect 427 47 483 67
rect 513 89 588 177
rect 513 55 534 89
rect 568 55 588 89
rect 513 47 588 55
rect 618 101 685 177
rect 618 67 629 101
rect 663 67 685 101
rect 618 47 685 67
rect 715 47 793 177
rect 823 161 891 177
rect 823 127 849 161
rect 883 127 891 161
rect 823 93 891 127
rect 823 59 849 93
rect 883 59 891 93
rect 823 47 891 59
<< pdiff >>
rect 33 485 86 497
rect 33 451 41 485
rect 75 451 86 485
rect 33 381 86 451
rect 33 347 41 381
rect 75 347 86 381
rect 33 297 86 347
rect 116 427 172 497
rect 116 393 127 427
rect 161 393 172 427
rect 116 359 172 393
rect 116 325 127 359
rect 161 325 172 359
rect 116 297 172 325
rect 202 485 255 497
rect 202 451 213 485
rect 247 451 255 485
rect 202 417 255 451
rect 202 383 213 417
rect 247 383 255 417
rect 202 349 255 383
rect 202 315 213 349
rect 247 315 255 349
rect 202 297 255 315
rect 315 477 397 497
rect 315 443 323 477
rect 357 443 397 477
rect 315 349 397 443
rect 315 315 323 349
rect 357 315 397 349
rect 315 297 397 315
rect 427 297 469 497
rect 499 297 577 497
rect 607 485 685 497
rect 607 451 630 485
rect 664 451 685 485
rect 607 417 685 451
rect 607 383 630 417
rect 664 383 685 417
rect 607 297 685 383
rect 715 485 793 497
rect 715 451 734 485
rect 768 451 793 485
rect 715 297 793 451
rect 823 485 876 497
rect 823 451 834 485
rect 868 451 876 485
rect 823 417 876 451
rect 823 383 834 417
rect 868 383 876 417
rect 823 297 876 383
<< ndiffc >>
rect 53 127 87 161
rect 53 59 87 93
rect 143 135 177 169
rect 143 67 177 101
rect 229 123 263 157
rect 229 55 263 89
rect 352 55 386 89
rect 438 67 472 101
rect 534 55 568 89
rect 629 67 663 101
rect 849 127 883 161
rect 849 59 883 93
<< pdiffc >>
rect 41 451 75 485
rect 41 347 75 381
rect 127 393 161 427
rect 127 325 161 359
rect 213 451 247 485
rect 213 383 247 417
rect 213 315 247 349
rect 323 443 357 477
rect 323 315 357 349
rect 630 451 664 485
rect 630 383 664 417
rect 734 451 768 485
rect 834 451 868 485
rect 834 383 868 417
<< poly >>
rect 86 497 116 523
rect 172 497 202 523
rect 397 497 427 523
rect 469 497 499 523
rect 577 497 607 523
rect 685 497 715 523
rect 793 497 823 523
rect 86 265 116 297
rect 172 265 202 297
rect 397 265 427 297
rect 86 249 283 265
rect 86 235 233 249
rect 102 215 233 235
rect 267 215 283 249
rect 102 199 283 215
rect 361 249 427 265
rect 361 215 377 249
rect 411 215 427 249
rect 361 199 427 215
rect 469 265 499 297
rect 577 265 607 297
rect 685 265 715 297
rect 793 265 823 297
rect 469 249 535 265
rect 469 215 485 249
rect 519 215 535 249
rect 469 199 535 215
rect 577 249 643 265
rect 577 215 593 249
rect 627 215 643 249
rect 577 199 643 215
rect 685 249 751 265
rect 685 215 701 249
rect 735 215 751 249
rect 102 177 132 199
rect 188 177 218 199
rect 397 177 427 199
rect 483 177 513 199
rect 588 177 618 199
rect 685 196 751 215
rect 793 249 859 265
rect 793 215 809 249
rect 843 215 859 249
rect 793 199 859 215
rect 685 177 715 196
rect 793 177 823 199
rect 102 21 132 47
rect 188 21 218 47
rect 397 21 427 47
rect 483 21 513 47
rect 588 21 618 47
rect 685 21 715 47
rect 793 21 823 47
<< polycont >>
rect 233 215 267 249
rect 377 215 411 249
rect 485 215 519 249
rect 593 215 627 249
rect 701 215 735 249
rect 809 215 843 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 17 485 87 527
rect 17 451 41 485
rect 75 451 87 485
rect 213 485 263 527
rect 17 381 87 451
rect 17 347 41 381
rect 75 347 87 381
rect 17 327 87 347
rect 121 427 179 478
rect 121 393 127 427
rect 161 393 179 427
rect 121 359 179 393
rect 121 325 127 359
rect 161 325 179 359
rect 17 161 87 177
rect 17 127 53 161
rect 17 93 87 127
rect 17 59 53 93
rect 17 17 87 59
rect 121 169 179 325
rect 247 451 263 485
rect 213 417 263 451
rect 247 383 263 417
rect 213 349 263 383
rect 247 315 263 349
rect 213 299 263 315
rect 299 477 357 493
rect 299 443 323 477
rect 614 485 680 493
rect 299 349 357 443
rect 299 315 323 349
rect 299 299 357 315
rect 299 265 341 299
rect 392 265 451 471
rect 213 249 341 265
rect 213 215 233 249
rect 267 215 341 249
rect 121 135 143 169
rect 177 135 179 169
rect 121 101 179 135
rect 121 67 143 101
rect 177 67 179 101
rect 121 51 179 67
rect 213 157 265 173
rect 213 123 229 157
rect 263 123 265 157
rect 299 157 341 215
rect 377 249 451 265
rect 411 215 451 249
rect 377 199 451 215
rect 485 249 547 471
rect 614 451 630 485
rect 664 451 680 485
rect 718 485 784 527
rect 718 451 734 485
rect 768 451 784 485
rect 818 485 903 493
rect 818 451 834 485
rect 868 451 903 485
rect 614 417 680 451
rect 818 417 903 451
rect 614 383 630 417
rect 664 383 834 417
rect 868 383 903 417
rect 519 215 547 249
rect 485 199 547 215
rect 581 249 639 348
rect 581 215 593 249
rect 627 215 639 249
rect 581 199 639 215
rect 673 249 755 348
rect 673 215 701 249
rect 735 215 755 249
rect 673 191 755 215
rect 789 249 903 348
rect 789 215 809 249
rect 843 215 903 249
rect 789 199 903 215
rect 701 165 755 191
rect 299 123 667 157
rect 213 89 265 123
rect 436 101 484 123
rect 213 55 229 89
rect 263 55 352 89
rect 386 55 402 89
rect 213 17 402 55
rect 436 67 438 101
rect 472 67 484 101
rect 618 101 667 123
rect 436 51 484 67
rect 518 55 534 89
rect 568 55 584 89
rect 518 17 584 55
rect 618 67 629 101
rect 663 67 667 101
rect 618 51 667 67
rect 701 58 799 165
rect 833 127 849 161
rect 883 127 903 161
rect 833 93 903 127
rect 833 59 849 93
rect 883 59 903 93
rect 833 17 903 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
flabel locali s 397 357 431 391 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 673 289 707 323 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 581 221 615 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 489 289 523 323 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 121 357 155 391 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 857 221 891 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 397 289 431 323 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 121 289 155 323 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 121 221 155 255 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 121 153 155 187 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 121 85 155 119 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 121 425 155 459 0 FreeSans 340 0 0 0 X
port 10 nsew signal output
flabel locali s 489 221 523 255 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 489 357 523 391 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 489 425 523 459 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 581 289 615 323 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 673 221 707 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 397 425 431 459 0 FreeSans 340 0 0 0 D1
port 5 nsew signal input
flabel locali s 765 85 799 119 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 857 289 891 323 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a2111o_2
rlabel metal1 s 0 -48 920 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 920 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 920 544
string GDS_END 3763378
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3754318
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 23.000 0.000 
<< end >>
