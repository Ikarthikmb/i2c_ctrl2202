magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 53 21 827 203
rect 53 17 64 21
rect 30 -17 64 17
<< scnmos >>
rect 131 47 161 177
rect 215 47 245 177
rect 299 47 329 177
rect 383 47 413 177
rect 467 47 497 177
rect 551 47 581 177
rect 635 47 665 177
rect 719 47 749 177
<< scpmoshvt >>
rect 131 297 161 497
rect 215 297 245 497
rect 299 297 329 497
rect 383 297 413 497
rect 467 297 497 497
rect 551 297 581 497
rect 635 297 665 497
rect 719 297 749 497
<< ndiff >>
rect 79 97 131 177
rect 79 63 87 97
rect 121 63 131 97
rect 79 47 131 63
rect 161 161 215 177
rect 161 127 171 161
rect 205 127 215 161
rect 161 93 215 127
rect 161 59 171 93
rect 205 59 215 93
rect 161 47 215 59
rect 245 97 299 177
rect 245 63 255 97
rect 289 63 299 97
rect 245 47 299 63
rect 329 129 383 177
rect 329 95 339 129
rect 373 95 383 129
rect 329 47 383 95
rect 413 97 467 177
rect 413 63 423 97
rect 457 63 467 97
rect 413 47 467 63
rect 497 129 551 177
rect 497 95 507 129
rect 541 95 551 129
rect 497 47 551 95
rect 581 97 635 177
rect 581 63 591 97
rect 625 63 635 97
rect 581 47 635 63
rect 665 129 719 177
rect 665 95 675 129
rect 709 95 719 129
rect 665 47 719 95
rect 749 161 801 177
rect 749 127 759 161
rect 793 127 801 161
rect 749 93 801 127
rect 749 59 759 93
rect 793 59 801 93
rect 749 47 801 59
<< pdiff >>
rect 79 485 131 497
rect 79 451 87 485
rect 121 451 131 485
rect 79 417 131 451
rect 79 383 87 417
rect 121 383 131 417
rect 79 349 131 383
rect 79 315 87 349
rect 121 315 131 349
rect 79 297 131 315
rect 161 479 215 497
rect 161 445 171 479
rect 205 445 215 479
rect 161 411 215 445
rect 161 377 171 411
rect 205 377 215 411
rect 161 343 215 377
rect 161 309 171 343
rect 205 309 215 343
rect 161 297 215 309
rect 245 485 299 497
rect 245 451 255 485
rect 289 451 299 485
rect 245 417 299 451
rect 245 383 255 417
rect 289 383 299 417
rect 245 297 299 383
rect 329 463 383 497
rect 329 429 339 463
rect 373 429 383 463
rect 329 368 383 429
rect 329 334 339 368
rect 373 334 383 368
rect 329 297 383 334
rect 413 485 467 497
rect 413 451 423 485
rect 457 451 467 485
rect 413 417 467 451
rect 413 383 423 417
rect 457 383 467 417
rect 413 297 467 383
rect 497 463 551 497
rect 497 429 507 463
rect 541 429 551 463
rect 497 368 551 429
rect 497 334 507 368
rect 541 334 551 368
rect 497 297 551 334
rect 581 485 635 497
rect 581 451 591 485
rect 625 451 635 485
rect 581 417 635 451
rect 581 383 591 417
rect 625 383 635 417
rect 581 297 635 383
rect 665 463 719 497
rect 665 429 675 463
rect 709 429 719 463
rect 665 368 719 429
rect 665 334 675 368
rect 709 334 719 368
rect 665 297 719 334
rect 749 485 801 497
rect 749 451 759 485
rect 793 451 801 485
rect 749 417 801 451
rect 749 383 759 417
rect 793 383 801 417
rect 749 349 801 383
rect 749 315 759 349
rect 793 315 801 349
rect 749 297 801 315
<< ndiffc >>
rect 87 63 121 97
rect 171 127 205 161
rect 171 59 205 93
rect 255 63 289 97
rect 339 95 373 129
rect 423 63 457 97
rect 507 95 541 129
rect 591 63 625 97
rect 675 95 709 129
rect 759 127 793 161
rect 759 59 793 93
<< pdiffc >>
rect 87 451 121 485
rect 87 383 121 417
rect 87 315 121 349
rect 171 445 205 479
rect 171 377 205 411
rect 171 309 205 343
rect 255 451 289 485
rect 255 383 289 417
rect 339 429 373 463
rect 339 334 373 368
rect 423 451 457 485
rect 423 383 457 417
rect 507 429 541 463
rect 507 334 541 368
rect 591 451 625 485
rect 591 383 625 417
rect 675 429 709 463
rect 675 334 709 368
rect 759 451 793 485
rect 759 383 793 417
rect 759 315 793 349
<< poly >>
rect 131 497 161 523
rect 215 497 245 523
rect 299 497 329 523
rect 383 497 413 523
rect 467 497 497 523
rect 551 497 581 523
rect 635 497 665 523
rect 719 497 749 523
rect 131 259 161 297
rect 215 259 245 297
rect 65 249 245 259
rect 65 215 92 249
rect 126 215 187 249
rect 221 215 245 249
rect 65 205 245 215
rect 131 177 161 205
rect 215 177 245 205
rect 299 259 329 297
rect 383 259 413 297
rect 467 259 497 297
rect 551 259 581 297
rect 635 259 665 297
rect 719 259 749 297
rect 299 249 749 259
rect 299 215 315 249
rect 349 215 749 249
rect 299 205 749 215
rect 299 177 329 205
rect 383 177 413 205
rect 467 177 497 205
rect 551 177 581 205
rect 635 177 665 205
rect 719 177 749 205
rect 131 21 161 47
rect 215 21 245 47
rect 299 21 329 47
rect 383 21 413 47
rect 467 21 497 47
rect 551 21 581 47
rect 635 21 665 47
rect 719 21 749 47
<< polycont >>
rect 92 215 126 249
rect 187 215 221 249
rect 315 215 349 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 87 485 121 527
rect 87 417 121 451
rect 87 349 121 383
rect 87 297 121 315
rect 155 479 221 493
rect 155 445 171 479
rect 205 445 221 479
rect 155 411 221 445
rect 155 377 171 411
rect 205 377 221 411
rect 155 343 221 377
rect 255 485 303 527
rect 289 451 303 485
rect 255 417 303 451
rect 289 383 303 417
rect 255 367 303 383
rect 339 463 373 493
rect 339 368 373 429
rect 155 309 171 343
rect 205 331 221 343
rect 407 485 473 527
rect 407 451 423 485
rect 457 451 473 485
rect 407 417 473 451
rect 407 383 423 417
rect 457 383 473 417
rect 407 367 473 383
rect 507 463 541 493
rect 507 368 541 429
rect 205 309 305 331
rect 155 297 305 309
rect 56 249 237 263
rect 56 215 92 249
rect 126 215 187 249
rect 221 215 237 249
rect 271 249 305 297
rect 339 323 373 334
rect 575 485 641 527
rect 575 451 591 485
rect 625 451 641 485
rect 575 417 641 451
rect 575 383 591 417
rect 625 383 641 417
rect 575 367 641 383
rect 675 463 709 493
rect 675 368 709 429
rect 507 323 541 334
rect 675 323 709 334
rect 339 289 709 323
rect 743 485 809 527
rect 743 451 759 485
rect 793 451 809 485
rect 743 417 809 451
rect 743 383 759 417
rect 793 383 809 417
rect 743 349 809 383
rect 743 315 759 349
rect 793 315 809 349
rect 743 297 809 315
rect 271 215 315 249
rect 349 215 365 249
rect 271 181 305 215
rect 442 181 709 289
rect 155 161 305 181
rect 155 127 171 161
rect 205 147 305 161
rect 339 147 709 181
rect 205 127 221 147
rect 87 97 121 113
rect 87 17 121 63
rect 155 93 221 127
rect 339 129 373 147
rect 155 59 171 93
rect 205 59 221 93
rect 155 51 221 59
rect 255 97 289 113
rect 255 17 289 63
rect 507 129 541 147
rect 339 51 373 95
rect 407 97 473 113
rect 407 63 423 97
rect 457 63 473 97
rect 407 17 473 63
rect 675 129 709 147
rect 507 51 541 95
rect 575 97 641 113
rect 575 63 591 97
rect 625 63 641 97
rect 575 17 641 63
rect 675 51 709 95
rect 743 161 809 177
rect 743 127 759 161
rect 793 127 809 161
rect 743 93 809 127
rect 743 59 759 93
rect 793 59 809 93
rect 743 17 809 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel locali s 442 221 476 255 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 442 289 476 323 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 442 153 476 187 0 FreeSans 200 0 0 0 X
port 6 nsew signal output
flabel locali s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 5 nsew power bidirectional abutment
flabel locali s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 2 nsew ground bidirectional abutment
flabel locali s 178 221 212 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 78 221 112 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 4 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 3 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 buf_6
rlabel metal1 s 0 -48 828 48 1 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 3104496
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3097518
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 20.700 13.600 
<< end >>
