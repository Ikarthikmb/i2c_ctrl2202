magic
tech sky130B
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__dfl1sd2__example_5595914180812  sky130_fd_pr__dfl1sd2__example_5595914180812_0
timestamp 1644511149
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180811  sky130_fd_pr__dfl1sd__example_5595914180811_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__dfl1sd__example_5595914180811  sky130_fd_pr__dfl1sd__example_5595914180811_1
timestamp 1644511149
transform 1 0 256 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 284 267 284 267 0 FreeSans 300 0 0 0 S
flabel comment s 128 267 128 267 0 FreeSans 300 0 0 0 D
flabel comment s -28 267 -28 267 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 35976956
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 35975392
<< end >>
