/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/rf_nfet_01v8_lvt/sky130_fd_pr__rf_nfet_01v8_lvt_bM02W3p00L0p18.spice