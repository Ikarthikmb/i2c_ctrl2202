/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/pfet_20v0/sky130_fd_pr__pfet_20v0__tt_discrete.corner.spice