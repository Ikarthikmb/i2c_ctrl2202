magic
tech sky130B
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__dfl1sd__example_5595914180815  sky130_fd_pr__dfl1sd__example_5595914180815_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_0
timestamp 1644511149
transform 1 0 180 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808100  sky130_fd_pr__hvdfl1sd__example_55959141808100_0
timestamp 1644511149
transform 1 0 416 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 444 97 444 97 0 FreeSans 300 0 0 0 D
flabel comment s 208 97 208 97 0 FreeSans 300 0 0 0 S
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 D
<< properties >>
string GDS_END 8098204
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8096698
<< end >>
