magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< labels >>
flabel comment s 125 300 125 300 0 FreeSans 300 0 0 0 D
flabel comment s -25 300 -25 300 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 7329348
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 7328580
<< end >>
