/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/npn_11v0/sky130_fd_pr__npn_11v0_W1p00L1p00.model.spice