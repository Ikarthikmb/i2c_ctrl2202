magic
tech sky130A
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdftpm1s2__example_55959141808649  sky130_fd_pr__hvdftpm1s2__example_55959141808649_0
timestamp 1644511149
transform -1 0 -91 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 145 500 145 500 0 FreeSans 300 0 0 0 D
flabel comment s -221 481 -221 481 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 3762036
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 3761178
<< end >>
