magic
tech sky130A
timestamp 1644511149
<< properties >>
string GDS_END 58740
string GDS_FILE $PDKPATH/libs.ref/sky130_sram_macros/gds/sky130_sram_1kbyte_1rw1r_8x1024_8.gds
string GDS_START 58416
<< end >>
