magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 1 21 911 203
rect 29 -17 63 21
<< locali >>
rect 17 199 75 394
rect 109 342 161 493
rect 295 342 333 493
rect 565 342 631 425
rect 109 308 631 342
rect 109 134 175 308
rect 209 215 381 273
rect 473 215 667 271
rect 712 249 891 259
rect 701 215 891 249
rect 823 153 891 215
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 23 435 75 527
rect 195 383 261 527
rect 367 383 433 527
rect 479 459 703 493
rect 479 420 531 459
rect 665 339 703 459
rect 737 373 803 527
rect 837 339 889 493
rect 665 305 889 339
rect 209 93 247 178
rect 281 127 789 169
rect 751 103 789 127
rect 209 89 433 93
rect 19 51 433 89
rect 479 17 545 89
rect 651 17 717 89
rect 823 17 889 89
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
<< metal1 >>
rect 0 561 920 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 920 561
rect 0 496 920 527
rect 0 17 920 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 920 17
rect 0 -48 920 -17
<< labels >>
rlabel locali s 823 153 891 215 6 A1
port 1 nsew signal input
rlabel locali s 701 215 891 249 6 A1
port 1 nsew signal input
rlabel locali s 712 249 891 259 6 A1
port 1 nsew signal input
rlabel locali s 473 215 667 271 6 A2
port 2 nsew signal input
rlabel locali s 209 215 381 273 6 B1
port 3 nsew signal input
rlabel locali s 17 199 75 394 6 C1
port 4 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 911 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 109 134 175 308 6 Y
port 9 nsew signal output
rlabel locali s 109 308 631 342 6 Y
port 9 nsew signal output
rlabel locali s 565 342 631 425 6 Y
port 9 nsew signal output
rlabel locali s 295 342 333 493 6 Y
port 9 nsew signal output
rlabel locali s 109 342 161 493 6 Y
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 920 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 792940
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 785544
<< end >>
