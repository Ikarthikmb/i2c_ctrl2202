magic
tech sky130B
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 1 21 1169 203
rect 29 -17 63 21
<< locali >>
rect 103 333 169 419
rect 555 333 621 417
rect 103 299 621 333
rect 18 215 169 265
rect 203 215 341 265
rect 375 221 434 299
rect 375 181 409 221
rect 481 215 613 265
rect 674 215 896 265
rect 950 215 1173 265
rect 103 131 409 181
<< obsli1 >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 18 459 253 493
rect 18 299 69 459
rect 203 401 253 459
rect 287 435 321 527
rect 355 401 421 491
rect 203 367 421 401
rect 467 451 877 489
rect 467 367 517 451
rect 655 299 689 451
rect 723 333 789 417
rect 827 367 877 451
rect 924 367 965 527
rect 999 333 1065 492
rect 723 299 1065 333
rect 1099 299 1143 527
rect 18 97 69 181
rect 447 143 1151 181
rect 447 97 481 143
rect 18 51 481 97
rect 524 17 590 109
rect 627 51 693 143
rect 727 17 761 109
rect 811 51 945 143
rect 981 17 1047 109
rect 1085 51 1151 143
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< obsli1c >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
rlabel locali s 950 215 1173 265 6 A1
port 1 nsew signal input
rlabel locali s 674 215 896 265 6 A2
port 2 nsew signal input
rlabel locali s 481 215 613 265 6 A3
port 3 nsew signal input
rlabel locali s 203 215 341 265 6 B1
port 4 nsew signal input
rlabel locali s 18 215 169 265 6 B2
port 5 nsew signal input
rlabel metal1 s 0 -48 1196 48 8 VGND
port 6 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 7 nsew ground bidirectional
rlabel pwell s 1 21 1169 203 6 VNB
port 7 nsew ground bidirectional
rlabel nwell s -38 261 1234 582 6 VPB
port 8 nsew power bidirectional
rlabel metal1 s 0 496 1196 592 6 VPWR
port 9 nsew power bidirectional abutment
rlabel locali s 103 131 409 181 6 Y
port 10 nsew signal output
rlabel locali s 375 181 409 221 6 Y
port 10 nsew signal output
rlabel locali s 375 221 434 299 6 Y
port 10 nsew signal output
rlabel locali s 103 299 621 333 6 Y
port 10 nsew signal output
rlabel locali s 555 333 621 417 6 Y
port 10 nsew signal output
rlabel locali s 103 333 169 419 6 Y
port 10 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1196 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1516096
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1506170
<< end >>
