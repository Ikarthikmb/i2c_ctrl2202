magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -66 377 450 897
<< pwell >>
rect 16 43 378 295
rect -26 -43 410 43
<< obsli1 >>
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 384 831
rect 50 746 340 751
rect 50 712 99 746
rect 133 712 172 746
rect 206 712 260 746
rect 294 712 340 746
rect 50 537 340 712
rect 95 250 161 406
rect 203 340 269 537
rect 95 169 356 250
rect 34 113 356 169
rect 34 79 43 113
rect 77 79 131 113
rect 165 79 219 113
rect 253 79 302 113
rect 336 79 356 113
rect 34 73 356 79
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
<< obsli1c >>
rect 31 797 65 831
rect 127 797 161 831
rect 223 797 257 831
rect 319 797 353 831
rect 99 712 133 746
rect 172 712 206 746
rect 260 712 294 746
rect 43 79 77 113
rect 131 79 165 113
rect 219 79 253 113
rect 302 79 336 113
rect 31 -17 65 17
rect 127 -17 161 17
rect 223 -17 257 17
rect 319 -17 353 17
<< metal1 >>
rect 0 831 384 837
rect 0 797 31 831
rect 65 797 127 831
rect 161 797 223 831
rect 257 797 319 831
rect 353 797 384 831
rect 0 791 384 797
rect 0 746 384 763
rect 0 712 99 746
rect 133 712 172 746
rect 206 712 260 746
rect 294 712 384 746
rect 0 689 384 712
rect 0 113 384 125
rect 0 79 43 113
rect 77 79 131 113
rect 165 79 219 113
rect 253 79 302 113
rect 336 79 384 113
rect 0 51 384 79
rect 0 17 384 23
rect 0 -17 31 17
rect 65 -17 127 17
rect 161 -17 223 17
rect 257 -17 319 17
rect 353 -17 384 17
rect 0 -23 384 -17
<< labels >>
rlabel metal1 s 0 51 384 125 6 VGND
port 1 nsew ground bidirectional
rlabel metal1 s 0 -23 384 23 8 VNB
port 2 nsew ground bidirectional
rlabel pwell s -26 -43 410 43 8 VNB
port 2 nsew ground bidirectional
rlabel pwell s 16 43 378 295 6 VNB
port 2 nsew ground bidirectional
rlabel metal1 s 0 791 384 837 6 VPB
port 3 nsew power bidirectional
rlabel nwell s -66 377 450 897 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 0 689 384 763 6 VPWR
port 4 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 384 814
string LEFclass CORE
string LEFsite unithv
string LEFsymmetry X Y
string LEFview TRUE
string GDS_END 959862
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hvl/gds/sky130_fd_sc_hvl.gds
string GDS_START 955112
<< end >>
