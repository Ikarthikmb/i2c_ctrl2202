/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/open_pdks/sources/sky130_sram_macros/sky130_sram_1kbyte_1rw1r_8x1024_8/sky130_sram_1kbyte_1rw1r_8x1024_8.lef