/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/open_pdks/sources/sky130_sram_macros/sky130_sram_2kbyte_1rw1r_32x512_8/sky130_sram_2kbyte_1rw1r_32x512_8.lef