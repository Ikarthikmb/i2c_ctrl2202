magic
tech sky130A
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__dfl1sd2__example_5595914180816  sky130_fd_pr__dfl1sd2__example_5595914180816_0
timestamp 1644511149
transform 1 0 50 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808140  sky130_fd_pr__hvdfl1sd2__example_55959141808140_1
timestamp 1644511149
transform 1 0 156 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 184 97 184 97 0 FreeSans 300 0 0 0 S
flabel comment s 78 97 78 97 0 FreeSans 300 0 0 0 D
flabel comment s -28 97 -28 97 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 6778292
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 6776912
<< end >>
