magic
tech sky130A
timestamp 1644511149
<< properties >>
string GDS_END 29783240
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 29774660
<< end >>
