magic
tech sky130A
magscale 1 2
timestamp 1644511149
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 1366 157 1839 203
rect 1 21 1839 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 258 47 288 119
rect 368 47 398 119
rect 464 47 494 131
rect 572 47 602 131
rect 762 47 792 131
rect 847 47 877 131
rect 1035 47 1065 131
rect 1142 47 1172 119
rect 1252 47 1282 119
rect 1347 47 1377 131
rect 1448 47 1478 177
rect 1532 47 1562 177
rect 1632 47 1662 177
rect 1716 47 1746 177
<< scpmoshvt >>
rect 79 369 109 497
rect 163 369 193 497
rect 259 413 289 497
rect 343 413 373 497
rect 487 345 517 473
rect 571 345 601 473
rect 759 316 789 424
rect 843 316 873 424
rect 1031 369 1061 497
rect 1166 413 1196 497
rect 1250 413 1280 497
rect 1351 369 1381 497
rect 1448 297 1478 497
rect 1532 297 1562 497
rect 1632 297 1662 497
rect 1716 297 1746 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 243 131
rect 413 119 464 131
rect 193 47 258 119
rect 288 107 368 119
rect 288 73 311 107
rect 345 73 368 107
rect 288 47 368 73
rect 398 47 464 119
rect 494 93 572 131
rect 494 59 515 93
rect 549 59 572 93
rect 494 47 572 59
rect 602 93 656 131
rect 602 59 614 93
rect 648 59 656 93
rect 602 47 656 59
rect 710 119 762 131
rect 710 85 718 119
rect 752 85 762 119
rect 710 47 762 85
rect 792 119 847 131
rect 792 85 803 119
rect 837 85 847 119
rect 792 47 847 85
rect 877 101 929 131
rect 877 67 887 101
rect 921 67 929 101
rect 877 47 929 67
rect 983 93 1035 131
rect 983 59 991 93
rect 1025 59 1035 93
rect 983 47 1035 59
rect 1065 119 1127 131
rect 1392 131 1448 177
rect 1297 119 1347 131
rect 1065 47 1142 119
rect 1172 93 1252 119
rect 1172 59 1195 93
rect 1229 59 1252 93
rect 1172 47 1252 59
rect 1282 47 1347 119
rect 1377 119 1448 131
rect 1377 85 1404 119
rect 1438 85 1448 119
rect 1377 47 1448 85
rect 1478 129 1532 177
rect 1478 95 1488 129
rect 1522 95 1532 129
rect 1478 47 1532 95
rect 1562 161 1632 177
rect 1562 127 1588 161
rect 1622 127 1632 161
rect 1562 93 1632 127
rect 1562 59 1588 93
rect 1622 59 1632 93
rect 1562 47 1632 59
rect 1662 129 1716 177
rect 1662 95 1672 129
rect 1706 95 1716 129
rect 1662 47 1716 95
rect 1746 161 1813 177
rect 1746 127 1771 161
rect 1805 127 1813 161
rect 1746 93 1813 127
rect 1746 59 1771 93
rect 1805 59 1813 93
rect 1746 47 1813 59
<< pdiff >>
rect 27 459 79 497
rect 27 425 35 459
rect 69 425 79 459
rect 27 369 79 425
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 369 163 451
rect 193 413 259 497
rect 289 459 343 497
rect 289 425 299 459
rect 333 425 343 459
rect 289 413 343 425
rect 373 473 472 497
rect 373 413 487 473
rect 193 369 244 413
rect 429 345 487 413
rect 517 461 571 473
rect 517 427 527 461
rect 561 427 571 461
rect 517 345 571 427
rect 601 391 653 473
rect 979 451 1031 497
rect 601 357 611 391
rect 645 357 653 391
rect 601 345 653 357
rect 707 412 759 424
rect 707 378 715 412
rect 749 378 759 412
rect 707 316 759 378
rect 789 362 843 424
rect 789 328 799 362
rect 833 328 843 362
rect 789 316 843 328
rect 873 363 925 424
rect 979 417 987 451
rect 1021 417 1031 451
rect 979 369 1031 417
rect 1061 413 1166 497
rect 1196 465 1250 497
rect 1196 431 1206 465
rect 1240 431 1250 465
rect 1196 413 1250 431
rect 1280 413 1351 497
rect 1061 369 1111 413
rect 873 329 883 363
rect 917 329 925 363
rect 873 316 925 329
rect 1295 369 1351 413
rect 1381 485 1448 497
rect 1381 451 1404 485
rect 1438 451 1448 485
rect 1381 417 1448 451
rect 1381 383 1404 417
rect 1438 383 1448 417
rect 1381 369 1448 383
rect 1396 297 1448 369
rect 1478 475 1532 497
rect 1478 441 1488 475
rect 1522 441 1532 475
rect 1478 401 1532 441
rect 1478 367 1488 401
rect 1522 367 1532 401
rect 1478 297 1532 367
rect 1562 485 1632 497
rect 1562 451 1588 485
rect 1622 451 1632 485
rect 1562 417 1632 451
rect 1562 383 1588 417
rect 1622 383 1632 417
rect 1562 349 1632 383
rect 1562 315 1588 349
rect 1622 315 1632 349
rect 1562 297 1632 315
rect 1662 475 1716 497
rect 1662 441 1672 475
rect 1706 441 1716 475
rect 1662 349 1716 441
rect 1662 315 1672 349
rect 1706 315 1716 349
rect 1662 297 1716 315
rect 1746 485 1813 497
rect 1746 451 1771 485
rect 1805 451 1813 485
rect 1746 417 1813 451
rect 1746 383 1771 417
rect 1805 383 1813 417
rect 1746 349 1813 383
rect 1746 315 1771 349
rect 1805 315 1813 349
rect 1746 297 1813 315
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 311 73 345 107
rect 515 59 549 93
rect 614 59 648 93
rect 718 85 752 119
rect 803 85 837 119
rect 887 67 921 101
rect 991 59 1025 93
rect 1195 59 1229 93
rect 1404 85 1438 119
rect 1488 95 1522 129
rect 1588 127 1622 161
rect 1588 59 1622 93
rect 1672 95 1706 129
rect 1771 127 1805 161
rect 1771 59 1805 93
<< pdiffc >>
rect 35 425 69 459
rect 119 451 153 485
rect 299 425 333 459
rect 527 427 561 461
rect 611 357 645 391
rect 715 378 749 412
rect 799 328 833 362
rect 987 417 1021 451
rect 1206 431 1240 465
rect 883 329 917 363
rect 1404 451 1438 485
rect 1404 383 1438 417
rect 1488 441 1522 475
rect 1488 367 1522 401
rect 1588 451 1622 485
rect 1588 383 1622 417
rect 1588 315 1622 349
rect 1672 441 1706 475
rect 1672 315 1706 349
rect 1771 451 1805 485
rect 1771 383 1805 417
rect 1771 315 1805 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 259 497 289 523
rect 343 497 373 523
rect 487 473 517 523
rect 571 493 873 523
rect 1031 497 1061 523
rect 1166 497 1196 523
rect 1250 497 1280 523
rect 1351 497 1381 523
rect 1448 497 1478 523
rect 1532 497 1562 523
rect 1632 497 1662 523
rect 1716 497 1746 523
rect 571 473 601 493
rect 79 265 109 369
rect 21 249 109 265
rect 21 215 32 249
rect 66 215 109 249
rect 163 219 193 369
rect 259 323 289 413
rect 343 375 373 413
rect 235 307 289 323
rect 331 365 397 375
rect 331 331 347 365
rect 381 331 397 365
rect 759 424 789 450
rect 843 424 873 493
rect 331 321 397 331
rect 487 330 517 345
rect 235 273 245 307
rect 279 279 289 307
rect 464 300 517 330
rect 279 273 398 279
rect 235 257 398 273
rect 259 249 398 257
rect 21 199 109 215
rect 79 131 109 199
rect 158 203 212 219
rect 158 169 168 203
rect 202 169 212 203
rect 158 153 212 169
rect 258 191 326 207
rect 258 157 282 191
rect 316 157 326 191
rect 163 131 193 153
rect 258 141 326 157
rect 258 119 288 141
rect 368 119 398 249
rect 464 219 494 300
rect 571 219 601 345
rect 1166 375 1196 413
rect 759 272 789 316
rect 843 290 873 316
rect 1031 279 1061 369
rect 1142 365 1208 375
rect 1142 331 1158 365
rect 1192 331 1208 365
rect 1142 321 1208 331
rect 1250 315 1280 413
rect 1250 299 1304 315
rect 1250 279 1260 299
rect 647 262 789 272
rect 647 228 663 262
rect 697 248 789 262
rect 980 263 1061 279
rect 697 228 877 248
rect 455 203 509 219
rect 455 169 465 203
rect 499 169 509 203
rect 455 153 509 169
rect 551 203 605 219
rect 647 218 877 228
rect 551 169 561 203
rect 595 176 605 203
rect 595 169 792 176
rect 551 153 792 169
rect 464 131 494 153
rect 570 146 792 153
rect 572 131 602 146
rect 762 131 792 146
rect 847 131 877 218
rect 980 229 990 263
rect 1024 243 1061 263
rect 1142 265 1260 279
rect 1294 265 1304 299
rect 1351 265 1381 369
rect 1448 265 1478 297
rect 1532 265 1562 297
rect 1632 265 1662 297
rect 1716 265 1746 297
rect 1142 249 1304 265
rect 1346 249 1400 265
rect 1024 229 1065 243
rect 980 213 1065 229
rect 1035 131 1065 213
rect 1142 119 1172 249
rect 1346 215 1356 249
rect 1390 215 1400 249
rect 1214 191 1282 207
rect 1346 199 1400 215
rect 1442 249 1746 265
rect 1442 215 1452 249
rect 1486 215 1746 249
rect 1442 199 1746 215
rect 1214 157 1224 191
rect 1258 157 1282 191
rect 1214 141 1282 157
rect 1252 119 1282 141
rect 1347 131 1377 199
rect 1448 177 1478 199
rect 1532 177 1562 199
rect 1632 177 1662 199
rect 1716 177 1746 199
rect 79 21 109 47
rect 163 21 193 47
rect 258 21 288 47
rect 368 21 398 47
rect 464 21 494 47
rect 572 21 602 47
rect 762 21 792 47
rect 847 21 877 47
rect 1035 21 1065 47
rect 1142 21 1172 47
rect 1252 21 1282 47
rect 1347 21 1377 47
rect 1448 21 1478 47
rect 1532 21 1562 47
rect 1632 21 1662 47
rect 1716 21 1746 47
<< polycont >>
rect 32 215 66 249
rect 347 331 381 365
rect 245 273 279 307
rect 168 169 202 203
rect 282 157 316 191
rect 1158 331 1192 365
rect 663 228 697 262
rect 465 169 499 203
rect 561 169 595 203
rect 990 229 1024 263
rect 1260 265 1294 299
rect 1356 215 1390 249
rect 1452 215 1486 249
rect 1224 157 1258 191
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 103 485 169 527
rect 27 459 69 475
rect 27 425 35 459
rect 103 451 119 485
rect 153 451 169 485
rect 520 461 566 527
rect 283 425 299 459
rect 333 425 398 459
rect 432 425 449 459
rect 27 417 69 425
rect 27 391 134 417
rect 27 383 306 391
rect 100 357 306 383
rect 340 365 381 391
rect 340 357 347 365
rect 30 323 66 349
rect 64 289 66 323
rect 30 249 66 289
rect 30 215 32 249
rect 30 195 66 215
rect 100 161 134 357
rect 313 331 347 357
rect 202 289 214 323
rect 248 307 279 323
rect 245 257 279 273
rect 313 315 381 331
rect 27 127 134 161
rect 168 203 248 219
rect 313 207 347 315
rect 415 281 449 425
rect 520 427 527 461
rect 561 427 566 461
rect 520 411 566 427
rect 662 425 674 459
rect 708 425 765 459
rect 715 412 765 425
rect 595 357 611 391
rect 645 357 664 391
rect 749 378 765 412
rect 715 362 765 378
rect 630 332 664 357
rect 630 298 684 332
rect 202 169 248 203
rect 168 153 248 169
rect 27 119 69 127
rect 27 85 35 119
rect 27 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 205 79 248 153
rect 282 191 347 207
rect 316 157 347 191
rect 282 141 347 157
rect 381 247 449 281
rect 650 278 684 298
rect 381 107 415 247
rect 483 203 524 264
rect 449 169 465 203
rect 499 169 524 203
rect 449 143 524 169
rect 558 203 616 264
rect 558 169 561 203
rect 595 169 616 203
rect 558 143 616 169
rect 650 262 697 278
rect 650 228 663 262
rect 650 212 697 228
rect 295 73 311 107
rect 345 73 415 107
rect 491 93 557 109
rect 650 93 684 212
rect 731 135 765 362
rect 103 17 169 59
rect 491 59 515 93
rect 549 59 557 93
rect 598 59 614 93
rect 648 59 684 93
rect 718 119 765 135
rect 752 85 765 119
rect 718 69 765 85
rect 799 425 858 459
rect 892 425 904 459
rect 952 451 1021 527
rect 1404 485 1438 527
rect 799 362 837 425
rect 952 417 987 451
rect 952 401 1021 417
rect 1066 431 1206 465
rect 1240 431 1256 465
rect 833 328 837 362
rect 799 119 837 328
rect 799 85 803 119
rect 799 69 837 85
rect 880 363 918 379
rect 880 329 883 363
rect 917 347 918 363
rect 1066 347 1100 431
rect 1306 425 1318 459
rect 1352 425 1370 459
rect 917 329 1100 347
rect 880 313 1100 329
rect 880 117 914 313
rect 950 263 1024 279
rect 950 229 990 263
rect 950 143 1024 229
rect 880 101 921 117
rect 880 67 887 101
rect 491 17 557 59
rect 880 51 921 67
rect 960 93 1026 109
rect 960 59 991 93
rect 1025 59 1026 93
rect 1066 93 1100 313
rect 1134 391 1192 397
rect 1168 365 1192 391
rect 1134 331 1158 357
rect 1134 207 1192 331
rect 1336 333 1370 425
rect 1404 417 1438 451
rect 1404 367 1438 383
rect 1472 475 1554 491
rect 1472 441 1488 475
rect 1522 441 1554 475
rect 1472 401 1554 441
rect 1472 367 1488 401
rect 1522 367 1554 401
rect 1226 323 1294 329
rect 1260 299 1294 323
rect 1336 299 1458 333
rect 1492 299 1554 367
rect 1588 485 1638 527
rect 1622 451 1638 485
rect 1588 417 1638 451
rect 1622 383 1638 417
rect 1588 349 1638 383
rect 1622 315 1638 349
rect 1588 299 1638 315
rect 1672 475 1737 491
rect 1706 441 1737 475
rect 1672 349 1737 441
rect 1706 315 1737 349
rect 1226 265 1260 289
rect 1424 265 1458 299
rect 1226 249 1294 265
rect 1328 249 1390 265
rect 1328 215 1356 249
rect 1134 191 1258 207
rect 1134 157 1224 191
rect 1134 141 1258 157
rect 1308 199 1390 215
rect 1424 249 1486 265
rect 1424 215 1452 249
rect 1424 199 1486 215
rect 1520 261 1554 299
rect 1672 261 1737 315
rect 1771 485 1821 527
rect 1805 451 1821 485
rect 1771 417 1821 451
rect 1805 383 1821 417
rect 1771 349 1821 383
rect 1805 315 1821 349
rect 1771 299 1821 315
rect 1520 213 1737 261
rect 1066 59 1195 93
rect 1229 59 1245 93
rect 1308 75 1370 199
rect 1404 119 1454 163
rect 1520 145 1554 213
rect 1438 85 1454 119
rect 960 17 1026 59
rect 1404 17 1454 85
rect 1488 129 1554 145
rect 1522 95 1554 129
rect 1488 53 1554 95
rect 1588 161 1638 177
rect 1622 127 1638 161
rect 1588 93 1638 127
rect 1622 59 1638 93
rect 1588 17 1638 59
rect 1672 129 1737 213
rect 1706 95 1737 129
rect 1672 53 1737 95
rect 1771 161 1821 177
rect 1805 127 1821 161
rect 1771 93 1821 127
rect 1805 59 1821 93
rect 1771 17 1821 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 398 425 432 459
rect 306 357 340 391
rect 30 289 64 323
rect 214 307 248 323
rect 214 289 245 307
rect 245 289 248 307
rect 674 425 708 459
rect 858 425 892 459
rect 1318 425 1352 459
rect 1134 365 1168 391
rect 1134 357 1158 365
rect 1158 357 1168 365
rect 1226 289 1260 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
<< metal1 >>
rect 0 561 1840 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1840 561
rect 0 496 1840 527
rect 386 459 444 465
rect 386 425 398 459
rect 432 456 444 459
rect 662 459 720 465
rect 662 456 674 459
rect 432 428 674 456
rect 432 425 444 428
rect 386 419 444 425
rect 662 425 674 428
rect 708 425 720 459
rect 662 419 720 425
rect 846 459 904 465
rect 846 425 858 459
rect 892 456 904 459
rect 1306 459 1364 465
rect 1306 456 1318 459
rect 892 428 1318 456
rect 892 425 904 428
rect 846 419 904 425
rect 1306 425 1318 428
rect 1352 425 1364 459
rect 1306 419 1364 425
rect 294 391 352 397
rect 294 357 306 391
rect 340 388 352 391
rect 1122 391 1180 397
rect 1122 388 1134 391
rect 340 360 1134 388
rect 340 357 352 360
rect 294 351 352 357
rect 1122 357 1134 360
rect 1168 357 1180 391
rect 1122 351 1180 357
rect 17 323 76 329
rect 17 289 30 323
rect 64 320 76 323
rect 202 323 260 329
rect 202 320 214 323
rect 64 292 214 320
rect 64 289 76 292
rect 17 283 76 289
rect 202 289 214 292
rect 248 320 260 323
rect 1214 323 1272 329
rect 1214 320 1226 323
rect 248 292 1226 320
rect 248 289 260 292
rect 202 283 260 289
rect 1214 289 1226 292
rect 1260 289 1272 323
rect 1214 283 1272 289
rect 0 17 1840 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1840 17
rect 0 -48 1840 -17
<< labels >>
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 8 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 9 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 7 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 10 nsew power bidirectional abutment
flabel locali s 1686 85 1720 119 0 FreeSans 400 0 0 0 X
port 11 nsew signal output
flabel locali s 1686 153 1720 187 0 FreeSans 400 0 0 0 X
port 11 nsew signal output
flabel locali s 1686 221 1720 255 0 FreeSans 400 0 0 0 X
port 11 nsew signal output
flabel locali s 1686 289 1720 323 0 FreeSans 400 0 0 0 X
port 11 nsew signal output
flabel locali s 1686 357 1720 391 0 FreeSans 400 0 0 0 X
port 11 nsew signal output
flabel locali s 1686 425 1720 459 0 FreeSans 400 0 0 0 X
port 11 nsew signal output
flabel locali s 30 221 64 255 0 FreeSans 400 0 0 0 S0
port 5 nsew signal input
flabel locali s 30 289 64 323 0 FreeSans 400 0 0 0 S0
port 5 nsew signal input
flabel locali s 214 153 248 187 0 FreeSans 400 0 0 0 A2
port 3 nsew signal input
flabel locali s 214 85 248 119 0 FreeSans 400 0 0 0 A2
port 3 nsew signal input
flabel locali s 490 153 524 187 0 FreeSans 400 0 0 0 A3
port 4 nsew signal input
flabel locali s 490 221 524 255 0 FreeSans 400 0 0 0 A3
port 4 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 400 0 0 0 S1
port 6 nsew signal input
flabel locali s 582 153 616 187 0 FreeSans 400 0 0 0 S1
port 6 nsew signal input
flabel locali s 950 221 984 255 0 FreeSans 400 0 0 0 A1
port 2 nsew signal input
flabel locali s 950 153 984 187 0 FreeSans 400 0 0 0 A1
port 2 nsew signal input
flabel locali s 1318 153 1352 187 0 FreeSans 400 0 0 0 A0
port 1 nsew signal input
flabel locali s 1318 85 1352 119 0 FreeSans 400 0 0 0 A0
port 1 nsew signal input
rlabel comment s 0 0 0 0 4 mux4_4
rlabel locali s 245 257 279 289 1 S0
port 5 nsew signal input
rlabel locali s 202 289 279 323 1 S0
port 5 nsew signal input
rlabel locali s 1226 249 1294 329 1 S0
port 5 nsew signal input
rlabel metal1 s 1214 320 1272 329 1 S0
port 5 nsew signal input
rlabel metal1 s 1214 283 1272 292 1 S0
port 5 nsew signal input
rlabel metal1 s 202 320 260 329 1 S0
port 5 nsew signal input
rlabel metal1 s 202 283 260 292 1 S0
port 5 nsew signal input
rlabel metal1 s 17 320 76 329 1 S0
port 5 nsew signal input
rlabel metal1 s 17 292 1272 320 1 S0
port 5 nsew signal input
rlabel metal1 s 17 283 76 292 1 S0
port 5 nsew signal input
rlabel metal1 s 0 -48 1840 48 1 VGND
port 7 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1840 592 1 VPWR
port 10 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1840 544
string GDS_END 1789346
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1773738
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 13.600 46.000 13.600 
<< end >>
