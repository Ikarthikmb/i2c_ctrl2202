magic
tech sky130A
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_0
timestamp 1644511149
transform -1 0 -7 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_1
timestamp 1644511149
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_2
timestamp 1644511149
transform 1 0 263 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_3
timestamp 1644511149
transform 1 0 426 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_4
timestamp 1644511149
transform 1 0 589 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_5
timestamp 1644511149
transform 1 0 752 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfm1sd2__example_55959141808563  sky130_fd_pr__hvdfm1sd2__example_55959141808563_6
timestamp 1644511149
transform 1 0 915 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 943 697 943 697 0 FreeSans 300 0 0 0 S
flabel comment s 780 697 780 697 0 FreeSans 300 0 0 0 D
flabel comment s 617 697 617 697 0 FreeSans 300 0 0 0 S
flabel comment s 454 697 454 697 0 FreeSans 300 0 0 0 D
flabel comment s 291 697 291 697 0 FreeSans 300 0 0 0 S
flabel comment s 128 697 128 697 0 FreeSans 300 0 0 0 D
flabel comment s -35 697 -35 697 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 8673962
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8669930
<< end >>
