magic
tech sky130B
magscale 1 2
timestamp 1644511149
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_0
timestamp 1644511149
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_1
timestamp 1644511149
transform 1 0 100 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_2
timestamp 1644511149
transform 1 0 256 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_3
timestamp 1644511149
transform 1 0 412 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_4
timestamp 1644511149
transform 1 0 568 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_5
timestamp 1644511149
transform 1 0 724 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_6
timestamp 1644511149
transform 1 0 880 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808178  sky130_fd_pr__hvdfl1sd2__example_55959141808178_7
timestamp 1644511149
transform 1 0 1036 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 1064 1491 1064 1491 0 FreeSans 300 0 0 0 D
flabel comment s 908 1491 908 1491 0 FreeSans 300 0 0 0 S
flabel comment s 752 1491 752 1491 0 FreeSans 300 0 0 0 D
flabel comment s 596 1491 596 1491 0 FreeSans 300 0 0 0 S
flabel comment s 440 1491 440 1491 0 FreeSans 300 0 0 0 D
flabel comment s 284 1491 284 1491 0 FreeSans 300 0 0 0 S
flabel comment s 128 1491 128 1491 0 FreeSans 300 0 0 0 D
flabel comment s -28 1491 -28 1491 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_END 8089926
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_START 8085760
<< end >>
