/home/drako/inventory/shuttle/caravel_tutorial/caravel_example/pdks/skywater-pdk/libraries/sky130_fd_pr/latest/cells/esd_rf_nfet_20v0_hbm/sky130_fd_pr__esd_rf_nfet_20v0_hbm_21vW60p00.spice